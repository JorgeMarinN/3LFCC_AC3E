magic
tech sky130A
timestamp 1668296084
<< metal5 >>
rect 3500 13500 6000 14000
rect 2500 13000 7000 13500
rect 1500 12500 3000 13000
rect 6500 12500 8000 13000
rect 1000 12000 2000 12500
rect 7500 12000 8500 12500
rect 1000 11500 1500 12000
rect 4500 11500 5000 12000
rect 8000 11500 8500 12000
rect 500 11000 1500 11500
rect 4000 11000 5500 11500
rect 8000 11000 9000 11500
rect 500 10000 1000 11000
rect 4500 10500 5000 11000
rect 0 7000 1000 10000
rect 8500 10000 9000 11000
rect 4000 8500 5500 9000
rect 3000 8000 6500 8500
rect 2000 7500 7500 8000
rect 8500 7000 9500 10000
rect 500 6000 1000 7000
rect 2000 6500 7500 7000
rect 2500 6000 7000 6500
rect 8500 6000 9000 7000
rect 11000 6500 12500 12500
rect 15500 6500 17000 12500
rect 19500 12000 23000 12500
rect 18500 11000 24000 12000
rect 11000 6000 13000 6500
rect 15000 6000 17000 6500
rect 18000 10500 20000 11000
rect 22500 10500 24500 11000
rect 18000 6500 19500 10500
rect 23000 10000 24500 10500
rect 23000 6500 24500 7000
rect 18000 6000 20000 6500
rect 22500 6000 24500 6500
rect 25500 6500 27000 12500
rect 30000 6500 31500 12500
rect 25500 6000 27500 6500
rect 29500 6000 31500 6500
rect 500 5500 1500 6000
rect 8000 5500 9000 6000
rect 1000 5000 1500 5500
rect 3000 5000 6500 5500
rect 8000 5000 8500 5500
rect 11500 5000 16500 6000
rect 18500 5000 24000 6000
rect 26000 5000 31000 6000
rect 1000 4500 2000 5000
rect 4000 4500 5500 5000
rect 7500 4500 8500 5000
rect 12500 4500 15500 5000
rect 19500 4500 23000 5000
rect 27000 4500 30000 5000
rect 1500 4000 3000 4500
rect 6500 4000 8000 4500
rect 2500 3500 7000 4000
rect 3500 3000 6000 3500
<< comment >>
rect -100 17000 32100 17100
rect -100 0 0 17000
rect 32000 0 32100 17000
rect -100 -100 32100 0
<< end >>
