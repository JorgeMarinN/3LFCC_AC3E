magic
tech sky130A
timestamp 1665354016
<< checkpaint >>
rect -1966 209166 39166 309166
rect -1966 168034 139166 209166
rect -1936 -1966 139166 168034
<< metal3 >>
rect 82000 173000 130000 174000
rect 82000 171300 82100 173000
rect 129900 171300 130000 173000
rect 82000 167000 130000 171300
<< via3 >>
rect 8100 171300 68900 173000
rect 82100 171300 129900 173000
<< metal4 >>
rect 8000 173000 69000 174000
rect 8000 171300 8100 173000
rect 68900 171300 69000 173000
rect 8000 167000 69000 171300
<< via4 >>
rect 8100 171300 68900 173000
rect 82100 171300 129900 173000
<< metal5 >>
rect 82000 173000 130000 174000
rect 82000 171300 82100 173000
rect 129900 171300 130000 173000
rect 82000 167000 130000 171300
use flying_cap  flying_cap_0
timestamp 1665353312
transform 1 0 30 0 1 0
box 0 0 137170 168000
use power_stage  power_stage_0
timestamp 1663434482
transform 0 -1 137200 1 0 170000
box 0 0 37200 137200
<< end >>
