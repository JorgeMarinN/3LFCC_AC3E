magic
tech sky130A
timestamp 1668306004
<< metal3 >>
rect 7000 36000 56000 42000
rect 7000 35000 7100 36000
rect 55900 35000 56000 36000
rect 7000 33000 56000 35000
<< via3 >>
rect 7100 35000 55900 36000
rect 69100 35000 129900 36000
<< metal4 >>
rect 69000 36000 130000 42000
rect 69000 35000 69100 36000
rect 129900 35000 130000 36000
rect 69000 33000 130000 35000
<< via4 >>
rect 7100 35000 55900 36000
rect 69100 35000 129900 36000
<< metal5 >>
rect 7000 36000 56000 42000
rect 7000 35000 7100 36000
rect 55900 35000 56000 36000
rect 7000 33000 56000 35000
use flying_cap  flying_cap_0
timestamp 1668303581
transform -1 0 137170 0 -1 209000
box -590 0 137170 168000
use power_stage  power_stage_0
timestamp 1663434482
transform 0 1 0 -1 0 37200
box 0 0 37200 137200
<< end >>
