magic
tech sky130A
magscale 1 2
timestamp 1665097055
<< nwell >>
rect -10 -6 1760 2244
<< mvpsubdiff >>
rect 128 -2526 152 -2458
rect 1590 -2526 1614 -2458
<< mvnsubdiff >>
rect 134 2126 164 2178
rect 1572 2126 1616 2178
<< mvpsubdiffcont >>
rect 152 -2526 1590 -2458
<< mvnsubdiffcont >>
rect 164 2126 1572 2178
<< poly >>
rect 134 -84 194 50
rect 292 -10 352 60
rect 450 -10 510 60
rect 292 -76 510 -10
rect 292 -78 352 -76
rect 450 -78 510 -76
rect 608 -10 668 60
rect 766 -10 826 60
rect 608 -76 826 -10
rect 608 -78 668 -76
rect 766 -78 826 -76
rect 924 -12 984 60
rect 1082 -12 1142 60
rect 924 -78 1142 -12
rect 1240 -12 1300 60
rect 1398 -12 1458 60
rect 1240 -78 1458 -12
rect 1556 -84 1616 60
rect 134 -486 194 -224
rect 292 -294 510 -228
rect 292 -496 352 -294
rect 450 -496 510 -294
rect 608 -294 826 -228
rect 608 -496 668 -294
rect 766 -496 826 -294
rect 924 -230 984 -228
rect 1082 -230 1142 -228
rect 924 -296 1142 -230
rect 924 -496 984 -296
rect 1082 -496 1142 -296
rect 1240 -230 1300 -228
rect 1398 -230 1458 -228
rect 1240 -296 1458 -230
rect 1240 -496 1300 -296
rect 1398 -496 1458 -296
rect 1556 -496 1616 -224
<< locali >>
rect 142 2126 164 2178
rect 1572 2126 1608 2178
rect 136 -2526 152 -2458
rect 1590 -2526 1606 -2458
<< viali >>
rect 164 2126 1572 2178
rect 152 -2524 1590 -2458
<< metal1 >>
rect 44 2178 1706 2184
rect 44 2126 164 2178
rect 1572 2126 1706 2178
rect 44 2120 1706 2126
rect 68 2048 102 2120
rect 384 2048 418 2120
rect 700 2048 734 2120
rect 1016 2048 1050 2120
rect 1332 2048 1366 2120
rect 1648 2048 1682 2120
rect 126 -70 136 -18
rect 188 -70 198 -18
rect 226 -128 260 72
rect 364 -70 374 -18
rect 426 -70 436 -18
rect 542 -128 576 72
rect 678 -70 688 -18
rect 740 -70 750 -18
rect 858 -128 892 72
rect 996 -70 1006 -18
rect 1058 -70 1068 -18
rect 1174 -128 1208 72
rect 1310 -70 1320 -18
rect 1372 -70 1382 -18
rect 1490 -128 1524 72
rect 1554 -70 1564 -18
rect 1616 -70 1626 -18
rect 206 -180 216 -128
rect 268 -180 278 -128
rect 522 -180 532 -128
rect 584 -180 594 -128
rect 840 -180 850 -128
rect 902 -180 912 -128
rect 1156 -180 1166 -128
rect 1218 -180 1228 -128
rect 1472 -180 1482 -128
rect 1534 -180 1544 -128
rect 126 -288 136 -236
rect 188 -288 198 -236
rect 226 -508 260 -180
rect 364 -288 374 -236
rect 426 -288 436 -236
rect 542 -508 576 -180
rect 678 -288 688 -236
rect 740 -288 750 -236
rect 858 -508 892 -180
rect 996 -288 1006 -236
rect 1058 -288 1068 -236
rect 1174 -508 1208 -180
rect 1310 -288 1320 -236
rect 1372 -288 1382 -236
rect 1490 -508 1524 -180
rect 1554 -288 1564 -236
rect 1616 -288 1626 -236
rect 68 -2426 102 -2352
rect 384 -2426 418 -2352
rect 700 -2426 734 -2352
rect 1016 -2426 1050 -2352
rect 1332 -2426 1366 -2352
rect 1648 -2426 1682 -2352
rect 68 -2458 1682 -2426
rect 68 -2524 152 -2458
rect 1590 -2524 1682 -2458
rect 68 -2532 1682 -2524
<< via1 >>
rect 136 -70 188 -18
rect 374 -70 426 -18
rect 688 -70 740 -18
rect 1006 -70 1058 -18
rect 1320 -70 1372 -18
rect 1564 -70 1616 -18
rect 216 -180 268 -128
rect 532 -180 584 -128
rect 850 -180 902 -128
rect 1166 -180 1218 -128
rect 1482 -180 1534 -128
rect 136 -288 188 -236
rect 374 -288 426 -236
rect 688 -288 740 -236
rect 1006 -288 1058 -236
rect 1320 -288 1372 -236
rect 1564 -288 1616 -236
<< metal2 >>
rect 136 -18 1758 -4
rect 188 -70 374 -18
rect 426 -70 688 -18
rect 740 -70 1006 -18
rect 1058 -70 1320 -18
rect 1372 -70 1564 -18
rect 1616 -70 1758 -18
rect 136 -84 1758 -70
rect -14 -128 1756 -114
rect -14 -180 216 -128
rect 268 -180 532 -128
rect 584 -180 850 -128
rect 902 -180 1166 -128
rect 1218 -180 1482 -128
rect 1534 -180 1756 -128
rect -14 -194 1756 -180
rect -12 -236 1758 -224
rect -12 -288 136 -236
rect 188 -288 374 -236
rect 426 -288 688 -236
rect 740 -288 1006 -236
rect 1058 -288 1320 -236
rect 1372 -288 1564 -236
rect 1616 -288 1758 -236
rect -12 -302 1758 -288
use cont_poly_min  cont_poly_min_0
timestamp 1663264347
transform 1 0 1591 0 1 -111
box -33 33 33 99
use cont_poly_min  cont_poly_min_1
timestamp 1663264347
transform 1 0 163 0 1 -111
box -33 33 33 99
use cont_poly_min  cont_poly_min_2
timestamp 1663264347
transform 1 0 401 0 1 -109
box -33 33 33 99
use cont_poly_min  cont_poly_min_3
timestamp 1663264347
transform 1 0 715 0 1 -109
box -33 33 33 99
use cont_poly_min  cont_poly_min_4
timestamp 1663264347
transform 1 0 1033 0 1 -111
box -33 33 33 99
use cont_poly_min  cont_poly_min_5
timestamp 1663264347
transform 1 0 1347 0 1 -111
box -33 33 33 99
use cont_poly_min  cont_poly_min_6
timestamp 1663264347
transform 1 0 163 0 1 -329
box -33 33 33 99
use cont_poly_min  cont_poly_min_7
timestamp 1663264347
transform 1 0 401 0 1 -327
box -33 33 33 99
use cont_poly_min  cont_poly_min_8
timestamp 1663264347
transform 1 0 715 0 1 -327
box -33 33 33 99
use cont_poly_min  cont_poly_min_9
timestamp 1663264347
transform 1 0 1033 0 1 -329
box -33 33 33 99
use cont_poly_min  cont_poly_min_10
timestamp 1663264347
transform 1 0 1347 0 1 -329
box -33 33 33 99
use cont_poly_min  cont_poly_min_11
timestamp 1663264347
transform 1 0 1591 0 1 -329
box -33 33 33 99
use sky130_fd_pr__nfet_g5v0d10v5_PVZBWB  sky130_fd_pr__nfet_g5v0d10v5_PVZBWB_0
timestamp 1663361110
transform 1 0 875 0 1 -1366
box -819 -1026 819 1026
use sky130_fd_pr__pfet_g5v0d10v5_VEZS85  sky130_fd_pr__pfet_g5v0d10v5_VEZS85_0
timestamp 1663361110
transform 1 0 875 0 1 1060
box -885 -1066 885 1066
<< labels >>
rlabel metal1 44 2178 1706 2184 1 VH
rlabel metal2 1534 -194 1756 -114 1 OUT
rlabel metal1 68 -2532 1682 -2526 1 GND
rlabel space -12 -84 136 -4 1 A
rlabel metal2 -12 -302 136 -224 1 B
<< end >>
