magic
tech sky130A
timestamp 1667696568
<< metal4 >>
rect 0 45759 28150 45779
rect 0 41449 20 45759
rect 4330 45743 28150 45759
rect 4330 41465 23836 45743
rect 28114 41465 28150 45743
rect 4330 41449 28150 41465
rect 0 41429 28150 41449
<< via4 >>
rect 20 41449 4330 45759
rect 23836 41465 28114 45743
<< metal5 >>
rect 0 65229 75529 69579
rect 5950 59279 69579 63629
rect 0 45759 4350 45779
rect 0 41449 20 45759
rect 4330 41449 4350 45759
rect 0 41429 4350 41449
rect 5950 4350 10300 59279
rect 11900 53329 63629 57679
rect 11900 10300 16250 53329
rect 17850 47379 57679 51729
rect 17850 16250 22200 47379
rect 23800 45743 28150 45779
rect 23800 41465 23836 45743
rect 28114 41465 28150 45743
rect 23800 22200 28150 41465
rect 53329 22200 57679 47379
rect 23800 17850 57679 22200
rect 59279 16250 63629 53329
rect 17850 11900 63629 16250
rect 65229 10300 69579 59279
rect 11900 5950 69579 10300
rect 71179 4350 75529 65229
rect 5950 0 75529 4350
<< end >>
