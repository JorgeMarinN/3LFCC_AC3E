magic
tech sky130A
timestamp 1666628647
<< metal4 >>
rect 92339 104019 105379 104080
rect 92339 91101 92400 104019
rect 105318 91101 105379 104019
rect 92339 36959 105379 91101
<< via4 >>
rect 92400 91101 105318 104019
<< metal5 >>
rect 50000 133380 146420 146420
rect 50000 119699 132740 132740
rect 50000 63040 63040 119699
rect 63680 106019 119059 119059
rect 63680 76720 76720 106019
rect 77360 104019 105379 105379
rect 77360 92339 92400 104019
rect 77360 90400 90400 92339
rect 92339 91101 92400 92339
rect 105318 91101 105379 104019
rect 92339 91040 105379 91101
rect 106019 90400 119059 106019
rect 77360 77360 119059 90400
rect 119699 76720 132740 119699
rect 63680 63680 132740 76720
rect 133380 63040 146420 133380
rect 50000 50000 146420 63040
<< end >>
