magic
tech sky130A
timestamp 1662490911
<< metal2 >>
rect 3000 131460 5200 132000
rect 3000 131270 4960 131460
rect 3000 130400 5200 131270
rect 3000 66960 5740 67200
rect 5930 66960 6800 67200
rect 3000 65600 6800 66960
rect 3000 56640 6800 58000
rect 3000 56400 5740 56640
rect 5930 56400 6800 56640
rect 3000 5749 4962 6000
rect 3000 5200 5300 5749
<< metal3 >>
rect 6000 133000 36000 136000
rect 3400 130100 4400 131039
rect 1000 104000 4000 130000
rect 33000 106000 36000 133000
rect 1000 95000 31000 104000
rect 1000 68000 4000 95000
rect 6161 66000 7100 66400
rect 33000 66000 36000 93000
rect 6161 65400 36000 66000
rect 7000 63000 36000 65400
rect 7000 61000 27000 63000
rect 7000 58200 30000 61000
rect 6161 58000 30000 58200
rect 6161 57200 7100 58000
rect 1000 35000 4000 56000
rect 27000 37000 30000 58000
rect 1000 27000 25000 35000
rect 1000 7100 4000 27000
rect 1000 7000 4400 7100
rect 3400 6161 4400 7000
rect 27000 4000 30000 25000
rect 6000 1000 30000 4000
<< metal4 >>
rect 6000 133000 36000 136000
rect 3400 130100 4400 131039
rect 1000 104000 4000 130000
rect 33000 106000 36000 133000
rect 1000 95000 31000 104000
rect 1000 68000 4000 95000
rect 6161 66000 7100 66400
rect 33000 66000 36000 93000
rect 6161 65400 36000 66000
rect 7000 63000 36000 65400
rect 7000 61000 27000 63000
rect 7000 58200 30000 61000
rect 6161 58000 30000 58200
rect 6161 57200 7100 58000
rect 1000 35000 4000 56000
rect 27000 37000 30000 58000
rect 1000 27000 25000 35000
rect 1000 7100 4000 27000
rect 1000 7000 4400 7100
rect 3400 6161 4400 7000
rect 27000 4000 30000 25000
rect 6000 1000 30000 4000
<< metal5 >>
rect 6000 133000 36000 136000
rect 3400 130100 4400 131039
rect 1000 104000 4000 130000
rect 33000 106000 36000 133000
rect 1000 95000 31000 104000
rect 1000 68000 4000 95000
rect 6161 66000 7100 66400
rect 33000 66000 36000 93000
rect 6161 65400 36000 66000
rect 7000 63000 36000 65400
rect 7000 61000 27000 63000
rect 7000 58200 30000 61000
rect 6161 58000 30000 58200
rect 6161 57200 7100 58000
rect 1000 35000 4000 56000
rect 27000 37000 30000 58000
rect 1000 27000 25000 35000
rect 1000 7100 4000 27000
rect 1000 7000 4400 7100
rect 3400 6161 4400 7000
rect 27000 4000 30000 25000
rect 6000 1000 30000 4000
use nmos_waffle_36x36  nmos_waffle_36x36_0
timestamp 1661896674
transform 1 0 5400 0 1 5400
box -5400 -5400 25200 25200
use nmos_waffle_36x36  nmos_waffle_36x36_1
timestamp 1661896674
transform 0 1 5400 -1 0 56200
box -5400 -5400 25200 25200
use pmos_waffle_48x48  pmos_waffle_48x48_0
timestamp 1661896674
transform 0 1 5400 1 0 67400
box -5400 -5400 31800 31800
use pmos_waffle_48x48  pmos_waffle_48x48_1
timestamp 1661896674
transform 1 0 5400 0 -1 131800
box -5400 -5400 31800 31800
<< end >>
