magic
tech sky130A
timestamp 1668197163
<< error_p >>
rect 496 19202 502 19217
rect 612 19202 1038 19204
rect 1148 19202 1154 19217
rect 1162 19202 1588 19204
rect 1596 19202 1602 19217
rect 1712 19202 2138 19204
rect 2248 19202 2254 19217
rect 2262 19202 2688 19204
rect 2696 19202 2702 19217
rect 2812 19202 3238 19204
rect 3348 19202 3354 19217
rect 3362 19202 3788 19204
rect 3796 19202 3802 19217
rect 3912 19202 4338 19204
rect 4448 19202 4454 19217
rect 4462 19202 4888 19204
rect 4896 19202 4902 19217
rect 5012 19202 5438 19204
rect 5548 19202 5554 19217
rect 5562 19202 5988 19204
rect 5996 19202 6002 19217
rect 6112 19202 6538 19204
rect 6648 19202 6654 19217
rect 6662 19202 7088 19204
rect 7096 19202 7102 19217
rect 7212 19202 7638 19204
rect 7748 19202 7754 19217
rect 7762 19202 8188 19204
rect 8196 19202 8202 19217
rect 8312 19202 8738 19204
rect 8848 19202 8854 19217
rect 8862 19202 9288 19204
rect 9296 19202 9302 19217
rect 9412 19202 9838 19204
rect 9948 19202 9954 19217
rect 9962 19202 10388 19204
rect 10396 19202 10402 19217
rect 10512 19202 10938 19204
rect 11048 19202 11054 19217
rect 11062 19202 11488 19204
rect 11496 19202 11502 19217
rect 11612 19202 12038 19204
rect 12148 19202 12154 19217
rect 12162 19202 12588 19204
rect 12596 19202 12602 19217
rect 12712 19202 13138 19204
rect 13248 19202 13254 19217
rect 13262 19202 13688 19204
rect 13696 19202 13702 19217
rect 13812 19202 14238 19204
rect 14348 19202 14354 19217
rect 14362 19202 14788 19204
rect 14796 19202 14802 19217
rect 14912 19202 15338 19204
rect 15448 19202 15454 19217
rect 15462 19202 15888 19204
rect 15896 19202 15902 19217
rect 16012 19202 16438 19204
rect 16548 19202 16554 19217
rect 16562 19202 16988 19204
rect 16996 19202 17002 19217
rect 17112 19202 17538 19204
rect 17648 19202 17654 19217
rect 17662 19202 18088 19204
rect 18096 19202 18102 19217
rect 18212 19202 18638 19204
rect 18748 19202 18754 19217
rect 19170 19204 19194 19224
rect 18762 19202 19194 19204
rect 19196 19202 19217 19217
rect 19170 19200 19194 19202
rect 19202 19196 19217 19202
rect 628 19172 885 19195
rect 1178 19172 1435 19195
rect 1728 19172 1985 19195
rect 2278 19172 2535 19195
rect 2828 19172 3085 19195
rect 3378 19172 3635 19195
rect 3928 19172 4185 19195
rect 4478 19172 4735 19195
rect 5028 19172 5285 19195
rect 5578 19172 5835 19195
rect 6128 19172 6385 19195
rect 6678 19172 6935 19195
rect 7228 19172 7485 19195
rect 7778 19172 8035 19195
rect 8328 19172 8585 19195
rect 8878 19172 9135 19195
rect 9428 19172 9685 19195
rect 9978 19172 10235 19195
rect 10528 19172 10785 19195
rect 11078 19172 11335 19195
rect 11628 19172 11885 19195
rect 12178 19172 12435 19195
rect 12728 19172 12985 19195
rect 13278 19172 13535 19195
rect 13828 19172 14085 19195
rect 14378 19172 14635 19195
rect 14928 19172 15185 19195
rect 15478 19172 15735 19195
rect 16028 19172 16285 19195
rect 16578 19172 16835 19195
rect 17128 19172 17385 19195
rect 17678 19172 17935 19195
rect 18228 19172 18485 19195
rect 18778 19172 19035 19195
rect 19200 19188 19208 19194
rect 19200 19186 19204 19188
rect 605 19035 609 19172
rect 784 19075 885 19172
rect 765 19035 885 19075
rect 1155 19035 1159 19172
rect 1334 19075 1435 19172
rect 1315 19035 1435 19075
rect 1705 19035 1709 19172
rect 1884 19075 1985 19172
rect 1865 19035 1985 19075
rect 2255 19035 2259 19172
rect 2434 19075 2535 19172
rect 2415 19035 2535 19075
rect 2805 19035 2809 19172
rect 2984 19075 3085 19172
rect 2965 19035 3085 19075
rect 3355 19035 3359 19172
rect 3534 19075 3635 19172
rect 3515 19035 3635 19075
rect 3905 19035 3909 19172
rect 4084 19075 4185 19172
rect 4065 19035 4185 19075
rect 4455 19035 4459 19172
rect 4634 19075 4735 19172
rect 4615 19035 4735 19075
rect 5005 19035 5009 19172
rect 5184 19075 5285 19172
rect 5165 19035 5285 19075
rect 5555 19035 5559 19172
rect 5734 19075 5835 19172
rect 5715 19035 5835 19075
rect 6105 19035 6109 19172
rect 6284 19075 6385 19172
rect 6265 19035 6385 19075
rect 6655 19035 6659 19172
rect 6834 19075 6935 19172
rect 6815 19035 6935 19075
rect 7205 19035 7209 19172
rect 7384 19075 7485 19172
rect 7365 19035 7485 19075
rect 7755 19035 7759 19172
rect 7934 19075 8035 19172
rect 7915 19035 8035 19075
rect 8305 19035 8309 19172
rect 8484 19075 8585 19172
rect 8465 19035 8585 19075
rect 8855 19035 8859 19172
rect 9034 19075 9135 19172
rect 9015 19035 9135 19075
rect 9405 19035 9409 19172
rect 9584 19075 9685 19172
rect 9565 19035 9685 19075
rect 9955 19035 9959 19172
rect 10134 19075 10235 19172
rect 10115 19035 10235 19075
rect 10505 19035 10509 19172
rect 10684 19075 10785 19172
rect 10665 19035 10785 19075
rect 11055 19035 11059 19172
rect 11234 19075 11335 19172
rect 11215 19035 11335 19075
rect 11605 19035 11609 19172
rect 11784 19075 11885 19172
rect 11765 19035 11885 19075
rect 12155 19035 12159 19172
rect 12334 19075 12435 19172
rect 12315 19035 12435 19075
rect 12705 19035 12709 19172
rect 12884 19075 12985 19172
rect 12865 19035 12985 19075
rect 13255 19035 13259 19172
rect 13434 19075 13535 19172
rect 13415 19035 13535 19075
rect 13805 19035 13809 19172
rect 13984 19075 14085 19172
rect 13965 19035 14085 19075
rect 14355 19035 14359 19172
rect 14534 19075 14635 19172
rect 14515 19035 14635 19075
rect 14905 19035 14909 19172
rect 15084 19075 15185 19172
rect 15065 19035 15185 19075
rect 15455 19035 15459 19172
rect 15634 19075 15735 19172
rect 15615 19035 15735 19075
rect 16005 19035 16009 19172
rect 16184 19075 16285 19172
rect 16165 19035 16285 19075
rect 16555 19035 16559 19172
rect 16734 19075 16835 19172
rect 16715 19035 16835 19075
rect 17105 19035 17109 19172
rect 17284 19075 17385 19172
rect 17265 19035 17385 19075
rect 17655 19035 17659 19172
rect 17834 19075 17935 19172
rect 17815 19035 17935 19075
rect 18205 19035 18209 19172
rect 18384 19075 18485 19172
rect 18365 19035 18485 19075
rect 18755 19035 18759 19172
rect 18934 19075 19035 19172
rect 18915 19035 19035 19075
rect 725 19028 842 19035
rect 885 19028 1045 19035
rect 725 18922 808 19028
rect 842 18922 1045 19028
rect 725 18915 765 18922
rect 808 18915 1045 18922
rect 1275 19028 1392 19035
rect 1435 19028 1595 19035
rect 1275 18922 1358 19028
rect 1392 18922 1595 19028
rect 1275 18915 1315 18922
rect 1358 18915 1595 18922
rect 1825 19028 1942 19035
rect 1985 19028 2145 19035
rect 1825 18922 1908 19028
rect 1942 18922 2145 19028
rect 1825 18915 1865 18922
rect 1908 18915 2145 18922
rect 2375 19028 2492 19035
rect 2535 19028 2695 19035
rect 2375 18922 2458 19028
rect 2492 18922 2695 19028
rect 2375 18915 2415 18922
rect 2458 18915 2695 18922
rect 2925 19028 3042 19035
rect 3085 19028 3245 19035
rect 2925 18922 3008 19028
rect 3042 18922 3245 19028
rect 2925 18915 2965 18922
rect 3008 18915 3245 18922
rect 3475 19028 3592 19035
rect 3635 19028 3795 19035
rect 3475 18922 3558 19028
rect 3592 18922 3795 19028
rect 3475 18915 3515 18922
rect 3558 18915 3795 18922
rect 4025 19028 4142 19035
rect 4185 19028 4345 19035
rect 4025 18922 4108 19028
rect 4142 18922 4345 19028
rect 4025 18915 4065 18922
rect 4108 18915 4345 18922
rect 4575 19028 4692 19035
rect 4735 19028 4895 19035
rect 4575 18922 4658 19028
rect 4692 18922 4895 19028
rect 4575 18915 4615 18922
rect 4658 18915 4895 18922
rect 5125 19028 5242 19035
rect 5285 19028 5445 19035
rect 5125 18922 5208 19028
rect 5242 18922 5445 19028
rect 5125 18915 5165 18922
rect 5208 18915 5445 18922
rect 5675 19028 5792 19035
rect 5835 19028 5995 19035
rect 5675 18922 5758 19028
rect 5792 18922 5995 19028
rect 5675 18915 5715 18922
rect 5758 18915 5995 18922
rect 6225 19028 6342 19035
rect 6385 19028 6545 19035
rect 6225 18922 6308 19028
rect 6342 18922 6545 19028
rect 6225 18915 6265 18922
rect 6308 18915 6545 18922
rect 6775 19028 6892 19035
rect 6935 19028 7095 19035
rect 6775 18922 6858 19028
rect 6892 18922 7095 19028
rect 6775 18915 6815 18922
rect 6858 18915 7095 18922
rect 7325 19028 7442 19035
rect 7485 19028 7645 19035
rect 7325 18922 7408 19028
rect 7442 18922 7645 19028
rect 7325 18915 7365 18922
rect 7408 18915 7645 18922
rect 7875 19028 7992 19035
rect 8035 19028 8195 19035
rect 7875 18922 7958 19028
rect 7992 18922 8195 19028
rect 7875 18915 7915 18922
rect 7958 18915 8195 18922
rect 8425 19028 8542 19035
rect 8585 19028 8745 19035
rect 8425 18922 8508 19028
rect 8542 18922 8745 19028
rect 8425 18915 8465 18922
rect 8508 18915 8745 18922
rect 8975 19028 9092 19035
rect 9135 19028 9295 19035
rect 8975 18922 9058 19028
rect 9092 18922 9295 19028
rect 8975 18915 9015 18922
rect 9058 18915 9295 18922
rect 9525 19028 9642 19035
rect 9685 19028 9845 19035
rect 9525 18922 9608 19028
rect 9642 18922 9845 19028
rect 9525 18915 9565 18922
rect 9608 18915 9845 18922
rect 10075 19028 10192 19035
rect 10235 19028 10395 19035
rect 10075 18922 10158 19028
rect 10192 18922 10395 19028
rect 10075 18915 10115 18922
rect 10158 18915 10395 18922
rect 10625 19028 10742 19035
rect 10785 19028 10945 19035
rect 10625 18922 10708 19028
rect 10742 18922 10945 19028
rect 10625 18915 10665 18922
rect 10708 18915 10945 18922
rect 11175 19028 11292 19035
rect 11335 19028 11495 19035
rect 11175 18922 11258 19028
rect 11292 18922 11495 19028
rect 11175 18915 11215 18922
rect 11258 18915 11495 18922
rect 11725 19028 11842 19035
rect 11885 19028 12045 19035
rect 11725 18922 11808 19028
rect 11842 18922 12045 19028
rect 11725 18915 11765 18922
rect 11808 18915 12045 18922
rect 12275 19028 12392 19035
rect 12435 19028 12595 19035
rect 12275 18922 12358 19028
rect 12392 18922 12595 19028
rect 12275 18915 12315 18922
rect 12358 18915 12595 18922
rect 12825 19028 12942 19035
rect 12985 19028 13145 19035
rect 12825 18922 12908 19028
rect 12942 18922 13145 19028
rect 12825 18915 12865 18922
rect 12908 18915 13145 18922
rect 13375 19028 13492 19035
rect 13535 19028 13695 19035
rect 13375 18922 13458 19028
rect 13492 18922 13695 19028
rect 13375 18915 13415 18922
rect 13458 18915 13695 18922
rect 13925 19028 14042 19035
rect 14085 19028 14245 19035
rect 13925 18922 14008 19028
rect 14042 18922 14245 19028
rect 13925 18915 13965 18922
rect 14008 18915 14245 18922
rect 14475 19028 14592 19035
rect 14635 19028 14795 19035
rect 14475 18922 14558 19028
rect 14592 18922 14795 19028
rect 14475 18915 14515 18922
rect 14558 18915 14795 18922
rect 15025 19028 15142 19035
rect 15185 19028 15345 19035
rect 15025 18922 15108 19028
rect 15142 18922 15345 19028
rect 15025 18915 15065 18922
rect 15108 18915 15345 18922
rect 15575 19028 15692 19035
rect 15735 19028 15895 19035
rect 15575 18922 15658 19028
rect 15692 18922 15895 19028
rect 15575 18915 15615 18922
rect 15658 18915 15895 18922
rect 16125 19028 16242 19035
rect 16285 19028 16445 19035
rect 16125 18922 16208 19028
rect 16242 18922 16445 19028
rect 16125 18915 16165 18922
rect 16208 18915 16445 18922
rect 16675 19028 16792 19035
rect 16835 19028 16995 19035
rect 16675 18922 16758 19028
rect 16792 18922 16995 19028
rect 16675 18915 16715 18922
rect 16758 18915 16995 18922
rect 17225 19028 17342 19035
rect 17385 19028 17545 19035
rect 17225 18922 17308 19028
rect 17342 18922 17545 19028
rect 17225 18915 17265 18922
rect 17308 18915 17545 18922
rect 17775 19028 17892 19035
rect 17935 19028 18095 19035
rect 17775 18922 17858 19028
rect 17892 18922 18095 19028
rect 17775 18915 17815 18922
rect 17858 18915 18095 18922
rect 18325 19028 18442 19035
rect 18485 19028 18645 19035
rect 18325 18922 18408 19028
rect 18442 18922 18645 19028
rect 18325 18915 18365 18922
rect 18408 18915 18645 18922
rect 18875 19028 18992 19035
rect 19035 19028 19195 19035
rect 18875 18922 18958 19028
rect 18992 18922 19195 19028
rect 18875 18915 18915 18922
rect 18958 18915 19195 18922
rect 765 18875 885 18915
rect 1315 18875 1435 18915
rect 1865 18875 1985 18915
rect 2415 18875 2535 18915
rect 2965 18875 3085 18915
rect 3515 18875 3635 18915
rect 4065 18875 4185 18915
rect 4615 18875 4735 18915
rect 5165 18875 5285 18915
rect 5715 18875 5835 18915
rect 6265 18875 6385 18915
rect 6815 18875 6935 18915
rect 7365 18875 7485 18915
rect 7915 18875 8035 18915
rect 8465 18875 8585 18915
rect 9015 18875 9135 18915
rect 9565 18875 9685 18915
rect 10115 18875 10235 18915
rect 10665 18875 10785 18915
rect 11215 18875 11335 18915
rect 11765 18875 11885 18915
rect 12315 18875 12435 18915
rect 12865 18875 12985 18915
rect 13415 18875 13535 18915
rect 13965 18875 14085 18915
rect 14515 18875 14635 18915
rect 15065 18875 15185 18915
rect 15615 18875 15735 18915
rect 16165 18875 16285 18915
rect 16715 18875 16835 18915
rect 17265 18875 17385 18915
rect 17815 18875 17935 18915
rect 18365 18875 18485 18915
rect 18915 18875 19035 18915
rect 19185 18754 19200 18771
rect 19202 18762 19204 19186
rect 19202 18748 19217 18754
rect 500 18675 507 18725
rect 500 18239 525 18640
rect 628 18622 885 18645
rect 1178 18622 1435 18645
rect 1728 18622 1985 18645
rect 2278 18622 2535 18645
rect 2828 18622 3085 18645
rect 3378 18622 3635 18645
rect 3928 18622 4185 18645
rect 4478 18622 4735 18645
rect 5028 18622 5285 18645
rect 5578 18622 5835 18645
rect 6128 18622 6385 18645
rect 6678 18622 6935 18645
rect 7228 18622 7485 18645
rect 7778 18622 8035 18645
rect 8328 18622 8585 18645
rect 8878 18622 9135 18645
rect 9428 18622 9685 18645
rect 9978 18622 10235 18645
rect 10528 18622 10785 18645
rect 11078 18622 11335 18645
rect 11628 18622 11885 18645
rect 12178 18622 12435 18645
rect 12728 18622 12985 18645
rect 13278 18622 13535 18645
rect 13828 18622 14085 18645
rect 14378 18622 14635 18645
rect 14928 18622 15185 18645
rect 15478 18622 15735 18645
rect 16028 18622 16285 18645
rect 16578 18622 16835 18645
rect 17128 18622 17385 18645
rect 17678 18622 17935 18645
rect 18228 18622 18485 18645
rect 18778 18622 19035 18645
rect 605 18485 609 18622
rect 784 18525 885 18622
rect 765 18485 885 18525
rect 1155 18485 1159 18622
rect 1334 18525 1435 18622
rect 1315 18485 1435 18525
rect 1705 18485 1709 18622
rect 1884 18525 1985 18622
rect 1865 18485 1985 18525
rect 2255 18485 2259 18622
rect 2434 18525 2535 18622
rect 2415 18485 2535 18525
rect 2805 18485 2809 18622
rect 2984 18525 3085 18622
rect 2965 18485 3085 18525
rect 3355 18485 3359 18622
rect 3534 18525 3635 18622
rect 3515 18485 3635 18525
rect 3905 18485 3909 18622
rect 4084 18525 4185 18622
rect 4065 18485 4185 18525
rect 4455 18485 4459 18622
rect 4634 18525 4735 18622
rect 4615 18485 4735 18525
rect 5005 18485 5009 18622
rect 5184 18525 5285 18622
rect 5165 18485 5285 18525
rect 5555 18485 5559 18622
rect 5734 18525 5835 18622
rect 5715 18485 5835 18525
rect 6105 18485 6109 18622
rect 6284 18525 6385 18622
rect 6265 18485 6385 18525
rect 6655 18485 6659 18622
rect 6834 18525 6935 18622
rect 6815 18485 6935 18525
rect 7205 18485 7209 18622
rect 7384 18525 7485 18622
rect 7365 18485 7485 18525
rect 7755 18485 7759 18622
rect 7934 18525 8035 18622
rect 7915 18485 8035 18525
rect 8305 18485 8309 18622
rect 8484 18525 8585 18622
rect 8465 18485 8585 18525
rect 8855 18485 8859 18622
rect 9034 18525 9135 18622
rect 9015 18485 9135 18525
rect 9405 18485 9409 18622
rect 9584 18525 9685 18622
rect 9565 18485 9685 18525
rect 9955 18485 9959 18622
rect 10134 18525 10235 18622
rect 10115 18485 10235 18525
rect 10505 18485 10509 18622
rect 10684 18525 10785 18622
rect 10665 18485 10785 18525
rect 11055 18485 11059 18622
rect 11234 18525 11335 18622
rect 11215 18485 11335 18525
rect 11605 18485 11609 18622
rect 11784 18525 11885 18622
rect 11765 18485 11885 18525
rect 12155 18485 12159 18622
rect 12334 18525 12435 18622
rect 12315 18485 12435 18525
rect 12705 18485 12709 18622
rect 12884 18525 12985 18622
rect 12865 18485 12985 18525
rect 13255 18485 13259 18622
rect 13434 18525 13535 18622
rect 13415 18485 13535 18525
rect 13805 18485 13809 18622
rect 13984 18525 14085 18622
rect 13965 18485 14085 18525
rect 14355 18485 14359 18622
rect 14534 18525 14635 18622
rect 14515 18485 14635 18525
rect 14905 18485 14909 18622
rect 15084 18525 15185 18622
rect 15065 18485 15185 18525
rect 15455 18485 15459 18622
rect 15634 18525 15735 18622
rect 15615 18485 15735 18525
rect 16005 18485 16009 18622
rect 16184 18525 16285 18622
rect 16165 18485 16285 18525
rect 16555 18485 16559 18622
rect 16734 18525 16835 18622
rect 16715 18485 16835 18525
rect 17105 18485 17109 18622
rect 17284 18525 17385 18622
rect 17265 18485 17385 18525
rect 17655 18485 17659 18622
rect 17834 18525 17935 18622
rect 17815 18485 17935 18525
rect 18205 18485 18209 18622
rect 18384 18525 18485 18622
rect 18365 18485 18485 18525
rect 18755 18485 18759 18622
rect 18934 18525 19035 18622
rect 18915 18485 19035 18525
rect 725 18478 842 18485
rect 885 18478 1045 18485
rect 725 18372 808 18478
rect 842 18372 1045 18478
rect 725 18365 765 18372
rect 808 18365 1045 18372
rect 1275 18478 1392 18485
rect 1435 18478 1595 18485
rect 1275 18372 1358 18478
rect 1392 18372 1595 18478
rect 1275 18365 1315 18372
rect 1358 18365 1595 18372
rect 1825 18478 1942 18485
rect 1985 18478 2145 18485
rect 1825 18372 1908 18478
rect 1942 18372 2145 18478
rect 1825 18365 1865 18372
rect 1908 18365 2145 18372
rect 2375 18478 2492 18485
rect 2535 18478 2695 18485
rect 2375 18372 2458 18478
rect 2492 18372 2695 18478
rect 2375 18365 2415 18372
rect 2458 18365 2695 18372
rect 2925 18478 3042 18485
rect 3085 18478 3245 18485
rect 2925 18372 3008 18478
rect 3042 18372 3245 18478
rect 2925 18365 2965 18372
rect 3008 18365 3245 18372
rect 3475 18478 3592 18485
rect 3635 18478 3795 18485
rect 3475 18372 3558 18478
rect 3592 18372 3795 18478
rect 3475 18365 3515 18372
rect 3558 18365 3795 18372
rect 4025 18478 4142 18485
rect 4185 18478 4345 18485
rect 4025 18372 4108 18478
rect 4142 18372 4345 18478
rect 4025 18365 4065 18372
rect 4108 18365 4345 18372
rect 4575 18478 4692 18485
rect 4735 18478 4895 18485
rect 4575 18372 4658 18478
rect 4692 18372 4895 18478
rect 4575 18365 4615 18372
rect 4658 18365 4895 18372
rect 5125 18478 5242 18485
rect 5285 18478 5445 18485
rect 5125 18372 5208 18478
rect 5242 18372 5445 18478
rect 5125 18365 5165 18372
rect 5208 18365 5445 18372
rect 5675 18478 5792 18485
rect 5835 18478 5995 18485
rect 5675 18372 5758 18478
rect 5792 18372 5995 18478
rect 5675 18365 5715 18372
rect 5758 18365 5995 18372
rect 6225 18478 6342 18485
rect 6385 18478 6545 18485
rect 6225 18372 6308 18478
rect 6342 18372 6545 18478
rect 6225 18365 6265 18372
rect 6308 18365 6545 18372
rect 6775 18478 6892 18485
rect 6935 18478 7095 18485
rect 6775 18372 6858 18478
rect 6892 18372 7095 18478
rect 6775 18365 6815 18372
rect 6858 18365 7095 18372
rect 7325 18478 7442 18485
rect 7485 18478 7645 18485
rect 7325 18372 7408 18478
rect 7442 18372 7645 18478
rect 7325 18365 7365 18372
rect 7408 18365 7645 18372
rect 7875 18478 7992 18485
rect 8035 18478 8195 18485
rect 7875 18372 7958 18478
rect 7992 18372 8195 18478
rect 7875 18365 7915 18372
rect 7958 18365 8195 18372
rect 8425 18478 8542 18485
rect 8585 18478 8745 18485
rect 8425 18372 8508 18478
rect 8542 18372 8745 18478
rect 8425 18365 8465 18372
rect 8508 18365 8745 18372
rect 8975 18478 9092 18485
rect 9135 18478 9295 18485
rect 8975 18372 9058 18478
rect 9092 18372 9295 18478
rect 8975 18365 9015 18372
rect 9058 18365 9295 18372
rect 9525 18478 9642 18485
rect 9685 18478 9845 18485
rect 9525 18372 9608 18478
rect 9642 18372 9845 18478
rect 9525 18365 9565 18372
rect 9608 18365 9845 18372
rect 10075 18478 10192 18485
rect 10235 18478 10395 18485
rect 10075 18372 10158 18478
rect 10192 18372 10395 18478
rect 10075 18365 10115 18372
rect 10158 18365 10395 18372
rect 10625 18478 10742 18485
rect 10785 18478 10945 18485
rect 10625 18372 10708 18478
rect 10742 18372 10945 18478
rect 10625 18365 10665 18372
rect 10708 18365 10945 18372
rect 11175 18478 11292 18485
rect 11335 18478 11495 18485
rect 11175 18372 11258 18478
rect 11292 18372 11495 18478
rect 11175 18365 11215 18372
rect 11258 18365 11495 18372
rect 11725 18478 11842 18485
rect 11885 18478 12045 18485
rect 11725 18372 11808 18478
rect 11842 18372 12045 18478
rect 11725 18365 11765 18372
rect 11808 18365 12045 18372
rect 12275 18478 12392 18485
rect 12435 18478 12595 18485
rect 12275 18372 12358 18478
rect 12392 18372 12595 18478
rect 12275 18365 12315 18372
rect 12358 18365 12595 18372
rect 12825 18478 12942 18485
rect 12985 18478 13145 18485
rect 12825 18372 12908 18478
rect 12942 18372 13145 18478
rect 12825 18365 12865 18372
rect 12908 18365 13145 18372
rect 13375 18478 13492 18485
rect 13535 18478 13695 18485
rect 13375 18372 13458 18478
rect 13492 18372 13695 18478
rect 13375 18365 13415 18372
rect 13458 18365 13695 18372
rect 13925 18478 14042 18485
rect 14085 18478 14245 18485
rect 13925 18372 14008 18478
rect 14042 18372 14245 18478
rect 13925 18365 13965 18372
rect 14008 18365 14245 18372
rect 14475 18478 14592 18485
rect 14635 18478 14795 18485
rect 14475 18372 14558 18478
rect 14592 18372 14795 18478
rect 14475 18365 14515 18372
rect 14558 18365 14795 18372
rect 15025 18478 15142 18485
rect 15185 18478 15345 18485
rect 15025 18372 15108 18478
rect 15142 18372 15345 18478
rect 15025 18365 15065 18372
rect 15108 18365 15345 18372
rect 15575 18478 15692 18485
rect 15735 18478 15895 18485
rect 15575 18372 15658 18478
rect 15692 18372 15895 18478
rect 15575 18365 15615 18372
rect 15658 18365 15895 18372
rect 16125 18478 16242 18485
rect 16285 18478 16445 18485
rect 16125 18372 16208 18478
rect 16242 18372 16445 18478
rect 16125 18365 16165 18372
rect 16208 18365 16445 18372
rect 16675 18478 16792 18485
rect 16835 18478 16995 18485
rect 16675 18372 16758 18478
rect 16792 18372 16995 18478
rect 16675 18365 16715 18372
rect 16758 18365 16995 18372
rect 17225 18478 17342 18485
rect 17385 18478 17545 18485
rect 17225 18372 17308 18478
rect 17342 18372 17545 18478
rect 17225 18365 17265 18372
rect 17308 18365 17545 18372
rect 17775 18478 17892 18485
rect 17935 18478 18095 18485
rect 17775 18372 17858 18478
rect 17892 18372 18095 18478
rect 17775 18365 17815 18372
rect 17858 18365 18095 18372
rect 18325 18478 18442 18485
rect 18485 18478 18645 18485
rect 18325 18372 18408 18478
rect 18442 18372 18645 18478
rect 18325 18365 18365 18372
rect 18408 18365 18645 18372
rect 18875 18478 18992 18485
rect 19035 18478 19195 18485
rect 18875 18372 18958 18478
rect 18992 18372 19195 18478
rect 18875 18365 18915 18372
rect 18958 18365 19195 18372
rect 765 18325 885 18365
rect 1315 18325 1435 18365
rect 1865 18325 1985 18365
rect 2415 18325 2535 18365
rect 2965 18325 3085 18365
rect 3515 18325 3635 18365
rect 4065 18325 4185 18365
rect 4615 18325 4735 18365
rect 5165 18325 5285 18365
rect 5715 18325 5835 18365
rect 6265 18325 6385 18365
rect 6815 18325 6935 18365
rect 7365 18325 7485 18365
rect 7915 18325 8035 18365
rect 8465 18325 8585 18365
rect 9015 18325 9135 18365
rect 9565 18325 9685 18365
rect 10115 18325 10235 18365
rect 10665 18325 10785 18365
rect 11215 18325 11335 18365
rect 11765 18325 11885 18365
rect 12315 18325 12435 18365
rect 12865 18325 12985 18365
rect 13415 18325 13535 18365
rect 13965 18325 14085 18365
rect 14515 18325 14635 18365
rect 15065 18325 15185 18365
rect 15615 18325 15735 18365
rect 16165 18325 16285 18365
rect 16715 18325 16835 18365
rect 17265 18325 17385 18365
rect 17815 18325 17935 18365
rect 18365 18325 18485 18365
rect 18915 18325 19035 18365
rect 19202 18212 19204 18638
rect 500 18125 507 18175
rect 19202 18096 19217 18102
rect 628 18072 885 18095
rect 1178 18072 1435 18095
rect 1728 18072 1985 18095
rect 2278 18072 2535 18095
rect 2828 18072 3085 18095
rect 3378 18072 3635 18095
rect 3928 18072 4185 18095
rect 4478 18072 4735 18095
rect 5028 18072 5285 18095
rect 5578 18072 5835 18095
rect 6128 18072 6385 18095
rect 6678 18072 6935 18095
rect 7228 18072 7485 18095
rect 7778 18072 8035 18095
rect 8328 18072 8585 18095
rect 8878 18072 9135 18095
rect 9428 18072 9685 18095
rect 9978 18072 10235 18095
rect 10528 18072 10785 18095
rect 11078 18072 11335 18095
rect 11628 18072 11885 18095
rect 12178 18072 12435 18095
rect 12728 18072 12985 18095
rect 13278 18072 13535 18095
rect 13828 18072 14085 18095
rect 14378 18072 14635 18095
rect 14928 18072 15185 18095
rect 15478 18072 15735 18095
rect 16028 18072 16285 18095
rect 16578 18072 16835 18095
rect 17128 18072 17385 18095
rect 17678 18072 17935 18095
rect 18228 18072 18485 18095
rect 18778 18072 19035 18095
rect 605 17935 609 18020
rect 784 17975 885 18072
rect 765 17935 885 17975
rect 1155 17935 1159 18020
rect 1334 17975 1435 18072
rect 1315 17935 1435 17975
rect 1705 17935 1709 18020
rect 1884 17975 1985 18072
rect 1865 17935 1985 17975
rect 2255 17935 2259 18020
rect 2434 17975 2535 18072
rect 2415 17935 2535 17975
rect 2805 17935 2809 18020
rect 2984 17975 3085 18072
rect 2965 17935 3085 17975
rect 3355 17935 3359 18020
rect 3534 17975 3635 18072
rect 3515 17935 3635 17975
rect 3905 17935 3909 18020
rect 4084 17975 4185 18072
rect 4065 17935 4185 17975
rect 4455 17935 4459 18020
rect 4634 17975 4735 18072
rect 4615 17935 4735 17975
rect 5005 17935 5009 18020
rect 5184 17975 5285 18072
rect 5165 17935 5285 17975
rect 5555 17935 5559 18020
rect 5734 17975 5835 18072
rect 5715 17935 5835 17975
rect 6105 17935 6109 18020
rect 6284 17975 6385 18072
rect 6265 17935 6385 17975
rect 6655 17935 6659 18020
rect 6834 17975 6935 18072
rect 6815 17935 6935 17975
rect 7205 17935 7209 18020
rect 7384 17975 7485 18072
rect 7365 17935 7485 17975
rect 7755 17935 7759 18020
rect 7934 17975 8035 18072
rect 7915 17935 8035 17975
rect 8305 17935 8309 18020
rect 8484 17975 8585 18072
rect 8465 17935 8585 17975
rect 8855 17935 8859 18020
rect 9034 17975 9135 18072
rect 9015 17935 9135 17975
rect 9405 17935 9409 18020
rect 9584 17975 9685 18072
rect 9565 17935 9685 17975
rect 9955 17935 9959 18020
rect 10134 17975 10235 18072
rect 10115 17935 10235 17975
rect 10505 17935 10509 18020
rect 10684 17975 10785 18072
rect 10665 17935 10785 17975
rect 11055 17935 11059 18020
rect 11234 17975 11335 18072
rect 11215 17935 11335 17975
rect 11605 17935 11609 18020
rect 11784 17975 11885 18072
rect 11765 17935 11885 17975
rect 12155 17935 12159 18020
rect 12334 17975 12435 18072
rect 12315 17935 12435 17975
rect 12705 17935 12709 18020
rect 12884 17975 12985 18072
rect 12865 17935 12985 17975
rect 13255 17935 13259 18020
rect 13434 17975 13535 18072
rect 13415 17935 13535 17975
rect 13805 17935 13809 18020
rect 13984 17975 14085 18072
rect 13965 17935 14085 17975
rect 14355 17935 14359 18020
rect 14534 17975 14635 18072
rect 14515 17935 14635 17975
rect 14905 17935 14909 18020
rect 15084 17975 15185 18072
rect 15065 17935 15185 17975
rect 15455 17935 15459 18020
rect 15634 17975 15735 18072
rect 15615 17935 15735 17975
rect 16005 17935 16009 18020
rect 16184 17975 16285 18072
rect 16165 17935 16285 17975
rect 16555 17935 16559 18020
rect 16734 17975 16835 18072
rect 16715 17935 16835 17975
rect 17105 17935 17109 18020
rect 17284 17975 17385 18072
rect 17265 17935 17385 17975
rect 17655 17935 17659 18020
rect 17834 17975 17935 18072
rect 17815 17935 17935 17975
rect 18205 17935 18209 18020
rect 18384 17975 18485 18072
rect 18365 17935 18485 17975
rect 18755 17935 18759 18020
rect 18934 17975 19035 18072
rect 18915 17935 19035 17975
rect 725 17928 842 17935
rect 885 17928 1045 17935
rect 725 17822 808 17928
rect 842 17822 1045 17928
rect 725 17815 765 17822
rect 808 17815 1045 17822
rect 1275 17928 1392 17935
rect 1435 17928 1595 17935
rect 1275 17822 1358 17928
rect 1392 17822 1595 17928
rect 1275 17815 1315 17822
rect 1358 17815 1595 17822
rect 1825 17928 1942 17935
rect 1985 17928 2145 17935
rect 1825 17822 1908 17928
rect 1942 17822 2145 17928
rect 1825 17815 1865 17822
rect 1908 17815 2145 17822
rect 2375 17928 2492 17935
rect 2535 17928 2695 17935
rect 2375 17822 2458 17928
rect 2492 17822 2695 17928
rect 2375 17815 2415 17822
rect 2458 17815 2695 17822
rect 2925 17928 3042 17935
rect 3085 17928 3245 17935
rect 2925 17822 3008 17928
rect 3042 17822 3245 17928
rect 2925 17815 2965 17822
rect 3008 17815 3245 17822
rect 3475 17928 3592 17935
rect 3635 17928 3795 17935
rect 3475 17822 3558 17928
rect 3592 17822 3795 17928
rect 3475 17815 3515 17822
rect 3558 17815 3795 17822
rect 4025 17928 4142 17935
rect 4185 17928 4345 17935
rect 4025 17822 4108 17928
rect 4142 17822 4345 17928
rect 4025 17815 4065 17822
rect 4108 17815 4345 17822
rect 4575 17928 4692 17935
rect 4735 17928 4895 17935
rect 4575 17822 4658 17928
rect 4692 17822 4895 17928
rect 4575 17815 4615 17822
rect 4658 17815 4895 17822
rect 5125 17928 5242 17935
rect 5285 17928 5445 17935
rect 5125 17822 5208 17928
rect 5242 17822 5445 17928
rect 5125 17815 5165 17822
rect 5208 17815 5445 17822
rect 5675 17928 5792 17935
rect 5835 17928 5995 17935
rect 5675 17822 5758 17928
rect 5792 17822 5995 17928
rect 5675 17815 5715 17822
rect 5758 17815 5995 17822
rect 6225 17928 6342 17935
rect 6385 17928 6545 17935
rect 6225 17822 6308 17928
rect 6342 17822 6545 17928
rect 6225 17815 6265 17822
rect 6308 17815 6545 17822
rect 6775 17928 6892 17935
rect 6935 17928 7095 17935
rect 6775 17822 6858 17928
rect 6892 17822 7095 17928
rect 6775 17815 6815 17822
rect 6858 17815 7095 17822
rect 7325 17928 7442 17935
rect 7485 17928 7645 17935
rect 7325 17822 7408 17928
rect 7442 17822 7645 17928
rect 7325 17815 7365 17822
rect 7408 17815 7645 17822
rect 7875 17928 7992 17935
rect 8035 17928 8195 17935
rect 7875 17822 7958 17928
rect 7992 17822 8195 17928
rect 7875 17815 7915 17822
rect 7958 17815 8195 17822
rect 8425 17928 8542 17935
rect 8585 17928 8745 17935
rect 8425 17822 8508 17928
rect 8542 17822 8745 17928
rect 8425 17815 8465 17822
rect 8508 17815 8745 17822
rect 8975 17928 9092 17935
rect 9135 17928 9295 17935
rect 8975 17822 9058 17928
rect 9092 17822 9295 17928
rect 8975 17815 9015 17822
rect 9058 17815 9295 17822
rect 9525 17928 9642 17935
rect 9685 17928 9845 17935
rect 9525 17822 9608 17928
rect 9642 17822 9845 17928
rect 9525 17815 9565 17822
rect 9608 17815 9845 17822
rect 10075 17928 10192 17935
rect 10235 17928 10395 17935
rect 10075 17822 10158 17928
rect 10192 17822 10395 17928
rect 10075 17815 10115 17822
rect 10158 17815 10395 17822
rect 10625 17928 10742 17935
rect 10785 17928 10945 17935
rect 10625 17822 10708 17928
rect 10742 17822 10945 17928
rect 10625 17815 10665 17822
rect 10708 17815 10945 17822
rect 11175 17928 11292 17935
rect 11335 17928 11495 17935
rect 11175 17822 11258 17928
rect 11292 17822 11495 17928
rect 11175 17815 11215 17822
rect 11258 17815 11495 17822
rect 11725 17928 11842 17935
rect 11885 17928 12045 17935
rect 11725 17822 11808 17928
rect 11842 17822 12045 17928
rect 11725 17815 11765 17822
rect 11808 17815 12045 17822
rect 12275 17928 12392 17935
rect 12435 17928 12595 17935
rect 12275 17822 12358 17928
rect 12392 17822 12595 17928
rect 12275 17815 12315 17822
rect 12358 17815 12595 17822
rect 12825 17928 12942 17935
rect 12985 17928 13145 17935
rect 12825 17822 12908 17928
rect 12942 17822 13145 17928
rect 12825 17815 12865 17822
rect 12908 17815 13145 17822
rect 13375 17928 13492 17935
rect 13535 17928 13695 17935
rect 13375 17822 13458 17928
rect 13492 17822 13695 17928
rect 13375 17815 13415 17822
rect 13458 17815 13695 17822
rect 13925 17928 14042 17935
rect 14085 17928 14245 17935
rect 13925 17822 14008 17928
rect 14042 17822 14245 17928
rect 13925 17815 13965 17822
rect 14008 17815 14245 17822
rect 14475 17928 14592 17935
rect 14635 17928 14795 17935
rect 14475 17822 14558 17928
rect 14592 17822 14795 17928
rect 14475 17815 14515 17822
rect 14558 17815 14795 17822
rect 15025 17928 15142 17935
rect 15185 17928 15345 17935
rect 15025 17822 15108 17928
rect 15142 17822 15345 17928
rect 15025 17815 15065 17822
rect 15108 17815 15345 17822
rect 15575 17928 15692 17935
rect 15735 17928 15895 17935
rect 15575 17822 15658 17928
rect 15692 17822 15895 17928
rect 15575 17815 15615 17822
rect 15658 17815 15895 17822
rect 16125 17928 16242 17935
rect 16285 17928 16445 17935
rect 16125 17822 16208 17928
rect 16242 17822 16445 17928
rect 16125 17815 16165 17822
rect 16208 17815 16445 17822
rect 16675 17928 16792 17935
rect 16835 17928 16995 17935
rect 16675 17822 16758 17928
rect 16792 17822 16995 17928
rect 16675 17815 16715 17822
rect 16758 17815 16995 17822
rect 17225 17928 17342 17935
rect 17385 17928 17545 17935
rect 17225 17822 17308 17928
rect 17342 17822 17545 17928
rect 17225 17815 17265 17822
rect 17308 17815 17545 17822
rect 17775 17928 17892 17935
rect 17935 17928 18095 17935
rect 17775 17822 17858 17928
rect 17892 17822 18095 17928
rect 17775 17815 17815 17822
rect 17858 17815 18095 17822
rect 18325 17928 18442 17935
rect 18485 17928 18645 17935
rect 18325 17822 18408 17928
rect 18442 17822 18645 17928
rect 18325 17815 18365 17822
rect 18408 17815 18645 17822
rect 18875 17928 18992 17935
rect 19035 17928 19195 17935
rect 18875 17822 18958 17928
rect 18992 17822 19195 17928
rect 18875 17815 18915 17822
rect 18958 17815 19195 17822
rect 765 17775 885 17815
rect 1315 17775 1435 17815
rect 1865 17775 1985 17815
rect 2415 17775 2535 17815
rect 2965 17775 3085 17815
rect 3515 17775 3635 17815
rect 4065 17775 4185 17815
rect 4615 17775 4735 17815
rect 5165 17775 5285 17815
rect 5715 17775 5835 17815
rect 6265 17775 6385 17815
rect 6815 17775 6935 17815
rect 7365 17775 7485 17815
rect 7915 17775 8035 17815
rect 8465 17775 8585 17815
rect 9015 17775 9135 17815
rect 9565 17775 9685 17815
rect 10115 17775 10235 17815
rect 10665 17775 10785 17815
rect 11215 17775 11335 17815
rect 11765 17775 11885 17815
rect 12315 17775 12435 17815
rect 12865 17775 12985 17815
rect 13415 17775 13535 17815
rect 13965 17775 14085 17815
rect 14515 17775 14635 17815
rect 15065 17775 15185 17815
rect 15615 17775 15735 17815
rect 16165 17775 16285 17815
rect 16715 17775 16835 17815
rect 17265 17775 17385 17815
rect 17815 17775 17935 17815
rect 18365 17775 18485 17815
rect 18915 17775 19035 17815
rect 19185 17654 19200 17671
rect 19202 17662 19204 18088
rect 19202 17648 19217 17654
rect 500 17575 507 17625
rect 500 17139 525 17540
rect 628 17522 885 17545
rect 1178 17522 1435 17545
rect 1728 17522 1985 17545
rect 2278 17522 2535 17545
rect 2828 17522 3085 17545
rect 3378 17522 3635 17545
rect 3928 17522 4185 17545
rect 4478 17522 4735 17545
rect 5028 17522 5285 17545
rect 5578 17522 5835 17545
rect 6128 17522 6385 17545
rect 6678 17522 6935 17545
rect 7228 17522 7485 17545
rect 7778 17522 8035 17545
rect 8328 17522 8585 17545
rect 8878 17522 9135 17545
rect 9428 17522 9685 17545
rect 9978 17522 10235 17545
rect 10528 17522 10785 17545
rect 11078 17522 11335 17545
rect 11628 17522 11885 17545
rect 12178 17522 12435 17545
rect 12728 17522 12985 17545
rect 13278 17522 13535 17545
rect 13828 17522 14085 17545
rect 14378 17522 14635 17545
rect 14928 17522 15185 17545
rect 15478 17522 15735 17545
rect 16028 17522 16285 17545
rect 16578 17522 16835 17545
rect 17128 17522 17385 17545
rect 17678 17522 17935 17545
rect 18228 17522 18485 17545
rect 18778 17522 19035 17545
rect 605 17385 609 17522
rect 784 17425 885 17522
rect 765 17385 885 17425
rect 1155 17385 1159 17522
rect 1334 17425 1435 17522
rect 1315 17385 1435 17425
rect 1705 17385 1709 17522
rect 1884 17425 1985 17522
rect 1865 17385 1985 17425
rect 2255 17385 2259 17522
rect 2434 17425 2535 17522
rect 2415 17385 2535 17425
rect 2805 17385 2809 17522
rect 2984 17425 3085 17522
rect 2965 17385 3085 17425
rect 3355 17385 3359 17522
rect 3534 17425 3635 17522
rect 3515 17385 3635 17425
rect 3905 17385 3909 17522
rect 4084 17425 4185 17522
rect 4065 17385 4185 17425
rect 4455 17385 4459 17522
rect 4634 17425 4735 17522
rect 4615 17385 4735 17425
rect 5005 17385 5009 17522
rect 5184 17425 5285 17522
rect 5165 17385 5285 17425
rect 5555 17385 5559 17522
rect 5734 17425 5835 17522
rect 5715 17385 5835 17425
rect 6105 17385 6109 17522
rect 6284 17425 6385 17522
rect 6265 17385 6385 17425
rect 6655 17385 6659 17522
rect 6834 17425 6935 17522
rect 6815 17385 6935 17425
rect 7205 17385 7209 17522
rect 7384 17425 7485 17522
rect 7365 17385 7485 17425
rect 7755 17385 7759 17522
rect 7934 17425 8035 17522
rect 7915 17385 8035 17425
rect 8305 17385 8309 17522
rect 8484 17425 8585 17522
rect 8465 17385 8585 17425
rect 8855 17385 8859 17522
rect 9034 17425 9135 17522
rect 9015 17385 9135 17425
rect 9405 17385 9409 17522
rect 9584 17425 9685 17522
rect 9565 17385 9685 17425
rect 9955 17385 9959 17522
rect 10134 17425 10235 17522
rect 10115 17385 10235 17425
rect 10505 17385 10509 17522
rect 10684 17425 10785 17522
rect 10665 17385 10785 17425
rect 11055 17385 11059 17522
rect 11234 17425 11335 17522
rect 11215 17385 11335 17425
rect 11605 17385 11609 17522
rect 11784 17425 11885 17522
rect 11765 17385 11885 17425
rect 12155 17385 12159 17522
rect 12334 17425 12435 17522
rect 12315 17385 12435 17425
rect 12705 17385 12709 17522
rect 12884 17425 12985 17522
rect 12865 17385 12985 17425
rect 13255 17385 13259 17522
rect 13434 17425 13535 17522
rect 13415 17385 13535 17425
rect 13805 17385 13809 17522
rect 13984 17425 14085 17522
rect 13965 17385 14085 17425
rect 14355 17385 14359 17522
rect 14534 17425 14635 17522
rect 14515 17385 14635 17425
rect 14905 17385 14909 17522
rect 15084 17425 15185 17522
rect 15065 17385 15185 17425
rect 15455 17385 15459 17522
rect 15634 17425 15735 17522
rect 15615 17385 15735 17425
rect 16005 17385 16009 17522
rect 16184 17425 16285 17522
rect 16165 17385 16285 17425
rect 16555 17385 16559 17522
rect 16734 17425 16835 17522
rect 16715 17385 16835 17425
rect 17105 17385 17109 17522
rect 17284 17425 17385 17522
rect 17265 17385 17385 17425
rect 17655 17385 17659 17522
rect 17834 17425 17935 17522
rect 17815 17385 17935 17425
rect 18205 17385 18209 17522
rect 18384 17425 18485 17522
rect 18365 17385 18485 17425
rect 18755 17385 18759 17522
rect 18934 17425 19035 17522
rect 18915 17385 19035 17425
rect 725 17378 842 17385
rect 885 17378 1045 17385
rect 725 17272 808 17378
rect 842 17272 1045 17378
rect 725 17265 765 17272
rect 808 17265 1045 17272
rect 1275 17378 1392 17385
rect 1435 17378 1595 17385
rect 1275 17272 1358 17378
rect 1392 17272 1595 17378
rect 1275 17265 1315 17272
rect 1358 17265 1595 17272
rect 1825 17378 1942 17385
rect 1985 17378 2145 17385
rect 1825 17272 1908 17378
rect 1942 17272 2145 17378
rect 1825 17265 1865 17272
rect 1908 17265 2145 17272
rect 2375 17378 2492 17385
rect 2535 17378 2695 17385
rect 2375 17272 2458 17378
rect 2492 17272 2695 17378
rect 2375 17265 2415 17272
rect 2458 17265 2695 17272
rect 2925 17378 3042 17385
rect 3085 17378 3245 17385
rect 2925 17272 3008 17378
rect 3042 17272 3245 17378
rect 2925 17265 2965 17272
rect 3008 17265 3245 17272
rect 3475 17378 3592 17385
rect 3635 17378 3795 17385
rect 3475 17272 3558 17378
rect 3592 17272 3795 17378
rect 3475 17265 3515 17272
rect 3558 17265 3795 17272
rect 4025 17378 4142 17385
rect 4185 17378 4345 17385
rect 4025 17272 4108 17378
rect 4142 17272 4345 17378
rect 4025 17265 4065 17272
rect 4108 17265 4345 17272
rect 4575 17378 4692 17385
rect 4735 17378 4895 17385
rect 4575 17272 4658 17378
rect 4692 17272 4895 17378
rect 4575 17265 4615 17272
rect 4658 17265 4895 17272
rect 5125 17378 5242 17385
rect 5285 17378 5445 17385
rect 5125 17272 5208 17378
rect 5242 17272 5445 17378
rect 5125 17265 5165 17272
rect 5208 17265 5445 17272
rect 5675 17378 5792 17385
rect 5835 17378 5995 17385
rect 5675 17272 5758 17378
rect 5792 17272 5995 17378
rect 5675 17265 5715 17272
rect 5758 17265 5995 17272
rect 6225 17378 6342 17385
rect 6385 17378 6545 17385
rect 6225 17272 6308 17378
rect 6342 17272 6545 17378
rect 6225 17265 6265 17272
rect 6308 17265 6545 17272
rect 6775 17378 6892 17385
rect 6935 17378 7095 17385
rect 6775 17272 6858 17378
rect 6892 17272 7095 17378
rect 6775 17265 6815 17272
rect 6858 17265 7095 17272
rect 7325 17378 7442 17385
rect 7485 17378 7645 17385
rect 7325 17272 7408 17378
rect 7442 17272 7645 17378
rect 7325 17265 7365 17272
rect 7408 17265 7645 17272
rect 7875 17378 7992 17385
rect 8035 17378 8195 17385
rect 7875 17272 7958 17378
rect 7992 17272 8195 17378
rect 7875 17265 7915 17272
rect 7958 17265 8195 17272
rect 8425 17378 8542 17385
rect 8585 17378 8745 17385
rect 8425 17272 8508 17378
rect 8542 17272 8745 17378
rect 8425 17265 8465 17272
rect 8508 17265 8745 17272
rect 8975 17378 9092 17385
rect 9135 17378 9295 17385
rect 8975 17272 9058 17378
rect 9092 17272 9295 17378
rect 8975 17265 9015 17272
rect 9058 17265 9295 17272
rect 9525 17378 9642 17385
rect 9685 17378 9845 17385
rect 9525 17272 9608 17378
rect 9642 17272 9845 17378
rect 9525 17265 9565 17272
rect 9608 17265 9845 17272
rect 10075 17378 10192 17385
rect 10235 17378 10395 17385
rect 10075 17272 10158 17378
rect 10192 17272 10395 17378
rect 10075 17265 10115 17272
rect 10158 17265 10395 17272
rect 10625 17378 10742 17385
rect 10785 17378 10945 17385
rect 10625 17272 10708 17378
rect 10742 17272 10945 17378
rect 10625 17265 10665 17272
rect 10708 17265 10945 17272
rect 11175 17378 11292 17385
rect 11335 17378 11495 17385
rect 11175 17272 11258 17378
rect 11292 17272 11495 17378
rect 11175 17265 11215 17272
rect 11258 17265 11495 17272
rect 11725 17378 11842 17385
rect 11885 17378 12045 17385
rect 11725 17272 11808 17378
rect 11842 17272 12045 17378
rect 11725 17265 11765 17272
rect 11808 17265 12045 17272
rect 12275 17378 12392 17385
rect 12435 17378 12595 17385
rect 12275 17272 12358 17378
rect 12392 17272 12595 17378
rect 12275 17265 12315 17272
rect 12358 17265 12595 17272
rect 12825 17378 12942 17385
rect 12985 17378 13145 17385
rect 12825 17272 12908 17378
rect 12942 17272 13145 17378
rect 12825 17265 12865 17272
rect 12908 17265 13145 17272
rect 13375 17378 13492 17385
rect 13535 17378 13695 17385
rect 13375 17272 13458 17378
rect 13492 17272 13695 17378
rect 13375 17265 13415 17272
rect 13458 17265 13695 17272
rect 13925 17378 14042 17385
rect 14085 17378 14245 17385
rect 13925 17272 14008 17378
rect 14042 17272 14245 17378
rect 13925 17265 13965 17272
rect 14008 17265 14245 17272
rect 14475 17378 14592 17385
rect 14635 17378 14795 17385
rect 14475 17272 14558 17378
rect 14592 17272 14795 17378
rect 14475 17265 14515 17272
rect 14558 17265 14795 17272
rect 15025 17378 15142 17385
rect 15185 17378 15345 17385
rect 15025 17272 15108 17378
rect 15142 17272 15345 17378
rect 15025 17265 15065 17272
rect 15108 17265 15345 17272
rect 15575 17378 15692 17385
rect 15735 17378 15895 17385
rect 15575 17272 15658 17378
rect 15692 17272 15895 17378
rect 15575 17265 15615 17272
rect 15658 17265 15895 17272
rect 16125 17378 16242 17385
rect 16285 17378 16445 17385
rect 16125 17272 16208 17378
rect 16242 17272 16445 17378
rect 16125 17265 16165 17272
rect 16208 17265 16445 17272
rect 16675 17378 16792 17385
rect 16835 17378 16995 17385
rect 16675 17272 16758 17378
rect 16792 17272 16995 17378
rect 16675 17265 16715 17272
rect 16758 17265 16995 17272
rect 17225 17378 17342 17385
rect 17385 17378 17545 17385
rect 17225 17272 17308 17378
rect 17342 17272 17545 17378
rect 17225 17265 17265 17272
rect 17308 17265 17545 17272
rect 17775 17378 17892 17385
rect 17935 17378 18095 17385
rect 17775 17272 17858 17378
rect 17892 17272 18095 17378
rect 17775 17265 17815 17272
rect 17858 17265 18095 17272
rect 18325 17378 18442 17385
rect 18485 17378 18645 17385
rect 18325 17272 18408 17378
rect 18442 17272 18645 17378
rect 18325 17265 18365 17272
rect 18408 17265 18645 17272
rect 18875 17378 18992 17385
rect 19035 17378 19195 17385
rect 18875 17272 18958 17378
rect 18992 17272 19195 17378
rect 18875 17265 18915 17272
rect 18958 17265 19195 17272
rect 765 17225 885 17265
rect 1315 17225 1435 17265
rect 1865 17225 1985 17265
rect 2415 17225 2535 17265
rect 2965 17225 3085 17265
rect 3515 17225 3635 17265
rect 4065 17225 4185 17265
rect 4615 17225 4735 17265
rect 5165 17225 5285 17265
rect 5715 17225 5835 17265
rect 6265 17225 6385 17265
rect 6815 17225 6935 17265
rect 7365 17225 7485 17265
rect 7915 17225 8035 17265
rect 8465 17225 8585 17265
rect 9015 17225 9135 17265
rect 9565 17225 9685 17265
rect 10115 17225 10235 17265
rect 10665 17225 10785 17265
rect 11215 17225 11335 17265
rect 11765 17225 11885 17265
rect 12315 17225 12435 17265
rect 12865 17225 12985 17265
rect 13415 17225 13535 17265
rect 13965 17225 14085 17265
rect 14515 17225 14635 17265
rect 15065 17225 15185 17265
rect 15615 17225 15735 17265
rect 16165 17225 16285 17265
rect 16715 17225 16835 17265
rect 17265 17225 17385 17265
rect 17815 17225 17935 17265
rect 18365 17225 18485 17265
rect 18915 17225 19035 17265
rect 19202 17112 19204 17538
rect 500 17025 507 17075
rect 19202 16996 19217 17002
rect 628 16972 885 16995
rect 1178 16972 1435 16995
rect 1728 16972 1985 16995
rect 2278 16972 2535 16995
rect 2828 16972 3085 16995
rect 3378 16972 3635 16995
rect 3928 16972 4185 16995
rect 4478 16972 4735 16995
rect 5028 16972 5285 16995
rect 5578 16972 5835 16995
rect 6128 16972 6385 16995
rect 6678 16972 6935 16995
rect 7228 16972 7485 16995
rect 7778 16972 8035 16995
rect 8328 16972 8585 16995
rect 8878 16972 9135 16995
rect 9428 16972 9685 16995
rect 9978 16972 10235 16995
rect 10528 16972 10785 16995
rect 11078 16972 11335 16995
rect 11628 16972 11885 16995
rect 12178 16972 12435 16995
rect 12728 16972 12985 16995
rect 13278 16972 13535 16995
rect 13828 16972 14085 16995
rect 14378 16972 14635 16995
rect 14928 16972 15185 16995
rect 15478 16972 15735 16995
rect 16028 16972 16285 16995
rect 16578 16972 16835 16995
rect 17128 16972 17385 16995
rect 17678 16972 17935 16995
rect 18228 16972 18485 16995
rect 18778 16972 19035 16995
rect 605 16835 609 16972
rect 784 16875 885 16972
rect 765 16835 885 16875
rect 1155 16835 1159 16972
rect 1334 16875 1435 16972
rect 1315 16835 1435 16875
rect 1705 16835 1709 16972
rect 1884 16875 1985 16972
rect 1865 16835 1985 16875
rect 2255 16835 2259 16972
rect 2434 16875 2535 16972
rect 2415 16835 2535 16875
rect 2805 16835 2809 16972
rect 2984 16875 3085 16972
rect 2965 16835 3085 16875
rect 3355 16835 3359 16972
rect 3534 16875 3635 16972
rect 3515 16835 3635 16875
rect 3905 16835 3909 16972
rect 4084 16875 4185 16972
rect 4065 16835 4185 16875
rect 4455 16835 4459 16972
rect 4634 16875 4735 16972
rect 4615 16835 4735 16875
rect 5005 16835 5009 16972
rect 5184 16875 5285 16972
rect 5165 16835 5285 16875
rect 5555 16835 5559 16972
rect 5734 16875 5835 16972
rect 5715 16835 5835 16875
rect 6105 16835 6109 16972
rect 6284 16875 6385 16972
rect 6265 16835 6385 16875
rect 6655 16835 6659 16972
rect 6834 16875 6935 16972
rect 6815 16835 6935 16875
rect 7205 16835 7209 16972
rect 7384 16875 7485 16972
rect 7365 16835 7485 16875
rect 7755 16835 7759 16972
rect 7934 16875 8035 16972
rect 7915 16835 8035 16875
rect 8305 16835 8309 16972
rect 8484 16875 8585 16972
rect 8465 16835 8585 16875
rect 8855 16835 8859 16972
rect 9034 16875 9135 16972
rect 9015 16835 9135 16875
rect 9405 16835 9409 16972
rect 9584 16875 9685 16972
rect 9565 16835 9685 16875
rect 9955 16835 9959 16972
rect 10134 16875 10235 16972
rect 10115 16835 10235 16875
rect 10505 16835 10509 16972
rect 10684 16875 10785 16972
rect 10665 16835 10785 16875
rect 11055 16835 11059 16972
rect 11234 16875 11335 16972
rect 11215 16835 11335 16875
rect 11605 16835 11609 16972
rect 11784 16875 11885 16972
rect 11765 16835 11885 16875
rect 12155 16835 12159 16972
rect 12334 16875 12435 16972
rect 12315 16835 12435 16875
rect 12705 16835 12709 16972
rect 12884 16875 12985 16972
rect 12865 16835 12985 16875
rect 13255 16835 13259 16972
rect 13434 16875 13535 16972
rect 13415 16835 13535 16875
rect 13805 16835 13809 16972
rect 13984 16875 14085 16972
rect 13965 16835 14085 16875
rect 14355 16835 14359 16972
rect 14534 16875 14635 16972
rect 14515 16835 14635 16875
rect 14905 16835 14909 16972
rect 15084 16875 15185 16972
rect 15065 16835 15185 16875
rect 15455 16835 15459 16972
rect 15634 16875 15735 16972
rect 15615 16835 15735 16875
rect 16005 16835 16009 16972
rect 16184 16875 16285 16972
rect 16165 16835 16285 16875
rect 16555 16835 16559 16972
rect 16734 16875 16835 16972
rect 16715 16835 16835 16875
rect 17105 16835 17109 16972
rect 17284 16875 17385 16972
rect 17265 16835 17385 16875
rect 17655 16835 17659 16972
rect 17834 16875 17935 16972
rect 17815 16835 17935 16875
rect 18205 16835 18209 16972
rect 18384 16875 18485 16972
rect 18365 16835 18485 16875
rect 18755 16835 18759 16972
rect 18934 16875 19035 16972
rect 18915 16835 19035 16875
rect 725 16828 842 16835
rect 885 16828 1045 16835
rect 725 16722 808 16828
rect 842 16722 1045 16828
rect 725 16715 765 16722
rect 808 16715 1045 16722
rect 1275 16828 1392 16835
rect 1435 16828 1595 16835
rect 1275 16722 1358 16828
rect 1392 16722 1595 16828
rect 1275 16715 1315 16722
rect 1358 16715 1595 16722
rect 1825 16828 1942 16835
rect 1985 16828 2145 16835
rect 1825 16722 1908 16828
rect 1942 16722 2145 16828
rect 1825 16715 1865 16722
rect 1908 16715 2145 16722
rect 2375 16828 2492 16835
rect 2535 16828 2695 16835
rect 2375 16722 2458 16828
rect 2492 16722 2695 16828
rect 2375 16715 2415 16722
rect 2458 16715 2695 16722
rect 2925 16828 3042 16835
rect 3085 16828 3245 16835
rect 2925 16722 3008 16828
rect 3042 16722 3245 16828
rect 2925 16715 2965 16722
rect 3008 16715 3245 16722
rect 3475 16828 3592 16835
rect 3635 16828 3795 16835
rect 3475 16722 3558 16828
rect 3592 16722 3795 16828
rect 3475 16715 3515 16722
rect 3558 16715 3795 16722
rect 4025 16828 4142 16835
rect 4185 16828 4345 16835
rect 4025 16722 4108 16828
rect 4142 16722 4345 16828
rect 4025 16715 4065 16722
rect 4108 16715 4345 16722
rect 4575 16828 4692 16835
rect 4735 16828 4895 16835
rect 4575 16722 4658 16828
rect 4692 16722 4895 16828
rect 4575 16715 4615 16722
rect 4658 16715 4895 16722
rect 5125 16828 5242 16835
rect 5285 16828 5445 16835
rect 5125 16722 5208 16828
rect 5242 16722 5445 16828
rect 5125 16715 5165 16722
rect 5208 16715 5445 16722
rect 5675 16828 5792 16835
rect 5835 16828 5995 16835
rect 5675 16722 5758 16828
rect 5792 16722 5995 16828
rect 5675 16715 5715 16722
rect 5758 16715 5995 16722
rect 6225 16828 6342 16835
rect 6385 16828 6545 16835
rect 6225 16722 6308 16828
rect 6342 16722 6545 16828
rect 6225 16715 6265 16722
rect 6308 16715 6545 16722
rect 6775 16828 6892 16835
rect 6935 16828 7095 16835
rect 6775 16722 6858 16828
rect 6892 16722 7095 16828
rect 6775 16715 6815 16722
rect 6858 16715 7095 16722
rect 7325 16828 7442 16835
rect 7485 16828 7645 16835
rect 7325 16722 7408 16828
rect 7442 16722 7645 16828
rect 7325 16715 7365 16722
rect 7408 16715 7645 16722
rect 7875 16828 7992 16835
rect 8035 16828 8195 16835
rect 7875 16722 7958 16828
rect 7992 16722 8195 16828
rect 7875 16715 7915 16722
rect 7958 16715 8195 16722
rect 8425 16828 8542 16835
rect 8585 16828 8745 16835
rect 8425 16722 8508 16828
rect 8542 16722 8745 16828
rect 8425 16715 8465 16722
rect 8508 16715 8745 16722
rect 8975 16828 9092 16835
rect 9135 16828 9295 16835
rect 8975 16722 9058 16828
rect 9092 16722 9295 16828
rect 8975 16715 9015 16722
rect 9058 16715 9295 16722
rect 9525 16828 9642 16835
rect 9685 16828 9845 16835
rect 9525 16722 9608 16828
rect 9642 16722 9845 16828
rect 9525 16715 9565 16722
rect 9608 16715 9845 16722
rect 10075 16828 10192 16835
rect 10235 16828 10395 16835
rect 10075 16722 10158 16828
rect 10192 16722 10395 16828
rect 10075 16715 10115 16722
rect 10158 16715 10395 16722
rect 10625 16828 10742 16835
rect 10785 16828 10945 16835
rect 10625 16722 10708 16828
rect 10742 16722 10945 16828
rect 10625 16715 10665 16722
rect 10708 16715 10945 16722
rect 11175 16828 11292 16835
rect 11335 16828 11495 16835
rect 11175 16722 11258 16828
rect 11292 16722 11495 16828
rect 11175 16715 11215 16722
rect 11258 16715 11495 16722
rect 11725 16828 11842 16835
rect 11885 16828 12045 16835
rect 11725 16722 11808 16828
rect 11842 16722 12045 16828
rect 11725 16715 11765 16722
rect 11808 16715 12045 16722
rect 12275 16828 12392 16835
rect 12435 16828 12595 16835
rect 12275 16722 12358 16828
rect 12392 16722 12595 16828
rect 12275 16715 12315 16722
rect 12358 16715 12595 16722
rect 12825 16828 12942 16835
rect 12985 16828 13145 16835
rect 12825 16722 12908 16828
rect 12942 16722 13145 16828
rect 12825 16715 12865 16722
rect 12908 16715 13145 16722
rect 13375 16828 13492 16835
rect 13535 16828 13695 16835
rect 13375 16722 13458 16828
rect 13492 16722 13695 16828
rect 13375 16715 13415 16722
rect 13458 16715 13695 16722
rect 13925 16828 14042 16835
rect 14085 16828 14245 16835
rect 13925 16722 14008 16828
rect 14042 16722 14245 16828
rect 13925 16715 13965 16722
rect 14008 16715 14245 16722
rect 14475 16828 14592 16835
rect 14635 16828 14795 16835
rect 14475 16722 14558 16828
rect 14592 16722 14795 16828
rect 14475 16715 14515 16722
rect 14558 16715 14795 16722
rect 15025 16828 15142 16835
rect 15185 16828 15345 16835
rect 15025 16722 15108 16828
rect 15142 16722 15345 16828
rect 15025 16715 15065 16722
rect 15108 16715 15345 16722
rect 15575 16828 15692 16835
rect 15735 16828 15895 16835
rect 15575 16722 15658 16828
rect 15692 16722 15895 16828
rect 15575 16715 15615 16722
rect 15658 16715 15895 16722
rect 16125 16828 16242 16835
rect 16285 16828 16445 16835
rect 16125 16722 16208 16828
rect 16242 16722 16445 16828
rect 16125 16715 16165 16722
rect 16208 16715 16445 16722
rect 16675 16828 16792 16835
rect 16835 16828 16995 16835
rect 16675 16722 16758 16828
rect 16792 16722 16995 16828
rect 16675 16715 16715 16722
rect 16758 16715 16995 16722
rect 17225 16828 17342 16835
rect 17385 16828 17545 16835
rect 17225 16722 17308 16828
rect 17342 16722 17545 16828
rect 17225 16715 17265 16722
rect 17308 16715 17545 16722
rect 17775 16828 17892 16835
rect 17935 16828 18095 16835
rect 17775 16722 17858 16828
rect 17892 16722 18095 16828
rect 17775 16715 17815 16722
rect 17858 16715 18095 16722
rect 18325 16828 18442 16835
rect 18485 16828 18645 16835
rect 18325 16722 18408 16828
rect 18442 16722 18645 16828
rect 18325 16715 18365 16722
rect 18408 16715 18645 16722
rect 18875 16828 18992 16835
rect 19035 16828 19195 16835
rect 18875 16722 18958 16828
rect 18992 16722 19195 16828
rect 18875 16715 18915 16722
rect 18958 16715 19195 16722
rect 765 16675 885 16715
rect 1315 16675 1435 16715
rect 1865 16675 1985 16715
rect 2415 16675 2535 16715
rect 2965 16675 3085 16715
rect 3515 16675 3635 16715
rect 4065 16675 4185 16715
rect 4615 16675 4735 16715
rect 5165 16675 5285 16715
rect 5715 16675 5835 16715
rect 6265 16675 6385 16715
rect 6815 16675 6935 16715
rect 7365 16675 7485 16715
rect 7915 16675 8035 16715
rect 8465 16675 8585 16715
rect 9015 16675 9135 16715
rect 9565 16675 9685 16715
rect 10115 16675 10235 16715
rect 10665 16675 10785 16715
rect 11215 16675 11335 16715
rect 11765 16675 11885 16715
rect 12315 16675 12435 16715
rect 12865 16675 12985 16715
rect 13415 16675 13535 16715
rect 13965 16675 14085 16715
rect 14515 16675 14635 16715
rect 15065 16675 15185 16715
rect 15615 16675 15735 16715
rect 16165 16675 16285 16715
rect 16715 16675 16835 16715
rect 17265 16675 17385 16715
rect 17815 16675 17935 16715
rect 18365 16675 18485 16715
rect 18915 16675 19035 16715
rect 19185 16554 19200 16571
rect 19202 16562 19204 16988
rect 19202 16548 19217 16554
rect 500 16475 507 16525
rect 500 16039 525 16440
rect 628 16422 885 16445
rect 1178 16422 1435 16445
rect 1728 16422 1985 16445
rect 2278 16422 2535 16445
rect 2828 16422 3085 16445
rect 3378 16422 3635 16445
rect 3928 16422 4185 16445
rect 4478 16422 4735 16445
rect 5028 16422 5285 16445
rect 5578 16422 5835 16445
rect 6128 16422 6385 16445
rect 6678 16422 6935 16445
rect 7228 16422 7485 16445
rect 7778 16422 8035 16445
rect 8328 16422 8585 16445
rect 8878 16422 9135 16445
rect 9428 16422 9685 16445
rect 9978 16422 10235 16445
rect 10528 16422 10785 16445
rect 11078 16422 11335 16445
rect 11628 16422 11885 16445
rect 12178 16422 12435 16445
rect 12728 16422 12985 16445
rect 13278 16422 13535 16445
rect 13828 16422 14085 16445
rect 14378 16422 14635 16445
rect 14928 16422 15185 16445
rect 15478 16422 15735 16445
rect 16028 16422 16285 16445
rect 16578 16422 16835 16445
rect 17128 16422 17385 16445
rect 17678 16422 17935 16445
rect 18228 16422 18485 16445
rect 18778 16422 19035 16445
rect 605 16285 609 16422
rect 784 16325 885 16422
rect 765 16285 885 16325
rect 1155 16285 1159 16422
rect 1334 16325 1435 16422
rect 1315 16285 1435 16325
rect 1705 16285 1709 16422
rect 1884 16325 1985 16422
rect 1865 16285 1985 16325
rect 2255 16285 2259 16422
rect 2434 16325 2535 16422
rect 2415 16285 2535 16325
rect 2805 16285 2809 16422
rect 2984 16325 3085 16422
rect 2965 16285 3085 16325
rect 3355 16285 3359 16422
rect 3534 16325 3635 16422
rect 3515 16285 3635 16325
rect 3905 16285 3909 16422
rect 4084 16325 4185 16422
rect 4065 16285 4185 16325
rect 4455 16285 4459 16422
rect 4634 16325 4735 16422
rect 4615 16285 4735 16325
rect 5005 16285 5009 16422
rect 5184 16325 5285 16422
rect 5165 16285 5285 16325
rect 5555 16285 5559 16422
rect 5734 16325 5835 16422
rect 5715 16285 5835 16325
rect 6105 16285 6109 16422
rect 6284 16325 6385 16422
rect 6265 16285 6385 16325
rect 6655 16285 6659 16422
rect 6834 16325 6935 16422
rect 6815 16285 6935 16325
rect 7205 16285 7209 16422
rect 7384 16325 7485 16422
rect 7365 16285 7485 16325
rect 7755 16285 7759 16422
rect 7934 16325 8035 16422
rect 7915 16285 8035 16325
rect 8305 16285 8309 16422
rect 8484 16325 8585 16422
rect 8465 16285 8585 16325
rect 8855 16285 8859 16422
rect 9034 16325 9135 16422
rect 9015 16285 9135 16325
rect 9405 16285 9409 16422
rect 9584 16325 9685 16422
rect 9565 16285 9685 16325
rect 9955 16285 9959 16422
rect 10134 16325 10235 16422
rect 10115 16285 10235 16325
rect 10505 16285 10509 16422
rect 10684 16325 10785 16422
rect 10665 16285 10785 16325
rect 11055 16285 11059 16422
rect 11234 16325 11335 16422
rect 11215 16285 11335 16325
rect 11605 16285 11609 16422
rect 11784 16325 11885 16422
rect 11765 16285 11885 16325
rect 12155 16285 12159 16422
rect 12334 16325 12435 16422
rect 12315 16285 12435 16325
rect 12705 16285 12709 16422
rect 12884 16325 12985 16422
rect 12865 16285 12985 16325
rect 13255 16285 13259 16422
rect 13434 16325 13535 16422
rect 13415 16285 13535 16325
rect 13805 16285 13809 16422
rect 13984 16325 14085 16422
rect 13965 16285 14085 16325
rect 14355 16285 14359 16422
rect 14534 16325 14635 16422
rect 14515 16285 14635 16325
rect 14905 16285 14909 16422
rect 15084 16325 15185 16422
rect 15065 16285 15185 16325
rect 15455 16285 15459 16422
rect 15634 16325 15735 16422
rect 15615 16285 15735 16325
rect 16005 16285 16009 16422
rect 16184 16325 16285 16422
rect 16165 16285 16285 16325
rect 16555 16285 16559 16422
rect 16734 16325 16835 16422
rect 16715 16285 16835 16325
rect 17105 16285 17109 16422
rect 17284 16325 17385 16422
rect 17265 16285 17385 16325
rect 17655 16285 17659 16422
rect 17834 16325 17935 16422
rect 17815 16285 17935 16325
rect 18205 16285 18209 16422
rect 18384 16325 18485 16422
rect 18365 16285 18485 16325
rect 18755 16285 18759 16422
rect 18934 16325 19035 16422
rect 18915 16285 19035 16325
rect 725 16278 842 16285
rect 885 16278 1045 16285
rect 725 16172 808 16278
rect 842 16172 1045 16278
rect 725 16165 765 16172
rect 808 16165 1045 16172
rect 1275 16278 1392 16285
rect 1435 16278 1595 16285
rect 1275 16172 1358 16278
rect 1392 16172 1595 16278
rect 1275 16165 1315 16172
rect 1358 16165 1595 16172
rect 1825 16278 1942 16285
rect 1985 16278 2145 16285
rect 1825 16172 1908 16278
rect 1942 16172 2145 16278
rect 1825 16165 1865 16172
rect 1908 16165 2145 16172
rect 2375 16278 2492 16285
rect 2535 16278 2695 16285
rect 2375 16172 2458 16278
rect 2492 16172 2695 16278
rect 2375 16165 2415 16172
rect 2458 16165 2695 16172
rect 2925 16278 3042 16285
rect 3085 16278 3245 16285
rect 2925 16172 3008 16278
rect 3042 16172 3245 16278
rect 2925 16165 2965 16172
rect 3008 16165 3245 16172
rect 3475 16278 3592 16285
rect 3635 16278 3795 16285
rect 3475 16172 3558 16278
rect 3592 16172 3795 16278
rect 3475 16165 3515 16172
rect 3558 16165 3795 16172
rect 4025 16278 4142 16285
rect 4185 16278 4345 16285
rect 4025 16172 4108 16278
rect 4142 16172 4345 16278
rect 4025 16165 4065 16172
rect 4108 16165 4345 16172
rect 4575 16278 4692 16285
rect 4735 16278 4895 16285
rect 4575 16172 4658 16278
rect 4692 16172 4895 16278
rect 4575 16165 4615 16172
rect 4658 16165 4895 16172
rect 5125 16278 5242 16285
rect 5285 16278 5445 16285
rect 5125 16172 5208 16278
rect 5242 16172 5445 16278
rect 5125 16165 5165 16172
rect 5208 16165 5445 16172
rect 5675 16278 5792 16285
rect 5835 16278 5995 16285
rect 5675 16172 5758 16278
rect 5792 16172 5995 16278
rect 5675 16165 5715 16172
rect 5758 16165 5995 16172
rect 6225 16278 6342 16285
rect 6385 16278 6545 16285
rect 6225 16172 6308 16278
rect 6342 16172 6545 16278
rect 6225 16165 6265 16172
rect 6308 16165 6545 16172
rect 6775 16278 6892 16285
rect 6935 16278 7095 16285
rect 6775 16172 6858 16278
rect 6892 16172 7095 16278
rect 6775 16165 6815 16172
rect 6858 16165 7095 16172
rect 7325 16278 7442 16285
rect 7485 16278 7645 16285
rect 7325 16172 7408 16278
rect 7442 16172 7645 16278
rect 7325 16165 7365 16172
rect 7408 16165 7645 16172
rect 7875 16278 7992 16285
rect 8035 16278 8195 16285
rect 7875 16172 7958 16278
rect 7992 16172 8195 16278
rect 7875 16165 7915 16172
rect 7958 16165 8195 16172
rect 8425 16278 8542 16285
rect 8585 16278 8745 16285
rect 8425 16172 8508 16278
rect 8542 16172 8745 16278
rect 8425 16165 8465 16172
rect 8508 16165 8745 16172
rect 8975 16278 9092 16285
rect 9135 16278 9295 16285
rect 8975 16172 9058 16278
rect 9092 16172 9295 16278
rect 8975 16165 9015 16172
rect 9058 16165 9295 16172
rect 9525 16278 9642 16285
rect 9685 16278 9845 16285
rect 9525 16172 9608 16278
rect 9642 16172 9845 16278
rect 9525 16165 9565 16172
rect 9608 16165 9845 16172
rect 10075 16278 10192 16285
rect 10235 16278 10395 16285
rect 10075 16172 10158 16278
rect 10192 16172 10395 16278
rect 10075 16165 10115 16172
rect 10158 16165 10395 16172
rect 10625 16278 10742 16285
rect 10785 16278 10945 16285
rect 10625 16172 10708 16278
rect 10742 16172 10945 16278
rect 10625 16165 10665 16172
rect 10708 16165 10945 16172
rect 11175 16278 11292 16285
rect 11335 16278 11495 16285
rect 11175 16172 11258 16278
rect 11292 16172 11495 16278
rect 11175 16165 11215 16172
rect 11258 16165 11495 16172
rect 11725 16278 11842 16285
rect 11885 16278 12045 16285
rect 11725 16172 11808 16278
rect 11842 16172 12045 16278
rect 11725 16165 11765 16172
rect 11808 16165 12045 16172
rect 12275 16278 12392 16285
rect 12435 16278 12595 16285
rect 12275 16172 12358 16278
rect 12392 16172 12595 16278
rect 12275 16165 12315 16172
rect 12358 16165 12595 16172
rect 12825 16278 12942 16285
rect 12985 16278 13145 16285
rect 12825 16172 12908 16278
rect 12942 16172 13145 16278
rect 12825 16165 12865 16172
rect 12908 16165 13145 16172
rect 13375 16278 13492 16285
rect 13535 16278 13695 16285
rect 13375 16172 13458 16278
rect 13492 16172 13695 16278
rect 13375 16165 13415 16172
rect 13458 16165 13695 16172
rect 13925 16278 14042 16285
rect 14085 16278 14245 16285
rect 13925 16172 14008 16278
rect 14042 16172 14245 16278
rect 13925 16165 13965 16172
rect 14008 16165 14245 16172
rect 14475 16278 14592 16285
rect 14635 16278 14795 16285
rect 14475 16172 14558 16278
rect 14592 16172 14795 16278
rect 14475 16165 14515 16172
rect 14558 16165 14795 16172
rect 15025 16278 15142 16285
rect 15185 16278 15345 16285
rect 15025 16172 15108 16278
rect 15142 16172 15345 16278
rect 15025 16165 15065 16172
rect 15108 16165 15345 16172
rect 15575 16278 15692 16285
rect 15735 16278 15895 16285
rect 15575 16172 15658 16278
rect 15692 16172 15895 16278
rect 15575 16165 15615 16172
rect 15658 16165 15895 16172
rect 16125 16278 16242 16285
rect 16285 16278 16445 16285
rect 16125 16172 16208 16278
rect 16242 16172 16445 16278
rect 16125 16165 16165 16172
rect 16208 16165 16445 16172
rect 16675 16278 16792 16285
rect 16835 16278 16995 16285
rect 16675 16172 16758 16278
rect 16792 16172 16995 16278
rect 16675 16165 16715 16172
rect 16758 16165 16995 16172
rect 17225 16278 17342 16285
rect 17385 16278 17545 16285
rect 17225 16172 17308 16278
rect 17342 16172 17545 16278
rect 17225 16165 17265 16172
rect 17308 16165 17545 16172
rect 17775 16278 17892 16285
rect 17935 16278 18095 16285
rect 17775 16172 17858 16278
rect 17892 16172 18095 16278
rect 17775 16165 17815 16172
rect 17858 16165 18095 16172
rect 18325 16278 18442 16285
rect 18485 16278 18645 16285
rect 18325 16172 18408 16278
rect 18442 16172 18645 16278
rect 18325 16165 18365 16172
rect 18408 16165 18645 16172
rect 18875 16278 18992 16285
rect 19035 16278 19195 16285
rect 18875 16172 18958 16278
rect 18992 16172 19195 16278
rect 18875 16165 18915 16172
rect 18958 16165 19195 16172
rect 765 16125 885 16165
rect 1315 16125 1435 16165
rect 1865 16125 1985 16165
rect 2415 16125 2535 16165
rect 2965 16125 3085 16165
rect 3515 16125 3635 16165
rect 4065 16125 4185 16165
rect 4615 16125 4735 16165
rect 5165 16125 5285 16165
rect 5715 16125 5835 16165
rect 6265 16125 6385 16165
rect 6815 16125 6935 16165
rect 7365 16125 7485 16165
rect 7915 16125 8035 16165
rect 8465 16125 8585 16165
rect 9015 16125 9135 16165
rect 9565 16125 9685 16165
rect 10115 16125 10235 16165
rect 10665 16125 10785 16165
rect 11215 16125 11335 16165
rect 11765 16125 11885 16165
rect 12315 16125 12435 16165
rect 12865 16125 12985 16165
rect 13415 16125 13535 16165
rect 13965 16125 14085 16165
rect 14515 16125 14635 16165
rect 15065 16125 15185 16165
rect 15615 16125 15735 16165
rect 16165 16125 16285 16165
rect 16715 16125 16835 16165
rect 17265 16125 17385 16165
rect 17815 16125 17935 16165
rect 18365 16125 18485 16165
rect 18915 16125 19035 16165
rect 19202 16012 19204 16438
rect 500 15925 507 15975
rect 19202 15896 19217 15902
rect 628 15872 885 15895
rect 1178 15872 1435 15895
rect 1728 15872 1985 15895
rect 2278 15872 2535 15895
rect 2828 15872 3085 15895
rect 3378 15872 3635 15895
rect 3928 15872 4185 15895
rect 4478 15872 4735 15895
rect 5028 15872 5285 15895
rect 5578 15872 5835 15895
rect 6128 15872 6385 15895
rect 6678 15872 6935 15895
rect 7228 15872 7485 15895
rect 7778 15872 8035 15895
rect 8328 15872 8585 15895
rect 8878 15872 9135 15895
rect 9428 15872 9685 15895
rect 9978 15872 10235 15895
rect 10528 15872 10785 15895
rect 11078 15872 11335 15895
rect 11628 15872 11885 15895
rect 12178 15872 12435 15895
rect 12728 15872 12985 15895
rect 13278 15872 13535 15895
rect 13828 15872 14085 15895
rect 14378 15872 14635 15895
rect 14928 15872 15185 15895
rect 15478 15872 15735 15895
rect 16028 15872 16285 15895
rect 16578 15872 16835 15895
rect 17128 15872 17385 15895
rect 17678 15872 17935 15895
rect 18228 15872 18485 15895
rect 18778 15872 19035 15895
rect 605 15735 609 15872
rect 784 15775 885 15872
rect 765 15735 885 15775
rect 1155 15735 1159 15872
rect 1334 15775 1435 15872
rect 1315 15735 1435 15775
rect 1705 15735 1709 15872
rect 1884 15775 1985 15872
rect 1865 15735 1985 15775
rect 2255 15735 2259 15872
rect 2434 15775 2535 15872
rect 2415 15735 2535 15775
rect 2805 15735 2809 15872
rect 2984 15775 3085 15872
rect 2965 15735 3085 15775
rect 3355 15735 3359 15872
rect 3534 15775 3635 15872
rect 3515 15735 3635 15775
rect 3905 15735 3909 15872
rect 4084 15775 4185 15872
rect 4065 15735 4185 15775
rect 4455 15735 4459 15872
rect 4634 15775 4735 15872
rect 4615 15735 4735 15775
rect 5005 15735 5009 15872
rect 5184 15775 5285 15872
rect 5165 15735 5285 15775
rect 5555 15735 5559 15872
rect 5734 15775 5835 15872
rect 5715 15735 5835 15775
rect 6105 15735 6109 15872
rect 6284 15775 6385 15872
rect 6265 15735 6385 15775
rect 6655 15735 6659 15872
rect 6834 15775 6935 15872
rect 6815 15735 6935 15775
rect 7205 15735 7209 15872
rect 7384 15775 7485 15872
rect 7365 15735 7485 15775
rect 7755 15735 7759 15872
rect 7934 15775 8035 15872
rect 7915 15735 8035 15775
rect 8305 15735 8309 15872
rect 8484 15775 8585 15872
rect 8465 15735 8585 15775
rect 8855 15735 8859 15872
rect 9034 15775 9135 15872
rect 9015 15735 9135 15775
rect 9405 15735 9409 15872
rect 9584 15775 9685 15872
rect 9565 15735 9685 15775
rect 9955 15735 9959 15872
rect 10134 15775 10235 15872
rect 10115 15735 10235 15775
rect 10505 15735 10509 15872
rect 10684 15775 10785 15872
rect 10665 15735 10785 15775
rect 11055 15735 11059 15872
rect 11234 15775 11335 15872
rect 11215 15735 11335 15775
rect 11605 15735 11609 15872
rect 11784 15775 11885 15872
rect 11765 15735 11885 15775
rect 12155 15735 12159 15872
rect 12334 15775 12435 15872
rect 12315 15735 12435 15775
rect 12705 15735 12709 15872
rect 12884 15775 12985 15872
rect 12865 15735 12985 15775
rect 13255 15735 13259 15872
rect 13434 15775 13535 15872
rect 13415 15735 13535 15775
rect 13805 15735 13809 15872
rect 13984 15775 14085 15872
rect 13965 15735 14085 15775
rect 14355 15735 14359 15872
rect 14534 15775 14635 15872
rect 14515 15735 14635 15775
rect 14905 15735 14909 15872
rect 15084 15775 15185 15872
rect 15065 15735 15185 15775
rect 15455 15735 15459 15872
rect 15634 15775 15735 15872
rect 15615 15735 15735 15775
rect 16005 15735 16009 15872
rect 16184 15775 16285 15872
rect 16165 15735 16285 15775
rect 16555 15735 16559 15872
rect 16734 15775 16835 15872
rect 16715 15735 16835 15775
rect 17105 15735 17109 15872
rect 17284 15775 17385 15872
rect 17265 15735 17385 15775
rect 17655 15735 17659 15872
rect 17834 15775 17935 15872
rect 17815 15735 17935 15775
rect 18205 15735 18209 15872
rect 18384 15775 18485 15872
rect 18365 15735 18485 15775
rect 18755 15735 18759 15872
rect 18934 15775 19035 15872
rect 18915 15735 19035 15775
rect 725 15728 842 15735
rect 885 15728 1045 15735
rect 725 15622 808 15728
rect 842 15622 1045 15728
rect 725 15615 765 15622
rect 808 15615 1045 15622
rect 1275 15728 1392 15735
rect 1435 15728 1595 15735
rect 1275 15622 1358 15728
rect 1392 15622 1595 15728
rect 1275 15615 1315 15622
rect 1358 15615 1595 15622
rect 1825 15728 1942 15735
rect 1985 15728 2145 15735
rect 1825 15622 1908 15728
rect 1942 15622 2145 15728
rect 1825 15615 1865 15622
rect 1908 15615 2145 15622
rect 2375 15728 2492 15735
rect 2535 15728 2695 15735
rect 2375 15622 2458 15728
rect 2492 15622 2695 15728
rect 2375 15615 2415 15622
rect 2458 15615 2695 15622
rect 2925 15728 3042 15735
rect 3085 15728 3245 15735
rect 2925 15622 3008 15728
rect 3042 15622 3245 15728
rect 2925 15615 2965 15622
rect 3008 15615 3245 15622
rect 3475 15728 3592 15735
rect 3635 15728 3795 15735
rect 3475 15622 3558 15728
rect 3592 15622 3795 15728
rect 3475 15615 3515 15622
rect 3558 15615 3795 15622
rect 4025 15728 4142 15735
rect 4185 15728 4345 15735
rect 4025 15622 4108 15728
rect 4142 15622 4345 15728
rect 4025 15615 4065 15622
rect 4108 15615 4345 15622
rect 4575 15728 4692 15735
rect 4735 15728 4895 15735
rect 4575 15622 4658 15728
rect 4692 15622 4895 15728
rect 4575 15615 4615 15622
rect 4658 15615 4895 15622
rect 5125 15728 5242 15735
rect 5285 15728 5445 15735
rect 5125 15622 5208 15728
rect 5242 15622 5445 15728
rect 5125 15615 5165 15622
rect 5208 15615 5445 15622
rect 5675 15728 5792 15735
rect 5835 15728 5995 15735
rect 5675 15622 5758 15728
rect 5792 15622 5995 15728
rect 5675 15615 5715 15622
rect 5758 15615 5995 15622
rect 6225 15728 6342 15735
rect 6385 15728 6545 15735
rect 6225 15622 6308 15728
rect 6342 15622 6545 15728
rect 6225 15615 6265 15622
rect 6308 15615 6545 15622
rect 6775 15728 6892 15735
rect 6935 15728 7095 15735
rect 6775 15622 6858 15728
rect 6892 15622 7095 15728
rect 6775 15615 6815 15622
rect 6858 15615 7095 15622
rect 7325 15728 7442 15735
rect 7485 15728 7645 15735
rect 7325 15622 7408 15728
rect 7442 15622 7645 15728
rect 7325 15615 7365 15622
rect 7408 15615 7645 15622
rect 7875 15728 7992 15735
rect 8035 15728 8195 15735
rect 7875 15622 7958 15728
rect 7992 15622 8195 15728
rect 7875 15615 7915 15622
rect 7958 15615 8195 15622
rect 8425 15728 8542 15735
rect 8585 15728 8745 15735
rect 8425 15622 8508 15728
rect 8542 15622 8745 15728
rect 8425 15615 8465 15622
rect 8508 15615 8745 15622
rect 8975 15728 9092 15735
rect 9135 15728 9295 15735
rect 8975 15622 9058 15728
rect 9092 15622 9295 15728
rect 8975 15615 9015 15622
rect 9058 15615 9295 15622
rect 9525 15728 9642 15735
rect 9685 15728 9845 15735
rect 9525 15622 9608 15728
rect 9642 15622 9845 15728
rect 9525 15615 9565 15622
rect 9608 15615 9845 15622
rect 10075 15728 10192 15735
rect 10235 15728 10395 15735
rect 10075 15622 10158 15728
rect 10192 15622 10395 15728
rect 10075 15615 10115 15622
rect 10158 15615 10395 15622
rect 10625 15728 10742 15735
rect 10785 15728 10945 15735
rect 10625 15622 10708 15728
rect 10742 15622 10945 15728
rect 10625 15615 10665 15622
rect 10708 15615 10945 15622
rect 11175 15728 11292 15735
rect 11335 15728 11495 15735
rect 11175 15622 11258 15728
rect 11292 15622 11495 15728
rect 11175 15615 11215 15622
rect 11258 15615 11495 15622
rect 11725 15728 11842 15735
rect 11885 15728 12045 15735
rect 11725 15622 11808 15728
rect 11842 15622 12045 15728
rect 11725 15615 11765 15622
rect 11808 15615 12045 15622
rect 12275 15728 12392 15735
rect 12435 15728 12595 15735
rect 12275 15622 12358 15728
rect 12392 15622 12595 15728
rect 12275 15615 12315 15622
rect 12358 15615 12595 15622
rect 12825 15728 12942 15735
rect 12985 15728 13145 15735
rect 12825 15622 12908 15728
rect 12942 15622 13145 15728
rect 12825 15615 12865 15622
rect 12908 15615 13145 15622
rect 13375 15728 13492 15735
rect 13535 15728 13695 15735
rect 13375 15622 13458 15728
rect 13492 15622 13695 15728
rect 13375 15615 13415 15622
rect 13458 15615 13695 15622
rect 13925 15728 14042 15735
rect 14085 15728 14245 15735
rect 13925 15622 14008 15728
rect 14042 15622 14245 15728
rect 13925 15615 13965 15622
rect 14008 15615 14245 15622
rect 14475 15728 14592 15735
rect 14635 15728 14795 15735
rect 14475 15622 14558 15728
rect 14592 15622 14795 15728
rect 14475 15615 14515 15622
rect 14558 15615 14795 15622
rect 15025 15728 15142 15735
rect 15185 15728 15345 15735
rect 15025 15622 15108 15728
rect 15142 15622 15345 15728
rect 15025 15615 15065 15622
rect 15108 15615 15345 15622
rect 15575 15728 15692 15735
rect 15735 15728 15895 15735
rect 15575 15622 15658 15728
rect 15692 15622 15895 15728
rect 15575 15615 15615 15622
rect 15658 15615 15895 15622
rect 16125 15728 16242 15735
rect 16285 15728 16445 15735
rect 16125 15622 16208 15728
rect 16242 15622 16445 15728
rect 16125 15615 16165 15622
rect 16208 15615 16445 15622
rect 16675 15728 16792 15735
rect 16835 15728 16995 15735
rect 16675 15622 16758 15728
rect 16792 15622 16995 15728
rect 16675 15615 16715 15622
rect 16758 15615 16995 15622
rect 17225 15728 17342 15735
rect 17385 15728 17545 15735
rect 17225 15622 17308 15728
rect 17342 15622 17545 15728
rect 17225 15615 17265 15622
rect 17308 15615 17545 15622
rect 17775 15728 17892 15735
rect 17935 15728 18095 15735
rect 17775 15622 17858 15728
rect 17892 15622 18095 15728
rect 17775 15615 17815 15622
rect 17858 15615 18095 15622
rect 18325 15728 18442 15735
rect 18485 15728 18645 15735
rect 18325 15622 18408 15728
rect 18442 15622 18645 15728
rect 18325 15615 18365 15622
rect 18408 15615 18645 15622
rect 18875 15728 18992 15735
rect 19035 15728 19195 15735
rect 18875 15622 18958 15728
rect 18992 15622 19195 15728
rect 18875 15615 18915 15622
rect 18958 15615 19195 15622
rect 765 15575 885 15615
rect 1315 15575 1435 15615
rect 1865 15575 1985 15615
rect 2415 15575 2535 15615
rect 2965 15575 3085 15615
rect 3515 15575 3635 15615
rect 4065 15575 4185 15615
rect 4615 15575 4735 15615
rect 5165 15575 5285 15615
rect 5715 15575 5835 15615
rect 6265 15575 6385 15615
rect 6815 15575 6935 15615
rect 7365 15575 7485 15615
rect 7915 15575 8035 15615
rect 8465 15575 8585 15615
rect 9015 15575 9135 15615
rect 9565 15575 9685 15615
rect 10115 15575 10235 15615
rect 10665 15575 10785 15615
rect 11215 15575 11335 15615
rect 11765 15575 11885 15615
rect 12315 15575 12435 15615
rect 12865 15575 12985 15615
rect 13415 15575 13535 15615
rect 13965 15575 14085 15615
rect 14515 15575 14635 15615
rect 15065 15575 15185 15615
rect 15615 15575 15735 15615
rect 16165 15575 16285 15615
rect 16715 15575 16835 15615
rect 17265 15575 17385 15615
rect 17815 15575 17935 15615
rect 18365 15575 18485 15615
rect 18915 15575 19035 15615
rect 19185 15454 19200 15471
rect 19202 15462 19204 15888
rect 19202 15448 19217 15454
rect 500 15375 507 15425
rect 500 14939 525 15340
rect 628 15322 885 15345
rect 1178 15322 1435 15345
rect 1728 15322 1985 15345
rect 2278 15322 2535 15345
rect 2828 15322 3085 15345
rect 3378 15322 3635 15345
rect 3928 15322 4185 15345
rect 4478 15322 4735 15345
rect 5028 15322 5285 15345
rect 5578 15322 5835 15345
rect 6128 15322 6385 15345
rect 6678 15322 6935 15345
rect 7228 15322 7485 15345
rect 7778 15322 8035 15345
rect 8328 15322 8585 15345
rect 8878 15322 9135 15345
rect 9428 15322 9685 15345
rect 9978 15322 10235 15345
rect 10528 15322 10785 15345
rect 11078 15322 11335 15345
rect 11628 15322 11885 15345
rect 12178 15322 12435 15345
rect 12728 15322 12985 15345
rect 13278 15322 13535 15345
rect 13828 15322 14085 15345
rect 14378 15322 14635 15345
rect 14928 15322 15185 15345
rect 15478 15322 15735 15345
rect 16028 15322 16285 15345
rect 16578 15322 16835 15345
rect 17128 15322 17385 15345
rect 17678 15322 17935 15345
rect 18228 15322 18485 15345
rect 18778 15322 19035 15345
rect 605 15185 609 15322
rect 784 15225 885 15322
rect 765 15185 885 15225
rect 1155 15185 1159 15322
rect 1334 15225 1435 15322
rect 1315 15185 1435 15225
rect 1705 15185 1709 15322
rect 1884 15225 1985 15322
rect 1865 15185 1985 15225
rect 2255 15185 2259 15322
rect 2434 15225 2535 15322
rect 2415 15185 2535 15225
rect 2805 15185 2809 15322
rect 2984 15225 3085 15322
rect 2965 15185 3085 15225
rect 3355 15185 3359 15322
rect 3534 15225 3635 15322
rect 3515 15185 3635 15225
rect 3905 15185 3909 15322
rect 4084 15225 4185 15322
rect 4065 15185 4185 15225
rect 4455 15185 4459 15322
rect 4634 15225 4735 15322
rect 4615 15185 4735 15225
rect 5005 15185 5009 15322
rect 5184 15225 5285 15322
rect 5165 15185 5285 15225
rect 5555 15185 5559 15322
rect 5734 15225 5835 15322
rect 5715 15185 5835 15225
rect 6105 15185 6109 15322
rect 6284 15225 6385 15322
rect 6265 15185 6385 15225
rect 6655 15185 6659 15322
rect 6834 15225 6935 15322
rect 6815 15185 6935 15225
rect 7205 15185 7209 15322
rect 7384 15225 7485 15322
rect 7365 15185 7485 15225
rect 7755 15185 7759 15322
rect 7934 15225 8035 15322
rect 7915 15185 8035 15225
rect 8305 15185 8309 15322
rect 8484 15225 8585 15322
rect 8465 15185 8585 15225
rect 8855 15185 8859 15322
rect 9034 15225 9135 15322
rect 9015 15185 9135 15225
rect 9405 15185 9409 15322
rect 9584 15225 9685 15322
rect 9565 15185 9685 15225
rect 9955 15185 9959 15322
rect 10134 15225 10235 15322
rect 10115 15185 10235 15225
rect 10505 15185 10509 15322
rect 10684 15225 10785 15322
rect 10665 15185 10785 15225
rect 11055 15185 11059 15322
rect 11234 15225 11335 15322
rect 11215 15185 11335 15225
rect 11605 15185 11609 15322
rect 11784 15225 11885 15322
rect 11765 15185 11885 15225
rect 12155 15185 12159 15322
rect 12334 15225 12435 15322
rect 12315 15185 12435 15225
rect 12705 15185 12709 15322
rect 12884 15225 12985 15322
rect 12865 15185 12985 15225
rect 13255 15185 13259 15322
rect 13434 15225 13535 15322
rect 13415 15185 13535 15225
rect 13805 15185 13809 15322
rect 13984 15225 14085 15322
rect 13965 15185 14085 15225
rect 14355 15185 14359 15322
rect 14534 15225 14635 15322
rect 14515 15185 14635 15225
rect 14905 15185 14909 15322
rect 15084 15225 15185 15322
rect 15065 15185 15185 15225
rect 15455 15185 15459 15322
rect 15634 15225 15735 15322
rect 15615 15185 15735 15225
rect 16005 15185 16009 15322
rect 16184 15225 16285 15322
rect 16165 15185 16285 15225
rect 16555 15185 16559 15322
rect 16734 15225 16835 15322
rect 16715 15185 16835 15225
rect 17105 15185 17109 15322
rect 17284 15225 17385 15322
rect 17265 15185 17385 15225
rect 17655 15185 17659 15322
rect 17834 15225 17935 15322
rect 17815 15185 17935 15225
rect 18205 15185 18209 15322
rect 18384 15225 18485 15322
rect 18365 15185 18485 15225
rect 18755 15185 18759 15322
rect 18934 15225 19035 15322
rect 18915 15185 19035 15225
rect 725 15178 842 15185
rect 885 15178 1045 15185
rect 725 15072 808 15178
rect 842 15072 1045 15178
rect 725 15065 765 15072
rect 808 15065 1045 15072
rect 1275 15178 1392 15185
rect 1435 15178 1595 15185
rect 1275 15072 1358 15178
rect 1392 15072 1595 15178
rect 1275 15065 1315 15072
rect 1358 15065 1595 15072
rect 1825 15178 1942 15185
rect 1985 15178 2145 15185
rect 1825 15072 1908 15178
rect 1942 15072 2145 15178
rect 1825 15065 1865 15072
rect 1908 15065 2145 15072
rect 2375 15178 2492 15185
rect 2535 15178 2695 15185
rect 2375 15072 2458 15178
rect 2492 15072 2695 15178
rect 2375 15065 2415 15072
rect 2458 15065 2695 15072
rect 2925 15178 3042 15185
rect 3085 15178 3245 15185
rect 2925 15072 3008 15178
rect 3042 15072 3245 15178
rect 2925 15065 2965 15072
rect 3008 15065 3245 15072
rect 3475 15178 3592 15185
rect 3635 15178 3795 15185
rect 3475 15072 3558 15178
rect 3592 15072 3795 15178
rect 3475 15065 3515 15072
rect 3558 15065 3795 15072
rect 4025 15178 4142 15185
rect 4185 15178 4345 15185
rect 4025 15072 4108 15178
rect 4142 15072 4345 15178
rect 4025 15065 4065 15072
rect 4108 15065 4345 15072
rect 4575 15178 4692 15185
rect 4735 15178 4895 15185
rect 4575 15072 4658 15178
rect 4692 15072 4895 15178
rect 4575 15065 4615 15072
rect 4658 15065 4895 15072
rect 5125 15178 5242 15185
rect 5285 15178 5445 15185
rect 5125 15072 5208 15178
rect 5242 15072 5445 15178
rect 5125 15065 5165 15072
rect 5208 15065 5445 15072
rect 5675 15178 5792 15185
rect 5835 15178 5995 15185
rect 5675 15072 5758 15178
rect 5792 15072 5995 15178
rect 5675 15065 5715 15072
rect 5758 15065 5995 15072
rect 6225 15178 6342 15185
rect 6385 15178 6545 15185
rect 6225 15072 6308 15178
rect 6342 15072 6545 15178
rect 6225 15065 6265 15072
rect 6308 15065 6545 15072
rect 6775 15178 6892 15185
rect 6935 15178 7095 15185
rect 6775 15072 6858 15178
rect 6892 15072 7095 15178
rect 6775 15065 6815 15072
rect 6858 15065 7095 15072
rect 7325 15178 7442 15185
rect 7485 15178 7645 15185
rect 7325 15072 7408 15178
rect 7442 15072 7645 15178
rect 7325 15065 7365 15072
rect 7408 15065 7645 15072
rect 7875 15178 7992 15185
rect 8035 15178 8195 15185
rect 7875 15072 7958 15178
rect 7992 15072 8195 15178
rect 7875 15065 7915 15072
rect 7958 15065 8195 15072
rect 8425 15178 8542 15185
rect 8585 15178 8745 15185
rect 8425 15072 8508 15178
rect 8542 15072 8745 15178
rect 8425 15065 8465 15072
rect 8508 15065 8745 15072
rect 8975 15178 9092 15185
rect 9135 15178 9295 15185
rect 8975 15072 9058 15178
rect 9092 15072 9295 15178
rect 8975 15065 9015 15072
rect 9058 15065 9295 15072
rect 9525 15178 9642 15185
rect 9685 15178 9845 15185
rect 9525 15072 9608 15178
rect 9642 15072 9845 15178
rect 9525 15065 9565 15072
rect 9608 15065 9845 15072
rect 10075 15178 10192 15185
rect 10235 15178 10395 15185
rect 10075 15072 10158 15178
rect 10192 15072 10395 15178
rect 10075 15065 10115 15072
rect 10158 15065 10395 15072
rect 10625 15178 10742 15185
rect 10785 15178 10945 15185
rect 10625 15072 10708 15178
rect 10742 15072 10945 15178
rect 10625 15065 10665 15072
rect 10708 15065 10945 15072
rect 11175 15178 11292 15185
rect 11335 15178 11495 15185
rect 11175 15072 11258 15178
rect 11292 15072 11495 15178
rect 11175 15065 11215 15072
rect 11258 15065 11495 15072
rect 11725 15178 11842 15185
rect 11885 15178 12045 15185
rect 11725 15072 11808 15178
rect 11842 15072 12045 15178
rect 11725 15065 11765 15072
rect 11808 15065 12045 15072
rect 12275 15178 12392 15185
rect 12435 15178 12595 15185
rect 12275 15072 12358 15178
rect 12392 15072 12595 15178
rect 12275 15065 12315 15072
rect 12358 15065 12595 15072
rect 12825 15178 12942 15185
rect 12985 15178 13145 15185
rect 12825 15072 12908 15178
rect 12942 15072 13145 15178
rect 12825 15065 12865 15072
rect 12908 15065 13145 15072
rect 13375 15178 13492 15185
rect 13535 15178 13695 15185
rect 13375 15072 13458 15178
rect 13492 15072 13695 15178
rect 13375 15065 13415 15072
rect 13458 15065 13695 15072
rect 13925 15178 14042 15185
rect 14085 15178 14245 15185
rect 13925 15072 14008 15178
rect 14042 15072 14245 15178
rect 13925 15065 13965 15072
rect 14008 15065 14245 15072
rect 14475 15178 14592 15185
rect 14635 15178 14795 15185
rect 14475 15072 14558 15178
rect 14592 15072 14795 15178
rect 14475 15065 14515 15072
rect 14558 15065 14795 15072
rect 15025 15178 15142 15185
rect 15185 15178 15345 15185
rect 15025 15072 15108 15178
rect 15142 15072 15345 15178
rect 15025 15065 15065 15072
rect 15108 15065 15345 15072
rect 15575 15178 15692 15185
rect 15735 15178 15895 15185
rect 15575 15072 15658 15178
rect 15692 15072 15895 15178
rect 15575 15065 15615 15072
rect 15658 15065 15895 15072
rect 16125 15178 16242 15185
rect 16285 15178 16445 15185
rect 16125 15072 16208 15178
rect 16242 15072 16445 15178
rect 16125 15065 16165 15072
rect 16208 15065 16445 15072
rect 16675 15178 16792 15185
rect 16835 15178 16995 15185
rect 16675 15072 16758 15178
rect 16792 15072 16995 15178
rect 16675 15065 16715 15072
rect 16758 15065 16995 15072
rect 17225 15178 17342 15185
rect 17385 15178 17545 15185
rect 17225 15072 17308 15178
rect 17342 15072 17545 15178
rect 17225 15065 17265 15072
rect 17308 15065 17545 15072
rect 17775 15178 17892 15185
rect 17935 15178 18095 15185
rect 17775 15072 17858 15178
rect 17892 15072 18095 15178
rect 17775 15065 17815 15072
rect 17858 15065 18095 15072
rect 18325 15178 18442 15185
rect 18485 15178 18645 15185
rect 18325 15072 18408 15178
rect 18442 15072 18645 15178
rect 18325 15065 18365 15072
rect 18408 15065 18645 15072
rect 18875 15178 18992 15185
rect 19035 15178 19195 15185
rect 18875 15072 18958 15178
rect 18992 15072 19195 15178
rect 18875 15065 18915 15072
rect 18958 15065 19195 15072
rect 765 15025 885 15065
rect 1315 15025 1435 15065
rect 1865 15025 1985 15065
rect 2415 15025 2535 15065
rect 2965 15025 3085 15065
rect 3515 15025 3635 15065
rect 4065 15025 4185 15065
rect 4615 15025 4735 15065
rect 5165 15025 5285 15065
rect 5715 15025 5835 15065
rect 6265 15025 6385 15065
rect 6815 15025 6935 15065
rect 7365 15025 7485 15065
rect 7915 15025 8035 15065
rect 8465 15025 8585 15065
rect 9015 15025 9135 15065
rect 9565 15025 9685 15065
rect 10115 15025 10235 15065
rect 10665 15025 10785 15065
rect 11215 15025 11335 15065
rect 11765 15025 11885 15065
rect 12315 15025 12435 15065
rect 12865 15025 12985 15065
rect 13415 15025 13535 15065
rect 13965 15025 14085 15065
rect 14515 15025 14635 15065
rect 15065 15025 15185 15065
rect 15615 15025 15735 15065
rect 16165 15025 16285 15065
rect 16715 15025 16835 15065
rect 17265 15025 17385 15065
rect 17815 15025 17935 15065
rect 18365 15025 18485 15065
rect 18915 15025 19035 15065
rect 19202 14912 19204 15338
rect 500 14825 507 14875
rect 19202 14796 19217 14802
rect 628 14772 885 14795
rect 1178 14772 1435 14795
rect 1728 14772 1985 14795
rect 2278 14772 2535 14795
rect 2828 14772 3085 14795
rect 3378 14772 3635 14795
rect 3928 14772 4185 14795
rect 4478 14772 4735 14795
rect 5028 14772 5285 14795
rect 5578 14772 5835 14795
rect 6128 14772 6385 14795
rect 6678 14772 6935 14795
rect 7228 14772 7485 14795
rect 7778 14772 8035 14795
rect 8328 14772 8585 14795
rect 8878 14772 9135 14795
rect 9428 14772 9685 14795
rect 9978 14772 10235 14795
rect 10528 14772 10785 14795
rect 11078 14772 11335 14795
rect 11628 14772 11885 14795
rect 12178 14772 12435 14795
rect 12728 14772 12985 14795
rect 13278 14772 13535 14795
rect 13828 14772 14085 14795
rect 14378 14772 14635 14795
rect 14928 14772 15185 14795
rect 15478 14772 15735 14795
rect 16028 14772 16285 14795
rect 16578 14772 16835 14795
rect 17128 14772 17385 14795
rect 17678 14772 17935 14795
rect 18228 14772 18485 14795
rect 18778 14772 19035 14795
rect 605 14635 609 14772
rect 784 14675 885 14772
rect 765 14635 885 14675
rect 1155 14635 1159 14772
rect 1334 14675 1435 14772
rect 1315 14635 1435 14675
rect 1705 14635 1709 14772
rect 1884 14675 1985 14772
rect 1865 14635 1985 14675
rect 2255 14635 2259 14772
rect 2434 14675 2535 14772
rect 2415 14635 2535 14675
rect 2805 14635 2809 14772
rect 2984 14675 3085 14772
rect 2965 14635 3085 14675
rect 3355 14635 3359 14772
rect 3534 14675 3635 14772
rect 3515 14635 3635 14675
rect 3905 14635 3909 14772
rect 4084 14675 4185 14772
rect 4065 14635 4185 14675
rect 4455 14635 4459 14772
rect 4634 14675 4735 14772
rect 4615 14635 4735 14675
rect 5005 14635 5009 14772
rect 5184 14675 5285 14772
rect 5165 14635 5285 14675
rect 5555 14635 5559 14772
rect 5734 14675 5835 14772
rect 5715 14635 5835 14675
rect 6105 14635 6109 14772
rect 6284 14675 6385 14772
rect 6265 14635 6385 14675
rect 6655 14635 6659 14772
rect 6834 14675 6935 14772
rect 6815 14635 6935 14675
rect 7205 14635 7209 14772
rect 7384 14675 7485 14772
rect 7365 14635 7485 14675
rect 7755 14635 7759 14772
rect 7934 14675 8035 14772
rect 7915 14635 8035 14675
rect 8305 14635 8309 14772
rect 8484 14675 8585 14772
rect 8465 14635 8585 14675
rect 8855 14635 8859 14772
rect 9034 14675 9135 14772
rect 9015 14635 9135 14675
rect 9405 14635 9409 14772
rect 9584 14675 9685 14772
rect 9565 14635 9685 14675
rect 9955 14635 9959 14772
rect 10134 14675 10235 14772
rect 10115 14635 10235 14675
rect 10505 14635 10509 14772
rect 10684 14675 10785 14772
rect 10665 14635 10785 14675
rect 11055 14635 11059 14772
rect 11234 14675 11335 14772
rect 11215 14635 11335 14675
rect 11605 14635 11609 14772
rect 11784 14675 11885 14772
rect 11765 14635 11885 14675
rect 12155 14635 12159 14772
rect 12334 14675 12435 14772
rect 12315 14635 12435 14675
rect 12705 14635 12709 14772
rect 12884 14675 12985 14772
rect 12865 14635 12985 14675
rect 13255 14635 13259 14772
rect 13434 14675 13535 14772
rect 13415 14635 13535 14675
rect 13805 14635 13809 14772
rect 13984 14675 14085 14772
rect 13965 14635 14085 14675
rect 14355 14635 14359 14772
rect 14534 14675 14635 14772
rect 14515 14635 14635 14675
rect 14905 14635 14909 14772
rect 15084 14675 15185 14772
rect 15065 14635 15185 14675
rect 15455 14635 15459 14772
rect 15634 14675 15735 14772
rect 15615 14635 15735 14675
rect 16005 14635 16009 14772
rect 16184 14675 16285 14772
rect 16165 14635 16285 14675
rect 16555 14635 16559 14772
rect 16734 14675 16835 14772
rect 16715 14635 16835 14675
rect 17105 14635 17109 14772
rect 17284 14675 17385 14772
rect 17265 14635 17385 14675
rect 17655 14635 17659 14772
rect 17834 14675 17935 14772
rect 17815 14635 17935 14675
rect 18205 14635 18209 14772
rect 18384 14675 18485 14772
rect 18365 14635 18485 14675
rect 18755 14635 18759 14772
rect 18934 14675 19035 14772
rect 18915 14635 19035 14675
rect 725 14628 842 14635
rect 885 14628 1045 14635
rect 725 14522 808 14628
rect 842 14522 1045 14628
rect 725 14515 765 14522
rect 808 14515 1045 14522
rect 1275 14628 1392 14635
rect 1435 14628 1595 14635
rect 1275 14522 1358 14628
rect 1392 14522 1595 14628
rect 1275 14515 1315 14522
rect 1358 14515 1595 14522
rect 1825 14628 1942 14635
rect 1985 14628 2145 14635
rect 1825 14522 1908 14628
rect 1942 14522 2145 14628
rect 1825 14515 1865 14522
rect 1908 14515 2145 14522
rect 2375 14628 2492 14635
rect 2535 14628 2695 14635
rect 2375 14522 2458 14628
rect 2492 14522 2695 14628
rect 2375 14515 2415 14522
rect 2458 14515 2695 14522
rect 2925 14628 3042 14635
rect 3085 14628 3245 14635
rect 2925 14522 3008 14628
rect 3042 14522 3245 14628
rect 2925 14515 2965 14522
rect 3008 14515 3245 14522
rect 3475 14628 3592 14635
rect 3635 14628 3795 14635
rect 3475 14522 3558 14628
rect 3592 14522 3795 14628
rect 3475 14515 3515 14522
rect 3558 14515 3795 14522
rect 4025 14628 4142 14635
rect 4185 14628 4345 14635
rect 4025 14522 4108 14628
rect 4142 14522 4345 14628
rect 4025 14515 4065 14522
rect 4108 14515 4345 14522
rect 4575 14628 4692 14635
rect 4735 14628 4895 14635
rect 4575 14522 4658 14628
rect 4692 14522 4895 14628
rect 4575 14515 4615 14522
rect 4658 14515 4895 14522
rect 5125 14628 5242 14635
rect 5285 14628 5445 14635
rect 5125 14522 5208 14628
rect 5242 14522 5445 14628
rect 5125 14515 5165 14522
rect 5208 14515 5445 14522
rect 5675 14628 5792 14635
rect 5835 14628 5995 14635
rect 5675 14522 5758 14628
rect 5792 14522 5995 14628
rect 5675 14515 5715 14522
rect 5758 14515 5995 14522
rect 6225 14628 6342 14635
rect 6385 14628 6545 14635
rect 6225 14522 6308 14628
rect 6342 14522 6545 14628
rect 6225 14515 6265 14522
rect 6308 14515 6545 14522
rect 6775 14628 6892 14635
rect 6935 14628 7095 14635
rect 6775 14522 6858 14628
rect 6892 14522 7095 14628
rect 6775 14515 6815 14522
rect 6858 14515 7095 14522
rect 7325 14628 7442 14635
rect 7485 14628 7645 14635
rect 7325 14522 7408 14628
rect 7442 14522 7645 14628
rect 7325 14515 7365 14522
rect 7408 14515 7645 14522
rect 7875 14628 7992 14635
rect 8035 14628 8195 14635
rect 7875 14522 7958 14628
rect 7992 14522 8195 14628
rect 7875 14515 7915 14522
rect 7958 14515 8195 14522
rect 8425 14628 8542 14635
rect 8585 14628 8745 14635
rect 8425 14522 8508 14628
rect 8542 14522 8745 14628
rect 8425 14515 8465 14522
rect 8508 14515 8745 14522
rect 8975 14628 9092 14635
rect 9135 14628 9295 14635
rect 8975 14522 9058 14628
rect 9092 14522 9295 14628
rect 8975 14515 9015 14522
rect 9058 14515 9295 14522
rect 9525 14628 9642 14635
rect 9685 14628 9845 14635
rect 9525 14522 9608 14628
rect 9642 14522 9845 14628
rect 9525 14515 9565 14522
rect 9608 14515 9845 14522
rect 10075 14628 10192 14635
rect 10235 14628 10395 14635
rect 10075 14522 10158 14628
rect 10192 14522 10395 14628
rect 10075 14515 10115 14522
rect 10158 14515 10395 14522
rect 10625 14628 10742 14635
rect 10785 14628 10945 14635
rect 10625 14522 10708 14628
rect 10742 14522 10945 14628
rect 10625 14515 10665 14522
rect 10708 14515 10945 14522
rect 11175 14628 11292 14635
rect 11335 14628 11495 14635
rect 11175 14522 11258 14628
rect 11292 14522 11495 14628
rect 11175 14515 11215 14522
rect 11258 14515 11495 14522
rect 11725 14628 11842 14635
rect 11885 14628 12045 14635
rect 11725 14522 11808 14628
rect 11842 14522 12045 14628
rect 11725 14515 11765 14522
rect 11808 14515 12045 14522
rect 12275 14628 12392 14635
rect 12435 14628 12595 14635
rect 12275 14522 12358 14628
rect 12392 14522 12595 14628
rect 12275 14515 12315 14522
rect 12358 14515 12595 14522
rect 12825 14628 12942 14635
rect 12985 14628 13145 14635
rect 12825 14522 12908 14628
rect 12942 14522 13145 14628
rect 12825 14515 12865 14522
rect 12908 14515 13145 14522
rect 13375 14628 13492 14635
rect 13535 14628 13695 14635
rect 13375 14522 13458 14628
rect 13492 14522 13695 14628
rect 13375 14515 13415 14522
rect 13458 14515 13695 14522
rect 13925 14628 14042 14635
rect 14085 14628 14245 14635
rect 13925 14522 14008 14628
rect 14042 14522 14245 14628
rect 13925 14515 13965 14522
rect 14008 14515 14245 14522
rect 14475 14628 14592 14635
rect 14635 14628 14795 14635
rect 14475 14522 14558 14628
rect 14592 14522 14795 14628
rect 14475 14515 14515 14522
rect 14558 14515 14795 14522
rect 15025 14628 15142 14635
rect 15185 14628 15345 14635
rect 15025 14522 15108 14628
rect 15142 14522 15345 14628
rect 15025 14515 15065 14522
rect 15108 14515 15345 14522
rect 15575 14628 15692 14635
rect 15735 14628 15895 14635
rect 15575 14522 15658 14628
rect 15692 14522 15895 14628
rect 15575 14515 15615 14522
rect 15658 14515 15895 14522
rect 16125 14628 16242 14635
rect 16285 14628 16445 14635
rect 16125 14522 16208 14628
rect 16242 14522 16445 14628
rect 16125 14515 16165 14522
rect 16208 14515 16445 14522
rect 16675 14628 16792 14635
rect 16835 14628 16995 14635
rect 16675 14522 16758 14628
rect 16792 14522 16995 14628
rect 16675 14515 16715 14522
rect 16758 14515 16995 14522
rect 17225 14628 17342 14635
rect 17385 14628 17545 14635
rect 17225 14522 17308 14628
rect 17342 14522 17545 14628
rect 17225 14515 17265 14522
rect 17308 14515 17545 14522
rect 17775 14628 17892 14635
rect 17935 14628 18095 14635
rect 17775 14522 17858 14628
rect 17892 14522 18095 14628
rect 17775 14515 17815 14522
rect 17858 14515 18095 14522
rect 18325 14628 18442 14635
rect 18485 14628 18645 14635
rect 18325 14522 18408 14628
rect 18442 14522 18645 14628
rect 18325 14515 18365 14522
rect 18408 14515 18645 14522
rect 18875 14628 18992 14635
rect 19035 14628 19195 14635
rect 18875 14522 18958 14628
rect 18992 14522 19195 14628
rect 18875 14515 18915 14522
rect 18958 14515 19195 14522
rect 765 14475 885 14515
rect 1315 14475 1435 14515
rect 1865 14475 1985 14515
rect 2415 14475 2535 14515
rect 2965 14475 3085 14515
rect 3515 14475 3635 14515
rect 4065 14475 4185 14515
rect 4615 14475 4735 14515
rect 5165 14475 5285 14515
rect 5715 14475 5835 14515
rect 6265 14475 6385 14515
rect 6815 14475 6935 14515
rect 7365 14475 7485 14515
rect 7915 14475 8035 14515
rect 8465 14475 8585 14515
rect 9015 14475 9135 14515
rect 9565 14475 9685 14515
rect 10115 14475 10235 14515
rect 10665 14475 10785 14515
rect 11215 14475 11335 14515
rect 11765 14475 11885 14515
rect 12315 14475 12435 14515
rect 12865 14475 12985 14515
rect 13415 14475 13535 14515
rect 13965 14475 14085 14515
rect 14515 14475 14635 14515
rect 15065 14475 15185 14515
rect 15615 14475 15735 14515
rect 16165 14475 16285 14515
rect 16715 14475 16835 14515
rect 17265 14475 17385 14515
rect 17815 14475 17935 14515
rect 18365 14475 18485 14515
rect 18915 14475 19035 14515
rect 19185 14354 19200 14371
rect 19202 14362 19204 14788
rect 19202 14348 19217 14354
rect 500 14275 507 14325
rect 500 13839 525 14240
rect 628 14222 885 14245
rect 1178 14222 1435 14245
rect 1728 14222 1985 14245
rect 2278 14222 2535 14245
rect 2828 14222 3085 14245
rect 3378 14222 3635 14245
rect 3928 14222 4185 14245
rect 4478 14222 4735 14245
rect 5028 14222 5285 14245
rect 5578 14222 5835 14245
rect 6128 14222 6385 14245
rect 6678 14222 6935 14245
rect 7228 14222 7485 14245
rect 7778 14222 8035 14245
rect 8328 14222 8585 14245
rect 8878 14222 9135 14245
rect 9428 14222 9685 14245
rect 9978 14222 10235 14245
rect 10528 14222 10785 14245
rect 11078 14222 11335 14245
rect 11628 14222 11885 14245
rect 12178 14222 12435 14245
rect 12728 14222 12985 14245
rect 13278 14222 13535 14245
rect 13828 14222 14085 14245
rect 14378 14222 14635 14245
rect 14928 14222 15185 14245
rect 15478 14222 15735 14245
rect 16028 14222 16285 14245
rect 16578 14222 16835 14245
rect 17128 14222 17385 14245
rect 17678 14222 17935 14245
rect 18228 14222 18485 14245
rect 18778 14222 19035 14245
rect 605 14085 609 14222
rect 784 14125 885 14222
rect 765 14085 885 14125
rect 1155 14085 1159 14222
rect 1334 14125 1435 14222
rect 1315 14085 1435 14125
rect 1705 14085 1709 14222
rect 1884 14125 1985 14222
rect 1865 14085 1985 14125
rect 2255 14085 2259 14222
rect 2434 14125 2535 14222
rect 2415 14085 2535 14125
rect 2805 14085 2809 14222
rect 2984 14125 3085 14222
rect 2965 14085 3085 14125
rect 3355 14085 3359 14222
rect 3534 14125 3635 14222
rect 3515 14085 3635 14125
rect 3905 14085 3909 14222
rect 4084 14125 4185 14222
rect 4065 14085 4185 14125
rect 4455 14085 4459 14222
rect 4634 14125 4735 14222
rect 4615 14085 4735 14125
rect 5005 14085 5009 14222
rect 5184 14125 5285 14222
rect 5165 14085 5285 14125
rect 5555 14085 5559 14222
rect 5734 14125 5835 14222
rect 5715 14085 5835 14125
rect 6105 14085 6109 14222
rect 6284 14125 6385 14222
rect 6265 14085 6385 14125
rect 6655 14085 6659 14222
rect 6834 14125 6935 14222
rect 6815 14085 6935 14125
rect 7205 14085 7209 14222
rect 7384 14125 7485 14222
rect 7365 14085 7485 14125
rect 7755 14085 7759 14222
rect 7934 14125 8035 14222
rect 7915 14085 8035 14125
rect 8305 14085 8309 14222
rect 8484 14125 8585 14222
rect 8465 14085 8585 14125
rect 8855 14085 8859 14222
rect 9034 14125 9135 14222
rect 9015 14085 9135 14125
rect 9405 14085 9409 14222
rect 9584 14125 9685 14222
rect 9565 14085 9685 14125
rect 9955 14085 9959 14222
rect 10134 14125 10235 14222
rect 10115 14085 10235 14125
rect 10505 14085 10509 14222
rect 10684 14125 10785 14222
rect 10665 14085 10785 14125
rect 11055 14085 11059 14222
rect 11234 14125 11335 14222
rect 11215 14085 11335 14125
rect 11605 14085 11609 14222
rect 11784 14125 11885 14222
rect 11765 14085 11885 14125
rect 12155 14085 12159 14222
rect 12334 14125 12435 14222
rect 12315 14085 12435 14125
rect 12705 14085 12709 14222
rect 12884 14125 12985 14222
rect 12865 14085 12985 14125
rect 13255 14085 13259 14222
rect 13434 14125 13535 14222
rect 13415 14085 13535 14125
rect 13805 14085 13809 14222
rect 13984 14125 14085 14222
rect 13965 14085 14085 14125
rect 14355 14085 14359 14222
rect 14534 14125 14635 14222
rect 14515 14085 14635 14125
rect 14905 14085 14909 14222
rect 15084 14125 15185 14222
rect 15065 14085 15185 14125
rect 15455 14085 15459 14222
rect 15634 14125 15735 14222
rect 15615 14085 15735 14125
rect 16005 14085 16009 14222
rect 16184 14125 16285 14222
rect 16165 14085 16285 14125
rect 16555 14085 16559 14222
rect 16734 14125 16835 14222
rect 16715 14085 16835 14125
rect 17105 14085 17109 14222
rect 17284 14125 17385 14222
rect 17265 14085 17385 14125
rect 17655 14085 17659 14222
rect 17834 14125 17935 14222
rect 17815 14085 17935 14125
rect 18205 14085 18209 14222
rect 18384 14125 18485 14222
rect 18365 14085 18485 14125
rect 18755 14085 18759 14222
rect 18934 14125 19035 14222
rect 18915 14085 19035 14125
rect 725 14078 842 14085
rect 885 14078 1045 14085
rect 725 13972 808 14078
rect 842 13972 1045 14078
rect 725 13965 765 13972
rect 808 13965 1045 13972
rect 1275 14078 1392 14085
rect 1435 14078 1595 14085
rect 1275 13972 1358 14078
rect 1392 13972 1595 14078
rect 1275 13965 1315 13972
rect 1358 13965 1595 13972
rect 1825 14078 1942 14085
rect 1985 14078 2145 14085
rect 1825 13972 1908 14078
rect 1942 13972 2145 14078
rect 1825 13965 1865 13972
rect 1908 13965 2145 13972
rect 2375 14078 2492 14085
rect 2535 14078 2695 14085
rect 2375 13972 2458 14078
rect 2492 13972 2695 14078
rect 2375 13965 2415 13972
rect 2458 13965 2695 13972
rect 2925 14078 3042 14085
rect 3085 14078 3245 14085
rect 2925 13972 3008 14078
rect 3042 13972 3245 14078
rect 2925 13965 2965 13972
rect 3008 13965 3245 13972
rect 3475 14078 3592 14085
rect 3635 14078 3795 14085
rect 3475 13972 3558 14078
rect 3592 13972 3795 14078
rect 3475 13965 3515 13972
rect 3558 13965 3795 13972
rect 4025 14078 4142 14085
rect 4185 14078 4345 14085
rect 4025 13972 4108 14078
rect 4142 13972 4345 14078
rect 4025 13965 4065 13972
rect 4108 13965 4345 13972
rect 4575 14078 4692 14085
rect 4735 14078 4895 14085
rect 4575 13972 4658 14078
rect 4692 13972 4895 14078
rect 4575 13965 4615 13972
rect 4658 13965 4895 13972
rect 5125 14078 5242 14085
rect 5285 14078 5445 14085
rect 5125 13972 5208 14078
rect 5242 13972 5445 14078
rect 5125 13965 5165 13972
rect 5208 13965 5445 13972
rect 5675 14078 5792 14085
rect 5835 14078 5995 14085
rect 5675 13972 5758 14078
rect 5792 13972 5995 14078
rect 5675 13965 5715 13972
rect 5758 13965 5995 13972
rect 6225 14078 6342 14085
rect 6385 14078 6545 14085
rect 6225 13972 6308 14078
rect 6342 13972 6545 14078
rect 6225 13965 6265 13972
rect 6308 13965 6545 13972
rect 6775 14078 6892 14085
rect 6935 14078 7095 14085
rect 6775 13972 6858 14078
rect 6892 13972 7095 14078
rect 6775 13965 6815 13972
rect 6858 13965 7095 13972
rect 7325 14078 7442 14085
rect 7485 14078 7645 14085
rect 7325 13972 7408 14078
rect 7442 13972 7645 14078
rect 7325 13965 7365 13972
rect 7408 13965 7645 13972
rect 7875 14078 7992 14085
rect 8035 14078 8195 14085
rect 7875 13972 7958 14078
rect 7992 13972 8195 14078
rect 7875 13965 7915 13972
rect 7958 13965 8195 13972
rect 8425 14078 8542 14085
rect 8585 14078 8745 14085
rect 8425 13972 8508 14078
rect 8542 13972 8745 14078
rect 8425 13965 8465 13972
rect 8508 13965 8745 13972
rect 8975 14078 9092 14085
rect 9135 14078 9295 14085
rect 8975 13972 9058 14078
rect 9092 13972 9295 14078
rect 8975 13965 9015 13972
rect 9058 13965 9295 13972
rect 9525 14078 9642 14085
rect 9685 14078 9845 14085
rect 9525 13972 9608 14078
rect 9642 13972 9845 14078
rect 9525 13965 9565 13972
rect 9608 13965 9845 13972
rect 10075 14078 10192 14085
rect 10235 14078 10395 14085
rect 10075 13972 10158 14078
rect 10192 13972 10395 14078
rect 10075 13965 10115 13972
rect 10158 13965 10395 13972
rect 10625 14078 10742 14085
rect 10785 14078 10945 14085
rect 10625 13972 10708 14078
rect 10742 13972 10945 14078
rect 10625 13965 10665 13972
rect 10708 13965 10945 13972
rect 11175 14078 11292 14085
rect 11335 14078 11495 14085
rect 11175 13972 11258 14078
rect 11292 13972 11495 14078
rect 11175 13965 11215 13972
rect 11258 13965 11495 13972
rect 11725 14078 11842 14085
rect 11885 14078 12045 14085
rect 11725 13972 11808 14078
rect 11842 13972 12045 14078
rect 11725 13965 11765 13972
rect 11808 13965 12045 13972
rect 12275 14078 12392 14085
rect 12435 14078 12595 14085
rect 12275 13972 12358 14078
rect 12392 13972 12595 14078
rect 12275 13965 12315 13972
rect 12358 13965 12595 13972
rect 12825 14078 12942 14085
rect 12985 14078 13145 14085
rect 12825 13972 12908 14078
rect 12942 13972 13145 14078
rect 12825 13965 12865 13972
rect 12908 13965 13145 13972
rect 13375 14078 13492 14085
rect 13535 14078 13695 14085
rect 13375 13972 13458 14078
rect 13492 13972 13695 14078
rect 13375 13965 13415 13972
rect 13458 13965 13695 13972
rect 13925 14078 14042 14085
rect 14085 14078 14245 14085
rect 13925 13972 14008 14078
rect 14042 13972 14245 14078
rect 13925 13965 13965 13972
rect 14008 13965 14245 13972
rect 14475 14078 14592 14085
rect 14635 14078 14795 14085
rect 14475 13972 14558 14078
rect 14592 13972 14795 14078
rect 14475 13965 14515 13972
rect 14558 13965 14795 13972
rect 15025 14078 15142 14085
rect 15185 14078 15345 14085
rect 15025 13972 15108 14078
rect 15142 13972 15345 14078
rect 15025 13965 15065 13972
rect 15108 13965 15345 13972
rect 15575 14078 15692 14085
rect 15735 14078 15895 14085
rect 15575 13972 15658 14078
rect 15692 13972 15895 14078
rect 15575 13965 15615 13972
rect 15658 13965 15895 13972
rect 16125 14078 16242 14085
rect 16285 14078 16445 14085
rect 16125 13972 16208 14078
rect 16242 13972 16445 14078
rect 16125 13965 16165 13972
rect 16208 13965 16445 13972
rect 16675 14078 16792 14085
rect 16835 14078 16995 14085
rect 16675 13972 16758 14078
rect 16792 13972 16995 14078
rect 16675 13965 16715 13972
rect 16758 13965 16995 13972
rect 17225 14078 17342 14085
rect 17385 14078 17545 14085
rect 17225 13972 17308 14078
rect 17342 13972 17545 14078
rect 17225 13965 17265 13972
rect 17308 13965 17545 13972
rect 17775 14078 17892 14085
rect 17935 14078 18095 14085
rect 17775 13972 17858 14078
rect 17892 13972 18095 14078
rect 17775 13965 17815 13972
rect 17858 13965 18095 13972
rect 18325 14078 18442 14085
rect 18485 14078 18645 14085
rect 18325 13972 18408 14078
rect 18442 13972 18645 14078
rect 18325 13965 18365 13972
rect 18408 13965 18645 13972
rect 18875 14078 18992 14085
rect 19035 14078 19195 14085
rect 18875 13972 18958 14078
rect 18992 13972 19195 14078
rect 18875 13965 18915 13972
rect 18958 13965 19195 13972
rect 765 13925 885 13965
rect 1315 13925 1435 13965
rect 1865 13925 1985 13965
rect 2415 13925 2535 13965
rect 2965 13925 3085 13965
rect 3515 13925 3635 13965
rect 4065 13925 4185 13965
rect 4615 13925 4735 13965
rect 5165 13925 5285 13965
rect 5715 13925 5835 13965
rect 6265 13925 6385 13965
rect 6815 13925 6935 13965
rect 7365 13925 7485 13965
rect 7915 13925 8035 13965
rect 8465 13925 8585 13965
rect 9015 13925 9135 13965
rect 9565 13925 9685 13965
rect 10115 13925 10235 13965
rect 10665 13925 10785 13965
rect 11215 13925 11335 13965
rect 11765 13925 11885 13965
rect 12315 13925 12435 13965
rect 12865 13925 12985 13965
rect 13415 13925 13535 13965
rect 13965 13925 14085 13965
rect 14515 13925 14635 13965
rect 15065 13925 15185 13965
rect 15615 13925 15735 13965
rect 16165 13925 16285 13965
rect 16715 13925 16835 13965
rect 17265 13925 17385 13965
rect 17815 13925 17935 13965
rect 18365 13925 18485 13965
rect 18915 13925 19035 13965
rect 19202 13812 19204 14238
rect 500 13725 507 13775
rect 19202 13696 19217 13702
rect 628 13672 885 13695
rect 1178 13672 1435 13695
rect 1728 13672 1985 13695
rect 2278 13672 2535 13695
rect 2828 13672 3085 13695
rect 3378 13672 3635 13695
rect 3928 13672 4185 13695
rect 4478 13672 4735 13695
rect 5028 13672 5285 13695
rect 5578 13672 5835 13695
rect 6128 13672 6385 13695
rect 6678 13672 6935 13695
rect 7228 13672 7485 13695
rect 7778 13672 8035 13695
rect 8328 13672 8585 13695
rect 8878 13672 9135 13695
rect 9428 13672 9685 13695
rect 9978 13672 10235 13695
rect 10528 13672 10785 13695
rect 11078 13672 11335 13695
rect 11628 13672 11885 13695
rect 12178 13672 12435 13695
rect 12728 13672 12985 13695
rect 13278 13672 13535 13695
rect 13828 13672 14085 13695
rect 14378 13672 14635 13695
rect 14928 13672 15185 13695
rect 15478 13672 15735 13695
rect 16028 13672 16285 13695
rect 16578 13672 16835 13695
rect 17128 13672 17385 13695
rect 17678 13672 17935 13695
rect 18228 13672 18485 13695
rect 18778 13672 19035 13695
rect 605 13535 609 13672
rect 784 13575 885 13672
rect 765 13535 885 13575
rect 1155 13535 1159 13672
rect 1334 13575 1435 13672
rect 1315 13535 1435 13575
rect 1705 13535 1709 13672
rect 1884 13575 1985 13672
rect 1865 13535 1985 13575
rect 2255 13535 2259 13672
rect 2434 13575 2535 13672
rect 2415 13535 2535 13575
rect 2805 13535 2809 13672
rect 2984 13575 3085 13672
rect 2965 13535 3085 13575
rect 3355 13535 3359 13672
rect 3534 13575 3635 13672
rect 3515 13535 3635 13575
rect 3905 13535 3909 13672
rect 4084 13575 4185 13672
rect 4065 13535 4185 13575
rect 4455 13535 4459 13672
rect 4634 13575 4735 13672
rect 4615 13535 4735 13575
rect 5005 13535 5009 13672
rect 5184 13575 5285 13672
rect 5165 13535 5285 13575
rect 5555 13535 5559 13672
rect 5734 13575 5835 13672
rect 5715 13535 5835 13575
rect 6105 13535 6109 13672
rect 6284 13575 6385 13672
rect 6265 13535 6385 13575
rect 6655 13535 6659 13672
rect 6834 13575 6935 13672
rect 6815 13535 6935 13575
rect 7205 13535 7209 13672
rect 7384 13575 7485 13672
rect 7365 13535 7485 13575
rect 7755 13535 7759 13672
rect 7934 13575 8035 13672
rect 7915 13535 8035 13575
rect 8305 13535 8309 13672
rect 8484 13575 8585 13672
rect 8465 13535 8585 13575
rect 8855 13535 8859 13672
rect 9034 13575 9135 13672
rect 9015 13535 9135 13575
rect 9405 13535 9409 13672
rect 9584 13575 9685 13672
rect 9565 13535 9685 13575
rect 9955 13535 9959 13672
rect 10134 13575 10235 13672
rect 10115 13535 10235 13575
rect 10505 13535 10509 13672
rect 10684 13575 10785 13672
rect 10665 13535 10785 13575
rect 11055 13535 11059 13672
rect 11234 13575 11335 13672
rect 11215 13535 11335 13575
rect 11605 13535 11609 13672
rect 11784 13575 11885 13672
rect 11765 13535 11885 13575
rect 12155 13535 12159 13672
rect 12334 13575 12435 13672
rect 12315 13535 12435 13575
rect 12705 13535 12709 13672
rect 12884 13575 12985 13672
rect 12865 13535 12985 13575
rect 13255 13535 13259 13672
rect 13434 13575 13535 13672
rect 13415 13535 13535 13575
rect 13805 13535 13809 13672
rect 13984 13575 14085 13672
rect 13965 13535 14085 13575
rect 14355 13535 14359 13672
rect 14534 13575 14635 13672
rect 14515 13535 14635 13575
rect 14905 13535 14909 13672
rect 15084 13575 15185 13672
rect 15065 13535 15185 13575
rect 15455 13535 15459 13672
rect 15634 13575 15735 13672
rect 15615 13535 15735 13575
rect 16005 13535 16009 13672
rect 16184 13575 16285 13672
rect 16165 13535 16285 13575
rect 16555 13535 16559 13672
rect 16734 13575 16835 13672
rect 16715 13535 16835 13575
rect 17105 13535 17109 13672
rect 17284 13575 17385 13672
rect 17265 13535 17385 13575
rect 17655 13535 17659 13672
rect 17834 13575 17935 13672
rect 17815 13535 17935 13575
rect 18205 13535 18209 13672
rect 18384 13575 18485 13672
rect 18365 13535 18485 13575
rect 18755 13535 18759 13672
rect 18934 13575 19035 13672
rect 18915 13535 19035 13575
rect 725 13528 842 13535
rect 885 13528 1045 13535
rect 725 13422 808 13528
rect 842 13422 1045 13528
rect 725 13415 765 13422
rect 808 13415 1045 13422
rect 1275 13528 1392 13535
rect 1435 13528 1595 13535
rect 1275 13422 1358 13528
rect 1392 13422 1595 13528
rect 1275 13415 1315 13422
rect 1358 13415 1595 13422
rect 1825 13528 1942 13535
rect 1985 13528 2145 13535
rect 1825 13422 1908 13528
rect 1942 13422 2145 13528
rect 1825 13415 1865 13422
rect 1908 13415 2145 13422
rect 2375 13528 2492 13535
rect 2535 13528 2695 13535
rect 2375 13422 2458 13528
rect 2492 13422 2695 13528
rect 2375 13415 2415 13422
rect 2458 13415 2695 13422
rect 2925 13528 3042 13535
rect 3085 13528 3245 13535
rect 2925 13422 3008 13528
rect 3042 13422 3245 13528
rect 2925 13415 2965 13422
rect 3008 13415 3245 13422
rect 3475 13528 3592 13535
rect 3635 13528 3795 13535
rect 3475 13422 3558 13528
rect 3592 13422 3795 13528
rect 3475 13415 3515 13422
rect 3558 13415 3795 13422
rect 4025 13528 4142 13535
rect 4185 13528 4345 13535
rect 4025 13422 4108 13528
rect 4142 13422 4345 13528
rect 4025 13415 4065 13422
rect 4108 13415 4345 13422
rect 4575 13528 4692 13535
rect 4735 13528 4895 13535
rect 4575 13422 4658 13528
rect 4692 13422 4895 13528
rect 4575 13415 4615 13422
rect 4658 13415 4895 13422
rect 5125 13528 5242 13535
rect 5285 13528 5445 13535
rect 5125 13422 5208 13528
rect 5242 13422 5445 13528
rect 5125 13415 5165 13422
rect 5208 13415 5445 13422
rect 5675 13528 5792 13535
rect 5835 13528 5995 13535
rect 5675 13422 5758 13528
rect 5792 13422 5995 13528
rect 5675 13415 5715 13422
rect 5758 13415 5995 13422
rect 6225 13528 6342 13535
rect 6385 13528 6545 13535
rect 6225 13422 6308 13528
rect 6342 13422 6545 13528
rect 6225 13415 6265 13422
rect 6308 13415 6545 13422
rect 6775 13528 6892 13535
rect 6935 13528 7095 13535
rect 6775 13422 6858 13528
rect 6892 13422 7095 13528
rect 6775 13415 6815 13422
rect 6858 13415 7095 13422
rect 7325 13528 7442 13535
rect 7485 13528 7645 13535
rect 7325 13422 7408 13528
rect 7442 13422 7645 13528
rect 7325 13415 7365 13422
rect 7408 13415 7645 13422
rect 7875 13528 7992 13535
rect 8035 13528 8195 13535
rect 7875 13422 7958 13528
rect 7992 13422 8195 13528
rect 7875 13415 7915 13422
rect 7958 13415 8195 13422
rect 8425 13528 8542 13535
rect 8585 13528 8745 13535
rect 8425 13422 8508 13528
rect 8542 13422 8745 13528
rect 8425 13415 8465 13422
rect 8508 13415 8745 13422
rect 8975 13528 9092 13535
rect 9135 13528 9295 13535
rect 8975 13422 9058 13528
rect 9092 13422 9295 13528
rect 8975 13415 9015 13422
rect 9058 13415 9295 13422
rect 9525 13528 9642 13535
rect 9685 13528 9845 13535
rect 9525 13422 9608 13528
rect 9642 13422 9845 13528
rect 9525 13415 9565 13422
rect 9608 13415 9845 13422
rect 10075 13528 10192 13535
rect 10235 13528 10395 13535
rect 10075 13422 10158 13528
rect 10192 13422 10395 13528
rect 10075 13415 10115 13422
rect 10158 13415 10395 13422
rect 10625 13528 10742 13535
rect 10785 13528 10945 13535
rect 10625 13422 10708 13528
rect 10742 13422 10945 13528
rect 10625 13415 10665 13422
rect 10708 13415 10945 13422
rect 11175 13528 11292 13535
rect 11335 13528 11495 13535
rect 11175 13422 11258 13528
rect 11292 13422 11495 13528
rect 11175 13415 11215 13422
rect 11258 13415 11495 13422
rect 11725 13528 11842 13535
rect 11885 13528 12045 13535
rect 11725 13422 11808 13528
rect 11842 13422 12045 13528
rect 11725 13415 11765 13422
rect 11808 13415 12045 13422
rect 12275 13528 12392 13535
rect 12435 13528 12595 13535
rect 12275 13422 12358 13528
rect 12392 13422 12595 13528
rect 12275 13415 12315 13422
rect 12358 13415 12595 13422
rect 12825 13528 12942 13535
rect 12985 13528 13145 13535
rect 12825 13422 12908 13528
rect 12942 13422 13145 13528
rect 12825 13415 12865 13422
rect 12908 13415 13145 13422
rect 13375 13528 13492 13535
rect 13535 13528 13695 13535
rect 13375 13422 13458 13528
rect 13492 13422 13695 13528
rect 13375 13415 13415 13422
rect 13458 13415 13695 13422
rect 13925 13528 14042 13535
rect 14085 13528 14245 13535
rect 13925 13422 14008 13528
rect 14042 13422 14245 13528
rect 13925 13415 13965 13422
rect 14008 13415 14245 13422
rect 14475 13528 14592 13535
rect 14635 13528 14795 13535
rect 14475 13422 14558 13528
rect 14592 13422 14795 13528
rect 14475 13415 14515 13422
rect 14558 13415 14795 13422
rect 15025 13528 15142 13535
rect 15185 13528 15345 13535
rect 15025 13422 15108 13528
rect 15142 13422 15345 13528
rect 15025 13415 15065 13422
rect 15108 13415 15345 13422
rect 15575 13528 15692 13535
rect 15735 13528 15895 13535
rect 15575 13422 15658 13528
rect 15692 13422 15895 13528
rect 15575 13415 15615 13422
rect 15658 13415 15895 13422
rect 16125 13528 16242 13535
rect 16285 13528 16445 13535
rect 16125 13422 16208 13528
rect 16242 13422 16445 13528
rect 16125 13415 16165 13422
rect 16208 13415 16445 13422
rect 16675 13528 16792 13535
rect 16835 13528 16995 13535
rect 16675 13422 16758 13528
rect 16792 13422 16995 13528
rect 16675 13415 16715 13422
rect 16758 13415 16995 13422
rect 17225 13528 17342 13535
rect 17385 13528 17545 13535
rect 17225 13422 17308 13528
rect 17342 13422 17545 13528
rect 17225 13415 17265 13422
rect 17308 13415 17545 13422
rect 17775 13528 17892 13535
rect 17935 13528 18095 13535
rect 17775 13422 17858 13528
rect 17892 13422 18095 13528
rect 17775 13415 17815 13422
rect 17858 13415 18095 13422
rect 18325 13528 18442 13535
rect 18485 13528 18645 13535
rect 18325 13422 18408 13528
rect 18442 13422 18645 13528
rect 18325 13415 18365 13422
rect 18408 13415 18645 13422
rect 18875 13528 18992 13535
rect 19035 13528 19195 13535
rect 18875 13422 18958 13528
rect 18992 13422 19195 13528
rect 18875 13415 18915 13422
rect 18958 13415 19195 13422
rect 765 13375 885 13415
rect 1315 13375 1435 13415
rect 1865 13375 1985 13415
rect 2415 13375 2535 13415
rect 2965 13375 3085 13415
rect 3515 13375 3635 13415
rect 4065 13375 4185 13415
rect 4615 13375 4735 13415
rect 5165 13375 5285 13415
rect 5715 13375 5835 13415
rect 6265 13375 6385 13415
rect 6815 13375 6935 13415
rect 7365 13375 7485 13415
rect 7915 13375 8035 13415
rect 8465 13375 8585 13415
rect 9015 13375 9135 13415
rect 9565 13375 9685 13415
rect 10115 13375 10235 13415
rect 10665 13375 10785 13415
rect 11215 13375 11335 13415
rect 11765 13375 11885 13415
rect 12315 13375 12435 13415
rect 12865 13375 12985 13415
rect 13415 13375 13535 13415
rect 13965 13375 14085 13415
rect 14515 13375 14635 13415
rect 15065 13375 15185 13415
rect 15615 13375 15735 13415
rect 16165 13375 16285 13415
rect 16715 13375 16835 13415
rect 17265 13375 17385 13415
rect 17815 13375 17935 13415
rect 18365 13375 18485 13415
rect 18915 13375 19035 13415
rect 19185 13254 19200 13271
rect 19202 13262 19204 13688
rect 19202 13248 19217 13254
rect 500 13175 507 13225
rect 500 12739 525 13140
rect 628 13122 885 13145
rect 1178 13122 1435 13145
rect 1728 13122 1985 13145
rect 2278 13122 2535 13145
rect 2828 13122 3085 13145
rect 3378 13122 3635 13145
rect 3928 13122 4185 13145
rect 4478 13122 4735 13145
rect 5028 13122 5285 13145
rect 5578 13122 5835 13145
rect 6128 13122 6385 13145
rect 6678 13122 6935 13145
rect 7228 13122 7485 13145
rect 7778 13122 8035 13145
rect 8328 13122 8585 13145
rect 8878 13122 9135 13145
rect 9428 13122 9685 13145
rect 9978 13122 10235 13145
rect 10528 13122 10785 13145
rect 11078 13122 11335 13145
rect 11628 13122 11885 13145
rect 12178 13122 12435 13145
rect 12728 13122 12985 13145
rect 13278 13122 13535 13145
rect 13828 13122 14085 13145
rect 14378 13122 14635 13145
rect 14928 13122 15185 13145
rect 15478 13122 15735 13145
rect 16028 13122 16285 13145
rect 16578 13122 16835 13145
rect 17128 13122 17385 13145
rect 17678 13122 17935 13145
rect 18228 13122 18485 13145
rect 18778 13122 19035 13145
rect 605 12985 609 13122
rect 784 13025 885 13122
rect 765 12985 885 13025
rect 1155 12985 1159 13122
rect 1334 13025 1435 13122
rect 1315 12985 1435 13025
rect 1705 12985 1709 13122
rect 1884 13025 1985 13122
rect 1865 12985 1985 13025
rect 2255 12985 2259 13122
rect 2434 13025 2535 13122
rect 2415 12985 2535 13025
rect 2805 12985 2809 13122
rect 2984 13025 3085 13122
rect 2965 12985 3085 13025
rect 3355 12985 3359 13122
rect 3534 13025 3635 13122
rect 3515 12985 3635 13025
rect 3905 12985 3909 13122
rect 4084 13025 4185 13122
rect 4065 12985 4185 13025
rect 4455 12985 4459 13122
rect 4634 13025 4735 13122
rect 4615 12985 4735 13025
rect 5005 12985 5009 13122
rect 5184 13025 5285 13122
rect 5165 12985 5285 13025
rect 5555 12985 5559 13122
rect 5734 13025 5835 13122
rect 5715 12985 5835 13025
rect 6105 12985 6109 13122
rect 6284 13025 6385 13122
rect 6265 12985 6385 13025
rect 6655 12985 6659 13122
rect 6834 13025 6935 13122
rect 6815 12985 6935 13025
rect 7205 12985 7209 13122
rect 7384 13025 7485 13122
rect 7365 12985 7485 13025
rect 7755 12985 7759 13122
rect 7934 13025 8035 13122
rect 7915 12985 8035 13025
rect 8305 12985 8309 13122
rect 8484 13025 8585 13122
rect 8465 12985 8585 13025
rect 8855 12985 8859 13122
rect 9034 13025 9135 13122
rect 9015 12985 9135 13025
rect 9405 12985 9409 13122
rect 9584 13025 9685 13122
rect 9565 12985 9685 13025
rect 9955 12985 9959 13122
rect 10134 13025 10235 13122
rect 10115 12985 10235 13025
rect 10505 12985 10509 13122
rect 10684 13025 10785 13122
rect 10665 12985 10785 13025
rect 11055 12985 11059 13122
rect 11234 13025 11335 13122
rect 11215 12985 11335 13025
rect 11605 12985 11609 13122
rect 11784 13025 11885 13122
rect 11765 12985 11885 13025
rect 12155 12985 12159 13122
rect 12334 13025 12435 13122
rect 12315 12985 12435 13025
rect 12705 12985 12709 13122
rect 12884 13025 12985 13122
rect 12865 12985 12985 13025
rect 13255 12985 13259 13122
rect 13434 13025 13535 13122
rect 13415 12985 13535 13025
rect 13805 12985 13809 13122
rect 13984 13025 14085 13122
rect 13965 12985 14085 13025
rect 14355 12985 14359 13122
rect 14534 13025 14635 13122
rect 14515 12985 14635 13025
rect 14905 12985 14909 13122
rect 15084 13025 15185 13122
rect 15065 12985 15185 13025
rect 15455 12985 15459 13122
rect 15634 13025 15735 13122
rect 15615 12985 15735 13025
rect 16005 12985 16009 13122
rect 16184 13025 16285 13122
rect 16165 12985 16285 13025
rect 16555 12985 16559 13122
rect 16734 13025 16835 13122
rect 16715 12985 16835 13025
rect 17105 12985 17109 13122
rect 17284 13025 17385 13122
rect 17265 12985 17385 13025
rect 17655 12985 17659 13122
rect 17834 13025 17935 13122
rect 17815 12985 17935 13025
rect 18205 12985 18209 13122
rect 18384 13025 18485 13122
rect 18365 12985 18485 13025
rect 18755 12985 18759 13122
rect 18934 13025 19035 13122
rect 18915 12985 19035 13025
rect 725 12978 842 12985
rect 885 12978 1045 12985
rect 725 12872 808 12978
rect 842 12872 1045 12978
rect 725 12865 765 12872
rect 808 12865 1045 12872
rect 1275 12978 1392 12985
rect 1435 12978 1595 12985
rect 1275 12872 1358 12978
rect 1392 12872 1595 12978
rect 1275 12865 1315 12872
rect 1358 12865 1595 12872
rect 1825 12978 1942 12985
rect 1985 12978 2145 12985
rect 1825 12872 1908 12978
rect 1942 12872 2145 12978
rect 1825 12865 1865 12872
rect 1908 12865 2145 12872
rect 2375 12978 2492 12985
rect 2535 12978 2695 12985
rect 2375 12872 2458 12978
rect 2492 12872 2695 12978
rect 2375 12865 2415 12872
rect 2458 12865 2695 12872
rect 2925 12978 3042 12985
rect 3085 12978 3245 12985
rect 2925 12872 3008 12978
rect 3042 12872 3245 12978
rect 2925 12865 2965 12872
rect 3008 12865 3245 12872
rect 3475 12978 3592 12985
rect 3635 12978 3795 12985
rect 3475 12872 3558 12978
rect 3592 12872 3795 12978
rect 3475 12865 3515 12872
rect 3558 12865 3795 12872
rect 4025 12978 4142 12985
rect 4185 12978 4345 12985
rect 4025 12872 4108 12978
rect 4142 12872 4345 12978
rect 4025 12865 4065 12872
rect 4108 12865 4345 12872
rect 4575 12978 4692 12985
rect 4735 12978 4895 12985
rect 4575 12872 4658 12978
rect 4692 12872 4895 12978
rect 4575 12865 4615 12872
rect 4658 12865 4895 12872
rect 5125 12978 5242 12985
rect 5285 12978 5445 12985
rect 5125 12872 5208 12978
rect 5242 12872 5445 12978
rect 5125 12865 5165 12872
rect 5208 12865 5445 12872
rect 5675 12978 5792 12985
rect 5835 12978 5995 12985
rect 5675 12872 5758 12978
rect 5792 12872 5995 12978
rect 5675 12865 5715 12872
rect 5758 12865 5995 12872
rect 6225 12978 6342 12985
rect 6385 12978 6545 12985
rect 6225 12872 6308 12978
rect 6342 12872 6545 12978
rect 6225 12865 6265 12872
rect 6308 12865 6545 12872
rect 6775 12978 6892 12985
rect 6935 12978 7095 12985
rect 6775 12872 6858 12978
rect 6892 12872 7095 12978
rect 6775 12865 6815 12872
rect 6858 12865 7095 12872
rect 7325 12978 7442 12985
rect 7485 12978 7645 12985
rect 7325 12872 7408 12978
rect 7442 12872 7645 12978
rect 7325 12865 7365 12872
rect 7408 12865 7645 12872
rect 7875 12978 7992 12985
rect 8035 12978 8195 12985
rect 7875 12872 7958 12978
rect 7992 12872 8195 12978
rect 7875 12865 7915 12872
rect 7958 12865 8195 12872
rect 8425 12978 8542 12985
rect 8585 12978 8745 12985
rect 8425 12872 8508 12978
rect 8542 12872 8745 12978
rect 8425 12865 8465 12872
rect 8508 12865 8745 12872
rect 8975 12978 9092 12985
rect 9135 12978 9295 12985
rect 8975 12872 9058 12978
rect 9092 12872 9295 12978
rect 8975 12865 9015 12872
rect 9058 12865 9295 12872
rect 9525 12978 9642 12985
rect 9685 12978 9845 12985
rect 9525 12872 9608 12978
rect 9642 12872 9845 12978
rect 9525 12865 9565 12872
rect 9608 12865 9845 12872
rect 10075 12978 10192 12985
rect 10235 12978 10395 12985
rect 10075 12872 10158 12978
rect 10192 12872 10395 12978
rect 10075 12865 10115 12872
rect 10158 12865 10395 12872
rect 10625 12978 10742 12985
rect 10785 12978 10945 12985
rect 10625 12872 10708 12978
rect 10742 12872 10945 12978
rect 10625 12865 10665 12872
rect 10708 12865 10945 12872
rect 11175 12978 11292 12985
rect 11335 12978 11495 12985
rect 11175 12872 11258 12978
rect 11292 12872 11495 12978
rect 11175 12865 11215 12872
rect 11258 12865 11495 12872
rect 11725 12978 11842 12985
rect 11885 12978 12045 12985
rect 11725 12872 11808 12978
rect 11842 12872 12045 12978
rect 11725 12865 11765 12872
rect 11808 12865 12045 12872
rect 12275 12978 12392 12985
rect 12435 12978 12595 12985
rect 12275 12872 12358 12978
rect 12392 12872 12595 12978
rect 12275 12865 12315 12872
rect 12358 12865 12595 12872
rect 12825 12978 12942 12985
rect 12985 12978 13145 12985
rect 12825 12872 12908 12978
rect 12942 12872 13145 12978
rect 12825 12865 12865 12872
rect 12908 12865 13145 12872
rect 13375 12978 13492 12985
rect 13535 12978 13695 12985
rect 13375 12872 13458 12978
rect 13492 12872 13695 12978
rect 13375 12865 13415 12872
rect 13458 12865 13695 12872
rect 13925 12978 14042 12985
rect 14085 12978 14245 12985
rect 13925 12872 14008 12978
rect 14042 12872 14245 12978
rect 13925 12865 13965 12872
rect 14008 12865 14245 12872
rect 14475 12978 14592 12985
rect 14635 12978 14795 12985
rect 14475 12872 14558 12978
rect 14592 12872 14795 12978
rect 14475 12865 14515 12872
rect 14558 12865 14795 12872
rect 15025 12978 15142 12985
rect 15185 12978 15345 12985
rect 15025 12872 15108 12978
rect 15142 12872 15345 12978
rect 15025 12865 15065 12872
rect 15108 12865 15345 12872
rect 15575 12978 15692 12985
rect 15735 12978 15895 12985
rect 15575 12872 15658 12978
rect 15692 12872 15895 12978
rect 15575 12865 15615 12872
rect 15658 12865 15895 12872
rect 16125 12978 16242 12985
rect 16285 12978 16445 12985
rect 16125 12872 16208 12978
rect 16242 12872 16445 12978
rect 16125 12865 16165 12872
rect 16208 12865 16445 12872
rect 16675 12978 16792 12985
rect 16835 12978 16995 12985
rect 16675 12872 16758 12978
rect 16792 12872 16995 12978
rect 16675 12865 16715 12872
rect 16758 12865 16995 12872
rect 17225 12978 17342 12985
rect 17385 12978 17545 12985
rect 17225 12872 17308 12978
rect 17342 12872 17545 12978
rect 17225 12865 17265 12872
rect 17308 12865 17545 12872
rect 17775 12978 17892 12985
rect 17935 12978 18095 12985
rect 17775 12872 17858 12978
rect 17892 12872 18095 12978
rect 17775 12865 17815 12872
rect 17858 12865 18095 12872
rect 18325 12978 18442 12985
rect 18485 12978 18645 12985
rect 18325 12872 18408 12978
rect 18442 12872 18645 12978
rect 18325 12865 18365 12872
rect 18408 12865 18645 12872
rect 18875 12978 18992 12985
rect 19035 12978 19195 12985
rect 18875 12872 18958 12978
rect 18992 12872 19195 12978
rect 18875 12865 18915 12872
rect 18958 12865 19195 12872
rect 765 12825 885 12865
rect 1315 12825 1435 12865
rect 1865 12825 1985 12865
rect 2415 12825 2535 12865
rect 2965 12825 3085 12865
rect 3515 12825 3635 12865
rect 4065 12825 4185 12865
rect 4615 12825 4735 12865
rect 5165 12825 5285 12865
rect 5715 12825 5835 12865
rect 6265 12825 6385 12865
rect 6815 12825 6935 12865
rect 7365 12825 7485 12865
rect 7915 12825 8035 12865
rect 8465 12825 8585 12865
rect 9015 12825 9135 12865
rect 9565 12825 9685 12865
rect 10115 12825 10235 12865
rect 10665 12825 10785 12865
rect 11215 12825 11335 12865
rect 11765 12825 11885 12865
rect 12315 12825 12435 12865
rect 12865 12825 12985 12865
rect 13415 12825 13535 12865
rect 13965 12825 14085 12865
rect 14515 12825 14635 12865
rect 15065 12825 15185 12865
rect 15615 12825 15735 12865
rect 16165 12825 16285 12865
rect 16715 12825 16835 12865
rect 17265 12825 17385 12865
rect 17815 12825 17935 12865
rect 18365 12825 18485 12865
rect 18915 12825 19035 12865
rect 19202 12712 19204 13138
rect 500 12625 507 12675
rect 19202 12596 19217 12602
rect 628 12572 885 12595
rect 1178 12572 1435 12595
rect 1728 12572 1985 12595
rect 2278 12572 2535 12595
rect 2828 12572 3085 12595
rect 3378 12572 3635 12595
rect 3928 12572 4185 12595
rect 4478 12572 4735 12595
rect 5028 12572 5285 12595
rect 5578 12572 5835 12595
rect 6128 12572 6385 12595
rect 6678 12572 6935 12595
rect 7228 12572 7485 12595
rect 7778 12572 8035 12595
rect 8328 12572 8585 12595
rect 8878 12572 9135 12595
rect 9428 12572 9685 12595
rect 9978 12572 10235 12595
rect 10528 12572 10785 12595
rect 11078 12572 11335 12595
rect 11628 12572 11885 12595
rect 12178 12572 12435 12595
rect 12728 12572 12985 12595
rect 13278 12572 13535 12595
rect 13828 12572 14085 12595
rect 14378 12572 14635 12595
rect 14928 12572 15185 12595
rect 15478 12572 15735 12595
rect 16028 12572 16285 12595
rect 16578 12572 16835 12595
rect 17128 12572 17385 12595
rect 17678 12572 17935 12595
rect 18228 12572 18485 12595
rect 18778 12572 19035 12595
rect 605 12435 609 12572
rect 784 12475 885 12572
rect 765 12435 885 12475
rect 1155 12435 1159 12572
rect 1334 12475 1435 12572
rect 1315 12435 1435 12475
rect 1705 12435 1709 12572
rect 1884 12475 1985 12572
rect 1865 12435 1985 12475
rect 2255 12435 2259 12572
rect 2434 12475 2535 12572
rect 2415 12435 2535 12475
rect 2805 12435 2809 12572
rect 2984 12475 3085 12572
rect 2965 12435 3085 12475
rect 3355 12435 3359 12572
rect 3534 12475 3635 12572
rect 3515 12435 3635 12475
rect 3905 12435 3909 12572
rect 4084 12475 4185 12572
rect 4065 12435 4185 12475
rect 4455 12435 4459 12572
rect 4634 12475 4735 12572
rect 4615 12435 4735 12475
rect 5005 12435 5009 12572
rect 5184 12475 5285 12572
rect 5165 12435 5285 12475
rect 5555 12435 5559 12572
rect 5734 12475 5835 12572
rect 5715 12435 5835 12475
rect 6105 12435 6109 12572
rect 6284 12475 6385 12572
rect 6265 12435 6385 12475
rect 6655 12435 6659 12572
rect 6834 12475 6935 12572
rect 6815 12435 6935 12475
rect 7205 12435 7209 12572
rect 7384 12475 7485 12572
rect 7365 12435 7485 12475
rect 7755 12435 7759 12572
rect 7934 12475 8035 12572
rect 7915 12435 8035 12475
rect 8305 12435 8309 12572
rect 8484 12475 8585 12572
rect 8465 12435 8585 12475
rect 8855 12435 8859 12572
rect 9034 12475 9135 12572
rect 9015 12435 9135 12475
rect 9405 12435 9409 12572
rect 9584 12475 9685 12572
rect 9565 12435 9685 12475
rect 9955 12435 9959 12572
rect 10134 12475 10235 12572
rect 10115 12435 10235 12475
rect 10505 12435 10509 12572
rect 10684 12475 10785 12572
rect 10665 12435 10785 12475
rect 11055 12435 11059 12572
rect 11234 12475 11335 12572
rect 11215 12435 11335 12475
rect 11605 12435 11609 12572
rect 11784 12475 11885 12572
rect 11765 12435 11885 12475
rect 12155 12435 12159 12572
rect 12334 12475 12435 12572
rect 12315 12435 12435 12475
rect 12705 12435 12709 12572
rect 12884 12475 12985 12572
rect 12865 12435 12985 12475
rect 13255 12435 13259 12572
rect 13434 12475 13535 12572
rect 13415 12435 13535 12475
rect 13805 12435 13809 12572
rect 13984 12475 14085 12572
rect 13965 12435 14085 12475
rect 14355 12435 14359 12572
rect 14534 12475 14635 12572
rect 14515 12435 14635 12475
rect 14905 12435 14909 12572
rect 15084 12475 15185 12572
rect 15065 12435 15185 12475
rect 15455 12435 15459 12572
rect 15634 12475 15735 12572
rect 15615 12435 15735 12475
rect 16005 12435 16009 12572
rect 16184 12475 16285 12572
rect 16165 12435 16285 12475
rect 16555 12435 16559 12572
rect 16734 12475 16835 12572
rect 16715 12435 16835 12475
rect 17105 12435 17109 12572
rect 17284 12475 17385 12572
rect 17265 12435 17385 12475
rect 17655 12435 17659 12572
rect 17834 12475 17935 12572
rect 17815 12435 17935 12475
rect 18205 12435 18209 12572
rect 18384 12475 18485 12572
rect 18365 12435 18485 12475
rect 18755 12435 18759 12572
rect 18934 12475 19035 12572
rect 18915 12435 19035 12475
rect 725 12428 842 12435
rect 885 12428 1045 12435
rect 725 12322 808 12428
rect 842 12322 1045 12428
rect 725 12315 765 12322
rect 808 12315 1045 12322
rect 1275 12428 1392 12435
rect 1435 12428 1595 12435
rect 1275 12322 1358 12428
rect 1392 12322 1595 12428
rect 1275 12315 1315 12322
rect 1358 12315 1595 12322
rect 1825 12428 1942 12435
rect 1985 12428 2145 12435
rect 1825 12322 1908 12428
rect 1942 12322 2145 12428
rect 1825 12315 1865 12322
rect 1908 12315 2145 12322
rect 2375 12428 2492 12435
rect 2535 12428 2695 12435
rect 2375 12322 2458 12428
rect 2492 12322 2695 12428
rect 2375 12315 2415 12322
rect 2458 12315 2695 12322
rect 2925 12428 3042 12435
rect 3085 12428 3245 12435
rect 2925 12322 3008 12428
rect 3042 12322 3245 12428
rect 2925 12315 2965 12322
rect 3008 12315 3245 12322
rect 3475 12428 3592 12435
rect 3635 12428 3795 12435
rect 3475 12322 3558 12428
rect 3592 12322 3795 12428
rect 3475 12315 3515 12322
rect 3558 12315 3795 12322
rect 4025 12428 4142 12435
rect 4185 12428 4345 12435
rect 4025 12322 4108 12428
rect 4142 12322 4345 12428
rect 4025 12315 4065 12322
rect 4108 12315 4345 12322
rect 4575 12428 4692 12435
rect 4735 12428 4895 12435
rect 4575 12322 4658 12428
rect 4692 12322 4895 12428
rect 4575 12315 4615 12322
rect 4658 12315 4895 12322
rect 5125 12428 5242 12435
rect 5285 12428 5445 12435
rect 5125 12322 5208 12428
rect 5242 12322 5445 12428
rect 5125 12315 5165 12322
rect 5208 12315 5445 12322
rect 5675 12428 5792 12435
rect 5835 12428 5995 12435
rect 5675 12322 5758 12428
rect 5792 12322 5995 12428
rect 5675 12315 5715 12322
rect 5758 12315 5995 12322
rect 6225 12428 6342 12435
rect 6385 12428 6545 12435
rect 6225 12322 6308 12428
rect 6342 12322 6545 12428
rect 6225 12315 6265 12322
rect 6308 12315 6545 12322
rect 6775 12428 6892 12435
rect 6935 12428 7095 12435
rect 6775 12322 6858 12428
rect 6892 12322 7095 12428
rect 6775 12315 6815 12322
rect 6858 12315 7095 12322
rect 7325 12428 7442 12435
rect 7485 12428 7645 12435
rect 7325 12322 7408 12428
rect 7442 12322 7645 12428
rect 7325 12315 7365 12322
rect 7408 12315 7645 12322
rect 7875 12428 7992 12435
rect 8035 12428 8195 12435
rect 7875 12322 7958 12428
rect 7992 12322 8195 12428
rect 7875 12315 7915 12322
rect 7958 12315 8195 12322
rect 8425 12428 8542 12435
rect 8585 12428 8745 12435
rect 8425 12322 8508 12428
rect 8542 12322 8745 12428
rect 8425 12315 8465 12322
rect 8508 12315 8745 12322
rect 8975 12428 9092 12435
rect 9135 12428 9295 12435
rect 8975 12322 9058 12428
rect 9092 12322 9295 12428
rect 8975 12315 9015 12322
rect 9058 12315 9295 12322
rect 9525 12428 9642 12435
rect 9685 12428 9845 12435
rect 9525 12322 9608 12428
rect 9642 12322 9845 12428
rect 9525 12315 9565 12322
rect 9608 12315 9845 12322
rect 10075 12428 10192 12435
rect 10235 12428 10395 12435
rect 10075 12322 10158 12428
rect 10192 12322 10395 12428
rect 10075 12315 10115 12322
rect 10158 12315 10395 12322
rect 10625 12428 10742 12435
rect 10785 12428 10945 12435
rect 10625 12322 10708 12428
rect 10742 12322 10945 12428
rect 10625 12315 10665 12322
rect 10708 12315 10945 12322
rect 11175 12428 11292 12435
rect 11335 12428 11495 12435
rect 11175 12322 11258 12428
rect 11292 12322 11495 12428
rect 11175 12315 11215 12322
rect 11258 12315 11495 12322
rect 11725 12428 11842 12435
rect 11885 12428 12045 12435
rect 11725 12322 11808 12428
rect 11842 12322 12045 12428
rect 11725 12315 11765 12322
rect 11808 12315 12045 12322
rect 12275 12428 12392 12435
rect 12435 12428 12595 12435
rect 12275 12322 12358 12428
rect 12392 12322 12595 12428
rect 12275 12315 12315 12322
rect 12358 12315 12595 12322
rect 12825 12428 12942 12435
rect 12985 12428 13145 12435
rect 12825 12322 12908 12428
rect 12942 12322 13145 12428
rect 12825 12315 12865 12322
rect 12908 12315 13145 12322
rect 13375 12428 13492 12435
rect 13535 12428 13695 12435
rect 13375 12322 13458 12428
rect 13492 12322 13695 12428
rect 13375 12315 13415 12322
rect 13458 12315 13695 12322
rect 13925 12428 14042 12435
rect 14085 12428 14245 12435
rect 13925 12322 14008 12428
rect 14042 12322 14245 12428
rect 13925 12315 13965 12322
rect 14008 12315 14245 12322
rect 14475 12428 14592 12435
rect 14635 12428 14795 12435
rect 14475 12322 14558 12428
rect 14592 12322 14795 12428
rect 14475 12315 14515 12322
rect 14558 12315 14795 12322
rect 15025 12428 15142 12435
rect 15185 12428 15345 12435
rect 15025 12322 15108 12428
rect 15142 12322 15345 12428
rect 15025 12315 15065 12322
rect 15108 12315 15345 12322
rect 15575 12428 15692 12435
rect 15735 12428 15895 12435
rect 15575 12322 15658 12428
rect 15692 12322 15895 12428
rect 15575 12315 15615 12322
rect 15658 12315 15895 12322
rect 16125 12428 16242 12435
rect 16285 12428 16445 12435
rect 16125 12322 16208 12428
rect 16242 12322 16445 12428
rect 16125 12315 16165 12322
rect 16208 12315 16445 12322
rect 16675 12428 16792 12435
rect 16835 12428 16995 12435
rect 16675 12322 16758 12428
rect 16792 12322 16995 12428
rect 16675 12315 16715 12322
rect 16758 12315 16995 12322
rect 17225 12428 17342 12435
rect 17385 12428 17545 12435
rect 17225 12322 17308 12428
rect 17342 12322 17545 12428
rect 17225 12315 17265 12322
rect 17308 12315 17545 12322
rect 17775 12428 17892 12435
rect 17935 12428 18095 12435
rect 17775 12322 17858 12428
rect 17892 12322 18095 12428
rect 17775 12315 17815 12322
rect 17858 12315 18095 12322
rect 18325 12428 18442 12435
rect 18485 12428 18645 12435
rect 18325 12322 18408 12428
rect 18442 12322 18645 12428
rect 18325 12315 18365 12322
rect 18408 12315 18645 12322
rect 18875 12428 18992 12435
rect 19035 12428 19195 12435
rect 18875 12322 18958 12428
rect 18992 12322 19195 12428
rect 18875 12315 18915 12322
rect 18958 12315 19195 12322
rect 765 12275 885 12315
rect 1315 12275 1435 12315
rect 1865 12275 1985 12315
rect 2415 12275 2535 12315
rect 2965 12275 3085 12315
rect 3515 12275 3635 12315
rect 4065 12275 4185 12315
rect 4615 12275 4735 12315
rect 5165 12275 5285 12315
rect 5715 12275 5835 12315
rect 6265 12275 6385 12315
rect 6815 12275 6935 12315
rect 7365 12275 7485 12315
rect 7915 12275 8035 12315
rect 8465 12275 8585 12315
rect 9015 12275 9135 12315
rect 9565 12275 9685 12315
rect 10115 12275 10235 12315
rect 10665 12275 10785 12315
rect 11215 12275 11335 12315
rect 11765 12275 11885 12315
rect 12315 12275 12435 12315
rect 12865 12275 12985 12315
rect 13415 12275 13535 12315
rect 13965 12275 14085 12315
rect 14515 12275 14635 12315
rect 15065 12275 15185 12315
rect 15615 12275 15735 12315
rect 16165 12275 16285 12315
rect 16715 12275 16835 12315
rect 17265 12275 17385 12315
rect 17815 12275 17935 12315
rect 18365 12275 18485 12315
rect 18915 12275 19035 12315
rect 19185 12154 19200 12171
rect 19202 12162 19204 12588
rect 19202 12148 19217 12154
rect 500 12075 507 12125
rect 500 11639 525 12040
rect 628 12022 885 12045
rect 1178 12022 1435 12045
rect 1728 12022 1985 12045
rect 2278 12022 2535 12045
rect 2828 12022 3085 12045
rect 3378 12022 3635 12045
rect 3928 12022 4185 12045
rect 4478 12022 4735 12045
rect 5028 12022 5285 12045
rect 5578 12022 5835 12045
rect 6128 12022 6385 12045
rect 6678 12022 6935 12045
rect 7228 12022 7485 12045
rect 7778 12022 8035 12045
rect 8328 12022 8585 12045
rect 8878 12022 9135 12045
rect 9428 12022 9685 12045
rect 9978 12022 10235 12045
rect 10528 12022 10785 12045
rect 11078 12022 11335 12045
rect 11628 12022 11885 12045
rect 12178 12022 12435 12045
rect 12728 12022 12985 12045
rect 13278 12022 13535 12045
rect 13828 12022 14085 12045
rect 14378 12022 14635 12045
rect 14928 12022 15185 12045
rect 15478 12022 15735 12045
rect 16028 12022 16285 12045
rect 16578 12022 16835 12045
rect 17128 12022 17385 12045
rect 17678 12022 17935 12045
rect 18228 12022 18485 12045
rect 18778 12022 19035 12045
rect 605 11885 609 12022
rect 784 11925 885 12022
rect 765 11885 885 11925
rect 1155 11885 1159 12022
rect 1334 11925 1435 12022
rect 1315 11885 1435 11925
rect 1705 11885 1709 12022
rect 1884 11925 1985 12022
rect 1865 11885 1985 11925
rect 2255 11885 2259 12022
rect 2434 11925 2535 12022
rect 2415 11885 2535 11925
rect 2805 11885 2809 12022
rect 2984 11925 3085 12022
rect 2965 11885 3085 11925
rect 3355 11885 3359 12022
rect 3534 11925 3635 12022
rect 3515 11885 3635 11925
rect 3905 11885 3909 12022
rect 4084 11925 4185 12022
rect 4065 11885 4185 11925
rect 4455 11885 4459 12022
rect 4634 11925 4735 12022
rect 4615 11885 4735 11925
rect 5005 11885 5009 12022
rect 5184 11925 5285 12022
rect 5165 11885 5285 11925
rect 5555 11885 5559 12022
rect 5734 11925 5835 12022
rect 5715 11885 5835 11925
rect 6105 11885 6109 12022
rect 6284 11925 6385 12022
rect 6265 11885 6385 11925
rect 6655 11885 6659 12022
rect 6834 11925 6935 12022
rect 6815 11885 6935 11925
rect 7205 11885 7209 12022
rect 7384 11925 7485 12022
rect 7365 11885 7485 11925
rect 7755 11885 7759 12022
rect 7934 11925 8035 12022
rect 7915 11885 8035 11925
rect 8305 11885 8309 12022
rect 8484 11925 8585 12022
rect 8465 11885 8585 11925
rect 8855 11885 8859 12022
rect 9034 11925 9135 12022
rect 9015 11885 9135 11925
rect 9405 11885 9409 12022
rect 9584 11925 9685 12022
rect 9565 11885 9685 11925
rect 9955 11885 9959 12022
rect 10134 11925 10235 12022
rect 10115 11885 10235 11925
rect 10505 11885 10509 12022
rect 10684 11925 10785 12022
rect 10665 11885 10785 11925
rect 11055 11885 11059 12022
rect 11234 11925 11335 12022
rect 11215 11885 11335 11925
rect 11605 11885 11609 12022
rect 11784 11925 11885 12022
rect 11765 11885 11885 11925
rect 12155 11885 12159 12022
rect 12334 11925 12435 12022
rect 12315 11885 12435 11925
rect 12705 11885 12709 12022
rect 12884 11925 12985 12022
rect 12865 11885 12985 11925
rect 13255 11885 13259 12022
rect 13434 11925 13535 12022
rect 13415 11885 13535 11925
rect 13805 11885 13809 12022
rect 13984 11925 14085 12022
rect 13965 11885 14085 11925
rect 14355 11885 14359 12022
rect 14534 11925 14635 12022
rect 14515 11885 14635 11925
rect 14905 11885 14909 12022
rect 15084 11925 15185 12022
rect 15065 11885 15185 11925
rect 15455 11885 15459 12022
rect 15634 11925 15735 12022
rect 15615 11885 15735 11925
rect 16005 11885 16009 12022
rect 16184 11925 16285 12022
rect 16165 11885 16285 11925
rect 16555 11885 16559 12022
rect 16734 11925 16835 12022
rect 16715 11885 16835 11925
rect 17105 11885 17109 12022
rect 17284 11925 17385 12022
rect 17265 11885 17385 11925
rect 17655 11885 17659 12022
rect 17834 11925 17935 12022
rect 17815 11885 17935 11925
rect 18205 11885 18209 12022
rect 18384 11925 18485 12022
rect 18365 11885 18485 11925
rect 18755 11885 18759 12022
rect 18934 11925 19035 12022
rect 18915 11885 19035 11925
rect 725 11878 842 11885
rect 885 11878 1045 11885
rect 725 11772 808 11878
rect 842 11772 1045 11878
rect 725 11765 765 11772
rect 808 11765 1045 11772
rect 1275 11878 1392 11885
rect 1435 11878 1595 11885
rect 1275 11772 1358 11878
rect 1392 11772 1595 11878
rect 1275 11765 1315 11772
rect 1358 11765 1595 11772
rect 1825 11878 1942 11885
rect 1985 11878 2145 11885
rect 1825 11772 1908 11878
rect 1942 11772 2145 11878
rect 1825 11765 1865 11772
rect 1908 11765 2145 11772
rect 2375 11878 2492 11885
rect 2535 11878 2695 11885
rect 2375 11772 2458 11878
rect 2492 11772 2695 11878
rect 2375 11765 2415 11772
rect 2458 11765 2695 11772
rect 2925 11878 3042 11885
rect 3085 11878 3245 11885
rect 2925 11772 3008 11878
rect 3042 11772 3245 11878
rect 2925 11765 2965 11772
rect 3008 11765 3245 11772
rect 3475 11878 3592 11885
rect 3635 11878 3795 11885
rect 3475 11772 3558 11878
rect 3592 11772 3795 11878
rect 3475 11765 3515 11772
rect 3558 11765 3795 11772
rect 4025 11878 4142 11885
rect 4185 11878 4345 11885
rect 4025 11772 4108 11878
rect 4142 11772 4345 11878
rect 4025 11765 4065 11772
rect 4108 11765 4345 11772
rect 4575 11878 4692 11885
rect 4735 11878 4895 11885
rect 4575 11772 4658 11878
rect 4692 11772 4895 11878
rect 4575 11765 4615 11772
rect 4658 11765 4895 11772
rect 5125 11878 5242 11885
rect 5285 11878 5445 11885
rect 5125 11772 5208 11878
rect 5242 11772 5445 11878
rect 5125 11765 5165 11772
rect 5208 11765 5445 11772
rect 5675 11878 5792 11885
rect 5835 11878 5995 11885
rect 5675 11772 5758 11878
rect 5792 11772 5995 11878
rect 5675 11765 5715 11772
rect 5758 11765 5995 11772
rect 6225 11878 6342 11885
rect 6385 11878 6545 11885
rect 6225 11772 6308 11878
rect 6342 11772 6545 11878
rect 6225 11765 6265 11772
rect 6308 11765 6545 11772
rect 6775 11878 6892 11885
rect 6935 11878 7095 11885
rect 6775 11772 6858 11878
rect 6892 11772 7095 11878
rect 6775 11765 6815 11772
rect 6858 11765 7095 11772
rect 7325 11878 7442 11885
rect 7485 11878 7645 11885
rect 7325 11772 7408 11878
rect 7442 11772 7645 11878
rect 7325 11765 7365 11772
rect 7408 11765 7645 11772
rect 7875 11878 7992 11885
rect 8035 11878 8195 11885
rect 7875 11772 7958 11878
rect 7992 11772 8195 11878
rect 7875 11765 7915 11772
rect 7958 11765 8195 11772
rect 8425 11878 8542 11885
rect 8585 11878 8745 11885
rect 8425 11772 8508 11878
rect 8542 11772 8745 11878
rect 8425 11765 8465 11772
rect 8508 11765 8745 11772
rect 8975 11878 9092 11885
rect 9135 11878 9295 11885
rect 8975 11772 9058 11878
rect 9092 11772 9295 11878
rect 8975 11765 9015 11772
rect 9058 11765 9295 11772
rect 9525 11878 9642 11885
rect 9685 11878 9845 11885
rect 9525 11772 9608 11878
rect 9642 11772 9845 11878
rect 9525 11765 9565 11772
rect 9608 11765 9845 11772
rect 10075 11878 10192 11885
rect 10235 11878 10395 11885
rect 10075 11772 10158 11878
rect 10192 11772 10395 11878
rect 10075 11765 10115 11772
rect 10158 11765 10395 11772
rect 10625 11878 10742 11885
rect 10785 11878 10945 11885
rect 10625 11772 10708 11878
rect 10742 11772 10945 11878
rect 10625 11765 10665 11772
rect 10708 11765 10945 11772
rect 11175 11878 11292 11885
rect 11335 11878 11495 11885
rect 11175 11772 11258 11878
rect 11292 11772 11495 11878
rect 11175 11765 11215 11772
rect 11258 11765 11495 11772
rect 11725 11878 11842 11885
rect 11885 11878 12045 11885
rect 11725 11772 11808 11878
rect 11842 11772 12045 11878
rect 11725 11765 11765 11772
rect 11808 11765 12045 11772
rect 12275 11878 12392 11885
rect 12435 11878 12595 11885
rect 12275 11772 12358 11878
rect 12392 11772 12595 11878
rect 12275 11765 12315 11772
rect 12358 11765 12595 11772
rect 12825 11878 12942 11885
rect 12985 11878 13145 11885
rect 12825 11772 12908 11878
rect 12942 11772 13145 11878
rect 12825 11765 12865 11772
rect 12908 11765 13145 11772
rect 13375 11878 13492 11885
rect 13535 11878 13695 11885
rect 13375 11772 13458 11878
rect 13492 11772 13695 11878
rect 13375 11765 13415 11772
rect 13458 11765 13695 11772
rect 13925 11878 14042 11885
rect 14085 11878 14245 11885
rect 13925 11772 14008 11878
rect 14042 11772 14245 11878
rect 13925 11765 13965 11772
rect 14008 11765 14245 11772
rect 14475 11878 14592 11885
rect 14635 11878 14795 11885
rect 14475 11772 14558 11878
rect 14592 11772 14795 11878
rect 14475 11765 14515 11772
rect 14558 11765 14795 11772
rect 15025 11878 15142 11885
rect 15185 11878 15345 11885
rect 15025 11772 15108 11878
rect 15142 11772 15345 11878
rect 15025 11765 15065 11772
rect 15108 11765 15345 11772
rect 15575 11878 15692 11885
rect 15735 11878 15895 11885
rect 15575 11772 15658 11878
rect 15692 11772 15895 11878
rect 15575 11765 15615 11772
rect 15658 11765 15895 11772
rect 16125 11878 16242 11885
rect 16285 11878 16445 11885
rect 16125 11772 16208 11878
rect 16242 11772 16445 11878
rect 16125 11765 16165 11772
rect 16208 11765 16445 11772
rect 16675 11878 16792 11885
rect 16835 11878 16995 11885
rect 16675 11772 16758 11878
rect 16792 11772 16995 11878
rect 16675 11765 16715 11772
rect 16758 11765 16995 11772
rect 17225 11878 17342 11885
rect 17385 11878 17545 11885
rect 17225 11772 17308 11878
rect 17342 11772 17545 11878
rect 17225 11765 17265 11772
rect 17308 11765 17545 11772
rect 17775 11878 17892 11885
rect 17935 11878 18095 11885
rect 17775 11772 17858 11878
rect 17892 11772 18095 11878
rect 17775 11765 17815 11772
rect 17858 11765 18095 11772
rect 18325 11878 18442 11885
rect 18485 11878 18645 11885
rect 18325 11772 18408 11878
rect 18442 11772 18645 11878
rect 18325 11765 18365 11772
rect 18408 11765 18645 11772
rect 18875 11878 18992 11885
rect 19035 11878 19195 11885
rect 18875 11772 18958 11878
rect 18992 11772 19195 11878
rect 18875 11765 18915 11772
rect 18958 11765 19195 11772
rect 765 11725 885 11765
rect 1315 11725 1435 11765
rect 1865 11725 1985 11765
rect 2415 11725 2535 11765
rect 2965 11725 3085 11765
rect 3515 11725 3635 11765
rect 4065 11725 4185 11765
rect 4615 11725 4735 11765
rect 5165 11725 5285 11765
rect 5715 11725 5835 11765
rect 6265 11725 6385 11765
rect 6815 11725 6935 11765
rect 7365 11725 7485 11765
rect 7915 11725 8035 11765
rect 8465 11725 8585 11765
rect 9015 11725 9135 11765
rect 9565 11725 9685 11765
rect 10115 11725 10235 11765
rect 10665 11725 10785 11765
rect 11215 11725 11335 11765
rect 11765 11725 11885 11765
rect 12315 11725 12435 11765
rect 12865 11725 12985 11765
rect 13415 11725 13535 11765
rect 13965 11725 14085 11765
rect 14515 11725 14635 11765
rect 15065 11725 15185 11765
rect 15615 11725 15735 11765
rect 16165 11725 16285 11765
rect 16715 11725 16835 11765
rect 17265 11725 17385 11765
rect 17815 11725 17935 11765
rect 18365 11725 18485 11765
rect 18915 11725 19035 11765
rect 19202 11612 19204 12038
rect 500 11525 507 11575
rect 19202 11496 19217 11502
rect 628 11472 885 11495
rect 1178 11472 1435 11495
rect 1728 11472 1985 11495
rect 2278 11472 2535 11495
rect 2828 11472 3085 11495
rect 3378 11472 3635 11495
rect 3928 11472 4185 11495
rect 4478 11472 4735 11495
rect 5028 11472 5285 11495
rect 5578 11472 5835 11495
rect 6128 11472 6385 11495
rect 6678 11472 6935 11495
rect 7228 11472 7485 11495
rect 7778 11472 8035 11495
rect 8328 11472 8585 11495
rect 8878 11472 9135 11495
rect 9428 11472 9685 11495
rect 9978 11472 10235 11495
rect 10528 11472 10785 11495
rect 11078 11472 11335 11495
rect 11628 11472 11885 11495
rect 12178 11472 12435 11495
rect 12728 11472 12985 11495
rect 13278 11472 13535 11495
rect 13828 11472 14085 11495
rect 14378 11472 14635 11495
rect 14928 11472 15185 11495
rect 15478 11472 15735 11495
rect 16028 11472 16285 11495
rect 16578 11472 16835 11495
rect 17128 11472 17385 11495
rect 17678 11472 17935 11495
rect 18228 11472 18485 11495
rect 18778 11472 19035 11495
rect 605 11335 609 11472
rect 784 11375 885 11472
rect 765 11335 885 11375
rect 1155 11335 1159 11472
rect 1334 11375 1435 11472
rect 1315 11335 1435 11375
rect 1705 11335 1709 11472
rect 1884 11375 1985 11472
rect 1865 11335 1985 11375
rect 2255 11335 2259 11472
rect 2434 11375 2535 11472
rect 2415 11335 2535 11375
rect 2805 11335 2809 11472
rect 2984 11375 3085 11472
rect 2965 11335 3085 11375
rect 3355 11335 3359 11472
rect 3534 11375 3635 11472
rect 3515 11335 3635 11375
rect 3905 11335 3909 11472
rect 4084 11375 4185 11472
rect 4065 11335 4185 11375
rect 4455 11335 4459 11472
rect 4634 11375 4735 11472
rect 4615 11335 4735 11375
rect 5005 11335 5009 11472
rect 5184 11375 5285 11472
rect 5165 11335 5285 11375
rect 5555 11335 5559 11472
rect 5734 11375 5835 11472
rect 5715 11335 5835 11375
rect 6105 11335 6109 11472
rect 6284 11375 6385 11472
rect 6265 11335 6385 11375
rect 6655 11335 6659 11472
rect 6834 11375 6935 11472
rect 6815 11335 6935 11375
rect 7205 11335 7209 11472
rect 7384 11375 7485 11472
rect 7365 11335 7485 11375
rect 7755 11335 7759 11472
rect 7934 11375 8035 11472
rect 7915 11335 8035 11375
rect 8305 11335 8309 11472
rect 8484 11375 8585 11472
rect 8465 11335 8585 11375
rect 8855 11335 8859 11472
rect 9034 11375 9135 11472
rect 9015 11335 9135 11375
rect 9405 11335 9409 11472
rect 9584 11375 9685 11472
rect 9565 11335 9685 11375
rect 9955 11335 9959 11472
rect 10134 11375 10235 11472
rect 10115 11335 10235 11375
rect 10505 11335 10509 11472
rect 10684 11375 10785 11472
rect 10665 11335 10785 11375
rect 11055 11335 11059 11472
rect 11234 11375 11335 11472
rect 11215 11335 11335 11375
rect 11605 11335 11609 11472
rect 11784 11375 11885 11472
rect 11765 11335 11885 11375
rect 12155 11335 12159 11472
rect 12334 11375 12435 11472
rect 12315 11335 12435 11375
rect 12705 11335 12709 11472
rect 12884 11375 12985 11472
rect 12865 11335 12985 11375
rect 13255 11335 13259 11472
rect 13434 11375 13535 11472
rect 13415 11335 13535 11375
rect 13805 11335 13809 11472
rect 13984 11375 14085 11472
rect 13965 11335 14085 11375
rect 14355 11335 14359 11472
rect 14534 11375 14635 11472
rect 14515 11335 14635 11375
rect 14905 11335 14909 11472
rect 15084 11375 15185 11472
rect 15065 11335 15185 11375
rect 15455 11335 15459 11472
rect 15634 11375 15735 11472
rect 15615 11335 15735 11375
rect 16005 11335 16009 11472
rect 16184 11375 16285 11472
rect 16165 11335 16285 11375
rect 16555 11335 16559 11472
rect 16734 11375 16835 11472
rect 16715 11335 16835 11375
rect 17105 11335 17109 11472
rect 17284 11375 17385 11472
rect 17265 11335 17385 11375
rect 17655 11335 17659 11472
rect 17834 11375 17935 11472
rect 17815 11335 17935 11375
rect 18205 11335 18209 11472
rect 18384 11375 18485 11472
rect 18365 11335 18485 11375
rect 18755 11335 18759 11472
rect 18934 11375 19035 11472
rect 18915 11335 19035 11375
rect 725 11328 842 11335
rect 885 11328 1045 11335
rect 725 11222 808 11328
rect 842 11222 1045 11328
rect 725 11215 765 11222
rect 808 11215 1045 11222
rect 1275 11328 1392 11335
rect 1435 11328 1595 11335
rect 1275 11222 1358 11328
rect 1392 11222 1595 11328
rect 1275 11215 1315 11222
rect 1358 11215 1595 11222
rect 1825 11328 1942 11335
rect 1985 11328 2145 11335
rect 1825 11222 1908 11328
rect 1942 11222 2145 11328
rect 1825 11215 1865 11222
rect 1908 11215 2145 11222
rect 2375 11328 2492 11335
rect 2535 11328 2695 11335
rect 2375 11222 2458 11328
rect 2492 11222 2695 11328
rect 2375 11215 2415 11222
rect 2458 11215 2695 11222
rect 2925 11328 3042 11335
rect 3085 11328 3245 11335
rect 2925 11222 3008 11328
rect 3042 11222 3245 11328
rect 2925 11215 2965 11222
rect 3008 11215 3245 11222
rect 3475 11328 3592 11335
rect 3635 11328 3795 11335
rect 3475 11222 3558 11328
rect 3592 11222 3795 11328
rect 3475 11215 3515 11222
rect 3558 11215 3795 11222
rect 4025 11328 4142 11335
rect 4185 11328 4345 11335
rect 4025 11222 4108 11328
rect 4142 11222 4345 11328
rect 4025 11215 4065 11222
rect 4108 11215 4345 11222
rect 4575 11328 4692 11335
rect 4735 11328 4895 11335
rect 4575 11222 4658 11328
rect 4692 11222 4895 11328
rect 4575 11215 4615 11222
rect 4658 11215 4895 11222
rect 5125 11328 5242 11335
rect 5285 11328 5445 11335
rect 5125 11222 5208 11328
rect 5242 11222 5445 11328
rect 5125 11215 5165 11222
rect 5208 11215 5445 11222
rect 5675 11328 5792 11335
rect 5835 11328 5995 11335
rect 5675 11222 5758 11328
rect 5792 11222 5995 11328
rect 5675 11215 5715 11222
rect 5758 11215 5995 11222
rect 6225 11328 6342 11335
rect 6385 11328 6545 11335
rect 6225 11222 6308 11328
rect 6342 11222 6545 11328
rect 6225 11215 6265 11222
rect 6308 11215 6545 11222
rect 6775 11328 6892 11335
rect 6935 11328 7095 11335
rect 6775 11222 6858 11328
rect 6892 11222 7095 11328
rect 6775 11215 6815 11222
rect 6858 11215 7095 11222
rect 7325 11328 7442 11335
rect 7485 11328 7645 11335
rect 7325 11222 7408 11328
rect 7442 11222 7645 11328
rect 7325 11215 7365 11222
rect 7408 11215 7645 11222
rect 7875 11328 7992 11335
rect 8035 11328 8195 11335
rect 7875 11222 7958 11328
rect 7992 11222 8195 11328
rect 7875 11215 7915 11222
rect 7958 11215 8195 11222
rect 8425 11328 8542 11335
rect 8585 11328 8745 11335
rect 8425 11222 8508 11328
rect 8542 11222 8745 11328
rect 8425 11215 8465 11222
rect 8508 11215 8745 11222
rect 8975 11328 9092 11335
rect 9135 11328 9295 11335
rect 8975 11222 9058 11328
rect 9092 11222 9295 11328
rect 8975 11215 9015 11222
rect 9058 11215 9295 11222
rect 9525 11328 9642 11335
rect 9685 11328 9845 11335
rect 9525 11222 9608 11328
rect 9642 11222 9845 11328
rect 9525 11215 9565 11222
rect 9608 11215 9845 11222
rect 10075 11328 10192 11335
rect 10235 11328 10395 11335
rect 10075 11222 10158 11328
rect 10192 11222 10395 11328
rect 10075 11215 10115 11222
rect 10158 11215 10395 11222
rect 10625 11328 10742 11335
rect 10785 11328 10945 11335
rect 10625 11222 10708 11328
rect 10742 11222 10945 11328
rect 10625 11215 10665 11222
rect 10708 11215 10945 11222
rect 11175 11328 11292 11335
rect 11335 11328 11495 11335
rect 11175 11222 11258 11328
rect 11292 11222 11495 11328
rect 11175 11215 11215 11222
rect 11258 11215 11495 11222
rect 11725 11328 11842 11335
rect 11885 11328 12045 11335
rect 11725 11222 11808 11328
rect 11842 11222 12045 11328
rect 11725 11215 11765 11222
rect 11808 11215 12045 11222
rect 12275 11328 12392 11335
rect 12435 11328 12595 11335
rect 12275 11222 12358 11328
rect 12392 11222 12595 11328
rect 12275 11215 12315 11222
rect 12358 11215 12595 11222
rect 12825 11328 12942 11335
rect 12985 11328 13145 11335
rect 12825 11222 12908 11328
rect 12942 11222 13145 11328
rect 12825 11215 12865 11222
rect 12908 11215 13145 11222
rect 13375 11328 13492 11335
rect 13535 11328 13695 11335
rect 13375 11222 13458 11328
rect 13492 11222 13695 11328
rect 13375 11215 13415 11222
rect 13458 11215 13695 11222
rect 13925 11328 14042 11335
rect 14085 11328 14245 11335
rect 13925 11222 14008 11328
rect 14042 11222 14245 11328
rect 13925 11215 13965 11222
rect 14008 11215 14245 11222
rect 14475 11328 14592 11335
rect 14635 11328 14795 11335
rect 14475 11222 14558 11328
rect 14592 11222 14795 11328
rect 14475 11215 14515 11222
rect 14558 11215 14795 11222
rect 15025 11328 15142 11335
rect 15185 11328 15345 11335
rect 15025 11222 15108 11328
rect 15142 11222 15345 11328
rect 15025 11215 15065 11222
rect 15108 11215 15345 11222
rect 15575 11328 15692 11335
rect 15735 11328 15895 11335
rect 15575 11222 15658 11328
rect 15692 11222 15895 11328
rect 15575 11215 15615 11222
rect 15658 11215 15895 11222
rect 16125 11328 16242 11335
rect 16285 11328 16445 11335
rect 16125 11222 16208 11328
rect 16242 11222 16445 11328
rect 16125 11215 16165 11222
rect 16208 11215 16445 11222
rect 16675 11328 16792 11335
rect 16835 11328 16995 11335
rect 16675 11222 16758 11328
rect 16792 11222 16995 11328
rect 16675 11215 16715 11222
rect 16758 11215 16995 11222
rect 17225 11328 17342 11335
rect 17385 11328 17545 11335
rect 17225 11222 17308 11328
rect 17342 11222 17545 11328
rect 17225 11215 17265 11222
rect 17308 11215 17545 11222
rect 17775 11328 17892 11335
rect 17935 11328 18095 11335
rect 17775 11222 17858 11328
rect 17892 11222 18095 11328
rect 17775 11215 17815 11222
rect 17858 11215 18095 11222
rect 18325 11328 18442 11335
rect 18485 11328 18645 11335
rect 18325 11222 18408 11328
rect 18442 11222 18645 11328
rect 18325 11215 18365 11222
rect 18408 11215 18645 11222
rect 18875 11328 18992 11335
rect 19035 11328 19195 11335
rect 18875 11222 18958 11328
rect 18992 11222 19195 11328
rect 18875 11215 18915 11222
rect 18958 11215 19195 11222
rect 765 11175 885 11215
rect 1315 11175 1435 11215
rect 1865 11175 1985 11215
rect 2415 11175 2535 11215
rect 2965 11175 3085 11215
rect 3515 11175 3635 11215
rect 4065 11175 4185 11215
rect 4615 11175 4735 11215
rect 5165 11175 5285 11215
rect 5715 11175 5835 11215
rect 6265 11175 6385 11215
rect 6815 11175 6935 11215
rect 7365 11175 7485 11215
rect 7915 11175 8035 11215
rect 8465 11175 8585 11215
rect 9015 11175 9135 11215
rect 9565 11175 9685 11215
rect 10115 11175 10235 11215
rect 10665 11175 10785 11215
rect 11215 11175 11335 11215
rect 11765 11175 11885 11215
rect 12315 11175 12435 11215
rect 12865 11175 12985 11215
rect 13415 11175 13535 11215
rect 13965 11175 14085 11215
rect 14515 11175 14635 11215
rect 15065 11175 15185 11215
rect 15615 11175 15735 11215
rect 16165 11175 16285 11215
rect 16715 11175 16835 11215
rect 17265 11175 17385 11215
rect 17815 11175 17935 11215
rect 18365 11175 18485 11215
rect 18915 11175 19035 11215
rect 19185 11054 19200 11071
rect 19202 11062 19204 11488
rect 19202 11048 19217 11054
rect 500 10975 507 11025
rect 500 10539 525 10940
rect 628 10922 885 10945
rect 1178 10922 1435 10945
rect 1728 10922 1985 10945
rect 2278 10922 2535 10945
rect 2828 10922 3085 10945
rect 3378 10922 3635 10945
rect 3928 10922 4185 10945
rect 4478 10922 4735 10945
rect 5028 10922 5285 10945
rect 5578 10922 5835 10945
rect 6128 10922 6385 10945
rect 6678 10922 6935 10945
rect 7228 10922 7485 10945
rect 7778 10922 8035 10945
rect 8328 10922 8585 10945
rect 8878 10922 9135 10945
rect 9428 10922 9685 10945
rect 9978 10922 10235 10945
rect 10528 10922 10785 10945
rect 11078 10922 11335 10945
rect 11628 10922 11885 10945
rect 12178 10922 12435 10945
rect 12728 10922 12985 10945
rect 13278 10922 13535 10945
rect 13828 10922 14085 10945
rect 14378 10922 14635 10945
rect 14928 10922 15185 10945
rect 15478 10922 15735 10945
rect 16028 10922 16285 10945
rect 16578 10922 16835 10945
rect 17128 10922 17385 10945
rect 17678 10922 17935 10945
rect 18228 10922 18485 10945
rect 18778 10922 19035 10945
rect 605 10785 609 10922
rect 784 10825 885 10922
rect 765 10785 885 10825
rect 1155 10785 1159 10922
rect 1334 10825 1435 10922
rect 1315 10785 1435 10825
rect 1705 10785 1709 10922
rect 1884 10825 1985 10922
rect 1865 10785 1985 10825
rect 2255 10785 2259 10922
rect 2434 10825 2535 10922
rect 2415 10785 2535 10825
rect 2805 10785 2809 10922
rect 2984 10825 3085 10922
rect 2965 10785 3085 10825
rect 3355 10785 3359 10922
rect 3534 10825 3635 10922
rect 3515 10785 3635 10825
rect 3905 10785 3909 10922
rect 4084 10825 4185 10922
rect 4065 10785 4185 10825
rect 4455 10785 4459 10922
rect 4634 10825 4735 10922
rect 4615 10785 4735 10825
rect 5005 10785 5009 10922
rect 5184 10825 5285 10922
rect 5165 10785 5285 10825
rect 5555 10785 5559 10922
rect 5734 10825 5835 10922
rect 5715 10785 5835 10825
rect 6105 10785 6109 10922
rect 6284 10825 6385 10922
rect 6265 10785 6385 10825
rect 6655 10785 6659 10922
rect 6834 10825 6935 10922
rect 6815 10785 6935 10825
rect 7205 10785 7209 10922
rect 7384 10825 7485 10922
rect 7365 10785 7485 10825
rect 7755 10785 7759 10922
rect 7934 10825 8035 10922
rect 7915 10785 8035 10825
rect 8305 10785 8309 10922
rect 8484 10825 8585 10922
rect 8465 10785 8585 10825
rect 8855 10785 8859 10922
rect 9034 10825 9135 10922
rect 9015 10785 9135 10825
rect 9405 10785 9409 10922
rect 9584 10825 9685 10922
rect 9565 10785 9685 10825
rect 9955 10785 9959 10922
rect 10134 10825 10235 10922
rect 10115 10785 10235 10825
rect 10505 10785 10509 10922
rect 10684 10825 10785 10922
rect 10665 10785 10785 10825
rect 11055 10785 11059 10922
rect 11234 10825 11335 10922
rect 11215 10785 11335 10825
rect 11605 10785 11609 10922
rect 11784 10825 11885 10922
rect 11765 10785 11885 10825
rect 12155 10785 12159 10922
rect 12334 10825 12435 10922
rect 12315 10785 12435 10825
rect 12705 10785 12709 10922
rect 12884 10825 12985 10922
rect 12865 10785 12985 10825
rect 13255 10785 13259 10922
rect 13434 10825 13535 10922
rect 13415 10785 13535 10825
rect 13805 10785 13809 10922
rect 13984 10825 14085 10922
rect 13965 10785 14085 10825
rect 14355 10785 14359 10922
rect 14534 10825 14635 10922
rect 14515 10785 14635 10825
rect 14905 10785 14909 10922
rect 15084 10825 15185 10922
rect 15065 10785 15185 10825
rect 15455 10785 15459 10922
rect 15634 10825 15735 10922
rect 15615 10785 15735 10825
rect 16005 10785 16009 10922
rect 16184 10825 16285 10922
rect 16165 10785 16285 10825
rect 16555 10785 16559 10922
rect 16734 10825 16835 10922
rect 16715 10785 16835 10825
rect 17105 10785 17109 10922
rect 17284 10825 17385 10922
rect 17265 10785 17385 10825
rect 17655 10785 17659 10922
rect 17834 10825 17935 10922
rect 17815 10785 17935 10825
rect 18205 10785 18209 10922
rect 18384 10825 18485 10922
rect 18365 10785 18485 10825
rect 18755 10785 18759 10922
rect 18934 10825 19035 10922
rect 18915 10785 19035 10825
rect 725 10778 842 10785
rect 885 10778 1045 10785
rect 725 10672 808 10778
rect 842 10672 1045 10778
rect 725 10665 765 10672
rect 808 10665 1045 10672
rect 1275 10778 1392 10785
rect 1435 10778 1595 10785
rect 1275 10672 1358 10778
rect 1392 10672 1595 10778
rect 1275 10665 1315 10672
rect 1358 10665 1595 10672
rect 1825 10778 1942 10785
rect 1985 10778 2145 10785
rect 1825 10672 1908 10778
rect 1942 10672 2145 10778
rect 1825 10665 1865 10672
rect 1908 10665 2145 10672
rect 2375 10778 2492 10785
rect 2535 10778 2695 10785
rect 2375 10672 2458 10778
rect 2492 10672 2695 10778
rect 2375 10665 2415 10672
rect 2458 10665 2695 10672
rect 2925 10778 3042 10785
rect 3085 10778 3245 10785
rect 2925 10672 3008 10778
rect 3042 10672 3245 10778
rect 2925 10665 2965 10672
rect 3008 10665 3245 10672
rect 3475 10778 3592 10785
rect 3635 10778 3795 10785
rect 3475 10672 3558 10778
rect 3592 10672 3795 10778
rect 3475 10665 3515 10672
rect 3558 10665 3795 10672
rect 4025 10778 4142 10785
rect 4185 10778 4345 10785
rect 4025 10672 4108 10778
rect 4142 10672 4345 10778
rect 4025 10665 4065 10672
rect 4108 10665 4345 10672
rect 4575 10778 4692 10785
rect 4735 10778 4895 10785
rect 4575 10672 4658 10778
rect 4692 10672 4895 10778
rect 4575 10665 4615 10672
rect 4658 10665 4895 10672
rect 5125 10778 5242 10785
rect 5285 10778 5445 10785
rect 5125 10672 5208 10778
rect 5242 10672 5445 10778
rect 5125 10665 5165 10672
rect 5208 10665 5445 10672
rect 5675 10778 5792 10785
rect 5835 10778 5995 10785
rect 5675 10672 5758 10778
rect 5792 10672 5995 10778
rect 5675 10665 5715 10672
rect 5758 10665 5995 10672
rect 6225 10778 6342 10785
rect 6385 10778 6545 10785
rect 6225 10672 6308 10778
rect 6342 10672 6545 10778
rect 6225 10665 6265 10672
rect 6308 10665 6545 10672
rect 6775 10778 6892 10785
rect 6935 10778 7095 10785
rect 6775 10672 6858 10778
rect 6892 10672 7095 10778
rect 6775 10665 6815 10672
rect 6858 10665 7095 10672
rect 7325 10778 7442 10785
rect 7485 10778 7645 10785
rect 7325 10672 7408 10778
rect 7442 10672 7645 10778
rect 7325 10665 7365 10672
rect 7408 10665 7645 10672
rect 7875 10778 7992 10785
rect 8035 10778 8195 10785
rect 7875 10672 7958 10778
rect 7992 10672 8195 10778
rect 7875 10665 7915 10672
rect 7958 10665 8195 10672
rect 8425 10778 8542 10785
rect 8585 10778 8745 10785
rect 8425 10672 8508 10778
rect 8542 10672 8745 10778
rect 8425 10665 8465 10672
rect 8508 10665 8745 10672
rect 8975 10778 9092 10785
rect 9135 10778 9295 10785
rect 8975 10672 9058 10778
rect 9092 10672 9295 10778
rect 8975 10665 9015 10672
rect 9058 10665 9295 10672
rect 9525 10778 9642 10785
rect 9685 10778 9845 10785
rect 9525 10672 9608 10778
rect 9642 10672 9845 10778
rect 9525 10665 9565 10672
rect 9608 10665 9845 10672
rect 10075 10778 10192 10785
rect 10235 10778 10395 10785
rect 10075 10672 10158 10778
rect 10192 10672 10395 10778
rect 10075 10665 10115 10672
rect 10158 10665 10395 10672
rect 10625 10778 10742 10785
rect 10785 10778 10945 10785
rect 10625 10672 10708 10778
rect 10742 10672 10945 10778
rect 10625 10665 10665 10672
rect 10708 10665 10945 10672
rect 11175 10778 11292 10785
rect 11335 10778 11495 10785
rect 11175 10672 11258 10778
rect 11292 10672 11495 10778
rect 11175 10665 11215 10672
rect 11258 10665 11495 10672
rect 11725 10778 11842 10785
rect 11885 10778 12045 10785
rect 11725 10672 11808 10778
rect 11842 10672 12045 10778
rect 11725 10665 11765 10672
rect 11808 10665 12045 10672
rect 12275 10778 12392 10785
rect 12435 10778 12595 10785
rect 12275 10672 12358 10778
rect 12392 10672 12595 10778
rect 12275 10665 12315 10672
rect 12358 10665 12595 10672
rect 12825 10778 12942 10785
rect 12985 10778 13145 10785
rect 12825 10672 12908 10778
rect 12942 10672 13145 10778
rect 12825 10665 12865 10672
rect 12908 10665 13145 10672
rect 13375 10778 13492 10785
rect 13535 10778 13695 10785
rect 13375 10672 13458 10778
rect 13492 10672 13695 10778
rect 13375 10665 13415 10672
rect 13458 10665 13695 10672
rect 13925 10778 14042 10785
rect 14085 10778 14245 10785
rect 13925 10672 14008 10778
rect 14042 10672 14245 10778
rect 13925 10665 13965 10672
rect 14008 10665 14245 10672
rect 14475 10778 14592 10785
rect 14635 10778 14795 10785
rect 14475 10672 14558 10778
rect 14592 10672 14795 10778
rect 14475 10665 14515 10672
rect 14558 10665 14795 10672
rect 15025 10778 15142 10785
rect 15185 10778 15345 10785
rect 15025 10672 15108 10778
rect 15142 10672 15345 10778
rect 15025 10665 15065 10672
rect 15108 10665 15345 10672
rect 15575 10778 15692 10785
rect 15735 10778 15895 10785
rect 15575 10672 15658 10778
rect 15692 10672 15895 10778
rect 15575 10665 15615 10672
rect 15658 10665 15895 10672
rect 16125 10778 16242 10785
rect 16285 10778 16445 10785
rect 16125 10672 16208 10778
rect 16242 10672 16445 10778
rect 16125 10665 16165 10672
rect 16208 10665 16445 10672
rect 16675 10778 16792 10785
rect 16835 10778 16995 10785
rect 16675 10672 16758 10778
rect 16792 10672 16995 10778
rect 16675 10665 16715 10672
rect 16758 10665 16995 10672
rect 17225 10778 17342 10785
rect 17385 10778 17545 10785
rect 17225 10672 17308 10778
rect 17342 10672 17545 10778
rect 17225 10665 17265 10672
rect 17308 10665 17545 10672
rect 17775 10778 17892 10785
rect 17935 10778 18095 10785
rect 17775 10672 17858 10778
rect 17892 10672 18095 10778
rect 17775 10665 17815 10672
rect 17858 10665 18095 10672
rect 18325 10778 18442 10785
rect 18485 10778 18645 10785
rect 18325 10672 18408 10778
rect 18442 10672 18645 10778
rect 18325 10665 18365 10672
rect 18408 10665 18645 10672
rect 18875 10778 18992 10785
rect 19035 10778 19195 10785
rect 18875 10672 18958 10778
rect 18992 10672 19195 10778
rect 18875 10665 18915 10672
rect 18958 10665 19195 10672
rect 765 10625 885 10665
rect 1315 10625 1435 10665
rect 1865 10625 1985 10665
rect 2415 10625 2535 10665
rect 2965 10625 3085 10665
rect 3515 10625 3635 10665
rect 4065 10625 4185 10665
rect 4615 10625 4735 10665
rect 5165 10625 5285 10665
rect 5715 10625 5835 10665
rect 6265 10625 6385 10665
rect 6815 10625 6935 10665
rect 7365 10625 7485 10665
rect 7915 10625 8035 10665
rect 8465 10625 8585 10665
rect 9015 10625 9135 10665
rect 9565 10625 9685 10665
rect 10115 10625 10235 10665
rect 10665 10625 10785 10665
rect 11215 10625 11335 10665
rect 11765 10625 11885 10665
rect 12315 10625 12435 10665
rect 12865 10625 12985 10665
rect 13415 10625 13535 10665
rect 13965 10625 14085 10665
rect 14515 10625 14635 10665
rect 15065 10625 15185 10665
rect 15615 10625 15735 10665
rect 16165 10625 16285 10665
rect 16715 10625 16835 10665
rect 17265 10625 17385 10665
rect 17815 10625 17935 10665
rect 18365 10625 18485 10665
rect 18915 10625 19035 10665
rect 19202 10512 19204 10938
rect 500 10425 507 10475
rect 19202 10396 19217 10402
rect 628 10372 885 10395
rect 1178 10372 1435 10395
rect 1728 10372 1985 10395
rect 2278 10372 2535 10395
rect 2828 10372 3085 10395
rect 3378 10372 3635 10395
rect 3928 10372 4185 10395
rect 4478 10372 4735 10395
rect 5028 10372 5285 10395
rect 5578 10372 5835 10395
rect 6128 10372 6385 10395
rect 6678 10372 6935 10395
rect 7228 10372 7485 10395
rect 7778 10372 8035 10395
rect 8328 10372 8585 10395
rect 8878 10372 9135 10395
rect 9428 10372 9685 10395
rect 9978 10372 10235 10395
rect 10528 10372 10785 10395
rect 11078 10372 11335 10395
rect 11628 10372 11885 10395
rect 12178 10372 12435 10395
rect 12728 10372 12985 10395
rect 13278 10372 13535 10395
rect 13828 10372 14085 10395
rect 14378 10372 14635 10395
rect 14928 10372 15185 10395
rect 15478 10372 15735 10395
rect 16028 10372 16285 10395
rect 16578 10372 16835 10395
rect 17128 10372 17385 10395
rect 17678 10372 17935 10395
rect 18228 10372 18485 10395
rect 18778 10372 19035 10395
rect 605 10235 609 10372
rect 784 10275 885 10372
rect 765 10235 885 10275
rect 1155 10235 1159 10372
rect 1334 10275 1435 10372
rect 1315 10235 1435 10275
rect 1705 10235 1709 10372
rect 1884 10275 1985 10372
rect 1865 10235 1985 10275
rect 2255 10235 2259 10372
rect 2434 10275 2535 10372
rect 2415 10235 2535 10275
rect 2805 10235 2809 10372
rect 2984 10275 3085 10372
rect 2965 10235 3085 10275
rect 3355 10235 3359 10372
rect 3534 10275 3635 10372
rect 3515 10235 3635 10275
rect 3905 10235 3909 10372
rect 4084 10275 4185 10372
rect 4065 10235 4185 10275
rect 4455 10235 4459 10372
rect 4634 10275 4735 10372
rect 4615 10235 4735 10275
rect 5005 10235 5009 10372
rect 5184 10275 5285 10372
rect 5165 10235 5285 10275
rect 5555 10235 5559 10372
rect 5734 10275 5835 10372
rect 5715 10235 5835 10275
rect 6105 10235 6109 10372
rect 6284 10275 6385 10372
rect 6265 10235 6385 10275
rect 6655 10235 6659 10372
rect 6834 10275 6935 10372
rect 6815 10235 6935 10275
rect 7205 10235 7209 10372
rect 7384 10275 7485 10372
rect 7365 10235 7485 10275
rect 7755 10235 7759 10372
rect 7934 10275 8035 10372
rect 7915 10235 8035 10275
rect 8305 10235 8309 10372
rect 8484 10275 8585 10372
rect 8465 10235 8585 10275
rect 8855 10235 8859 10372
rect 9034 10275 9135 10372
rect 9015 10235 9135 10275
rect 9405 10235 9409 10372
rect 9584 10275 9685 10372
rect 9565 10235 9685 10275
rect 9955 10235 9959 10372
rect 10134 10275 10235 10372
rect 10115 10235 10235 10275
rect 10505 10235 10509 10372
rect 10684 10275 10785 10372
rect 10665 10235 10785 10275
rect 11055 10235 11059 10372
rect 11234 10275 11335 10372
rect 11215 10235 11335 10275
rect 11605 10235 11609 10372
rect 11784 10275 11885 10372
rect 11765 10235 11885 10275
rect 12155 10235 12159 10372
rect 12334 10275 12435 10372
rect 12315 10235 12435 10275
rect 12705 10235 12709 10372
rect 12884 10275 12985 10372
rect 12865 10235 12985 10275
rect 13255 10235 13259 10372
rect 13434 10275 13535 10372
rect 13415 10235 13535 10275
rect 13805 10235 13809 10372
rect 13984 10275 14085 10372
rect 13965 10235 14085 10275
rect 14355 10235 14359 10372
rect 14534 10275 14635 10372
rect 14515 10235 14635 10275
rect 14905 10235 14909 10372
rect 15084 10275 15185 10372
rect 15065 10235 15185 10275
rect 15455 10235 15459 10372
rect 15634 10275 15735 10372
rect 15615 10235 15735 10275
rect 16005 10235 16009 10372
rect 16184 10275 16285 10372
rect 16165 10235 16285 10275
rect 16555 10235 16559 10372
rect 16734 10275 16835 10372
rect 16715 10235 16835 10275
rect 17105 10235 17109 10372
rect 17284 10275 17385 10372
rect 17265 10235 17385 10275
rect 17655 10235 17659 10372
rect 17834 10275 17935 10372
rect 17815 10235 17935 10275
rect 18205 10235 18209 10372
rect 18384 10275 18485 10372
rect 18365 10235 18485 10275
rect 18755 10235 18759 10372
rect 18934 10275 19035 10372
rect 18915 10235 19035 10275
rect 725 10228 842 10235
rect 885 10228 1045 10235
rect 725 10122 808 10228
rect 842 10122 1045 10228
rect 725 10115 765 10122
rect 808 10115 1045 10122
rect 1275 10228 1392 10235
rect 1435 10228 1595 10235
rect 1275 10122 1358 10228
rect 1392 10122 1595 10228
rect 1275 10115 1315 10122
rect 1358 10115 1595 10122
rect 1825 10228 1942 10235
rect 1985 10228 2145 10235
rect 1825 10122 1908 10228
rect 1942 10122 2145 10228
rect 1825 10115 1865 10122
rect 1908 10115 2145 10122
rect 2375 10228 2492 10235
rect 2535 10228 2695 10235
rect 2375 10122 2458 10228
rect 2492 10122 2695 10228
rect 2375 10115 2415 10122
rect 2458 10115 2695 10122
rect 2925 10228 3042 10235
rect 3085 10228 3245 10235
rect 2925 10122 3008 10228
rect 3042 10122 3245 10228
rect 2925 10115 2965 10122
rect 3008 10115 3245 10122
rect 3475 10228 3592 10235
rect 3635 10228 3795 10235
rect 3475 10122 3558 10228
rect 3592 10122 3795 10228
rect 3475 10115 3515 10122
rect 3558 10115 3795 10122
rect 4025 10228 4142 10235
rect 4185 10228 4345 10235
rect 4025 10122 4108 10228
rect 4142 10122 4345 10228
rect 4025 10115 4065 10122
rect 4108 10115 4345 10122
rect 4575 10228 4692 10235
rect 4735 10228 4895 10235
rect 4575 10122 4658 10228
rect 4692 10122 4895 10228
rect 4575 10115 4615 10122
rect 4658 10115 4895 10122
rect 5125 10228 5242 10235
rect 5285 10228 5445 10235
rect 5125 10122 5208 10228
rect 5242 10122 5445 10228
rect 5125 10115 5165 10122
rect 5208 10115 5445 10122
rect 5675 10228 5792 10235
rect 5835 10228 5995 10235
rect 5675 10122 5758 10228
rect 5792 10122 5995 10228
rect 5675 10115 5715 10122
rect 5758 10115 5995 10122
rect 6225 10228 6342 10235
rect 6385 10228 6545 10235
rect 6225 10122 6308 10228
rect 6342 10122 6545 10228
rect 6225 10115 6265 10122
rect 6308 10115 6545 10122
rect 6775 10228 6892 10235
rect 6935 10228 7095 10235
rect 6775 10122 6858 10228
rect 6892 10122 7095 10228
rect 6775 10115 6815 10122
rect 6858 10115 7095 10122
rect 7325 10228 7442 10235
rect 7485 10228 7645 10235
rect 7325 10122 7408 10228
rect 7442 10122 7645 10228
rect 7325 10115 7365 10122
rect 7408 10115 7645 10122
rect 7875 10228 7992 10235
rect 8035 10228 8195 10235
rect 7875 10122 7958 10228
rect 7992 10122 8195 10228
rect 7875 10115 7915 10122
rect 7958 10115 8195 10122
rect 8425 10228 8542 10235
rect 8585 10228 8745 10235
rect 8425 10122 8508 10228
rect 8542 10122 8745 10228
rect 8425 10115 8465 10122
rect 8508 10115 8745 10122
rect 8975 10228 9092 10235
rect 9135 10228 9295 10235
rect 8975 10122 9058 10228
rect 9092 10122 9295 10228
rect 8975 10115 9015 10122
rect 9058 10115 9295 10122
rect 9525 10228 9642 10235
rect 9685 10228 9845 10235
rect 9525 10122 9608 10228
rect 9642 10122 9845 10228
rect 9525 10115 9565 10122
rect 9608 10115 9845 10122
rect 10075 10228 10192 10235
rect 10235 10228 10395 10235
rect 10075 10122 10158 10228
rect 10192 10122 10395 10228
rect 10075 10115 10115 10122
rect 10158 10115 10395 10122
rect 10625 10228 10742 10235
rect 10785 10228 10945 10235
rect 10625 10122 10708 10228
rect 10742 10122 10945 10228
rect 10625 10115 10665 10122
rect 10708 10115 10945 10122
rect 11175 10228 11292 10235
rect 11335 10228 11495 10235
rect 11175 10122 11258 10228
rect 11292 10122 11495 10228
rect 11175 10115 11215 10122
rect 11258 10115 11495 10122
rect 11725 10228 11842 10235
rect 11885 10228 12045 10235
rect 11725 10122 11808 10228
rect 11842 10122 12045 10228
rect 11725 10115 11765 10122
rect 11808 10115 12045 10122
rect 12275 10228 12392 10235
rect 12435 10228 12595 10235
rect 12275 10122 12358 10228
rect 12392 10122 12595 10228
rect 12275 10115 12315 10122
rect 12358 10115 12595 10122
rect 12825 10228 12942 10235
rect 12985 10228 13145 10235
rect 12825 10122 12908 10228
rect 12942 10122 13145 10228
rect 12825 10115 12865 10122
rect 12908 10115 13145 10122
rect 13375 10228 13492 10235
rect 13535 10228 13695 10235
rect 13375 10122 13458 10228
rect 13492 10122 13695 10228
rect 13375 10115 13415 10122
rect 13458 10115 13695 10122
rect 13925 10228 14042 10235
rect 14085 10228 14245 10235
rect 13925 10122 14008 10228
rect 14042 10122 14245 10228
rect 13925 10115 13965 10122
rect 14008 10115 14245 10122
rect 14475 10228 14592 10235
rect 14635 10228 14795 10235
rect 14475 10122 14558 10228
rect 14592 10122 14795 10228
rect 14475 10115 14515 10122
rect 14558 10115 14795 10122
rect 15025 10228 15142 10235
rect 15185 10228 15345 10235
rect 15025 10122 15108 10228
rect 15142 10122 15345 10228
rect 15025 10115 15065 10122
rect 15108 10115 15345 10122
rect 15575 10228 15692 10235
rect 15735 10228 15895 10235
rect 15575 10122 15658 10228
rect 15692 10122 15895 10228
rect 15575 10115 15615 10122
rect 15658 10115 15895 10122
rect 16125 10228 16242 10235
rect 16285 10228 16445 10235
rect 16125 10122 16208 10228
rect 16242 10122 16445 10228
rect 16125 10115 16165 10122
rect 16208 10115 16445 10122
rect 16675 10228 16792 10235
rect 16835 10228 16995 10235
rect 16675 10122 16758 10228
rect 16792 10122 16995 10228
rect 16675 10115 16715 10122
rect 16758 10115 16995 10122
rect 17225 10228 17342 10235
rect 17385 10228 17545 10235
rect 17225 10122 17308 10228
rect 17342 10122 17545 10228
rect 17225 10115 17265 10122
rect 17308 10115 17545 10122
rect 17775 10228 17892 10235
rect 17935 10228 18095 10235
rect 17775 10122 17858 10228
rect 17892 10122 18095 10228
rect 17775 10115 17815 10122
rect 17858 10115 18095 10122
rect 18325 10228 18442 10235
rect 18485 10228 18645 10235
rect 18325 10122 18408 10228
rect 18442 10122 18645 10228
rect 18325 10115 18365 10122
rect 18408 10115 18645 10122
rect 18875 10228 18992 10235
rect 19035 10228 19195 10235
rect 18875 10122 18958 10228
rect 18992 10122 19195 10228
rect 18875 10115 18915 10122
rect 18958 10115 19195 10122
rect 765 10075 885 10115
rect 1315 10075 1435 10115
rect 1865 10075 1985 10115
rect 2415 10075 2535 10115
rect 2965 10075 3085 10115
rect 3515 10075 3635 10115
rect 4065 10075 4185 10115
rect 4615 10075 4735 10115
rect 5165 10075 5285 10115
rect 5715 10075 5835 10115
rect 6265 10075 6385 10115
rect 6815 10075 6935 10115
rect 7365 10075 7485 10115
rect 7915 10075 8035 10115
rect 8465 10075 8585 10115
rect 9015 10075 9135 10115
rect 9565 10075 9685 10115
rect 10115 10075 10235 10115
rect 10665 10075 10785 10115
rect 11215 10075 11335 10115
rect 11765 10075 11885 10115
rect 12315 10075 12435 10115
rect 12865 10075 12985 10115
rect 13415 10075 13535 10115
rect 13965 10075 14085 10115
rect 14515 10075 14635 10115
rect 15065 10075 15185 10115
rect 15615 10075 15735 10115
rect 16165 10075 16285 10115
rect 16715 10075 16835 10115
rect 17265 10075 17385 10115
rect 17815 10075 17935 10115
rect 18365 10075 18485 10115
rect 18915 10075 19035 10115
rect 19185 9954 19200 9971
rect 19202 9962 19204 10388
rect 19202 9948 19217 9954
rect 500 9875 507 9925
rect 500 9439 525 9840
rect 628 9822 885 9845
rect 1178 9822 1435 9845
rect 1728 9822 1985 9845
rect 2278 9822 2535 9845
rect 2828 9822 3085 9845
rect 3378 9822 3635 9845
rect 3928 9822 4185 9845
rect 4478 9822 4735 9845
rect 5028 9822 5285 9845
rect 5578 9822 5835 9845
rect 6128 9822 6385 9845
rect 6678 9822 6935 9845
rect 7228 9822 7485 9845
rect 7778 9822 8035 9845
rect 8328 9822 8585 9845
rect 8878 9822 9135 9845
rect 9428 9822 9685 9845
rect 9978 9822 10235 9845
rect 10528 9822 10785 9845
rect 11078 9822 11335 9845
rect 11628 9822 11885 9845
rect 12178 9822 12435 9845
rect 12728 9822 12985 9845
rect 13278 9822 13535 9845
rect 13828 9822 14085 9845
rect 14378 9822 14635 9845
rect 14928 9822 15185 9845
rect 15478 9822 15735 9845
rect 16028 9822 16285 9845
rect 16578 9822 16835 9845
rect 17128 9822 17385 9845
rect 17678 9822 17935 9845
rect 18228 9822 18485 9845
rect 18778 9822 19035 9845
rect 605 9685 609 9822
rect 784 9725 885 9822
rect 765 9685 885 9725
rect 1155 9685 1159 9822
rect 1334 9725 1435 9822
rect 1315 9685 1435 9725
rect 1705 9685 1709 9822
rect 1884 9725 1985 9822
rect 1865 9685 1985 9725
rect 2255 9685 2259 9822
rect 2434 9725 2535 9822
rect 2415 9685 2535 9725
rect 2805 9685 2809 9822
rect 2984 9725 3085 9822
rect 2965 9685 3085 9725
rect 3355 9685 3359 9822
rect 3534 9725 3635 9822
rect 3515 9685 3635 9725
rect 3905 9685 3909 9822
rect 4084 9725 4185 9822
rect 4065 9685 4185 9725
rect 4455 9685 4459 9822
rect 4634 9725 4735 9822
rect 4615 9685 4735 9725
rect 5005 9685 5009 9822
rect 5184 9725 5285 9822
rect 5165 9685 5285 9725
rect 5555 9685 5559 9822
rect 5734 9725 5835 9822
rect 5715 9685 5835 9725
rect 6105 9685 6109 9822
rect 6284 9725 6385 9822
rect 6265 9685 6385 9725
rect 6655 9685 6659 9822
rect 6834 9725 6935 9822
rect 6815 9685 6935 9725
rect 7205 9685 7209 9822
rect 7384 9725 7485 9822
rect 7365 9685 7485 9725
rect 7755 9685 7759 9822
rect 7934 9725 8035 9822
rect 7915 9685 8035 9725
rect 8305 9685 8309 9822
rect 8484 9725 8585 9822
rect 8465 9685 8585 9725
rect 8855 9685 8859 9822
rect 9034 9725 9135 9822
rect 9015 9685 9135 9725
rect 9405 9685 9409 9822
rect 9584 9725 9685 9822
rect 9565 9685 9685 9725
rect 9955 9685 9959 9822
rect 10134 9725 10235 9822
rect 10115 9685 10235 9725
rect 10505 9685 10509 9822
rect 10684 9725 10785 9822
rect 10665 9685 10785 9725
rect 11055 9685 11059 9822
rect 11234 9725 11335 9822
rect 11215 9685 11335 9725
rect 11605 9685 11609 9822
rect 11784 9725 11885 9822
rect 11765 9685 11885 9725
rect 12155 9685 12159 9822
rect 12334 9725 12435 9822
rect 12315 9685 12435 9725
rect 12705 9685 12709 9822
rect 12884 9725 12985 9822
rect 12865 9685 12985 9725
rect 13255 9685 13259 9822
rect 13434 9725 13535 9822
rect 13415 9685 13535 9725
rect 13805 9685 13809 9822
rect 13984 9725 14085 9822
rect 13965 9685 14085 9725
rect 14355 9685 14359 9822
rect 14534 9725 14635 9822
rect 14515 9685 14635 9725
rect 14905 9685 14909 9822
rect 15084 9725 15185 9822
rect 15065 9685 15185 9725
rect 15455 9685 15459 9822
rect 15634 9725 15735 9822
rect 15615 9685 15735 9725
rect 16005 9685 16009 9822
rect 16184 9725 16285 9822
rect 16165 9685 16285 9725
rect 16555 9685 16559 9822
rect 16734 9725 16835 9822
rect 16715 9685 16835 9725
rect 17105 9685 17109 9822
rect 17284 9725 17385 9822
rect 17265 9685 17385 9725
rect 17655 9685 17659 9822
rect 17834 9725 17935 9822
rect 17815 9685 17935 9725
rect 18205 9685 18209 9822
rect 18384 9725 18485 9822
rect 18365 9685 18485 9725
rect 18755 9685 18759 9822
rect 18934 9725 19035 9822
rect 18915 9685 19035 9725
rect 725 9678 842 9685
rect 885 9678 1045 9685
rect 725 9572 808 9678
rect 842 9572 1045 9678
rect 725 9565 765 9572
rect 808 9565 1045 9572
rect 1275 9678 1392 9685
rect 1435 9678 1595 9685
rect 1275 9572 1358 9678
rect 1392 9572 1595 9678
rect 1275 9565 1315 9572
rect 1358 9565 1595 9572
rect 1825 9678 1942 9685
rect 1985 9678 2145 9685
rect 1825 9572 1908 9678
rect 1942 9572 2145 9678
rect 1825 9565 1865 9572
rect 1908 9565 2145 9572
rect 2375 9678 2492 9685
rect 2535 9678 2695 9685
rect 2375 9572 2458 9678
rect 2492 9572 2695 9678
rect 2375 9565 2415 9572
rect 2458 9565 2695 9572
rect 2925 9678 3042 9685
rect 3085 9678 3245 9685
rect 2925 9572 3008 9678
rect 3042 9572 3245 9678
rect 2925 9565 2965 9572
rect 3008 9565 3245 9572
rect 3475 9678 3592 9685
rect 3635 9678 3795 9685
rect 3475 9572 3558 9678
rect 3592 9572 3795 9678
rect 3475 9565 3515 9572
rect 3558 9565 3795 9572
rect 4025 9678 4142 9685
rect 4185 9678 4345 9685
rect 4025 9572 4108 9678
rect 4142 9572 4345 9678
rect 4025 9565 4065 9572
rect 4108 9565 4345 9572
rect 4575 9678 4692 9685
rect 4735 9678 4895 9685
rect 4575 9572 4658 9678
rect 4692 9572 4895 9678
rect 4575 9565 4615 9572
rect 4658 9565 4895 9572
rect 5125 9678 5242 9685
rect 5285 9678 5445 9685
rect 5125 9572 5208 9678
rect 5242 9572 5445 9678
rect 5125 9565 5165 9572
rect 5208 9565 5445 9572
rect 5675 9678 5792 9685
rect 5835 9678 5995 9685
rect 5675 9572 5758 9678
rect 5792 9572 5995 9678
rect 5675 9565 5715 9572
rect 5758 9565 5995 9572
rect 6225 9678 6342 9685
rect 6385 9678 6545 9685
rect 6225 9572 6308 9678
rect 6342 9572 6545 9678
rect 6225 9565 6265 9572
rect 6308 9565 6545 9572
rect 6775 9678 6892 9685
rect 6935 9678 7095 9685
rect 6775 9572 6858 9678
rect 6892 9572 7095 9678
rect 6775 9565 6815 9572
rect 6858 9565 7095 9572
rect 7325 9678 7442 9685
rect 7485 9678 7645 9685
rect 7325 9572 7408 9678
rect 7442 9572 7645 9678
rect 7325 9565 7365 9572
rect 7408 9565 7645 9572
rect 7875 9678 7992 9685
rect 8035 9678 8195 9685
rect 7875 9572 7958 9678
rect 7992 9572 8195 9678
rect 7875 9565 7915 9572
rect 7958 9565 8195 9572
rect 8425 9678 8542 9685
rect 8585 9678 8745 9685
rect 8425 9572 8508 9678
rect 8542 9572 8745 9678
rect 8425 9565 8465 9572
rect 8508 9565 8745 9572
rect 8975 9678 9092 9685
rect 9135 9678 9295 9685
rect 8975 9572 9058 9678
rect 9092 9572 9295 9678
rect 8975 9565 9015 9572
rect 9058 9565 9295 9572
rect 9525 9678 9642 9685
rect 9685 9678 9845 9685
rect 9525 9572 9608 9678
rect 9642 9572 9845 9678
rect 9525 9565 9565 9572
rect 9608 9565 9845 9572
rect 10075 9678 10192 9685
rect 10235 9678 10395 9685
rect 10075 9572 10158 9678
rect 10192 9572 10395 9678
rect 10075 9565 10115 9572
rect 10158 9565 10395 9572
rect 10625 9678 10742 9685
rect 10785 9678 10945 9685
rect 10625 9572 10708 9678
rect 10742 9572 10945 9678
rect 10625 9565 10665 9572
rect 10708 9565 10945 9572
rect 11175 9678 11292 9685
rect 11335 9678 11495 9685
rect 11175 9572 11258 9678
rect 11292 9572 11495 9678
rect 11175 9565 11215 9572
rect 11258 9565 11495 9572
rect 11725 9678 11842 9685
rect 11885 9678 12045 9685
rect 11725 9572 11808 9678
rect 11842 9572 12045 9678
rect 11725 9565 11765 9572
rect 11808 9565 12045 9572
rect 12275 9678 12392 9685
rect 12435 9678 12595 9685
rect 12275 9572 12358 9678
rect 12392 9572 12595 9678
rect 12275 9565 12315 9572
rect 12358 9565 12595 9572
rect 12825 9678 12942 9685
rect 12985 9678 13145 9685
rect 12825 9572 12908 9678
rect 12942 9572 13145 9678
rect 12825 9565 12865 9572
rect 12908 9565 13145 9572
rect 13375 9678 13492 9685
rect 13535 9678 13695 9685
rect 13375 9572 13458 9678
rect 13492 9572 13695 9678
rect 13375 9565 13415 9572
rect 13458 9565 13695 9572
rect 13925 9678 14042 9685
rect 14085 9678 14245 9685
rect 13925 9572 14008 9678
rect 14042 9572 14245 9678
rect 13925 9565 13965 9572
rect 14008 9565 14245 9572
rect 14475 9678 14592 9685
rect 14635 9678 14795 9685
rect 14475 9572 14558 9678
rect 14592 9572 14795 9678
rect 14475 9565 14515 9572
rect 14558 9565 14795 9572
rect 15025 9678 15142 9685
rect 15185 9678 15345 9685
rect 15025 9572 15108 9678
rect 15142 9572 15345 9678
rect 15025 9565 15065 9572
rect 15108 9565 15345 9572
rect 15575 9678 15692 9685
rect 15735 9678 15895 9685
rect 15575 9572 15658 9678
rect 15692 9572 15895 9678
rect 15575 9565 15615 9572
rect 15658 9565 15895 9572
rect 16125 9678 16242 9685
rect 16285 9678 16445 9685
rect 16125 9572 16208 9678
rect 16242 9572 16445 9678
rect 16125 9565 16165 9572
rect 16208 9565 16445 9572
rect 16675 9678 16792 9685
rect 16835 9678 16995 9685
rect 16675 9572 16758 9678
rect 16792 9572 16995 9678
rect 16675 9565 16715 9572
rect 16758 9565 16995 9572
rect 17225 9678 17342 9685
rect 17385 9678 17545 9685
rect 17225 9572 17308 9678
rect 17342 9572 17545 9678
rect 17225 9565 17265 9572
rect 17308 9565 17545 9572
rect 17775 9678 17892 9685
rect 17935 9678 18095 9685
rect 17775 9572 17858 9678
rect 17892 9572 18095 9678
rect 17775 9565 17815 9572
rect 17858 9565 18095 9572
rect 18325 9678 18442 9685
rect 18485 9678 18645 9685
rect 18325 9572 18408 9678
rect 18442 9572 18645 9678
rect 18325 9565 18365 9572
rect 18408 9565 18645 9572
rect 18875 9678 18992 9685
rect 19035 9678 19195 9685
rect 18875 9572 18958 9678
rect 18992 9572 19195 9678
rect 18875 9565 18915 9572
rect 18958 9565 19195 9572
rect 765 9525 885 9565
rect 1315 9525 1435 9565
rect 1865 9525 1985 9565
rect 2415 9525 2535 9565
rect 2965 9525 3085 9565
rect 3515 9525 3635 9565
rect 4065 9525 4185 9565
rect 4615 9525 4735 9565
rect 5165 9525 5285 9565
rect 5715 9525 5835 9565
rect 6265 9525 6385 9565
rect 6815 9525 6935 9565
rect 7365 9525 7485 9565
rect 7915 9525 8035 9565
rect 8465 9525 8585 9565
rect 9015 9525 9135 9565
rect 9565 9525 9685 9565
rect 10115 9525 10235 9565
rect 10665 9525 10785 9565
rect 11215 9525 11335 9565
rect 11765 9525 11885 9565
rect 12315 9525 12435 9565
rect 12865 9525 12985 9565
rect 13415 9525 13535 9565
rect 13965 9525 14085 9565
rect 14515 9525 14635 9565
rect 15065 9525 15185 9565
rect 15615 9525 15735 9565
rect 16165 9525 16285 9565
rect 16715 9525 16835 9565
rect 17265 9525 17385 9565
rect 17815 9525 17935 9565
rect 18365 9525 18485 9565
rect 18915 9525 19035 9565
rect 19202 9412 19204 9838
rect 500 9325 507 9375
rect 19202 9296 19217 9302
rect 628 9272 885 9295
rect 1178 9272 1435 9295
rect 1728 9272 1985 9295
rect 2278 9272 2535 9295
rect 2828 9272 3085 9295
rect 3378 9272 3635 9295
rect 3928 9272 4185 9295
rect 4478 9272 4735 9295
rect 5028 9272 5285 9295
rect 5578 9272 5835 9295
rect 6128 9272 6385 9295
rect 6678 9272 6935 9295
rect 7228 9272 7485 9295
rect 7778 9272 8035 9295
rect 8328 9272 8585 9295
rect 8878 9272 9135 9295
rect 9428 9272 9685 9295
rect 9978 9272 10235 9295
rect 10528 9272 10785 9295
rect 11078 9272 11335 9295
rect 11628 9272 11885 9295
rect 12178 9272 12435 9295
rect 12728 9272 12985 9295
rect 13278 9272 13535 9295
rect 13828 9272 14085 9295
rect 14378 9272 14635 9295
rect 14928 9272 15185 9295
rect 15478 9272 15735 9295
rect 16028 9272 16285 9295
rect 16578 9272 16835 9295
rect 17128 9272 17385 9295
rect 17678 9272 17935 9295
rect 18228 9272 18485 9295
rect 18778 9272 19035 9295
rect 605 9135 609 9272
rect 784 9175 885 9272
rect 765 9135 885 9175
rect 1155 9135 1159 9272
rect 1334 9175 1435 9272
rect 1315 9135 1435 9175
rect 1705 9135 1709 9272
rect 1884 9175 1985 9272
rect 1865 9135 1985 9175
rect 2255 9135 2259 9272
rect 2434 9175 2535 9272
rect 2415 9135 2535 9175
rect 2805 9135 2809 9272
rect 2984 9175 3085 9272
rect 2965 9135 3085 9175
rect 3355 9135 3359 9272
rect 3534 9175 3635 9272
rect 3515 9135 3635 9175
rect 3905 9135 3909 9272
rect 4084 9175 4185 9272
rect 4065 9135 4185 9175
rect 4455 9135 4459 9272
rect 4634 9175 4735 9272
rect 4615 9135 4735 9175
rect 5005 9135 5009 9272
rect 5184 9175 5285 9272
rect 5165 9135 5285 9175
rect 5555 9135 5559 9272
rect 5734 9175 5835 9272
rect 5715 9135 5835 9175
rect 6105 9135 6109 9272
rect 6284 9175 6385 9272
rect 6265 9135 6385 9175
rect 6655 9135 6659 9272
rect 6834 9175 6935 9272
rect 6815 9135 6935 9175
rect 7205 9135 7209 9272
rect 7384 9175 7485 9272
rect 7365 9135 7485 9175
rect 7755 9135 7759 9272
rect 7934 9175 8035 9272
rect 7915 9135 8035 9175
rect 8305 9135 8309 9272
rect 8484 9175 8585 9272
rect 8465 9135 8585 9175
rect 8855 9135 8859 9272
rect 9034 9175 9135 9272
rect 9015 9135 9135 9175
rect 9405 9135 9409 9272
rect 9584 9175 9685 9272
rect 9565 9135 9685 9175
rect 9955 9135 9959 9272
rect 10134 9175 10235 9272
rect 10115 9135 10235 9175
rect 10505 9135 10509 9272
rect 10684 9175 10785 9272
rect 10665 9135 10785 9175
rect 11055 9135 11059 9272
rect 11234 9175 11335 9272
rect 11215 9135 11335 9175
rect 11605 9135 11609 9272
rect 11784 9175 11885 9272
rect 11765 9135 11885 9175
rect 12155 9135 12159 9272
rect 12334 9175 12435 9272
rect 12315 9135 12435 9175
rect 12705 9135 12709 9272
rect 12884 9175 12985 9272
rect 12865 9135 12985 9175
rect 13255 9135 13259 9272
rect 13434 9175 13535 9272
rect 13415 9135 13535 9175
rect 13805 9135 13809 9272
rect 13984 9175 14085 9272
rect 13965 9135 14085 9175
rect 14355 9135 14359 9272
rect 14534 9175 14635 9272
rect 14515 9135 14635 9175
rect 14905 9135 14909 9272
rect 15084 9175 15185 9272
rect 15065 9135 15185 9175
rect 15455 9135 15459 9272
rect 15634 9175 15735 9272
rect 15615 9135 15735 9175
rect 16005 9135 16009 9272
rect 16184 9175 16285 9272
rect 16165 9135 16285 9175
rect 16555 9135 16559 9272
rect 16734 9175 16835 9272
rect 16715 9135 16835 9175
rect 17105 9135 17109 9272
rect 17284 9175 17385 9272
rect 17265 9135 17385 9175
rect 17655 9135 17659 9272
rect 17834 9175 17935 9272
rect 17815 9135 17935 9175
rect 18205 9135 18209 9272
rect 18384 9175 18485 9272
rect 18365 9135 18485 9175
rect 18755 9135 18759 9272
rect 18934 9175 19035 9272
rect 18915 9135 19035 9175
rect 725 9128 842 9135
rect 885 9128 1045 9135
rect 725 9022 808 9128
rect 842 9022 1045 9128
rect 725 9015 765 9022
rect 808 9015 1045 9022
rect 1275 9128 1392 9135
rect 1435 9128 1595 9135
rect 1275 9022 1358 9128
rect 1392 9022 1595 9128
rect 1275 9015 1315 9022
rect 1358 9015 1595 9022
rect 1825 9128 1942 9135
rect 1985 9128 2145 9135
rect 1825 9022 1908 9128
rect 1942 9022 2145 9128
rect 1825 9015 1865 9022
rect 1908 9015 2145 9022
rect 2375 9128 2492 9135
rect 2535 9128 2695 9135
rect 2375 9022 2458 9128
rect 2492 9022 2695 9128
rect 2375 9015 2415 9022
rect 2458 9015 2695 9022
rect 2925 9128 3042 9135
rect 3085 9128 3245 9135
rect 2925 9022 3008 9128
rect 3042 9022 3245 9128
rect 2925 9015 2965 9022
rect 3008 9015 3245 9022
rect 3475 9128 3592 9135
rect 3635 9128 3795 9135
rect 3475 9022 3558 9128
rect 3592 9022 3795 9128
rect 3475 9015 3515 9022
rect 3558 9015 3795 9022
rect 4025 9128 4142 9135
rect 4185 9128 4345 9135
rect 4025 9022 4108 9128
rect 4142 9022 4345 9128
rect 4025 9015 4065 9022
rect 4108 9015 4345 9022
rect 4575 9128 4692 9135
rect 4735 9128 4895 9135
rect 4575 9022 4658 9128
rect 4692 9022 4895 9128
rect 4575 9015 4615 9022
rect 4658 9015 4895 9022
rect 5125 9128 5242 9135
rect 5285 9128 5445 9135
rect 5125 9022 5208 9128
rect 5242 9022 5445 9128
rect 5125 9015 5165 9022
rect 5208 9015 5445 9022
rect 5675 9128 5792 9135
rect 5835 9128 5995 9135
rect 5675 9022 5758 9128
rect 5792 9022 5995 9128
rect 5675 9015 5715 9022
rect 5758 9015 5995 9022
rect 6225 9128 6342 9135
rect 6385 9128 6545 9135
rect 6225 9022 6308 9128
rect 6342 9022 6545 9128
rect 6225 9015 6265 9022
rect 6308 9015 6545 9022
rect 6775 9128 6892 9135
rect 6935 9128 7095 9135
rect 6775 9022 6858 9128
rect 6892 9022 7095 9128
rect 6775 9015 6815 9022
rect 6858 9015 7095 9022
rect 7325 9128 7442 9135
rect 7485 9128 7645 9135
rect 7325 9022 7408 9128
rect 7442 9022 7645 9128
rect 7325 9015 7365 9022
rect 7408 9015 7645 9022
rect 7875 9128 7992 9135
rect 8035 9128 8195 9135
rect 7875 9022 7958 9128
rect 7992 9022 8195 9128
rect 7875 9015 7915 9022
rect 7958 9015 8195 9022
rect 8425 9128 8542 9135
rect 8585 9128 8745 9135
rect 8425 9022 8508 9128
rect 8542 9022 8745 9128
rect 8425 9015 8465 9022
rect 8508 9015 8745 9022
rect 8975 9128 9092 9135
rect 9135 9128 9295 9135
rect 8975 9022 9058 9128
rect 9092 9022 9295 9128
rect 8975 9015 9015 9022
rect 9058 9015 9295 9022
rect 9525 9128 9642 9135
rect 9685 9128 9845 9135
rect 9525 9022 9608 9128
rect 9642 9022 9845 9128
rect 9525 9015 9565 9022
rect 9608 9015 9845 9022
rect 10075 9128 10192 9135
rect 10235 9128 10395 9135
rect 10075 9022 10158 9128
rect 10192 9022 10395 9128
rect 10075 9015 10115 9022
rect 10158 9015 10395 9022
rect 10625 9128 10742 9135
rect 10785 9128 10945 9135
rect 10625 9022 10708 9128
rect 10742 9022 10945 9128
rect 10625 9015 10665 9022
rect 10708 9015 10945 9022
rect 11175 9128 11292 9135
rect 11335 9128 11495 9135
rect 11175 9022 11258 9128
rect 11292 9022 11495 9128
rect 11175 9015 11215 9022
rect 11258 9015 11495 9022
rect 11725 9128 11842 9135
rect 11885 9128 12045 9135
rect 11725 9022 11808 9128
rect 11842 9022 12045 9128
rect 11725 9015 11765 9022
rect 11808 9015 12045 9022
rect 12275 9128 12392 9135
rect 12435 9128 12595 9135
rect 12275 9022 12358 9128
rect 12392 9022 12595 9128
rect 12275 9015 12315 9022
rect 12358 9015 12595 9022
rect 12825 9128 12942 9135
rect 12985 9128 13145 9135
rect 12825 9022 12908 9128
rect 12942 9022 13145 9128
rect 12825 9015 12865 9022
rect 12908 9015 13145 9022
rect 13375 9128 13492 9135
rect 13535 9128 13695 9135
rect 13375 9022 13458 9128
rect 13492 9022 13695 9128
rect 13375 9015 13415 9022
rect 13458 9015 13695 9022
rect 13925 9128 14042 9135
rect 14085 9128 14245 9135
rect 13925 9022 14008 9128
rect 14042 9022 14245 9128
rect 13925 9015 13965 9022
rect 14008 9015 14245 9022
rect 14475 9128 14592 9135
rect 14635 9128 14795 9135
rect 14475 9022 14558 9128
rect 14592 9022 14795 9128
rect 14475 9015 14515 9022
rect 14558 9015 14795 9022
rect 15025 9128 15142 9135
rect 15185 9128 15345 9135
rect 15025 9022 15108 9128
rect 15142 9022 15345 9128
rect 15025 9015 15065 9022
rect 15108 9015 15345 9022
rect 15575 9128 15692 9135
rect 15735 9128 15895 9135
rect 15575 9022 15658 9128
rect 15692 9022 15895 9128
rect 15575 9015 15615 9022
rect 15658 9015 15895 9022
rect 16125 9128 16242 9135
rect 16285 9128 16445 9135
rect 16125 9022 16208 9128
rect 16242 9022 16445 9128
rect 16125 9015 16165 9022
rect 16208 9015 16445 9022
rect 16675 9128 16792 9135
rect 16835 9128 16995 9135
rect 16675 9022 16758 9128
rect 16792 9022 16995 9128
rect 16675 9015 16715 9022
rect 16758 9015 16995 9022
rect 17225 9128 17342 9135
rect 17385 9128 17545 9135
rect 17225 9022 17308 9128
rect 17342 9022 17545 9128
rect 17225 9015 17265 9022
rect 17308 9015 17545 9022
rect 17775 9128 17892 9135
rect 17935 9128 18095 9135
rect 17775 9022 17858 9128
rect 17892 9022 18095 9128
rect 17775 9015 17815 9022
rect 17858 9015 18095 9022
rect 18325 9128 18442 9135
rect 18485 9128 18645 9135
rect 18325 9022 18408 9128
rect 18442 9022 18645 9128
rect 18325 9015 18365 9022
rect 18408 9015 18645 9022
rect 18875 9128 18992 9135
rect 19035 9128 19195 9135
rect 18875 9022 18958 9128
rect 18992 9022 19195 9128
rect 18875 9015 18915 9022
rect 18958 9015 19195 9022
rect 765 8975 885 9015
rect 1315 8975 1435 9015
rect 1865 8975 1985 9015
rect 2415 8975 2535 9015
rect 2965 8975 3085 9015
rect 3515 8975 3635 9015
rect 4065 8975 4185 9015
rect 4615 8975 4735 9015
rect 5165 8975 5285 9015
rect 5715 8975 5835 9015
rect 6265 8975 6385 9015
rect 6815 8975 6935 9015
rect 7365 8975 7485 9015
rect 7915 8975 8035 9015
rect 8465 8975 8585 9015
rect 9015 8975 9135 9015
rect 9565 8975 9685 9015
rect 10115 8975 10235 9015
rect 10665 8975 10785 9015
rect 11215 8975 11335 9015
rect 11765 8975 11885 9015
rect 12315 8975 12435 9015
rect 12865 8975 12985 9015
rect 13415 8975 13535 9015
rect 13965 8975 14085 9015
rect 14515 8975 14635 9015
rect 15065 8975 15185 9015
rect 15615 8975 15735 9015
rect 16165 8975 16285 9015
rect 16715 8975 16835 9015
rect 17265 8975 17385 9015
rect 17815 8975 17935 9015
rect 18365 8975 18485 9015
rect 18915 8975 19035 9015
rect 19185 8854 19200 8871
rect 19202 8862 19204 9288
rect 19202 8848 19217 8854
rect 500 8775 507 8825
rect 500 8339 525 8740
rect 628 8722 885 8745
rect 1178 8722 1435 8745
rect 1728 8722 1985 8745
rect 2278 8722 2535 8745
rect 2828 8722 3085 8745
rect 3378 8722 3635 8745
rect 3928 8722 4185 8745
rect 4478 8722 4735 8745
rect 5028 8722 5285 8745
rect 5578 8722 5835 8745
rect 6128 8722 6385 8745
rect 6678 8722 6935 8745
rect 7228 8722 7485 8745
rect 7778 8722 8035 8745
rect 8328 8722 8585 8745
rect 8878 8722 9135 8745
rect 9428 8722 9685 8745
rect 9978 8722 10235 8745
rect 10528 8722 10785 8745
rect 11078 8722 11335 8745
rect 11628 8722 11885 8745
rect 12178 8722 12435 8745
rect 12728 8722 12985 8745
rect 13278 8722 13535 8745
rect 13828 8722 14085 8745
rect 14378 8722 14635 8745
rect 14928 8722 15185 8745
rect 15478 8722 15735 8745
rect 16028 8722 16285 8745
rect 16578 8722 16835 8745
rect 17128 8722 17385 8745
rect 17678 8722 17935 8745
rect 18228 8722 18485 8745
rect 18778 8722 19035 8745
rect 605 8585 609 8722
rect 784 8625 885 8722
rect 765 8585 885 8625
rect 1155 8585 1159 8722
rect 1334 8625 1435 8722
rect 1315 8585 1435 8625
rect 1705 8585 1709 8722
rect 1884 8625 1985 8722
rect 1865 8585 1985 8625
rect 2255 8585 2259 8722
rect 2434 8625 2535 8722
rect 2415 8585 2535 8625
rect 2805 8585 2809 8722
rect 2984 8625 3085 8722
rect 2965 8585 3085 8625
rect 3355 8585 3359 8722
rect 3534 8625 3635 8722
rect 3515 8585 3635 8625
rect 3905 8585 3909 8722
rect 4084 8625 4185 8722
rect 4065 8585 4185 8625
rect 4455 8585 4459 8722
rect 4634 8625 4735 8722
rect 4615 8585 4735 8625
rect 5005 8585 5009 8722
rect 5184 8625 5285 8722
rect 5165 8585 5285 8625
rect 5555 8585 5559 8722
rect 5734 8625 5835 8722
rect 5715 8585 5835 8625
rect 6105 8585 6109 8722
rect 6284 8625 6385 8722
rect 6265 8585 6385 8625
rect 6655 8585 6659 8722
rect 6834 8625 6935 8722
rect 6815 8585 6935 8625
rect 7205 8585 7209 8722
rect 7384 8625 7485 8722
rect 7365 8585 7485 8625
rect 7755 8585 7759 8722
rect 7934 8625 8035 8722
rect 7915 8585 8035 8625
rect 8305 8585 8309 8722
rect 8484 8625 8585 8722
rect 8465 8585 8585 8625
rect 8855 8585 8859 8722
rect 9034 8625 9135 8722
rect 9015 8585 9135 8625
rect 9405 8585 9409 8722
rect 9584 8625 9685 8722
rect 9565 8585 9685 8625
rect 9955 8585 9959 8722
rect 10134 8625 10235 8722
rect 10115 8585 10235 8625
rect 10505 8585 10509 8722
rect 10684 8625 10785 8722
rect 10665 8585 10785 8625
rect 11055 8585 11059 8722
rect 11234 8625 11335 8722
rect 11215 8585 11335 8625
rect 11605 8585 11609 8722
rect 11784 8625 11885 8722
rect 11765 8585 11885 8625
rect 12155 8585 12159 8722
rect 12334 8625 12435 8722
rect 12315 8585 12435 8625
rect 12705 8585 12709 8722
rect 12884 8625 12985 8722
rect 12865 8585 12985 8625
rect 13255 8585 13259 8722
rect 13434 8625 13535 8722
rect 13415 8585 13535 8625
rect 13805 8585 13809 8722
rect 13984 8625 14085 8722
rect 13965 8585 14085 8625
rect 14355 8585 14359 8722
rect 14534 8625 14635 8722
rect 14515 8585 14635 8625
rect 14905 8585 14909 8722
rect 15084 8625 15185 8722
rect 15065 8585 15185 8625
rect 15455 8585 15459 8722
rect 15634 8625 15735 8722
rect 15615 8585 15735 8625
rect 16005 8585 16009 8722
rect 16184 8625 16285 8722
rect 16165 8585 16285 8625
rect 16555 8585 16559 8722
rect 16734 8625 16835 8722
rect 16715 8585 16835 8625
rect 17105 8585 17109 8722
rect 17284 8625 17385 8722
rect 17265 8585 17385 8625
rect 17655 8585 17659 8722
rect 17834 8625 17935 8722
rect 17815 8585 17935 8625
rect 18205 8585 18209 8722
rect 18384 8625 18485 8722
rect 18365 8585 18485 8625
rect 18755 8585 18759 8722
rect 18934 8625 19035 8722
rect 18915 8585 19035 8625
rect 725 8578 842 8585
rect 885 8578 1045 8585
rect 725 8472 808 8578
rect 842 8472 1045 8578
rect 725 8465 765 8472
rect 808 8465 1045 8472
rect 1275 8578 1392 8585
rect 1435 8578 1595 8585
rect 1275 8472 1358 8578
rect 1392 8472 1595 8578
rect 1275 8465 1315 8472
rect 1358 8465 1595 8472
rect 1825 8578 1942 8585
rect 1985 8578 2145 8585
rect 1825 8472 1908 8578
rect 1942 8472 2145 8578
rect 1825 8465 1865 8472
rect 1908 8465 2145 8472
rect 2375 8578 2492 8585
rect 2535 8578 2695 8585
rect 2375 8472 2458 8578
rect 2492 8472 2695 8578
rect 2375 8465 2415 8472
rect 2458 8465 2695 8472
rect 2925 8578 3042 8585
rect 3085 8578 3245 8585
rect 2925 8472 3008 8578
rect 3042 8472 3245 8578
rect 2925 8465 2965 8472
rect 3008 8465 3245 8472
rect 3475 8578 3592 8585
rect 3635 8578 3795 8585
rect 3475 8472 3558 8578
rect 3592 8472 3795 8578
rect 3475 8465 3515 8472
rect 3558 8465 3795 8472
rect 4025 8578 4142 8585
rect 4185 8578 4345 8585
rect 4025 8472 4108 8578
rect 4142 8472 4345 8578
rect 4025 8465 4065 8472
rect 4108 8465 4345 8472
rect 4575 8578 4692 8585
rect 4735 8578 4895 8585
rect 4575 8472 4658 8578
rect 4692 8472 4895 8578
rect 4575 8465 4615 8472
rect 4658 8465 4895 8472
rect 5125 8578 5242 8585
rect 5285 8578 5445 8585
rect 5125 8472 5208 8578
rect 5242 8472 5445 8578
rect 5125 8465 5165 8472
rect 5208 8465 5445 8472
rect 5675 8578 5792 8585
rect 5835 8578 5995 8585
rect 5675 8472 5758 8578
rect 5792 8472 5995 8578
rect 5675 8465 5715 8472
rect 5758 8465 5995 8472
rect 6225 8578 6342 8585
rect 6385 8578 6545 8585
rect 6225 8472 6308 8578
rect 6342 8472 6545 8578
rect 6225 8465 6265 8472
rect 6308 8465 6545 8472
rect 6775 8578 6892 8585
rect 6935 8578 7095 8585
rect 6775 8472 6858 8578
rect 6892 8472 7095 8578
rect 6775 8465 6815 8472
rect 6858 8465 7095 8472
rect 7325 8578 7442 8585
rect 7485 8578 7645 8585
rect 7325 8472 7408 8578
rect 7442 8472 7645 8578
rect 7325 8465 7365 8472
rect 7408 8465 7645 8472
rect 7875 8578 7992 8585
rect 8035 8578 8195 8585
rect 7875 8472 7958 8578
rect 7992 8472 8195 8578
rect 7875 8465 7915 8472
rect 7958 8465 8195 8472
rect 8425 8578 8542 8585
rect 8585 8578 8745 8585
rect 8425 8472 8508 8578
rect 8542 8472 8745 8578
rect 8425 8465 8465 8472
rect 8508 8465 8745 8472
rect 8975 8578 9092 8585
rect 9135 8578 9295 8585
rect 8975 8472 9058 8578
rect 9092 8472 9295 8578
rect 8975 8465 9015 8472
rect 9058 8465 9295 8472
rect 9525 8578 9642 8585
rect 9685 8578 9845 8585
rect 9525 8472 9608 8578
rect 9642 8472 9845 8578
rect 9525 8465 9565 8472
rect 9608 8465 9845 8472
rect 10075 8578 10192 8585
rect 10235 8578 10395 8585
rect 10075 8472 10158 8578
rect 10192 8472 10395 8578
rect 10075 8465 10115 8472
rect 10158 8465 10395 8472
rect 10625 8578 10742 8585
rect 10785 8578 10945 8585
rect 10625 8472 10708 8578
rect 10742 8472 10945 8578
rect 10625 8465 10665 8472
rect 10708 8465 10945 8472
rect 11175 8578 11292 8585
rect 11335 8578 11495 8585
rect 11175 8472 11258 8578
rect 11292 8472 11495 8578
rect 11175 8465 11215 8472
rect 11258 8465 11495 8472
rect 11725 8578 11842 8585
rect 11885 8578 12045 8585
rect 11725 8472 11808 8578
rect 11842 8472 12045 8578
rect 11725 8465 11765 8472
rect 11808 8465 12045 8472
rect 12275 8578 12392 8585
rect 12435 8578 12595 8585
rect 12275 8472 12358 8578
rect 12392 8472 12595 8578
rect 12275 8465 12315 8472
rect 12358 8465 12595 8472
rect 12825 8578 12942 8585
rect 12985 8578 13145 8585
rect 12825 8472 12908 8578
rect 12942 8472 13145 8578
rect 12825 8465 12865 8472
rect 12908 8465 13145 8472
rect 13375 8578 13492 8585
rect 13535 8578 13695 8585
rect 13375 8472 13458 8578
rect 13492 8472 13695 8578
rect 13375 8465 13415 8472
rect 13458 8465 13695 8472
rect 13925 8578 14042 8585
rect 14085 8578 14245 8585
rect 13925 8472 14008 8578
rect 14042 8472 14245 8578
rect 13925 8465 13965 8472
rect 14008 8465 14245 8472
rect 14475 8578 14592 8585
rect 14635 8578 14795 8585
rect 14475 8472 14558 8578
rect 14592 8472 14795 8578
rect 14475 8465 14515 8472
rect 14558 8465 14795 8472
rect 15025 8578 15142 8585
rect 15185 8578 15345 8585
rect 15025 8472 15108 8578
rect 15142 8472 15345 8578
rect 15025 8465 15065 8472
rect 15108 8465 15345 8472
rect 15575 8578 15692 8585
rect 15735 8578 15895 8585
rect 15575 8472 15658 8578
rect 15692 8472 15895 8578
rect 15575 8465 15615 8472
rect 15658 8465 15895 8472
rect 16125 8578 16242 8585
rect 16285 8578 16445 8585
rect 16125 8472 16208 8578
rect 16242 8472 16445 8578
rect 16125 8465 16165 8472
rect 16208 8465 16445 8472
rect 16675 8578 16792 8585
rect 16835 8578 16995 8585
rect 16675 8472 16758 8578
rect 16792 8472 16995 8578
rect 16675 8465 16715 8472
rect 16758 8465 16995 8472
rect 17225 8578 17342 8585
rect 17385 8578 17545 8585
rect 17225 8472 17308 8578
rect 17342 8472 17545 8578
rect 17225 8465 17265 8472
rect 17308 8465 17545 8472
rect 17775 8578 17892 8585
rect 17935 8578 18095 8585
rect 17775 8472 17858 8578
rect 17892 8472 18095 8578
rect 17775 8465 17815 8472
rect 17858 8465 18095 8472
rect 18325 8578 18442 8585
rect 18485 8578 18645 8585
rect 18325 8472 18408 8578
rect 18442 8472 18645 8578
rect 18325 8465 18365 8472
rect 18408 8465 18645 8472
rect 18875 8578 18992 8585
rect 19035 8578 19195 8585
rect 18875 8472 18958 8578
rect 18992 8472 19195 8578
rect 18875 8465 18915 8472
rect 18958 8465 19195 8472
rect 765 8425 885 8465
rect 1315 8425 1435 8465
rect 1865 8425 1985 8465
rect 2415 8425 2535 8465
rect 2965 8425 3085 8465
rect 3515 8425 3635 8465
rect 4065 8425 4185 8465
rect 4615 8425 4735 8465
rect 5165 8425 5285 8465
rect 5715 8425 5835 8465
rect 6265 8425 6385 8465
rect 6815 8425 6935 8465
rect 7365 8425 7485 8465
rect 7915 8425 8035 8465
rect 8465 8425 8585 8465
rect 9015 8425 9135 8465
rect 9565 8425 9685 8465
rect 10115 8425 10235 8465
rect 10665 8425 10785 8465
rect 11215 8425 11335 8465
rect 11765 8425 11885 8465
rect 12315 8425 12435 8465
rect 12865 8425 12985 8465
rect 13415 8425 13535 8465
rect 13965 8425 14085 8465
rect 14515 8425 14635 8465
rect 15065 8425 15185 8465
rect 15615 8425 15735 8465
rect 16165 8425 16285 8465
rect 16715 8425 16835 8465
rect 17265 8425 17385 8465
rect 17815 8425 17935 8465
rect 18365 8425 18485 8465
rect 18915 8425 19035 8465
rect 19202 8312 19204 8738
rect 500 8225 507 8275
rect 19202 8196 19217 8202
rect 628 8172 885 8195
rect 1178 8172 1435 8195
rect 1728 8172 1985 8195
rect 2278 8172 2535 8195
rect 2828 8172 3085 8195
rect 3378 8172 3635 8195
rect 3928 8172 4185 8195
rect 4478 8172 4735 8195
rect 5028 8172 5285 8195
rect 5578 8172 5835 8195
rect 6128 8172 6385 8195
rect 6678 8172 6935 8195
rect 7228 8172 7485 8195
rect 7778 8172 8035 8195
rect 8328 8172 8585 8195
rect 8878 8172 9135 8195
rect 9428 8172 9685 8195
rect 9978 8172 10235 8195
rect 10528 8172 10785 8195
rect 11078 8172 11335 8195
rect 11628 8172 11885 8195
rect 12178 8172 12435 8195
rect 12728 8172 12985 8195
rect 13278 8172 13535 8195
rect 13828 8172 14085 8195
rect 14378 8172 14635 8195
rect 14928 8172 15185 8195
rect 15478 8172 15735 8195
rect 16028 8172 16285 8195
rect 16578 8172 16835 8195
rect 17128 8172 17385 8195
rect 17678 8172 17935 8195
rect 18228 8172 18485 8195
rect 18778 8172 19035 8195
rect 605 8035 609 8172
rect 784 8075 885 8172
rect 765 8035 885 8075
rect 1155 8035 1159 8172
rect 1334 8075 1435 8172
rect 1315 8035 1435 8075
rect 1705 8035 1709 8172
rect 1884 8075 1985 8172
rect 1865 8035 1985 8075
rect 2255 8035 2259 8172
rect 2434 8075 2535 8172
rect 2415 8035 2535 8075
rect 2805 8035 2809 8172
rect 2984 8075 3085 8172
rect 2965 8035 3085 8075
rect 3355 8035 3359 8172
rect 3534 8075 3635 8172
rect 3515 8035 3635 8075
rect 3905 8035 3909 8172
rect 4084 8075 4185 8172
rect 4065 8035 4185 8075
rect 4455 8035 4459 8172
rect 4634 8075 4735 8172
rect 4615 8035 4735 8075
rect 5005 8035 5009 8172
rect 5184 8075 5285 8172
rect 5165 8035 5285 8075
rect 5555 8035 5559 8172
rect 5734 8075 5835 8172
rect 5715 8035 5835 8075
rect 6105 8035 6109 8172
rect 6284 8075 6385 8172
rect 6265 8035 6385 8075
rect 6655 8035 6659 8172
rect 6834 8075 6935 8172
rect 6815 8035 6935 8075
rect 7205 8035 7209 8172
rect 7384 8075 7485 8172
rect 7365 8035 7485 8075
rect 7755 8035 7759 8172
rect 7934 8075 8035 8172
rect 7915 8035 8035 8075
rect 8305 8035 8309 8172
rect 8484 8075 8585 8172
rect 8465 8035 8585 8075
rect 8855 8035 8859 8172
rect 9034 8075 9135 8172
rect 9015 8035 9135 8075
rect 9405 8035 9409 8172
rect 9584 8075 9685 8172
rect 9565 8035 9685 8075
rect 9955 8035 9959 8172
rect 10134 8075 10235 8172
rect 10115 8035 10235 8075
rect 10505 8035 10509 8172
rect 10684 8075 10785 8172
rect 10665 8035 10785 8075
rect 11055 8035 11059 8172
rect 11234 8075 11335 8172
rect 11215 8035 11335 8075
rect 11605 8035 11609 8172
rect 11784 8075 11885 8172
rect 11765 8035 11885 8075
rect 12155 8035 12159 8172
rect 12334 8075 12435 8172
rect 12315 8035 12435 8075
rect 12705 8035 12709 8172
rect 12884 8075 12985 8172
rect 12865 8035 12985 8075
rect 13255 8035 13259 8172
rect 13434 8075 13535 8172
rect 13415 8035 13535 8075
rect 13805 8035 13809 8172
rect 13984 8075 14085 8172
rect 13965 8035 14085 8075
rect 14355 8035 14359 8172
rect 14534 8075 14635 8172
rect 14515 8035 14635 8075
rect 14905 8035 14909 8172
rect 15084 8075 15185 8172
rect 15065 8035 15185 8075
rect 15455 8035 15459 8172
rect 15634 8075 15735 8172
rect 15615 8035 15735 8075
rect 16005 8035 16009 8172
rect 16184 8075 16285 8172
rect 16165 8035 16285 8075
rect 16555 8035 16559 8172
rect 16734 8075 16835 8172
rect 16715 8035 16835 8075
rect 17105 8035 17109 8172
rect 17284 8075 17385 8172
rect 17265 8035 17385 8075
rect 17655 8035 17659 8172
rect 17834 8075 17935 8172
rect 17815 8035 17935 8075
rect 18205 8035 18209 8172
rect 18384 8075 18485 8172
rect 18365 8035 18485 8075
rect 18755 8035 18759 8172
rect 18934 8075 19035 8172
rect 18915 8035 19035 8075
rect 725 8028 842 8035
rect 885 8028 1045 8035
rect 725 7922 808 8028
rect 842 7922 1045 8028
rect 725 7915 765 7922
rect 808 7915 1045 7922
rect 1275 8028 1392 8035
rect 1435 8028 1595 8035
rect 1275 7922 1358 8028
rect 1392 7922 1595 8028
rect 1275 7915 1315 7922
rect 1358 7915 1595 7922
rect 1825 8028 1942 8035
rect 1985 8028 2145 8035
rect 1825 7922 1908 8028
rect 1942 7922 2145 8028
rect 1825 7915 1865 7922
rect 1908 7915 2145 7922
rect 2375 8028 2492 8035
rect 2535 8028 2695 8035
rect 2375 7922 2458 8028
rect 2492 7922 2695 8028
rect 2375 7915 2415 7922
rect 2458 7915 2695 7922
rect 2925 8028 3042 8035
rect 3085 8028 3245 8035
rect 2925 7922 3008 8028
rect 3042 7922 3245 8028
rect 2925 7915 2965 7922
rect 3008 7915 3245 7922
rect 3475 8028 3592 8035
rect 3635 8028 3795 8035
rect 3475 7922 3558 8028
rect 3592 7922 3795 8028
rect 3475 7915 3515 7922
rect 3558 7915 3795 7922
rect 4025 8028 4142 8035
rect 4185 8028 4345 8035
rect 4025 7922 4108 8028
rect 4142 7922 4345 8028
rect 4025 7915 4065 7922
rect 4108 7915 4345 7922
rect 4575 8028 4692 8035
rect 4735 8028 4895 8035
rect 4575 7922 4658 8028
rect 4692 7922 4895 8028
rect 4575 7915 4615 7922
rect 4658 7915 4895 7922
rect 5125 8028 5242 8035
rect 5285 8028 5445 8035
rect 5125 7922 5208 8028
rect 5242 7922 5445 8028
rect 5125 7915 5165 7922
rect 5208 7915 5445 7922
rect 5675 8028 5792 8035
rect 5835 8028 5995 8035
rect 5675 7922 5758 8028
rect 5792 7922 5995 8028
rect 5675 7915 5715 7922
rect 5758 7915 5995 7922
rect 6225 8028 6342 8035
rect 6385 8028 6545 8035
rect 6225 7922 6308 8028
rect 6342 7922 6545 8028
rect 6225 7915 6265 7922
rect 6308 7915 6545 7922
rect 6775 8028 6892 8035
rect 6935 8028 7095 8035
rect 6775 7922 6858 8028
rect 6892 7922 7095 8028
rect 6775 7915 6815 7922
rect 6858 7915 7095 7922
rect 7325 8028 7442 8035
rect 7485 8028 7645 8035
rect 7325 7922 7408 8028
rect 7442 7922 7645 8028
rect 7325 7915 7365 7922
rect 7408 7915 7645 7922
rect 7875 8028 7992 8035
rect 8035 8028 8195 8035
rect 7875 7922 7958 8028
rect 7992 7922 8195 8028
rect 7875 7915 7915 7922
rect 7958 7915 8195 7922
rect 8425 8028 8542 8035
rect 8585 8028 8745 8035
rect 8425 7922 8508 8028
rect 8542 7922 8745 8028
rect 8425 7915 8465 7922
rect 8508 7915 8745 7922
rect 8975 8028 9092 8035
rect 9135 8028 9295 8035
rect 8975 7922 9058 8028
rect 9092 7922 9295 8028
rect 8975 7915 9015 7922
rect 9058 7915 9295 7922
rect 9525 8028 9642 8035
rect 9685 8028 9845 8035
rect 9525 7922 9608 8028
rect 9642 7922 9845 8028
rect 9525 7915 9565 7922
rect 9608 7915 9845 7922
rect 10075 8028 10192 8035
rect 10235 8028 10395 8035
rect 10075 7922 10158 8028
rect 10192 7922 10395 8028
rect 10075 7915 10115 7922
rect 10158 7915 10395 7922
rect 10625 8028 10742 8035
rect 10785 8028 10945 8035
rect 10625 7922 10708 8028
rect 10742 7922 10945 8028
rect 10625 7915 10665 7922
rect 10708 7915 10945 7922
rect 11175 8028 11292 8035
rect 11335 8028 11495 8035
rect 11175 7922 11258 8028
rect 11292 7922 11495 8028
rect 11175 7915 11215 7922
rect 11258 7915 11495 7922
rect 11725 8028 11842 8035
rect 11885 8028 12045 8035
rect 11725 7922 11808 8028
rect 11842 7922 12045 8028
rect 11725 7915 11765 7922
rect 11808 7915 12045 7922
rect 12275 8028 12392 8035
rect 12435 8028 12595 8035
rect 12275 7922 12358 8028
rect 12392 7922 12595 8028
rect 12275 7915 12315 7922
rect 12358 7915 12595 7922
rect 12825 8028 12942 8035
rect 12985 8028 13145 8035
rect 12825 7922 12908 8028
rect 12942 7922 13145 8028
rect 12825 7915 12865 7922
rect 12908 7915 13145 7922
rect 13375 8028 13492 8035
rect 13535 8028 13695 8035
rect 13375 7922 13458 8028
rect 13492 7922 13695 8028
rect 13375 7915 13415 7922
rect 13458 7915 13695 7922
rect 13925 8028 14042 8035
rect 14085 8028 14245 8035
rect 13925 7922 14008 8028
rect 14042 7922 14245 8028
rect 13925 7915 13965 7922
rect 14008 7915 14245 7922
rect 14475 8028 14592 8035
rect 14635 8028 14795 8035
rect 14475 7922 14558 8028
rect 14592 7922 14795 8028
rect 14475 7915 14515 7922
rect 14558 7915 14795 7922
rect 15025 8028 15142 8035
rect 15185 8028 15345 8035
rect 15025 7922 15108 8028
rect 15142 7922 15345 8028
rect 15025 7915 15065 7922
rect 15108 7915 15345 7922
rect 15575 8028 15692 8035
rect 15735 8028 15895 8035
rect 15575 7922 15658 8028
rect 15692 7922 15895 8028
rect 15575 7915 15615 7922
rect 15658 7915 15895 7922
rect 16125 8028 16242 8035
rect 16285 8028 16445 8035
rect 16125 7922 16208 8028
rect 16242 7922 16445 8028
rect 16125 7915 16165 7922
rect 16208 7915 16445 7922
rect 16675 8028 16792 8035
rect 16835 8028 16995 8035
rect 16675 7922 16758 8028
rect 16792 7922 16995 8028
rect 16675 7915 16715 7922
rect 16758 7915 16995 7922
rect 17225 8028 17342 8035
rect 17385 8028 17545 8035
rect 17225 7922 17308 8028
rect 17342 7922 17545 8028
rect 17225 7915 17265 7922
rect 17308 7915 17545 7922
rect 17775 8028 17892 8035
rect 17935 8028 18095 8035
rect 17775 7922 17858 8028
rect 17892 7922 18095 8028
rect 17775 7915 17815 7922
rect 17858 7915 18095 7922
rect 18325 8028 18442 8035
rect 18485 8028 18645 8035
rect 18325 7922 18408 8028
rect 18442 7922 18645 8028
rect 18325 7915 18365 7922
rect 18408 7915 18645 7922
rect 18875 8028 18992 8035
rect 19035 8028 19195 8035
rect 18875 7922 18958 8028
rect 18992 7922 19195 8028
rect 18875 7915 18915 7922
rect 18958 7915 19195 7922
rect 765 7875 885 7915
rect 1315 7875 1435 7915
rect 1865 7875 1985 7915
rect 2415 7875 2535 7915
rect 2965 7875 3085 7915
rect 3515 7875 3635 7915
rect 4065 7875 4185 7915
rect 4615 7875 4735 7915
rect 5165 7875 5285 7915
rect 5715 7875 5835 7915
rect 6265 7875 6385 7915
rect 6815 7875 6935 7915
rect 7365 7875 7485 7915
rect 7915 7875 8035 7915
rect 8465 7875 8585 7915
rect 9015 7875 9135 7915
rect 9565 7875 9685 7915
rect 10115 7875 10235 7915
rect 10665 7875 10785 7915
rect 11215 7875 11335 7915
rect 11765 7875 11885 7915
rect 12315 7875 12435 7915
rect 12865 7875 12985 7915
rect 13415 7875 13535 7915
rect 13965 7875 14085 7915
rect 14515 7875 14635 7915
rect 15065 7875 15185 7915
rect 15615 7875 15735 7915
rect 16165 7875 16285 7915
rect 16715 7875 16835 7915
rect 17265 7875 17385 7915
rect 17815 7875 17935 7915
rect 18365 7875 18485 7915
rect 18915 7875 19035 7915
rect 19185 7754 19200 7771
rect 19202 7762 19204 8188
rect 19202 7748 19217 7754
rect 500 7675 507 7725
rect 500 7239 525 7640
rect 628 7622 885 7645
rect 1178 7622 1435 7645
rect 1728 7622 1985 7645
rect 2278 7622 2535 7645
rect 2828 7622 3085 7645
rect 3378 7622 3635 7645
rect 3928 7622 4185 7645
rect 4478 7622 4735 7645
rect 5028 7622 5285 7645
rect 5578 7622 5835 7645
rect 6128 7622 6385 7645
rect 6678 7622 6935 7645
rect 7228 7622 7485 7645
rect 7778 7622 8035 7645
rect 8328 7622 8585 7645
rect 8878 7622 9135 7645
rect 9428 7622 9685 7645
rect 9978 7622 10235 7645
rect 10528 7622 10785 7645
rect 11078 7622 11335 7645
rect 11628 7622 11885 7645
rect 12178 7622 12435 7645
rect 12728 7622 12985 7645
rect 13278 7622 13535 7645
rect 13828 7622 14085 7645
rect 14378 7622 14635 7645
rect 14928 7622 15185 7645
rect 15478 7622 15735 7645
rect 16028 7622 16285 7645
rect 16578 7622 16835 7645
rect 17128 7622 17385 7645
rect 17678 7622 17935 7645
rect 18228 7622 18485 7645
rect 18778 7622 19035 7645
rect 605 7485 609 7622
rect 784 7525 885 7622
rect 765 7485 885 7525
rect 1155 7485 1159 7622
rect 1334 7525 1435 7622
rect 1315 7485 1435 7525
rect 1705 7485 1709 7622
rect 1884 7525 1985 7622
rect 1865 7485 1985 7525
rect 2255 7485 2259 7622
rect 2434 7525 2535 7622
rect 2415 7485 2535 7525
rect 2805 7485 2809 7622
rect 2984 7525 3085 7622
rect 2965 7485 3085 7525
rect 3355 7485 3359 7622
rect 3534 7525 3635 7622
rect 3515 7485 3635 7525
rect 3905 7485 3909 7622
rect 4084 7525 4185 7622
rect 4065 7485 4185 7525
rect 4455 7485 4459 7622
rect 4634 7525 4735 7622
rect 4615 7485 4735 7525
rect 5005 7485 5009 7622
rect 5184 7525 5285 7622
rect 5165 7485 5285 7525
rect 5555 7485 5559 7622
rect 5734 7525 5835 7622
rect 5715 7485 5835 7525
rect 6105 7485 6109 7622
rect 6284 7525 6385 7622
rect 6265 7485 6385 7525
rect 6655 7485 6659 7622
rect 6834 7525 6935 7622
rect 6815 7485 6935 7525
rect 7205 7485 7209 7622
rect 7384 7525 7485 7622
rect 7365 7485 7485 7525
rect 7755 7485 7759 7622
rect 7934 7525 8035 7622
rect 7915 7485 8035 7525
rect 8305 7485 8309 7622
rect 8484 7525 8585 7622
rect 8465 7485 8585 7525
rect 8855 7485 8859 7622
rect 9034 7525 9135 7622
rect 9015 7485 9135 7525
rect 9405 7485 9409 7622
rect 9584 7525 9685 7622
rect 9565 7485 9685 7525
rect 9955 7485 9959 7622
rect 10134 7525 10235 7622
rect 10115 7485 10235 7525
rect 10505 7485 10509 7622
rect 10684 7525 10785 7622
rect 10665 7485 10785 7525
rect 11055 7485 11059 7622
rect 11234 7525 11335 7622
rect 11215 7485 11335 7525
rect 11605 7485 11609 7622
rect 11784 7525 11885 7622
rect 11765 7485 11885 7525
rect 12155 7485 12159 7622
rect 12334 7525 12435 7622
rect 12315 7485 12435 7525
rect 12705 7485 12709 7622
rect 12884 7525 12985 7622
rect 12865 7485 12985 7525
rect 13255 7485 13259 7622
rect 13434 7525 13535 7622
rect 13415 7485 13535 7525
rect 13805 7485 13809 7622
rect 13984 7525 14085 7622
rect 13965 7485 14085 7525
rect 14355 7485 14359 7622
rect 14534 7525 14635 7622
rect 14515 7485 14635 7525
rect 14905 7485 14909 7622
rect 15084 7525 15185 7622
rect 15065 7485 15185 7525
rect 15455 7485 15459 7622
rect 15634 7525 15735 7622
rect 15615 7485 15735 7525
rect 16005 7485 16009 7622
rect 16184 7525 16285 7622
rect 16165 7485 16285 7525
rect 16555 7485 16559 7622
rect 16734 7525 16835 7622
rect 16715 7485 16835 7525
rect 17105 7485 17109 7622
rect 17284 7525 17385 7622
rect 17265 7485 17385 7525
rect 17655 7485 17659 7622
rect 17834 7525 17935 7622
rect 17815 7485 17935 7525
rect 18205 7485 18209 7622
rect 18384 7525 18485 7622
rect 18365 7485 18485 7525
rect 18755 7485 18759 7622
rect 18934 7525 19035 7622
rect 18915 7485 19035 7525
rect 725 7478 842 7485
rect 885 7478 1045 7485
rect 725 7372 808 7478
rect 842 7372 1045 7478
rect 725 7365 765 7372
rect 808 7365 1045 7372
rect 1275 7478 1392 7485
rect 1435 7478 1595 7485
rect 1275 7372 1358 7478
rect 1392 7372 1595 7478
rect 1275 7365 1315 7372
rect 1358 7365 1595 7372
rect 1825 7478 1942 7485
rect 1985 7478 2145 7485
rect 1825 7372 1908 7478
rect 1942 7372 2145 7478
rect 1825 7365 1865 7372
rect 1908 7365 2145 7372
rect 2375 7478 2492 7485
rect 2535 7478 2695 7485
rect 2375 7372 2458 7478
rect 2492 7372 2695 7478
rect 2375 7365 2415 7372
rect 2458 7365 2695 7372
rect 2925 7478 3042 7485
rect 3085 7478 3245 7485
rect 2925 7372 3008 7478
rect 3042 7372 3245 7478
rect 2925 7365 2965 7372
rect 3008 7365 3245 7372
rect 3475 7478 3592 7485
rect 3635 7478 3795 7485
rect 3475 7372 3558 7478
rect 3592 7372 3795 7478
rect 3475 7365 3515 7372
rect 3558 7365 3795 7372
rect 4025 7478 4142 7485
rect 4185 7478 4345 7485
rect 4025 7372 4108 7478
rect 4142 7372 4345 7478
rect 4025 7365 4065 7372
rect 4108 7365 4345 7372
rect 4575 7478 4692 7485
rect 4735 7478 4895 7485
rect 4575 7372 4658 7478
rect 4692 7372 4895 7478
rect 4575 7365 4615 7372
rect 4658 7365 4895 7372
rect 5125 7478 5242 7485
rect 5285 7478 5445 7485
rect 5125 7372 5208 7478
rect 5242 7372 5445 7478
rect 5125 7365 5165 7372
rect 5208 7365 5445 7372
rect 5675 7478 5792 7485
rect 5835 7478 5995 7485
rect 5675 7372 5758 7478
rect 5792 7372 5995 7478
rect 5675 7365 5715 7372
rect 5758 7365 5995 7372
rect 6225 7478 6342 7485
rect 6385 7478 6545 7485
rect 6225 7372 6308 7478
rect 6342 7372 6545 7478
rect 6225 7365 6265 7372
rect 6308 7365 6545 7372
rect 6775 7478 6892 7485
rect 6935 7478 7095 7485
rect 6775 7372 6858 7478
rect 6892 7372 7095 7478
rect 6775 7365 6815 7372
rect 6858 7365 7095 7372
rect 7325 7478 7442 7485
rect 7485 7478 7645 7485
rect 7325 7372 7408 7478
rect 7442 7372 7645 7478
rect 7325 7365 7365 7372
rect 7408 7365 7645 7372
rect 7875 7478 7992 7485
rect 8035 7478 8195 7485
rect 7875 7372 7958 7478
rect 7992 7372 8195 7478
rect 7875 7365 7915 7372
rect 7958 7365 8195 7372
rect 8425 7478 8542 7485
rect 8585 7478 8745 7485
rect 8425 7372 8508 7478
rect 8542 7372 8745 7478
rect 8425 7365 8465 7372
rect 8508 7365 8745 7372
rect 8975 7478 9092 7485
rect 9135 7478 9295 7485
rect 8975 7372 9058 7478
rect 9092 7372 9295 7478
rect 8975 7365 9015 7372
rect 9058 7365 9295 7372
rect 9525 7478 9642 7485
rect 9685 7478 9845 7485
rect 9525 7372 9608 7478
rect 9642 7372 9845 7478
rect 9525 7365 9565 7372
rect 9608 7365 9845 7372
rect 10075 7478 10192 7485
rect 10235 7478 10395 7485
rect 10075 7372 10158 7478
rect 10192 7372 10395 7478
rect 10075 7365 10115 7372
rect 10158 7365 10395 7372
rect 10625 7478 10742 7485
rect 10785 7478 10945 7485
rect 10625 7372 10708 7478
rect 10742 7372 10945 7478
rect 10625 7365 10665 7372
rect 10708 7365 10945 7372
rect 11175 7478 11292 7485
rect 11335 7478 11495 7485
rect 11175 7372 11258 7478
rect 11292 7372 11495 7478
rect 11175 7365 11215 7372
rect 11258 7365 11495 7372
rect 11725 7478 11842 7485
rect 11885 7478 12045 7485
rect 11725 7372 11808 7478
rect 11842 7372 12045 7478
rect 11725 7365 11765 7372
rect 11808 7365 12045 7372
rect 12275 7478 12392 7485
rect 12435 7478 12595 7485
rect 12275 7372 12358 7478
rect 12392 7372 12595 7478
rect 12275 7365 12315 7372
rect 12358 7365 12595 7372
rect 12825 7478 12942 7485
rect 12985 7478 13145 7485
rect 12825 7372 12908 7478
rect 12942 7372 13145 7478
rect 12825 7365 12865 7372
rect 12908 7365 13145 7372
rect 13375 7478 13492 7485
rect 13535 7478 13695 7485
rect 13375 7372 13458 7478
rect 13492 7372 13695 7478
rect 13375 7365 13415 7372
rect 13458 7365 13695 7372
rect 13925 7478 14042 7485
rect 14085 7478 14245 7485
rect 13925 7372 14008 7478
rect 14042 7372 14245 7478
rect 13925 7365 13965 7372
rect 14008 7365 14245 7372
rect 14475 7478 14592 7485
rect 14635 7478 14795 7485
rect 14475 7372 14558 7478
rect 14592 7372 14795 7478
rect 14475 7365 14515 7372
rect 14558 7365 14795 7372
rect 15025 7478 15142 7485
rect 15185 7478 15345 7485
rect 15025 7372 15108 7478
rect 15142 7372 15345 7478
rect 15025 7365 15065 7372
rect 15108 7365 15345 7372
rect 15575 7478 15692 7485
rect 15735 7478 15895 7485
rect 15575 7372 15658 7478
rect 15692 7372 15895 7478
rect 15575 7365 15615 7372
rect 15658 7365 15895 7372
rect 16125 7478 16242 7485
rect 16285 7478 16445 7485
rect 16125 7372 16208 7478
rect 16242 7372 16445 7478
rect 16125 7365 16165 7372
rect 16208 7365 16445 7372
rect 16675 7478 16792 7485
rect 16835 7478 16995 7485
rect 16675 7372 16758 7478
rect 16792 7372 16995 7478
rect 16675 7365 16715 7372
rect 16758 7365 16995 7372
rect 17225 7478 17342 7485
rect 17385 7478 17545 7485
rect 17225 7372 17308 7478
rect 17342 7372 17545 7478
rect 17225 7365 17265 7372
rect 17308 7365 17545 7372
rect 17775 7478 17892 7485
rect 17935 7478 18095 7485
rect 17775 7372 17858 7478
rect 17892 7372 18095 7478
rect 17775 7365 17815 7372
rect 17858 7365 18095 7372
rect 18325 7478 18442 7485
rect 18485 7478 18645 7485
rect 18325 7372 18408 7478
rect 18442 7372 18645 7478
rect 18325 7365 18365 7372
rect 18408 7365 18645 7372
rect 18875 7478 18992 7485
rect 19035 7478 19195 7485
rect 18875 7372 18958 7478
rect 18992 7372 19195 7478
rect 18875 7365 18915 7372
rect 18958 7365 19195 7372
rect 765 7325 885 7365
rect 1315 7325 1435 7365
rect 1865 7325 1985 7365
rect 2415 7325 2535 7365
rect 2965 7325 3085 7365
rect 3515 7325 3635 7365
rect 4065 7325 4185 7365
rect 4615 7325 4735 7365
rect 5165 7325 5285 7365
rect 5715 7325 5835 7365
rect 6265 7325 6385 7365
rect 6815 7325 6935 7365
rect 7365 7325 7485 7365
rect 7915 7325 8035 7365
rect 8465 7325 8585 7365
rect 9015 7325 9135 7365
rect 9565 7325 9685 7365
rect 10115 7325 10235 7365
rect 10665 7325 10785 7365
rect 11215 7325 11335 7365
rect 11765 7325 11885 7365
rect 12315 7325 12435 7365
rect 12865 7325 12985 7365
rect 13415 7325 13535 7365
rect 13965 7325 14085 7365
rect 14515 7325 14635 7365
rect 15065 7325 15185 7365
rect 15615 7325 15735 7365
rect 16165 7325 16285 7365
rect 16715 7325 16835 7365
rect 17265 7325 17385 7365
rect 17815 7325 17935 7365
rect 18365 7325 18485 7365
rect 18915 7325 19035 7365
rect 19202 7212 19204 7638
rect 500 7125 507 7175
rect 19202 7096 19217 7102
rect 628 7072 885 7095
rect 1178 7072 1435 7095
rect 1728 7072 1985 7095
rect 2278 7072 2535 7095
rect 2828 7072 3085 7095
rect 3378 7072 3635 7095
rect 3928 7072 4185 7095
rect 4478 7072 4735 7095
rect 5028 7072 5285 7095
rect 5578 7072 5835 7095
rect 6128 7072 6385 7095
rect 6678 7072 6935 7095
rect 7228 7072 7485 7095
rect 7778 7072 8035 7095
rect 8328 7072 8585 7095
rect 8878 7072 9135 7095
rect 9428 7072 9685 7095
rect 9978 7072 10235 7095
rect 10528 7072 10785 7095
rect 11078 7072 11335 7095
rect 11628 7072 11885 7095
rect 12178 7072 12435 7095
rect 12728 7072 12985 7095
rect 13278 7072 13535 7095
rect 13828 7072 14085 7095
rect 14378 7072 14635 7095
rect 14928 7072 15185 7095
rect 15478 7072 15735 7095
rect 16028 7072 16285 7095
rect 16578 7072 16835 7095
rect 17128 7072 17385 7095
rect 17678 7072 17935 7095
rect 18228 7072 18485 7095
rect 18778 7072 19035 7095
rect 605 6935 609 7072
rect 784 6975 885 7072
rect 765 6935 885 6975
rect 1155 6935 1159 7072
rect 1334 6975 1435 7072
rect 1315 6935 1435 6975
rect 1705 6935 1709 7072
rect 1884 6975 1985 7072
rect 1865 6935 1985 6975
rect 2255 6935 2259 7072
rect 2434 6975 2535 7072
rect 2415 6935 2535 6975
rect 2805 6935 2809 7072
rect 2984 6975 3085 7072
rect 2965 6935 3085 6975
rect 3355 6935 3359 7072
rect 3534 6975 3635 7072
rect 3515 6935 3635 6975
rect 3905 6935 3909 7072
rect 4084 6975 4185 7072
rect 4065 6935 4185 6975
rect 4455 6935 4459 7072
rect 4634 6975 4735 7072
rect 4615 6935 4735 6975
rect 5005 6935 5009 7072
rect 5184 6975 5285 7072
rect 5165 6935 5285 6975
rect 5555 6935 5559 7072
rect 5734 6975 5835 7072
rect 5715 6935 5835 6975
rect 6105 6935 6109 7072
rect 6284 6975 6385 7072
rect 6265 6935 6385 6975
rect 6655 6935 6659 7072
rect 6834 6975 6935 7072
rect 6815 6935 6935 6975
rect 7205 6935 7209 7072
rect 7384 6975 7485 7072
rect 7365 6935 7485 6975
rect 7755 6935 7759 7072
rect 7934 6975 8035 7072
rect 7915 6935 8035 6975
rect 8305 6935 8309 7072
rect 8484 6975 8585 7072
rect 8465 6935 8585 6975
rect 8855 6935 8859 7072
rect 9034 6975 9135 7072
rect 9015 6935 9135 6975
rect 9405 6935 9409 7072
rect 9584 6975 9685 7072
rect 9565 6935 9685 6975
rect 9955 6935 9959 7072
rect 10134 6975 10235 7072
rect 10115 6935 10235 6975
rect 10505 6935 10509 7072
rect 10684 6975 10785 7072
rect 10665 6935 10785 6975
rect 11055 6935 11059 7072
rect 11234 6975 11335 7072
rect 11215 6935 11335 6975
rect 11605 6935 11609 7072
rect 11784 6975 11885 7072
rect 11765 6935 11885 6975
rect 12155 6935 12159 7072
rect 12334 6975 12435 7072
rect 12315 6935 12435 6975
rect 12705 6935 12709 7072
rect 12884 6975 12985 7072
rect 12865 6935 12985 6975
rect 13255 6935 13259 7072
rect 13434 6975 13535 7072
rect 13415 6935 13535 6975
rect 13805 6935 13809 7072
rect 13984 6975 14085 7072
rect 13965 6935 14085 6975
rect 14355 6935 14359 7072
rect 14534 6975 14635 7072
rect 14515 6935 14635 6975
rect 14905 6935 14909 7072
rect 15084 6975 15185 7072
rect 15065 6935 15185 6975
rect 15455 6935 15459 7072
rect 15634 6975 15735 7072
rect 15615 6935 15735 6975
rect 16005 6935 16009 7072
rect 16184 6975 16285 7072
rect 16165 6935 16285 6975
rect 16555 6935 16559 7072
rect 16734 6975 16835 7072
rect 16715 6935 16835 6975
rect 17105 6935 17109 7072
rect 17284 6975 17385 7072
rect 17265 6935 17385 6975
rect 17655 6935 17659 7072
rect 17834 6975 17935 7072
rect 17815 6935 17935 6975
rect 18205 6935 18209 7072
rect 18384 6975 18485 7072
rect 18365 6935 18485 6975
rect 18755 6935 18759 7072
rect 18934 6975 19035 7072
rect 18915 6935 19035 6975
rect 725 6928 842 6935
rect 885 6928 1045 6935
rect 725 6822 808 6928
rect 842 6822 1045 6928
rect 725 6815 765 6822
rect 808 6815 1045 6822
rect 1275 6928 1392 6935
rect 1435 6928 1595 6935
rect 1275 6822 1358 6928
rect 1392 6822 1595 6928
rect 1275 6815 1315 6822
rect 1358 6815 1595 6822
rect 1825 6928 1942 6935
rect 1985 6928 2145 6935
rect 1825 6822 1908 6928
rect 1942 6822 2145 6928
rect 1825 6815 1865 6822
rect 1908 6815 2145 6822
rect 2375 6928 2492 6935
rect 2535 6928 2695 6935
rect 2375 6822 2458 6928
rect 2492 6822 2695 6928
rect 2375 6815 2415 6822
rect 2458 6815 2695 6822
rect 2925 6928 3042 6935
rect 3085 6928 3245 6935
rect 2925 6822 3008 6928
rect 3042 6822 3245 6928
rect 2925 6815 2965 6822
rect 3008 6815 3245 6822
rect 3475 6928 3592 6935
rect 3635 6928 3795 6935
rect 3475 6822 3558 6928
rect 3592 6822 3795 6928
rect 3475 6815 3515 6822
rect 3558 6815 3795 6822
rect 4025 6928 4142 6935
rect 4185 6928 4345 6935
rect 4025 6822 4108 6928
rect 4142 6822 4345 6928
rect 4025 6815 4065 6822
rect 4108 6815 4345 6822
rect 4575 6928 4692 6935
rect 4735 6928 4895 6935
rect 4575 6822 4658 6928
rect 4692 6822 4895 6928
rect 4575 6815 4615 6822
rect 4658 6815 4895 6822
rect 5125 6928 5242 6935
rect 5285 6928 5445 6935
rect 5125 6822 5208 6928
rect 5242 6822 5445 6928
rect 5125 6815 5165 6822
rect 5208 6815 5445 6822
rect 5675 6928 5792 6935
rect 5835 6928 5995 6935
rect 5675 6822 5758 6928
rect 5792 6822 5995 6928
rect 5675 6815 5715 6822
rect 5758 6815 5995 6822
rect 6225 6928 6342 6935
rect 6385 6928 6545 6935
rect 6225 6822 6308 6928
rect 6342 6822 6545 6928
rect 6225 6815 6265 6822
rect 6308 6815 6545 6822
rect 6775 6928 6892 6935
rect 6935 6928 7095 6935
rect 6775 6822 6858 6928
rect 6892 6822 7095 6928
rect 6775 6815 6815 6822
rect 6858 6815 7095 6822
rect 7325 6928 7442 6935
rect 7485 6928 7645 6935
rect 7325 6822 7408 6928
rect 7442 6822 7645 6928
rect 7325 6815 7365 6822
rect 7408 6815 7645 6822
rect 7875 6928 7992 6935
rect 8035 6928 8195 6935
rect 7875 6822 7958 6928
rect 7992 6822 8195 6928
rect 7875 6815 7915 6822
rect 7958 6815 8195 6822
rect 8425 6928 8542 6935
rect 8585 6928 8745 6935
rect 8425 6822 8508 6928
rect 8542 6822 8745 6928
rect 8425 6815 8465 6822
rect 8508 6815 8745 6822
rect 8975 6928 9092 6935
rect 9135 6928 9295 6935
rect 8975 6822 9058 6928
rect 9092 6822 9295 6928
rect 8975 6815 9015 6822
rect 9058 6815 9295 6822
rect 9525 6928 9642 6935
rect 9685 6928 9845 6935
rect 9525 6822 9608 6928
rect 9642 6822 9845 6928
rect 9525 6815 9565 6822
rect 9608 6815 9845 6822
rect 10075 6928 10192 6935
rect 10235 6928 10395 6935
rect 10075 6822 10158 6928
rect 10192 6822 10395 6928
rect 10075 6815 10115 6822
rect 10158 6815 10395 6822
rect 10625 6928 10742 6935
rect 10785 6928 10945 6935
rect 10625 6822 10708 6928
rect 10742 6822 10945 6928
rect 10625 6815 10665 6822
rect 10708 6815 10945 6822
rect 11175 6928 11292 6935
rect 11335 6928 11495 6935
rect 11175 6822 11258 6928
rect 11292 6822 11495 6928
rect 11175 6815 11215 6822
rect 11258 6815 11495 6822
rect 11725 6928 11842 6935
rect 11885 6928 12045 6935
rect 11725 6822 11808 6928
rect 11842 6822 12045 6928
rect 11725 6815 11765 6822
rect 11808 6815 12045 6822
rect 12275 6928 12392 6935
rect 12435 6928 12595 6935
rect 12275 6822 12358 6928
rect 12392 6822 12595 6928
rect 12275 6815 12315 6822
rect 12358 6815 12595 6822
rect 12825 6928 12942 6935
rect 12985 6928 13145 6935
rect 12825 6822 12908 6928
rect 12942 6822 13145 6928
rect 12825 6815 12865 6822
rect 12908 6815 13145 6822
rect 13375 6928 13492 6935
rect 13535 6928 13695 6935
rect 13375 6822 13458 6928
rect 13492 6822 13695 6928
rect 13375 6815 13415 6822
rect 13458 6815 13695 6822
rect 13925 6928 14042 6935
rect 14085 6928 14245 6935
rect 13925 6822 14008 6928
rect 14042 6822 14245 6928
rect 13925 6815 13965 6822
rect 14008 6815 14245 6822
rect 14475 6928 14592 6935
rect 14635 6928 14795 6935
rect 14475 6822 14558 6928
rect 14592 6822 14795 6928
rect 14475 6815 14515 6822
rect 14558 6815 14795 6822
rect 15025 6928 15142 6935
rect 15185 6928 15345 6935
rect 15025 6822 15108 6928
rect 15142 6822 15345 6928
rect 15025 6815 15065 6822
rect 15108 6815 15345 6822
rect 15575 6928 15692 6935
rect 15735 6928 15895 6935
rect 15575 6822 15658 6928
rect 15692 6822 15895 6928
rect 15575 6815 15615 6822
rect 15658 6815 15895 6822
rect 16125 6928 16242 6935
rect 16285 6928 16445 6935
rect 16125 6822 16208 6928
rect 16242 6822 16445 6928
rect 16125 6815 16165 6822
rect 16208 6815 16445 6822
rect 16675 6928 16792 6935
rect 16835 6928 16995 6935
rect 16675 6822 16758 6928
rect 16792 6822 16995 6928
rect 16675 6815 16715 6822
rect 16758 6815 16995 6822
rect 17225 6928 17342 6935
rect 17385 6928 17545 6935
rect 17225 6822 17308 6928
rect 17342 6822 17545 6928
rect 17225 6815 17265 6822
rect 17308 6815 17545 6822
rect 17775 6928 17892 6935
rect 17935 6928 18095 6935
rect 17775 6822 17858 6928
rect 17892 6822 18095 6928
rect 17775 6815 17815 6822
rect 17858 6815 18095 6822
rect 18325 6928 18442 6935
rect 18485 6928 18645 6935
rect 18325 6822 18408 6928
rect 18442 6822 18645 6928
rect 18325 6815 18365 6822
rect 18408 6815 18645 6822
rect 18875 6928 18992 6935
rect 19035 6928 19195 6935
rect 18875 6822 18958 6928
rect 18992 6822 19195 6928
rect 18875 6815 18915 6822
rect 18958 6815 19195 6822
rect 765 6775 885 6815
rect 1315 6775 1435 6815
rect 1865 6775 1985 6815
rect 2415 6775 2535 6815
rect 2965 6775 3085 6815
rect 3515 6775 3635 6815
rect 4065 6775 4185 6815
rect 4615 6775 4735 6815
rect 5165 6775 5285 6815
rect 5715 6775 5835 6815
rect 6265 6775 6385 6815
rect 6815 6775 6935 6815
rect 7365 6775 7485 6815
rect 7915 6775 8035 6815
rect 8465 6775 8585 6815
rect 9015 6775 9135 6815
rect 9565 6775 9685 6815
rect 10115 6775 10235 6815
rect 10665 6775 10785 6815
rect 11215 6775 11335 6815
rect 11765 6775 11885 6815
rect 12315 6775 12435 6815
rect 12865 6775 12985 6815
rect 13415 6775 13535 6815
rect 13965 6775 14085 6815
rect 14515 6775 14635 6815
rect 15065 6775 15185 6815
rect 15615 6775 15735 6815
rect 16165 6775 16285 6815
rect 16715 6775 16835 6815
rect 17265 6775 17385 6815
rect 17815 6775 17935 6815
rect 18365 6775 18485 6815
rect 18915 6775 19035 6815
rect 19185 6654 19200 6671
rect 19202 6662 19204 7088
rect 19202 6648 19217 6654
rect 500 6575 507 6625
rect 500 6139 525 6540
rect 628 6522 885 6545
rect 1178 6522 1435 6545
rect 1728 6522 1985 6545
rect 2278 6522 2535 6545
rect 2828 6522 3085 6545
rect 3378 6522 3635 6545
rect 3928 6522 4185 6545
rect 4478 6522 4735 6545
rect 5028 6522 5285 6545
rect 5578 6522 5835 6545
rect 6128 6522 6385 6545
rect 6678 6522 6935 6545
rect 7228 6522 7485 6545
rect 7778 6522 8035 6545
rect 8328 6522 8585 6545
rect 8878 6522 9135 6545
rect 9428 6522 9685 6545
rect 9978 6522 10235 6545
rect 10528 6522 10785 6545
rect 11078 6522 11335 6545
rect 11628 6522 11885 6545
rect 12178 6522 12435 6545
rect 12728 6522 12985 6545
rect 13278 6522 13535 6545
rect 13828 6522 14085 6545
rect 14378 6522 14635 6545
rect 14928 6522 15185 6545
rect 15478 6522 15735 6545
rect 16028 6522 16285 6545
rect 16578 6522 16835 6545
rect 17128 6522 17385 6545
rect 17678 6522 17935 6545
rect 18228 6522 18485 6545
rect 18778 6522 19035 6545
rect 605 6385 609 6522
rect 784 6425 885 6522
rect 765 6385 885 6425
rect 1155 6385 1159 6522
rect 1334 6425 1435 6522
rect 1315 6385 1435 6425
rect 1705 6385 1709 6522
rect 1884 6425 1985 6522
rect 1865 6385 1985 6425
rect 2255 6385 2259 6522
rect 2434 6425 2535 6522
rect 2415 6385 2535 6425
rect 2805 6385 2809 6522
rect 2984 6425 3085 6522
rect 2965 6385 3085 6425
rect 3355 6385 3359 6522
rect 3534 6425 3635 6522
rect 3515 6385 3635 6425
rect 3905 6385 3909 6522
rect 4084 6425 4185 6522
rect 4065 6385 4185 6425
rect 4455 6385 4459 6522
rect 4634 6425 4735 6522
rect 4615 6385 4735 6425
rect 5005 6385 5009 6522
rect 5184 6425 5285 6522
rect 5165 6385 5285 6425
rect 5555 6385 5559 6522
rect 5734 6425 5835 6522
rect 5715 6385 5835 6425
rect 6105 6385 6109 6522
rect 6284 6425 6385 6522
rect 6265 6385 6385 6425
rect 6655 6385 6659 6522
rect 6834 6425 6935 6522
rect 6815 6385 6935 6425
rect 7205 6385 7209 6522
rect 7384 6425 7485 6522
rect 7365 6385 7485 6425
rect 7755 6385 7759 6522
rect 7934 6425 8035 6522
rect 7915 6385 8035 6425
rect 8305 6385 8309 6522
rect 8484 6425 8585 6522
rect 8465 6385 8585 6425
rect 8855 6385 8859 6522
rect 9034 6425 9135 6522
rect 9015 6385 9135 6425
rect 9405 6385 9409 6522
rect 9584 6425 9685 6522
rect 9565 6385 9685 6425
rect 9955 6385 9959 6522
rect 10134 6425 10235 6522
rect 10115 6385 10235 6425
rect 10505 6385 10509 6522
rect 10684 6425 10785 6522
rect 10665 6385 10785 6425
rect 11055 6385 11059 6522
rect 11234 6425 11335 6522
rect 11215 6385 11335 6425
rect 11605 6385 11609 6522
rect 11784 6425 11885 6522
rect 11765 6385 11885 6425
rect 12155 6385 12159 6522
rect 12334 6425 12435 6522
rect 12315 6385 12435 6425
rect 12705 6385 12709 6522
rect 12884 6425 12985 6522
rect 12865 6385 12985 6425
rect 13255 6385 13259 6522
rect 13434 6425 13535 6522
rect 13415 6385 13535 6425
rect 13805 6385 13809 6522
rect 13984 6425 14085 6522
rect 13965 6385 14085 6425
rect 14355 6385 14359 6522
rect 14534 6425 14635 6522
rect 14515 6385 14635 6425
rect 14905 6385 14909 6522
rect 15084 6425 15185 6522
rect 15065 6385 15185 6425
rect 15455 6385 15459 6522
rect 15634 6425 15735 6522
rect 15615 6385 15735 6425
rect 16005 6385 16009 6522
rect 16184 6425 16285 6522
rect 16165 6385 16285 6425
rect 16555 6385 16559 6522
rect 16734 6425 16835 6522
rect 16715 6385 16835 6425
rect 17105 6385 17109 6522
rect 17284 6425 17385 6522
rect 17265 6385 17385 6425
rect 17655 6385 17659 6522
rect 17834 6425 17935 6522
rect 17815 6385 17935 6425
rect 18205 6385 18209 6522
rect 18384 6425 18485 6522
rect 18365 6385 18485 6425
rect 18755 6385 18759 6522
rect 18934 6425 19035 6522
rect 18915 6385 19035 6425
rect 725 6378 842 6385
rect 885 6378 1045 6385
rect 725 6272 808 6378
rect 842 6272 1045 6378
rect 725 6265 765 6272
rect 808 6265 1045 6272
rect 1275 6378 1392 6385
rect 1435 6378 1595 6385
rect 1275 6272 1358 6378
rect 1392 6272 1595 6378
rect 1275 6265 1315 6272
rect 1358 6265 1595 6272
rect 1825 6378 1942 6385
rect 1985 6378 2145 6385
rect 1825 6272 1908 6378
rect 1942 6272 2145 6378
rect 1825 6265 1865 6272
rect 1908 6265 2145 6272
rect 2375 6378 2492 6385
rect 2535 6378 2695 6385
rect 2375 6272 2458 6378
rect 2492 6272 2695 6378
rect 2375 6265 2415 6272
rect 2458 6265 2695 6272
rect 2925 6378 3042 6385
rect 3085 6378 3245 6385
rect 2925 6272 3008 6378
rect 3042 6272 3245 6378
rect 2925 6265 2965 6272
rect 3008 6265 3245 6272
rect 3475 6378 3592 6385
rect 3635 6378 3795 6385
rect 3475 6272 3558 6378
rect 3592 6272 3795 6378
rect 3475 6265 3515 6272
rect 3558 6265 3795 6272
rect 4025 6378 4142 6385
rect 4185 6378 4345 6385
rect 4025 6272 4108 6378
rect 4142 6272 4345 6378
rect 4025 6265 4065 6272
rect 4108 6265 4345 6272
rect 4575 6378 4692 6385
rect 4735 6378 4895 6385
rect 4575 6272 4658 6378
rect 4692 6272 4895 6378
rect 4575 6265 4615 6272
rect 4658 6265 4895 6272
rect 5125 6378 5242 6385
rect 5285 6378 5445 6385
rect 5125 6272 5208 6378
rect 5242 6272 5445 6378
rect 5125 6265 5165 6272
rect 5208 6265 5445 6272
rect 5675 6378 5792 6385
rect 5835 6378 5995 6385
rect 5675 6272 5758 6378
rect 5792 6272 5995 6378
rect 5675 6265 5715 6272
rect 5758 6265 5995 6272
rect 6225 6378 6342 6385
rect 6385 6378 6545 6385
rect 6225 6272 6308 6378
rect 6342 6272 6545 6378
rect 6225 6265 6265 6272
rect 6308 6265 6545 6272
rect 6775 6378 6892 6385
rect 6935 6378 7095 6385
rect 6775 6272 6858 6378
rect 6892 6272 7095 6378
rect 6775 6265 6815 6272
rect 6858 6265 7095 6272
rect 7325 6378 7442 6385
rect 7485 6378 7645 6385
rect 7325 6272 7408 6378
rect 7442 6272 7645 6378
rect 7325 6265 7365 6272
rect 7408 6265 7645 6272
rect 7875 6378 7992 6385
rect 8035 6378 8195 6385
rect 7875 6272 7958 6378
rect 7992 6272 8195 6378
rect 7875 6265 7915 6272
rect 7958 6265 8195 6272
rect 8425 6378 8542 6385
rect 8585 6378 8745 6385
rect 8425 6272 8508 6378
rect 8542 6272 8745 6378
rect 8425 6265 8465 6272
rect 8508 6265 8745 6272
rect 8975 6378 9092 6385
rect 9135 6378 9295 6385
rect 8975 6272 9058 6378
rect 9092 6272 9295 6378
rect 8975 6265 9015 6272
rect 9058 6265 9295 6272
rect 9525 6378 9642 6385
rect 9685 6378 9845 6385
rect 9525 6272 9608 6378
rect 9642 6272 9845 6378
rect 9525 6265 9565 6272
rect 9608 6265 9845 6272
rect 10075 6378 10192 6385
rect 10235 6378 10395 6385
rect 10075 6272 10158 6378
rect 10192 6272 10395 6378
rect 10075 6265 10115 6272
rect 10158 6265 10395 6272
rect 10625 6378 10742 6385
rect 10785 6378 10945 6385
rect 10625 6272 10708 6378
rect 10742 6272 10945 6378
rect 10625 6265 10665 6272
rect 10708 6265 10945 6272
rect 11175 6378 11292 6385
rect 11335 6378 11495 6385
rect 11175 6272 11258 6378
rect 11292 6272 11495 6378
rect 11175 6265 11215 6272
rect 11258 6265 11495 6272
rect 11725 6378 11842 6385
rect 11885 6378 12045 6385
rect 11725 6272 11808 6378
rect 11842 6272 12045 6378
rect 11725 6265 11765 6272
rect 11808 6265 12045 6272
rect 12275 6378 12392 6385
rect 12435 6378 12595 6385
rect 12275 6272 12358 6378
rect 12392 6272 12595 6378
rect 12275 6265 12315 6272
rect 12358 6265 12595 6272
rect 12825 6378 12942 6385
rect 12985 6378 13145 6385
rect 12825 6272 12908 6378
rect 12942 6272 13145 6378
rect 12825 6265 12865 6272
rect 12908 6265 13145 6272
rect 13375 6378 13492 6385
rect 13535 6378 13695 6385
rect 13375 6272 13458 6378
rect 13492 6272 13695 6378
rect 13375 6265 13415 6272
rect 13458 6265 13695 6272
rect 13925 6378 14042 6385
rect 14085 6378 14245 6385
rect 13925 6272 14008 6378
rect 14042 6272 14245 6378
rect 13925 6265 13965 6272
rect 14008 6265 14245 6272
rect 14475 6378 14592 6385
rect 14635 6378 14795 6385
rect 14475 6272 14558 6378
rect 14592 6272 14795 6378
rect 14475 6265 14515 6272
rect 14558 6265 14795 6272
rect 15025 6378 15142 6385
rect 15185 6378 15345 6385
rect 15025 6272 15108 6378
rect 15142 6272 15345 6378
rect 15025 6265 15065 6272
rect 15108 6265 15345 6272
rect 15575 6378 15692 6385
rect 15735 6378 15895 6385
rect 15575 6272 15658 6378
rect 15692 6272 15895 6378
rect 15575 6265 15615 6272
rect 15658 6265 15895 6272
rect 16125 6378 16242 6385
rect 16285 6378 16445 6385
rect 16125 6272 16208 6378
rect 16242 6272 16445 6378
rect 16125 6265 16165 6272
rect 16208 6265 16445 6272
rect 16675 6378 16792 6385
rect 16835 6378 16995 6385
rect 16675 6272 16758 6378
rect 16792 6272 16995 6378
rect 16675 6265 16715 6272
rect 16758 6265 16995 6272
rect 17225 6378 17342 6385
rect 17385 6378 17545 6385
rect 17225 6272 17308 6378
rect 17342 6272 17545 6378
rect 17225 6265 17265 6272
rect 17308 6265 17545 6272
rect 17775 6378 17892 6385
rect 17935 6378 18095 6385
rect 17775 6272 17858 6378
rect 17892 6272 18095 6378
rect 17775 6265 17815 6272
rect 17858 6265 18095 6272
rect 18325 6378 18442 6385
rect 18485 6378 18645 6385
rect 18325 6272 18408 6378
rect 18442 6272 18645 6378
rect 18325 6265 18365 6272
rect 18408 6265 18645 6272
rect 18875 6378 18992 6385
rect 19035 6378 19195 6385
rect 18875 6272 18958 6378
rect 18992 6272 19195 6378
rect 18875 6265 18915 6272
rect 18958 6265 19195 6272
rect 765 6225 885 6265
rect 1315 6225 1435 6265
rect 1865 6225 1985 6265
rect 2415 6225 2535 6265
rect 2965 6225 3085 6265
rect 3515 6225 3635 6265
rect 4065 6225 4185 6265
rect 4615 6225 4735 6265
rect 5165 6225 5285 6265
rect 5715 6225 5835 6265
rect 6265 6225 6385 6265
rect 6815 6225 6935 6265
rect 7365 6225 7485 6265
rect 7915 6225 8035 6265
rect 8465 6225 8585 6265
rect 9015 6225 9135 6265
rect 9565 6225 9685 6265
rect 10115 6225 10235 6265
rect 10665 6225 10785 6265
rect 11215 6225 11335 6265
rect 11765 6225 11885 6265
rect 12315 6225 12435 6265
rect 12865 6225 12985 6265
rect 13415 6225 13535 6265
rect 13965 6225 14085 6265
rect 14515 6225 14635 6265
rect 15065 6225 15185 6265
rect 15615 6225 15735 6265
rect 16165 6225 16285 6265
rect 16715 6225 16835 6265
rect 17265 6225 17385 6265
rect 17815 6225 17935 6265
rect 18365 6225 18485 6265
rect 18915 6225 19035 6265
rect 19202 6112 19204 6538
rect 500 6025 507 6075
rect 19202 5996 19217 6002
rect 628 5972 885 5995
rect 1178 5972 1435 5995
rect 1728 5972 1985 5995
rect 2278 5972 2535 5995
rect 2828 5972 3085 5995
rect 3378 5972 3635 5995
rect 3928 5972 4185 5995
rect 4478 5972 4735 5995
rect 5028 5972 5285 5995
rect 5578 5972 5835 5995
rect 6128 5972 6385 5995
rect 6678 5972 6935 5995
rect 7228 5972 7485 5995
rect 7778 5972 8035 5995
rect 8328 5972 8585 5995
rect 8878 5972 9135 5995
rect 9428 5972 9685 5995
rect 9978 5972 10235 5995
rect 10528 5972 10785 5995
rect 11078 5972 11335 5995
rect 11628 5972 11885 5995
rect 12178 5972 12435 5995
rect 12728 5972 12985 5995
rect 13278 5972 13535 5995
rect 13828 5972 14085 5995
rect 14378 5972 14635 5995
rect 14928 5972 15185 5995
rect 15478 5972 15735 5995
rect 16028 5972 16285 5995
rect 16578 5972 16835 5995
rect 17128 5972 17385 5995
rect 17678 5972 17935 5995
rect 18228 5972 18485 5995
rect 18778 5972 19035 5995
rect 605 5835 609 5972
rect 784 5875 885 5972
rect 765 5835 885 5875
rect 1155 5835 1159 5972
rect 1334 5875 1435 5972
rect 1315 5835 1435 5875
rect 1705 5835 1709 5972
rect 1884 5875 1985 5972
rect 1865 5835 1985 5875
rect 2255 5835 2259 5972
rect 2434 5875 2535 5972
rect 2415 5835 2535 5875
rect 2805 5835 2809 5972
rect 2984 5875 3085 5972
rect 2965 5835 3085 5875
rect 3355 5835 3359 5972
rect 3534 5875 3635 5972
rect 3515 5835 3635 5875
rect 3905 5835 3909 5972
rect 4084 5875 4185 5972
rect 4065 5835 4185 5875
rect 4455 5835 4459 5972
rect 4634 5875 4735 5972
rect 4615 5835 4735 5875
rect 5005 5835 5009 5972
rect 5184 5875 5285 5972
rect 5165 5835 5285 5875
rect 5555 5835 5559 5972
rect 5734 5875 5835 5972
rect 5715 5835 5835 5875
rect 6105 5835 6109 5972
rect 6284 5875 6385 5972
rect 6265 5835 6385 5875
rect 6655 5835 6659 5972
rect 6834 5875 6935 5972
rect 6815 5835 6935 5875
rect 7205 5835 7209 5972
rect 7384 5875 7485 5972
rect 7365 5835 7485 5875
rect 7755 5835 7759 5972
rect 7934 5875 8035 5972
rect 7915 5835 8035 5875
rect 8305 5835 8309 5972
rect 8484 5875 8585 5972
rect 8465 5835 8585 5875
rect 8855 5835 8859 5972
rect 9034 5875 9135 5972
rect 9015 5835 9135 5875
rect 9405 5835 9409 5972
rect 9584 5875 9685 5972
rect 9565 5835 9685 5875
rect 9955 5835 9959 5972
rect 10134 5875 10235 5972
rect 10115 5835 10235 5875
rect 10505 5835 10509 5972
rect 10684 5875 10785 5972
rect 10665 5835 10785 5875
rect 11055 5835 11059 5972
rect 11234 5875 11335 5972
rect 11215 5835 11335 5875
rect 11605 5835 11609 5972
rect 11784 5875 11885 5972
rect 11765 5835 11885 5875
rect 12155 5835 12159 5972
rect 12334 5875 12435 5972
rect 12315 5835 12435 5875
rect 12705 5835 12709 5972
rect 12884 5875 12985 5972
rect 12865 5835 12985 5875
rect 13255 5835 13259 5972
rect 13434 5875 13535 5972
rect 13415 5835 13535 5875
rect 13805 5835 13809 5972
rect 13984 5875 14085 5972
rect 13965 5835 14085 5875
rect 14355 5835 14359 5972
rect 14534 5875 14635 5972
rect 14515 5835 14635 5875
rect 14905 5835 14909 5972
rect 15084 5875 15185 5972
rect 15065 5835 15185 5875
rect 15455 5835 15459 5972
rect 15634 5875 15735 5972
rect 15615 5835 15735 5875
rect 16005 5835 16009 5972
rect 16184 5875 16285 5972
rect 16165 5835 16285 5875
rect 16555 5835 16559 5972
rect 16734 5875 16835 5972
rect 16715 5835 16835 5875
rect 17105 5835 17109 5972
rect 17284 5875 17385 5972
rect 17265 5835 17385 5875
rect 17655 5835 17659 5972
rect 17834 5875 17935 5972
rect 17815 5835 17935 5875
rect 18205 5835 18209 5972
rect 18384 5875 18485 5972
rect 18365 5835 18485 5875
rect 18755 5835 18759 5972
rect 18934 5875 19035 5972
rect 18915 5835 19035 5875
rect 725 5828 842 5835
rect 885 5828 1045 5835
rect 725 5722 808 5828
rect 842 5722 1045 5828
rect 725 5715 765 5722
rect 808 5715 1045 5722
rect 1275 5828 1392 5835
rect 1435 5828 1595 5835
rect 1275 5722 1358 5828
rect 1392 5722 1595 5828
rect 1275 5715 1315 5722
rect 1358 5715 1595 5722
rect 1825 5828 1942 5835
rect 1985 5828 2145 5835
rect 1825 5722 1908 5828
rect 1942 5722 2145 5828
rect 1825 5715 1865 5722
rect 1908 5715 2145 5722
rect 2375 5828 2492 5835
rect 2535 5828 2695 5835
rect 2375 5722 2458 5828
rect 2492 5722 2695 5828
rect 2375 5715 2415 5722
rect 2458 5715 2695 5722
rect 2925 5828 3042 5835
rect 3085 5828 3245 5835
rect 2925 5722 3008 5828
rect 3042 5722 3245 5828
rect 2925 5715 2965 5722
rect 3008 5715 3245 5722
rect 3475 5828 3592 5835
rect 3635 5828 3795 5835
rect 3475 5722 3558 5828
rect 3592 5722 3795 5828
rect 3475 5715 3515 5722
rect 3558 5715 3795 5722
rect 4025 5828 4142 5835
rect 4185 5828 4345 5835
rect 4025 5722 4108 5828
rect 4142 5722 4345 5828
rect 4025 5715 4065 5722
rect 4108 5715 4345 5722
rect 4575 5828 4692 5835
rect 4735 5828 4895 5835
rect 4575 5722 4658 5828
rect 4692 5722 4895 5828
rect 4575 5715 4615 5722
rect 4658 5715 4895 5722
rect 5125 5828 5242 5835
rect 5285 5828 5445 5835
rect 5125 5722 5208 5828
rect 5242 5722 5445 5828
rect 5125 5715 5165 5722
rect 5208 5715 5445 5722
rect 5675 5828 5792 5835
rect 5835 5828 5995 5835
rect 5675 5722 5758 5828
rect 5792 5722 5995 5828
rect 5675 5715 5715 5722
rect 5758 5715 5995 5722
rect 6225 5828 6342 5835
rect 6385 5828 6545 5835
rect 6225 5722 6308 5828
rect 6342 5722 6545 5828
rect 6225 5715 6265 5722
rect 6308 5715 6545 5722
rect 6775 5828 6892 5835
rect 6935 5828 7095 5835
rect 6775 5722 6858 5828
rect 6892 5722 7095 5828
rect 6775 5715 6815 5722
rect 6858 5715 7095 5722
rect 7325 5828 7442 5835
rect 7485 5828 7645 5835
rect 7325 5722 7408 5828
rect 7442 5722 7645 5828
rect 7325 5715 7365 5722
rect 7408 5715 7645 5722
rect 7875 5828 7992 5835
rect 8035 5828 8195 5835
rect 7875 5722 7958 5828
rect 7992 5722 8195 5828
rect 7875 5715 7915 5722
rect 7958 5715 8195 5722
rect 8425 5828 8542 5835
rect 8585 5828 8745 5835
rect 8425 5722 8508 5828
rect 8542 5722 8745 5828
rect 8425 5715 8465 5722
rect 8508 5715 8745 5722
rect 8975 5828 9092 5835
rect 9135 5828 9295 5835
rect 8975 5722 9058 5828
rect 9092 5722 9295 5828
rect 8975 5715 9015 5722
rect 9058 5715 9295 5722
rect 9525 5828 9642 5835
rect 9685 5828 9845 5835
rect 9525 5722 9608 5828
rect 9642 5722 9845 5828
rect 9525 5715 9565 5722
rect 9608 5715 9845 5722
rect 10075 5828 10192 5835
rect 10235 5828 10395 5835
rect 10075 5722 10158 5828
rect 10192 5722 10395 5828
rect 10075 5715 10115 5722
rect 10158 5715 10395 5722
rect 10625 5828 10742 5835
rect 10785 5828 10945 5835
rect 10625 5722 10708 5828
rect 10742 5722 10945 5828
rect 10625 5715 10665 5722
rect 10708 5715 10945 5722
rect 11175 5828 11292 5835
rect 11335 5828 11495 5835
rect 11175 5722 11258 5828
rect 11292 5722 11495 5828
rect 11175 5715 11215 5722
rect 11258 5715 11495 5722
rect 11725 5828 11842 5835
rect 11885 5828 12045 5835
rect 11725 5722 11808 5828
rect 11842 5722 12045 5828
rect 11725 5715 11765 5722
rect 11808 5715 12045 5722
rect 12275 5828 12392 5835
rect 12435 5828 12595 5835
rect 12275 5722 12358 5828
rect 12392 5722 12595 5828
rect 12275 5715 12315 5722
rect 12358 5715 12595 5722
rect 12825 5828 12942 5835
rect 12985 5828 13145 5835
rect 12825 5722 12908 5828
rect 12942 5722 13145 5828
rect 12825 5715 12865 5722
rect 12908 5715 13145 5722
rect 13375 5828 13492 5835
rect 13535 5828 13695 5835
rect 13375 5722 13458 5828
rect 13492 5722 13695 5828
rect 13375 5715 13415 5722
rect 13458 5715 13695 5722
rect 13925 5828 14042 5835
rect 14085 5828 14245 5835
rect 13925 5722 14008 5828
rect 14042 5722 14245 5828
rect 13925 5715 13965 5722
rect 14008 5715 14245 5722
rect 14475 5828 14592 5835
rect 14635 5828 14795 5835
rect 14475 5722 14558 5828
rect 14592 5722 14795 5828
rect 14475 5715 14515 5722
rect 14558 5715 14795 5722
rect 15025 5828 15142 5835
rect 15185 5828 15345 5835
rect 15025 5722 15108 5828
rect 15142 5722 15345 5828
rect 15025 5715 15065 5722
rect 15108 5715 15345 5722
rect 15575 5828 15692 5835
rect 15735 5828 15895 5835
rect 15575 5722 15658 5828
rect 15692 5722 15895 5828
rect 15575 5715 15615 5722
rect 15658 5715 15895 5722
rect 16125 5828 16242 5835
rect 16285 5828 16445 5835
rect 16125 5722 16208 5828
rect 16242 5722 16445 5828
rect 16125 5715 16165 5722
rect 16208 5715 16445 5722
rect 16675 5828 16792 5835
rect 16835 5828 16995 5835
rect 16675 5722 16758 5828
rect 16792 5722 16995 5828
rect 16675 5715 16715 5722
rect 16758 5715 16995 5722
rect 17225 5828 17342 5835
rect 17385 5828 17545 5835
rect 17225 5722 17308 5828
rect 17342 5722 17545 5828
rect 17225 5715 17265 5722
rect 17308 5715 17545 5722
rect 17775 5828 17892 5835
rect 17935 5828 18095 5835
rect 17775 5722 17858 5828
rect 17892 5722 18095 5828
rect 17775 5715 17815 5722
rect 17858 5715 18095 5722
rect 18325 5828 18442 5835
rect 18485 5828 18645 5835
rect 18325 5722 18408 5828
rect 18442 5722 18645 5828
rect 18325 5715 18365 5722
rect 18408 5715 18645 5722
rect 18875 5828 18992 5835
rect 19035 5828 19195 5835
rect 18875 5722 18958 5828
rect 18992 5722 19195 5828
rect 18875 5715 18915 5722
rect 18958 5715 19195 5722
rect 765 5675 885 5715
rect 1315 5675 1435 5715
rect 1865 5675 1985 5715
rect 2415 5675 2535 5715
rect 2965 5675 3085 5715
rect 3515 5675 3635 5715
rect 4065 5675 4185 5715
rect 4615 5675 4735 5715
rect 5165 5675 5285 5715
rect 5715 5675 5835 5715
rect 6265 5675 6385 5715
rect 6815 5675 6935 5715
rect 7365 5675 7485 5715
rect 7915 5675 8035 5715
rect 8465 5675 8585 5715
rect 9015 5675 9135 5715
rect 9565 5675 9685 5715
rect 10115 5675 10235 5715
rect 10665 5675 10785 5715
rect 11215 5675 11335 5715
rect 11765 5675 11885 5715
rect 12315 5675 12435 5715
rect 12865 5675 12985 5715
rect 13415 5675 13535 5715
rect 13965 5675 14085 5715
rect 14515 5675 14635 5715
rect 15065 5675 15185 5715
rect 15615 5675 15735 5715
rect 16165 5675 16285 5715
rect 16715 5675 16835 5715
rect 17265 5675 17385 5715
rect 17815 5675 17935 5715
rect 18365 5675 18485 5715
rect 18915 5675 19035 5715
rect 19185 5554 19200 5571
rect 19202 5562 19204 5988
rect 19202 5548 19217 5554
rect 500 5475 507 5525
rect 500 5039 525 5440
rect 628 5422 885 5445
rect 1178 5422 1435 5445
rect 1728 5422 1985 5445
rect 2278 5422 2535 5445
rect 2828 5422 3085 5445
rect 3378 5422 3635 5445
rect 3928 5422 4185 5445
rect 4478 5422 4735 5445
rect 5028 5422 5285 5445
rect 5578 5422 5835 5445
rect 6128 5422 6385 5445
rect 6678 5422 6935 5445
rect 7228 5422 7485 5445
rect 7778 5422 8035 5445
rect 8328 5422 8585 5445
rect 8878 5422 9135 5445
rect 9428 5422 9685 5445
rect 9978 5422 10235 5445
rect 10528 5422 10785 5445
rect 11078 5422 11335 5445
rect 11628 5422 11885 5445
rect 12178 5422 12435 5445
rect 12728 5422 12985 5445
rect 13278 5422 13535 5445
rect 13828 5422 14085 5445
rect 14378 5422 14635 5445
rect 14928 5422 15185 5445
rect 15478 5422 15735 5445
rect 16028 5422 16285 5445
rect 16578 5422 16835 5445
rect 17128 5422 17385 5445
rect 17678 5422 17935 5445
rect 18228 5422 18485 5445
rect 18778 5422 19035 5445
rect 605 5285 609 5422
rect 784 5325 885 5422
rect 765 5285 885 5325
rect 1155 5285 1159 5422
rect 1334 5325 1435 5422
rect 1315 5285 1435 5325
rect 1705 5285 1709 5422
rect 1884 5325 1985 5422
rect 1865 5285 1985 5325
rect 2255 5285 2259 5422
rect 2434 5325 2535 5422
rect 2415 5285 2535 5325
rect 2805 5285 2809 5422
rect 2984 5325 3085 5422
rect 2965 5285 3085 5325
rect 3355 5285 3359 5422
rect 3534 5325 3635 5422
rect 3515 5285 3635 5325
rect 3905 5285 3909 5422
rect 4084 5325 4185 5422
rect 4065 5285 4185 5325
rect 4455 5285 4459 5422
rect 4634 5325 4735 5422
rect 4615 5285 4735 5325
rect 5005 5285 5009 5422
rect 5184 5325 5285 5422
rect 5165 5285 5285 5325
rect 5555 5285 5559 5422
rect 5734 5325 5835 5422
rect 5715 5285 5835 5325
rect 6105 5285 6109 5422
rect 6284 5325 6385 5422
rect 6265 5285 6385 5325
rect 6655 5285 6659 5422
rect 6834 5325 6935 5422
rect 6815 5285 6935 5325
rect 7205 5285 7209 5422
rect 7384 5325 7485 5422
rect 7365 5285 7485 5325
rect 7755 5285 7759 5422
rect 7934 5325 8035 5422
rect 7915 5285 8035 5325
rect 8305 5285 8309 5422
rect 8484 5325 8585 5422
rect 8465 5285 8585 5325
rect 8855 5285 8859 5422
rect 9034 5325 9135 5422
rect 9015 5285 9135 5325
rect 9405 5285 9409 5422
rect 9584 5325 9685 5422
rect 9565 5285 9685 5325
rect 9955 5285 9959 5422
rect 10134 5325 10235 5422
rect 10115 5285 10235 5325
rect 10505 5285 10509 5422
rect 10684 5325 10785 5422
rect 10665 5285 10785 5325
rect 11055 5285 11059 5422
rect 11234 5325 11335 5422
rect 11215 5285 11335 5325
rect 11605 5285 11609 5422
rect 11784 5325 11885 5422
rect 11765 5285 11885 5325
rect 12155 5285 12159 5422
rect 12334 5325 12435 5422
rect 12315 5285 12435 5325
rect 12705 5285 12709 5422
rect 12884 5325 12985 5422
rect 12865 5285 12985 5325
rect 13255 5285 13259 5422
rect 13434 5325 13535 5422
rect 13415 5285 13535 5325
rect 13805 5285 13809 5422
rect 13984 5325 14085 5422
rect 13965 5285 14085 5325
rect 14355 5285 14359 5422
rect 14534 5325 14635 5422
rect 14515 5285 14635 5325
rect 14905 5285 14909 5422
rect 15084 5325 15185 5422
rect 15065 5285 15185 5325
rect 15455 5285 15459 5422
rect 15634 5325 15735 5422
rect 15615 5285 15735 5325
rect 16005 5285 16009 5422
rect 16184 5325 16285 5422
rect 16165 5285 16285 5325
rect 16555 5285 16559 5422
rect 16734 5325 16835 5422
rect 16715 5285 16835 5325
rect 17105 5285 17109 5422
rect 17284 5325 17385 5422
rect 17265 5285 17385 5325
rect 17655 5285 17659 5422
rect 17834 5325 17935 5422
rect 17815 5285 17935 5325
rect 18205 5285 18209 5422
rect 18384 5325 18485 5422
rect 18365 5285 18485 5325
rect 18755 5285 18759 5422
rect 18934 5325 19035 5422
rect 18915 5285 19035 5325
rect 725 5278 842 5285
rect 885 5278 1045 5285
rect 725 5172 808 5278
rect 842 5172 1045 5278
rect 725 5165 765 5172
rect 808 5165 1045 5172
rect 1275 5278 1392 5285
rect 1435 5278 1595 5285
rect 1275 5172 1358 5278
rect 1392 5172 1595 5278
rect 1275 5165 1315 5172
rect 1358 5165 1595 5172
rect 1825 5278 1942 5285
rect 1985 5278 2145 5285
rect 1825 5172 1908 5278
rect 1942 5172 2145 5278
rect 1825 5165 1865 5172
rect 1908 5165 2145 5172
rect 2375 5278 2492 5285
rect 2535 5278 2695 5285
rect 2375 5172 2458 5278
rect 2492 5172 2695 5278
rect 2375 5165 2415 5172
rect 2458 5165 2695 5172
rect 2925 5278 3042 5285
rect 3085 5278 3245 5285
rect 2925 5172 3008 5278
rect 3042 5172 3245 5278
rect 2925 5165 2965 5172
rect 3008 5165 3245 5172
rect 3475 5278 3592 5285
rect 3635 5278 3795 5285
rect 3475 5172 3558 5278
rect 3592 5172 3795 5278
rect 3475 5165 3515 5172
rect 3558 5165 3795 5172
rect 4025 5278 4142 5285
rect 4185 5278 4345 5285
rect 4025 5172 4108 5278
rect 4142 5172 4345 5278
rect 4025 5165 4065 5172
rect 4108 5165 4345 5172
rect 4575 5278 4692 5285
rect 4735 5278 4895 5285
rect 4575 5172 4658 5278
rect 4692 5172 4895 5278
rect 4575 5165 4615 5172
rect 4658 5165 4895 5172
rect 5125 5278 5242 5285
rect 5285 5278 5445 5285
rect 5125 5172 5208 5278
rect 5242 5172 5445 5278
rect 5125 5165 5165 5172
rect 5208 5165 5445 5172
rect 5675 5278 5792 5285
rect 5835 5278 5995 5285
rect 5675 5172 5758 5278
rect 5792 5172 5995 5278
rect 5675 5165 5715 5172
rect 5758 5165 5995 5172
rect 6225 5278 6342 5285
rect 6385 5278 6545 5285
rect 6225 5172 6308 5278
rect 6342 5172 6545 5278
rect 6225 5165 6265 5172
rect 6308 5165 6545 5172
rect 6775 5278 6892 5285
rect 6935 5278 7095 5285
rect 6775 5172 6858 5278
rect 6892 5172 7095 5278
rect 6775 5165 6815 5172
rect 6858 5165 7095 5172
rect 7325 5278 7442 5285
rect 7485 5278 7645 5285
rect 7325 5172 7408 5278
rect 7442 5172 7645 5278
rect 7325 5165 7365 5172
rect 7408 5165 7645 5172
rect 7875 5278 7992 5285
rect 8035 5278 8195 5285
rect 7875 5172 7958 5278
rect 7992 5172 8195 5278
rect 7875 5165 7915 5172
rect 7958 5165 8195 5172
rect 8425 5278 8542 5285
rect 8585 5278 8745 5285
rect 8425 5172 8508 5278
rect 8542 5172 8745 5278
rect 8425 5165 8465 5172
rect 8508 5165 8745 5172
rect 8975 5278 9092 5285
rect 9135 5278 9295 5285
rect 8975 5172 9058 5278
rect 9092 5172 9295 5278
rect 8975 5165 9015 5172
rect 9058 5165 9295 5172
rect 9525 5278 9642 5285
rect 9685 5278 9845 5285
rect 9525 5172 9608 5278
rect 9642 5172 9845 5278
rect 9525 5165 9565 5172
rect 9608 5165 9845 5172
rect 10075 5278 10192 5285
rect 10235 5278 10395 5285
rect 10075 5172 10158 5278
rect 10192 5172 10395 5278
rect 10075 5165 10115 5172
rect 10158 5165 10395 5172
rect 10625 5278 10742 5285
rect 10785 5278 10945 5285
rect 10625 5172 10708 5278
rect 10742 5172 10945 5278
rect 10625 5165 10665 5172
rect 10708 5165 10945 5172
rect 11175 5278 11292 5285
rect 11335 5278 11495 5285
rect 11175 5172 11258 5278
rect 11292 5172 11495 5278
rect 11175 5165 11215 5172
rect 11258 5165 11495 5172
rect 11725 5278 11842 5285
rect 11885 5278 12045 5285
rect 11725 5172 11808 5278
rect 11842 5172 12045 5278
rect 11725 5165 11765 5172
rect 11808 5165 12045 5172
rect 12275 5278 12392 5285
rect 12435 5278 12595 5285
rect 12275 5172 12358 5278
rect 12392 5172 12595 5278
rect 12275 5165 12315 5172
rect 12358 5165 12595 5172
rect 12825 5278 12942 5285
rect 12985 5278 13145 5285
rect 12825 5172 12908 5278
rect 12942 5172 13145 5278
rect 12825 5165 12865 5172
rect 12908 5165 13145 5172
rect 13375 5278 13492 5285
rect 13535 5278 13695 5285
rect 13375 5172 13458 5278
rect 13492 5172 13695 5278
rect 13375 5165 13415 5172
rect 13458 5165 13695 5172
rect 13925 5278 14042 5285
rect 14085 5278 14245 5285
rect 13925 5172 14008 5278
rect 14042 5172 14245 5278
rect 13925 5165 13965 5172
rect 14008 5165 14245 5172
rect 14475 5278 14592 5285
rect 14635 5278 14795 5285
rect 14475 5172 14558 5278
rect 14592 5172 14795 5278
rect 14475 5165 14515 5172
rect 14558 5165 14795 5172
rect 15025 5278 15142 5285
rect 15185 5278 15345 5285
rect 15025 5172 15108 5278
rect 15142 5172 15345 5278
rect 15025 5165 15065 5172
rect 15108 5165 15345 5172
rect 15575 5278 15692 5285
rect 15735 5278 15895 5285
rect 15575 5172 15658 5278
rect 15692 5172 15895 5278
rect 15575 5165 15615 5172
rect 15658 5165 15895 5172
rect 16125 5278 16242 5285
rect 16285 5278 16445 5285
rect 16125 5172 16208 5278
rect 16242 5172 16445 5278
rect 16125 5165 16165 5172
rect 16208 5165 16445 5172
rect 16675 5278 16792 5285
rect 16835 5278 16995 5285
rect 16675 5172 16758 5278
rect 16792 5172 16995 5278
rect 16675 5165 16715 5172
rect 16758 5165 16995 5172
rect 17225 5278 17342 5285
rect 17385 5278 17545 5285
rect 17225 5172 17308 5278
rect 17342 5172 17545 5278
rect 17225 5165 17265 5172
rect 17308 5165 17545 5172
rect 17775 5278 17892 5285
rect 17935 5278 18095 5285
rect 17775 5172 17858 5278
rect 17892 5172 18095 5278
rect 17775 5165 17815 5172
rect 17858 5165 18095 5172
rect 18325 5278 18442 5285
rect 18485 5278 18645 5285
rect 18325 5172 18408 5278
rect 18442 5172 18645 5278
rect 18325 5165 18365 5172
rect 18408 5165 18645 5172
rect 18875 5278 18992 5285
rect 19035 5278 19195 5285
rect 18875 5172 18958 5278
rect 18992 5172 19195 5278
rect 18875 5165 18915 5172
rect 18958 5165 19195 5172
rect 765 5125 885 5165
rect 1315 5125 1435 5165
rect 1865 5125 1985 5165
rect 2415 5125 2535 5165
rect 2965 5125 3085 5165
rect 3515 5125 3635 5165
rect 4065 5125 4185 5165
rect 4615 5125 4735 5165
rect 5165 5125 5285 5165
rect 5715 5125 5835 5165
rect 6265 5125 6385 5165
rect 6815 5125 6935 5165
rect 7365 5125 7485 5165
rect 7915 5125 8035 5165
rect 8465 5125 8585 5165
rect 9015 5125 9135 5165
rect 9565 5125 9685 5165
rect 10115 5125 10235 5165
rect 10665 5125 10785 5165
rect 11215 5125 11335 5165
rect 11765 5125 11885 5165
rect 12315 5125 12435 5165
rect 12865 5125 12985 5165
rect 13415 5125 13535 5165
rect 13965 5125 14085 5165
rect 14515 5125 14635 5165
rect 15065 5125 15185 5165
rect 15615 5125 15735 5165
rect 16165 5125 16285 5165
rect 16715 5125 16835 5165
rect 17265 5125 17385 5165
rect 17815 5125 17935 5165
rect 18365 5125 18485 5165
rect 18915 5125 19035 5165
rect 19202 5012 19204 5438
rect 500 4925 507 4975
rect 19202 4896 19217 4902
rect 628 4872 885 4895
rect 1178 4872 1435 4895
rect 1728 4872 1985 4895
rect 2278 4872 2535 4895
rect 2828 4872 3085 4895
rect 3378 4872 3635 4895
rect 3928 4872 4185 4895
rect 4478 4872 4735 4895
rect 5028 4872 5285 4895
rect 5578 4872 5835 4895
rect 6128 4872 6385 4895
rect 6678 4872 6935 4895
rect 7228 4872 7485 4895
rect 7778 4872 8035 4895
rect 8328 4872 8585 4895
rect 8878 4872 9135 4895
rect 9428 4872 9685 4895
rect 9978 4872 10235 4895
rect 10528 4872 10785 4895
rect 11078 4872 11335 4895
rect 11628 4872 11885 4895
rect 12178 4872 12435 4895
rect 12728 4872 12985 4895
rect 13278 4872 13535 4895
rect 13828 4872 14085 4895
rect 14378 4872 14635 4895
rect 14928 4872 15185 4895
rect 15478 4872 15735 4895
rect 16028 4872 16285 4895
rect 16578 4872 16835 4895
rect 17128 4872 17385 4895
rect 17678 4872 17935 4895
rect 18228 4872 18485 4895
rect 18778 4872 19035 4895
rect 605 4735 609 4872
rect 784 4775 885 4872
rect 765 4735 885 4775
rect 1155 4735 1159 4872
rect 1334 4775 1435 4872
rect 1315 4735 1435 4775
rect 1705 4735 1709 4872
rect 1884 4775 1985 4872
rect 1865 4735 1985 4775
rect 2255 4735 2259 4872
rect 2434 4775 2535 4872
rect 2415 4735 2535 4775
rect 2805 4735 2809 4872
rect 2984 4775 3085 4872
rect 2965 4735 3085 4775
rect 3355 4735 3359 4872
rect 3534 4775 3635 4872
rect 3515 4735 3635 4775
rect 3905 4735 3909 4872
rect 4084 4775 4185 4872
rect 4065 4735 4185 4775
rect 4455 4735 4459 4872
rect 4634 4775 4735 4872
rect 4615 4735 4735 4775
rect 5005 4735 5009 4872
rect 5184 4775 5285 4872
rect 5165 4735 5285 4775
rect 5555 4735 5559 4872
rect 5734 4775 5835 4872
rect 5715 4735 5835 4775
rect 6105 4735 6109 4872
rect 6284 4775 6385 4872
rect 6265 4735 6385 4775
rect 6655 4735 6659 4872
rect 6834 4775 6935 4872
rect 6815 4735 6935 4775
rect 7205 4735 7209 4872
rect 7384 4775 7485 4872
rect 7365 4735 7485 4775
rect 7755 4735 7759 4872
rect 7934 4775 8035 4872
rect 7915 4735 8035 4775
rect 8305 4735 8309 4872
rect 8484 4775 8585 4872
rect 8465 4735 8585 4775
rect 8855 4735 8859 4872
rect 9034 4775 9135 4872
rect 9015 4735 9135 4775
rect 9405 4735 9409 4872
rect 9584 4775 9685 4872
rect 9565 4735 9685 4775
rect 9955 4735 9959 4872
rect 10134 4775 10235 4872
rect 10115 4735 10235 4775
rect 10505 4735 10509 4872
rect 10684 4775 10785 4872
rect 10665 4735 10785 4775
rect 11055 4735 11059 4872
rect 11234 4775 11335 4872
rect 11215 4735 11335 4775
rect 11605 4735 11609 4872
rect 11784 4775 11885 4872
rect 11765 4735 11885 4775
rect 12155 4735 12159 4872
rect 12334 4775 12435 4872
rect 12315 4735 12435 4775
rect 12705 4735 12709 4872
rect 12884 4775 12985 4872
rect 12865 4735 12985 4775
rect 13255 4735 13259 4872
rect 13434 4775 13535 4872
rect 13415 4735 13535 4775
rect 13805 4735 13809 4872
rect 13984 4775 14085 4872
rect 13965 4735 14085 4775
rect 14355 4735 14359 4872
rect 14534 4775 14635 4872
rect 14515 4735 14635 4775
rect 14905 4735 14909 4872
rect 15084 4775 15185 4872
rect 15065 4735 15185 4775
rect 15455 4735 15459 4872
rect 15634 4775 15735 4872
rect 15615 4735 15735 4775
rect 16005 4735 16009 4872
rect 16184 4775 16285 4872
rect 16165 4735 16285 4775
rect 16555 4735 16559 4872
rect 16734 4775 16835 4872
rect 16715 4735 16835 4775
rect 17105 4735 17109 4872
rect 17284 4775 17385 4872
rect 17265 4735 17385 4775
rect 17655 4735 17659 4872
rect 17834 4775 17935 4872
rect 17815 4735 17935 4775
rect 18205 4735 18209 4872
rect 18384 4775 18485 4872
rect 18365 4735 18485 4775
rect 18755 4735 18759 4872
rect 18934 4775 19035 4872
rect 18915 4735 19035 4775
rect 725 4728 842 4735
rect 885 4728 1045 4735
rect 725 4622 808 4728
rect 842 4622 1045 4728
rect 725 4615 765 4622
rect 808 4615 1045 4622
rect 1275 4728 1392 4735
rect 1435 4728 1595 4735
rect 1275 4622 1358 4728
rect 1392 4622 1595 4728
rect 1275 4615 1315 4622
rect 1358 4615 1595 4622
rect 1825 4728 1942 4735
rect 1985 4728 2145 4735
rect 1825 4622 1908 4728
rect 1942 4622 2145 4728
rect 1825 4615 1865 4622
rect 1908 4615 2145 4622
rect 2375 4728 2492 4735
rect 2535 4728 2695 4735
rect 2375 4622 2458 4728
rect 2492 4622 2695 4728
rect 2375 4615 2415 4622
rect 2458 4615 2695 4622
rect 2925 4728 3042 4735
rect 3085 4728 3245 4735
rect 2925 4622 3008 4728
rect 3042 4622 3245 4728
rect 2925 4615 2965 4622
rect 3008 4615 3245 4622
rect 3475 4728 3592 4735
rect 3635 4728 3795 4735
rect 3475 4622 3558 4728
rect 3592 4622 3795 4728
rect 3475 4615 3515 4622
rect 3558 4615 3795 4622
rect 4025 4728 4142 4735
rect 4185 4728 4345 4735
rect 4025 4622 4108 4728
rect 4142 4622 4345 4728
rect 4025 4615 4065 4622
rect 4108 4615 4345 4622
rect 4575 4728 4692 4735
rect 4735 4728 4895 4735
rect 4575 4622 4658 4728
rect 4692 4622 4895 4728
rect 4575 4615 4615 4622
rect 4658 4615 4895 4622
rect 5125 4728 5242 4735
rect 5285 4728 5445 4735
rect 5125 4622 5208 4728
rect 5242 4622 5445 4728
rect 5125 4615 5165 4622
rect 5208 4615 5445 4622
rect 5675 4728 5792 4735
rect 5835 4728 5995 4735
rect 5675 4622 5758 4728
rect 5792 4622 5995 4728
rect 5675 4615 5715 4622
rect 5758 4615 5995 4622
rect 6225 4728 6342 4735
rect 6385 4728 6545 4735
rect 6225 4622 6308 4728
rect 6342 4622 6545 4728
rect 6225 4615 6265 4622
rect 6308 4615 6545 4622
rect 6775 4728 6892 4735
rect 6935 4728 7095 4735
rect 6775 4622 6858 4728
rect 6892 4622 7095 4728
rect 6775 4615 6815 4622
rect 6858 4615 7095 4622
rect 7325 4728 7442 4735
rect 7485 4728 7645 4735
rect 7325 4622 7408 4728
rect 7442 4622 7645 4728
rect 7325 4615 7365 4622
rect 7408 4615 7645 4622
rect 7875 4728 7992 4735
rect 8035 4728 8195 4735
rect 7875 4622 7958 4728
rect 7992 4622 8195 4728
rect 7875 4615 7915 4622
rect 7958 4615 8195 4622
rect 8425 4728 8542 4735
rect 8585 4728 8745 4735
rect 8425 4622 8508 4728
rect 8542 4622 8745 4728
rect 8425 4615 8465 4622
rect 8508 4615 8745 4622
rect 8975 4728 9092 4735
rect 9135 4728 9295 4735
rect 8975 4622 9058 4728
rect 9092 4622 9295 4728
rect 8975 4615 9015 4622
rect 9058 4615 9295 4622
rect 9525 4728 9642 4735
rect 9685 4728 9845 4735
rect 9525 4622 9608 4728
rect 9642 4622 9845 4728
rect 9525 4615 9565 4622
rect 9608 4615 9845 4622
rect 10075 4728 10192 4735
rect 10235 4728 10395 4735
rect 10075 4622 10158 4728
rect 10192 4622 10395 4728
rect 10075 4615 10115 4622
rect 10158 4615 10395 4622
rect 10625 4728 10742 4735
rect 10785 4728 10945 4735
rect 10625 4622 10708 4728
rect 10742 4622 10945 4728
rect 10625 4615 10665 4622
rect 10708 4615 10945 4622
rect 11175 4728 11292 4735
rect 11335 4728 11495 4735
rect 11175 4622 11258 4728
rect 11292 4622 11495 4728
rect 11175 4615 11215 4622
rect 11258 4615 11495 4622
rect 11725 4728 11842 4735
rect 11885 4728 12045 4735
rect 11725 4622 11808 4728
rect 11842 4622 12045 4728
rect 11725 4615 11765 4622
rect 11808 4615 12045 4622
rect 12275 4728 12392 4735
rect 12435 4728 12595 4735
rect 12275 4622 12358 4728
rect 12392 4622 12595 4728
rect 12275 4615 12315 4622
rect 12358 4615 12595 4622
rect 12825 4728 12942 4735
rect 12985 4728 13145 4735
rect 12825 4622 12908 4728
rect 12942 4622 13145 4728
rect 12825 4615 12865 4622
rect 12908 4615 13145 4622
rect 13375 4728 13492 4735
rect 13535 4728 13695 4735
rect 13375 4622 13458 4728
rect 13492 4622 13695 4728
rect 13375 4615 13415 4622
rect 13458 4615 13695 4622
rect 13925 4728 14042 4735
rect 14085 4728 14245 4735
rect 13925 4622 14008 4728
rect 14042 4622 14245 4728
rect 13925 4615 13965 4622
rect 14008 4615 14245 4622
rect 14475 4728 14592 4735
rect 14635 4728 14795 4735
rect 14475 4622 14558 4728
rect 14592 4622 14795 4728
rect 14475 4615 14515 4622
rect 14558 4615 14795 4622
rect 15025 4728 15142 4735
rect 15185 4728 15345 4735
rect 15025 4622 15108 4728
rect 15142 4622 15345 4728
rect 15025 4615 15065 4622
rect 15108 4615 15345 4622
rect 15575 4728 15692 4735
rect 15735 4728 15895 4735
rect 15575 4622 15658 4728
rect 15692 4622 15895 4728
rect 15575 4615 15615 4622
rect 15658 4615 15895 4622
rect 16125 4728 16242 4735
rect 16285 4728 16445 4735
rect 16125 4622 16208 4728
rect 16242 4622 16445 4728
rect 16125 4615 16165 4622
rect 16208 4615 16445 4622
rect 16675 4728 16792 4735
rect 16835 4728 16995 4735
rect 16675 4622 16758 4728
rect 16792 4622 16995 4728
rect 16675 4615 16715 4622
rect 16758 4615 16995 4622
rect 17225 4728 17342 4735
rect 17385 4728 17545 4735
rect 17225 4622 17308 4728
rect 17342 4622 17545 4728
rect 17225 4615 17265 4622
rect 17308 4615 17545 4622
rect 17775 4728 17892 4735
rect 17935 4728 18095 4735
rect 17775 4622 17858 4728
rect 17892 4622 18095 4728
rect 17775 4615 17815 4622
rect 17858 4615 18095 4622
rect 18325 4728 18442 4735
rect 18485 4728 18645 4735
rect 18325 4622 18408 4728
rect 18442 4622 18645 4728
rect 18325 4615 18365 4622
rect 18408 4615 18645 4622
rect 18875 4728 18992 4735
rect 19035 4728 19195 4735
rect 18875 4622 18958 4728
rect 18992 4622 19195 4728
rect 18875 4615 18915 4622
rect 18958 4615 19195 4622
rect 765 4575 885 4615
rect 1315 4575 1435 4615
rect 1865 4575 1985 4615
rect 2415 4575 2535 4615
rect 2965 4575 3085 4615
rect 3515 4575 3635 4615
rect 4065 4575 4185 4615
rect 4615 4575 4735 4615
rect 5165 4575 5285 4615
rect 5715 4575 5835 4615
rect 6265 4575 6385 4615
rect 6815 4575 6935 4615
rect 7365 4575 7485 4615
rect 7915 4575 8035 4615
rect 8465 4575 8585 4615
rect 9015 4575 9135 4615
rect 9565 4575 9685 4615
rect 10115 4575 10235 4615
rect 10665 4575 10785 4615
rect 11215 4575 11335 4615
rect 11765 4575 11885 4615
rect 12315 4575 12435 4615
rect 12865 4575 12985 4615
rect 13415 4575 13535 4615
rect 13965 4575 14085 4615
rect 14515 4575 14635 4615
rect 15065 4575 15185 4615
rect 15615 4575 15735 4615
rect 16165 4575 16285 4615
rect 16715 4575 16835 4615
rect 17265 4575 17385 4615
rect 17815 4575 17935 4615
rect 18365 4575 18485 4615
rect 18915 4575 19035 4615
rect 19185 4454 19200 4471
rect 19202 4462 19204 4888
rect 19202 4448 19217 4454
rect 500 4375 507 4425
rect 500 3939 525 4340
rect 628 4322 885 4345
rect 1178 4322 1435 4345
rect 1728 4322 1985 4345
rect 2278 4322 2535 4345
rect 2828 4322 3085 4345
rect 3378 4322 3635 4345
rect 3928 4322 4185 4345
rect 4478 4322 4735 4345
rect 5028 4322 5285 4345
rect 5578 4322 5835 4345
rect 6128 4322 6385 4345
rect 6678 4322 6935 4345
rect 7228 4322 7485 4345
rect 7778 4322 8035 4345
rect 8328 4322 8585 4345
rect 8878 4322 9135 4345
rect 9428 4322 9685 4345
rect 9978 4322 10235 4345
rect 10528 4322 10785 4345
rect 11078 4322 11335 4345
rect 11628 4322 11885 4345
rect 12178 4322 12435 4345
rect 12728 4322 12985 4345
rect 13278 4322 13535 4345
rect 13828 4322 14085 4345
rect 14378 4322 14635 4345
rect 14928 4322 15185 4345
rect 15478 4322 15735 4345
rect 16028 4322 16285 4345
rect 16578 4322 16835 4345
rect 17128 4322 17385 4345
rect 17678 4322 17935 4345
rect 18228 4322 18485 4345
rect 18778 4322 19035 4345
rect 605 4185 609 4322
rect 784 4225 885 4322
rect 765 4185 885 4225
rect 1155 4185 1159 4322
rect 1334 4225 1435 4322
rect 1315 4185 1435 4225
rect 1705 4185 1709 4322
rect 1884 4225 1985 4322
rect 1865 4185 1985 4225
rect 2255 4185 2259 4322
rect 2434 4225 2535 4322
rect 2415 4185 2535 4225
rect 2805 4185 2809 4322
rect 2984 4225 3085 4322
rect 2965 4185 3085 4225
rect 3355 4185 3359 4322
rect 3534 4225 3635 4322
rect 3515 4185 3635 4225
rect 3905 4185 3909 4322
rect 4084 4225 4185 4322
rect 4065 4185 4185 4225
rect 4455 4185 4459 4322
rect 4634 4225 4735 4322
rect 4615 4185 4735 4225
rect 5005 4185 5009 4322
rect 5184 4225 5285 4322
rect 5165 4185 5285 4225
rect 5555 4185 5559 4322
rect 5734 4225 5835 4322
rect 5715 4185 5835 4225
rect 6105 4185 6109 4322
rect 6284 4225 6385 4322
rect 6265 4185 6385 4225
rect 6655 4185 6659 4322
rect 6834 4225 6935 4322
rect 6815 4185 6935 4225
rect 7205 4185 7209 4322
rect 7384 4225 7485 4322
rect 7365 4185 7485 4225
rect 7755 4185 7759 4322
rect 7934 4225 8035 4322
rect 7915 4185 8035 4225
rect 8305 4185 8309 4322
rect 8484 4225 8585 4322
rect 8465 4185 8585 4225
rect 8855 4185 8859 4322
rect 9034 4225 9135 4322
rect 9015 4185 9135 4225
rect 9405 4185 9409 4322
rect 9584 4225 9685 4322
rect 9565 4185 9685 4225
rect 9955 4185 9959 4322
rect 10134 4225 10235 4322
rect 10115 4185 10235 4225
rect 10505 4185 10509 4322
rect 10684 4225 10785 4322
rect 10665 4185 10785 4225
rect 11055 4185 11059 4322
rect 11234 4225 11335 4322
rect 11215 4185 11335 4225
rect 11605 4185 11609 4322
rect 11784 4225 11885 4322
rect 11765 4185 11885 4225
rect 12155 4185 12159 4322
rect 12334 4225 12435 4322
rect 12315 4185 12435 4225
rect 12705 4185 12709 4322
rect 12884 4225 12985 4322
rect 12865 4185 12985 4225
rect 13255 4185 13259 4322
rect 13434 4225 13535 4322
rect 13415 4185 13535 4225
rect 13805 4185 13809 4322
rect 13984 4225 14085 4322
rect 13965 4185 14085 4225
rect 14355 4185 14359 4322
rect 14534 4225 14635 4322
rect 14515 4185 14635 4225
rect 14905 4185 14909 4322
rect 15084 4225 15185 4322
rect 15065 4185 15185 4225
rect 15455 4185 15459 4322
rect 15634 4225 15735 4322
rect 15615 4185 15735 4225
rect 16005 4185 16009 4322
rect 16184 4225 16285 4322
rect 16165 4185 16285 4225
rect 16555 4185 16559 4322
rect 16734 4225 16835 4322
rect 16715 4185 16835 4225
rect 17105 4185 17109 4322
rect 17284 4225 17385 4322
rect 17265 4185 17385 4225
rect 17655 4185 17659 4322
rect 17834 4225 17935 4322
rect 17815 4185 17935 4225
rect 18205 4185 18209 4322
rect 18384 4225 18485 4322
rect 18365 4185 18485 4225
rect 18755 4185 18759 4322
rect 18934 4225 19035 4322
rect 18915 4185 19035 4225
rect 725 4178 842 4185
rect 885 4178 1045 4185
rect 725 4072 808 4178
rect 842 4072 1045 4178
rect 725 4065 765 4072
rect 808 4065 1045 4072
rect 1275 4178 1392 4185
rect 1435 4178 1595 4185
rect 1275 4072 1358 4178
rect 1392 4072 1595 4178
rect 1275 4065 1315 4072
rect 1358 4065 1595 4072
rect 1825 4178 1942 4185
rect 1985 4178 2145 4185
rect 1825 4072 1908 4178
rect 1942 4072 2145 4178
rect 1825 4065 1865 4072
rect 1908 4065 2145 4072
rect 2375 4178 2492 4185
rect 2535 4178 2695 4185
rect 2375 4072 2458 4178
rect 2492 4072 2695 4178
rect 2375 4065 2415 4072
rect 2458 4065 2695 4072
rect 2925 4178 3042 4185
rect 3085 4178 3245 4185
rect 2925 4072 3008 4178
rect 3042 4072 3245 4178
rect 2925 4065 2965 4072
rect 3008 4065 3245 4072
rect 3475 4178 3592 4185
rect 3635 4178 3795 4185
rect 3475 4072 3558 4178
rect 3592 4072 3795 4178
rect 3475 4065 3515 4072
rect 3558 4065 3795 4072
rect 4025 4178 4142 4185
rect 4185 4178 4345 4185
rect 4025 4072 4108 4178
rect 4142 4072 4345 4178
rect 4025 4065 4065 4072
rect 4108 4065 4345 4072
rect 4575 4178 4692 4185
rect 4735 4178 4895 4185
rect 4575 4072 4658 4178
rect 4692 4072 4895 4178
rect 4575 4065 4615 4072
rect 4658 4065 4895 4072
rect 5125 4178 5242 4185
rect 5285 4178 5445 4185
rect 5125 4072 5208 4178
rect 5242 4072 5445 4178
rect 5125 4065 5165 4072
rect 5208 4065 5445 4072
rect 5675 4178 5792 4185
rect 5835 4178 5995 4185
rect 5675 4072 5758 4178
rect 5792 4072 5995 4178
rect 5675 4065 5715 4072
rect 5758 4065 5995 4072
rect 6225 4178 6342 4185
rect 6385 4178 6545 4185
rect 6225 4072 6308 4178
rect 6342 4072 6545 4178
rect 6225 4065 6265 4072
rect 6308 4065 6545 4072
rect 6775 4178 6892 4185
rect 6935 4178 7095 4185
rect 6775 4072 6858 4178
rect 6892 4072 7095 4178
rect 6775 4065 6815 4072
rect 6858 4065 7095 4072
rect 7325 4178 7442 4185
rect 7485 4178 7645 4185
rect 7325 4072 7408 4178
rect 7442 4072 7645 4178
rect 7325 4065 7365 4072
rect 7408 4065 7645 4072
rect 7875 4178 7992 4185
rect 8035 4178 8195 4185
rect 7875 4072 7958 4178
rect 7992 4072 8195 4178
rect 7875 4065 7915 4072
rect 7958 4065 8195 4072
rect 8425 4178 8542 4185
rect 8585 4178 8745 4185
rect 8425 4072 8508 4178
rect 8542 4072 8745 4178
rect 8425 4065 8465 4072
rect 8508 4065 8745 4072
rect 8975 4178 9092 4185
rect 9135 4178 9295 4185
rect 8975 4072 9058 4178
rect 9092 4072 9295 4178
rect 8975 4065 9015 4072
rect 9058 4065 9295 4072
rect 9525 4178 9642 4185
rect 9685 4178 9845 4185
rect 9525 4072 9608 4178
rect 9642 4072 9845 4178
rect 9525 4065 9565 4072
rect 9608 4065 9845 4072
rect 10075 4178 10192 4185
rect 10235 4178 10395 4185
rect 10075 4072 10158 4178
rect 10192 4072 10395 4178
rect 10075 4065 10115 4072
rect 10158 4065 10395 4072
rect 10625 4178 10742 4185
rect 10785 4178 10945 4185
rect 10625 4072 10708 4178
rect 10742 4072 10945 4178
rect 10625 4065 10665 4072
rect 10708 4065 10945 4072
rect 11175 4178 11292 4185
rect 11335 4178 11495 4185
rect 11175 4072 11258 4178
rect 11292 4072 11495 4178
rect 11175 4065 11215 4072
rect 11258 4065 11495 4072
rect 11725 4178 11842 4185
rect 11885 4178 12045 4185
rect 11725 4072 11808 4178
rect 11842 4072 12045 4178
rect 11725 4065 11765 4072
rect 11808 4065 12045 4072
rect 12275 4178 12392 4185
rect 12435 4178 12595 4185
rect 12275 4072 12358 4178
rect 12392 4072 12595 4178
rect 12275 4065 12315 4072
rect 12358 4065 12595 4072
rect 12825 4178 12942 4185
rect 12985 4178 13145 4185
rect 12825 4072 12908 4178
rect 12942 4072 13145 4178
rect 12825 4065 12865 4072
rect 12908 4065 13145 4072
rect 13375 4178 13492 4185
rect 13535 4178 13695 4185
rect 13375 4072 13458 4178
rect 13492 4072 13695 4178
rect 13375 4065 13415 4072
rect 13458 4065 13695 4072
rect 13925 4178 14042 4185
rect 14085 4178 14245 4185
rect 13925 4072 14008 4178
rect 14042 4072 14245 4178
rect 13925 4065 13965 4072
rect 14008 4065 14245 4072
rect 14475 4178 14592 4185
rect 14635 4178 14795 4185
rect 14475 4072 14558 4178
rect 14592 4072 14795 4178
rect 14475 4065 14515 4072
rect 14558 4065 14795 4072
rect 15025 4178 15142 4185
rect 15185 4178 15345 4185
rect 15025 4072 15108 4178
rect 15142 4072 15345 4178
rect 15025 4065 15065 4072
rect 15108 4065 15345 4072
rect 15575 4178 15692 4185
rect 15735 4178 15895 4185
rect 15575 4072 15658 4178
rect 15692 4072 15895 4178
rect 15575 4065 15615 4072
rect 15658 4065 15895 4072
rect 16125 4178 16242 4185
rect 16285 4178 16445 4185
rect 16125 4072 16208 4178
rect 16242 4072 16445 4178
rect 16125 4065 16165 4072
rect 16208 4065 16445 4072
rect 16675 4178 16792 4185
rect 16835 4178 16995 4185
rect 16675 4072 16758 4178
rect 16792 4072 16995 4178
rect 16675 4065 16715 4072
rect 16758 4065 16995 4072
rect 17225 4178 17342 4185
rect 17385 4178 17545 4185
rect 17225 4072 17308 4178
rect 17342 4072 17545 4178
rect 17225 4065 17265 4072
rect 17308 4065 17545 4072
rect 17775 4178 17892 4185
rect 17935 4178 18095 4185
rect 17775 4072 17858 4178
rect 17892 4072 18095 4178
rect 17775 4065 17815 4072
rect 17858 4065 18095 4072
rect 18325 4178 18442 4185
rect 18485 4178 18645 4185
rect 18325 4072 18408 4178
rect 18442 4072 18645 4178
rect 18325 4065 18365 4072
rect 18408 4065 18645 4072
rect 18875 4178 18992 4185
rect 19035 4178 19195 4185
rect 18875 4072 18958 4178
rect 18992 4072 19195 4178
rect 18875 4065 18915 4072
rect 18958 4065 19195 4072
rect 765 4025 885 4065
rect 1315 4025 1435 4065
rect 1865 4025 1985 4065
rect 2415 4025 2535 4065
rect 2965 4025 3085 4065
rect 3515 4025 3635 4065
rect 4065 4025 4185 4065
rect 4615 4025 4735 4065
rect 5165 4025 5285 4065
rect 5715 4025 5835 4065
rect 6265 4025 6385 4065
rect 6815 4025 6935 4065
rect 7365 4025 7485 4065
rect 7915 4025 8035 4065
rect 8465 4025 8585 4065
rect 9015 4025 9135 4065
rect 9565 4025 9685 4065
rect 10115 4025 10235 4065
rect 10665 4025 10785 4065
rect 11215 4025 11335 4065
rect 11765 4025 11885 4065
rect 12315 4025 12435 4065
rect 12865 4025 12985 4065
rect 13415 4025 13535 4065
rect 13965 4025 14085 4065
rect 14515 4025 14635 4065
rect 15065 4025 15185 4065
rect 15615 4025 15735 4065
rect 16165 4025 16285 4065
rect 16715 4025 16835 4065
rect 17265 4025 17385 4065
rect 17815 4025 17935 4065
rect 18365 4025 18485 4065
rect 18915 4025 19035 4065
rect 19202 3912 19204 4338
rect 500 3825 507 3875
rect 19202 3796 19217 3802
rect 628 3772 885 3795
rect 1178 3772 1435 3795
rect 1728 3772 1985 3795
rect 2278 3772 2535 3795
rect 2828 3772 3085 3795
rect 3378 3772 3635 3795
rect 3928 3772 4185 3795
rect 4478 3772 4735 3795
rect 5028 3772 5285 3795
rect 5578 3772 5835 3795
rect 6128 3772 6385 3795
rect 6678 3772 6935 3795
rect 7228 3772 7485 3795
rect 7778 3772 8035 3795
rect 8328 3772 8585 3795
rect 8878 3772 9135 3795
rect 9428 3772 9685 3795
rect 9978 3772 10235 3795
rect 10528 3772 10785 3795
rect 11078 3772 11335 3795
rect 11628 3772 11885 3795
rect 12178 3772 12435 3795
rect 12728 3772 12985 3795
rect 13278 3772 13535 3795
rect 13828 3772 14085 3795
rect 14378 3772 14635 3795
rect 14928 3772 15185 3795
rect 15478 3772 15735 3795
rect 16028 3772 16285 3795
rect 16578 3772 16835 3795
rect 17128 3772 17385 3795
rect 17678 3772 17935 3795
rect 18228 3772 18485 3795
rect 18778 3772 19035 3795
rect 605 3635 609 3772
rect 784 3675 885 3772
rect 765 3635 885 3675
rect 1155 3635 1159 3772
rect 1334 3675 1435 3772
rect 1315 3635 1435 3675
rect 1705 3635 1709 3772
rect 1884 3675 1985 3772
rect 1865 3635 1985 3675
rect 2255 3635 2259 3772
rect 2434 3675 2535 3772
rect 2415 3635 2535 3675
rect 2805 3635 2809 3772
rect 2984 3675 3085 3772
rect 2965 3635 3085 3675
rect 3355 3635 3359 3772
rect 3534 3675 3635 3772
rect 3515 3635 3635 3675
rect 3905 3635 3909 3772
rect 4084 3675 4185 3772
rect 4065 3635 4185 3675
rect 4455 3635 4459 3772
rect 4634 3675 4735 3772
rect 4615 3635 4735 3675
rect 5005 3635 5009 3772
rect 5184 3675 5285 3772
rect 5165 3635 5285 3675
rect 5555 3635 5559 3772
rect 5734 3675 5835 3772
rect 5715 3635 5835 3675
rect 6105 3635 6109 3772
rect 6284 3675 6385 3772
rect 6265 3635 6385 3675
rect 6655 3635 6659 3772
rect 6834 3675 6935 3772
rect 6815 3635 6935 3675
rect 7205 3635 7209 3772
rect 7384 3675 7485 3772
rect 7365 3635 7485 3675
rect 7755 3635 7759 3772
rect 7934 3675 8035 3772
rect 7915 3635 8035 3675
rect 8305 3635 8309 3772
rect 8484 3675 8585 3772
rect 8465 3635 8585 3675
rect 8855 3635 8859 3772
rect 9034 3675 9135 3772
rect 9015 3635 9135 3675
rect 9405 3635 9409 3772
rect 9584 3675 9685 3772
rect 9565 3635 9685 3675
rect 9955 3635 9959 3772
rect 10134 3675 10235 3772
rect 10115 3635 10235 3675
rect 10505 3635 10509 3772
rect 10684 3675 10785 3772
rect 10665 3635 10785 3675
rect 11055 3635 11059 3772
rect 11234 3675 11335 3772
rect 11215 3635 11335 3675
rect 11605 3635 11609 3772
rect 11784 3675 11885 3772
rect 11765 3635 11885 3675
rect 12155 3635 12159 3772
rect 12334 3675 12435 3772
rect 12315 3635 12435 3675
rect 12705 3635 12709 3772
rect 12884 3675 12985 3772
rect 12865 3635 12985 3675
rect 13255 3635 13259 3772
rect 13434 3675 13535 3772
rect 13415 3635 13535 3675
rect 13805 3635 13809 3772
rect 13984 3675 14085 3772
rect 13965 3635 14085 3675
rect 14355 3635 14359 3772
rect 14534 3675 14635 3772
rect 14515 3635 14635 3675
rect 14905 3635 14909 3772
rect 15084 3675 15185 3772
rect 15065 3635 15185 3675
rect 15455 3635 15459 3772
rect 15634 3675 15735 3772
rect 15615 3635 15735 3675
rect 16005 3635 16009 3772
rect 16184 3675 16285 3772
rect 16165 3635 16285 3675
rect 16555 3635 16559 3772
rect 16734 3675 16835 3772
rect 16715 3635 16835 3675
rect 17105 3635 17109 3772
rect 17284 3675 17385 3772
rect 17265 3635 17385 3675
rect 17655 3635 17659 3772
rect 17834 3675 17935 3772
rect 17815 3635 17935 3675
rect 18205 3635 18209 3772
rect 18384 3675 18485 3772
rect 18365 3635 18485 3675
rect 18755 3635 18759 3772
rect 18934 3675 19035 3772
rect 18915 3635 19035 3675
rect 725 3628 842 3635
rect 885 3628 1045 3635
rect 725 3522 808 3628
rect 842 3522 1045 3628
rect 725 3515 765 3522
rect 808 3515 1045 3522
rect 1275 3628 1392 3635
rect 1435 3628 1595 3635
rect 1275 3522 1358 3628
rect 1392 3522 1595 3628
rect 1275 3515 1315 3522
rect 1358 3515 1595 3522
rect 1825 3628 1942 3635
rect 1985 3628 2145 3635
rect 1825 3522 1908 3628
rect 1942 3522 2145 3628
rect 1825 3515 1865 3522
rect 1908 3515 2145 3522
rect 2375 3628 2492 3635
rect 2535 3628 2695 3635
rect 2375 3522 2458 3628
rect 2492 3522 2695 3628
rect 2375 3515 2415 3522
rect 2458 3515 2695 3522
rect 2925 3628 3042 3635
rect 3085 3628 3245 3635
rect 2925 3522 3008 3628
rect 3042 3522 3245 3628
rect 2925 3515 2965 3522
rect 3008 3515 3245 3522
rect 3475 3628 3592 3635
rect 3635 3628 3795 3635
rect 3475 3522 3558 3628
rect 3592 3522 3795 3628
rect 3475 3515 3515 3522
rect 3558 3515 3795 3522
rect 4025 3628 4142 3635
rect 4185 3628 4345 3635
rect 4025 3522 4108 3628
rect 4142 3522 4345 3628
rect 4025 3515 4065 3522
rect 4108 3515 4345 3522
rect 4575 3628 4692 3635
rect 4735 3628 4895 3635
rect 4575 3522 4658 3628
rect 4692 3522 4895 3628
rect 4575 3515 4615 3522
rect 4658 3515 4895 3522
rect 5125 3628 5242 3635
rect 5285 3628 5445 3635
rect 5125 3522 5208 3628
rect 5242 3522 5445 3628
rect 5125 3515 5165 3522
rect 5208 3515 5445 3522
rect 5675 3628 5792 3635
rect 5835 3628 5995 3635
rect 5675 3522 5758 3628
rect 5792 3522 5995 3628
rect 5675 3515 5715 3522
rect 5758 3515 5995 3522
rect 6225 3628 6342 3635
rect 6385 3628 6545 3635
rect 6225 3522 6308 3628
rect 6342 3522 6545 3628
rect 6225 3515 6265 3522
rect 6308 3515 6545 3522
rect 6775 3628 6892 3635
rect 6935 3628 7095 3635
rect 6775 3522 6858 3628
rect 6892 3522 7095 3628
rect 6775 3515 6815 3522
rect 6858 3515 7095 3522
rect 7325 3628 7442 3635
rect 7485 3628 7645 3635
rect 7325 3522 7408 3628
rect 7442 3522 7645 3628
rect 7325 3515 7365 3522
rect 7408 3515 7645 3522
rect 7875 3628 7992 3635
rect 8035 3628 8195 3635
rect 7875 3522 7958 3628
rect 7992 3522 8195 3628
rect 7875 3515 7915 3522
rect 7958 3515 8195 3522
rect 8425 3628 8542 3635
rect 8585 3628 8745 3635
rect 8425 3522 8508 3628
rect 8542 3522 8745 3628
rect 8425 3515 8465 3522
rect 8508 3515 8745 3522
rect 8975 3628 9092 3635
rect 9135 3628 9295 3635
rect 8975 3522 9058 3628
rect 9092 3522 9295 3628
rect 8975 3515 9015 3522
rect 9058 3515 9295 3522
rect 9525 3628 9642 3635
rect 9685 3628 9845 3635
rect 9525 3522 9608 3628
rect 9642 3522 9845 3628
rect 9525 3515 9565 3522
rect 9608 3515 9845 3522
rect 10075 3628 10192 3635
rect 10235 3628 10395 3635
rect 10075 3522 10158 3628
rect 10192 3522 10395 3628
rect 10075 3515 10115 3522
rect 10158 3515 10395 3522
rect 10625 3628 10742 3635
rect 10785 3628 10945 3635
rect 10625 3522 10708 3628
rect 10742 3522 10945 3628
rect 10625 3515 10665 3522
rect 10708 3515 10945 3522
rect 11175 3628 11292 3635
rect 11335 3628 11495 3635
rect 11175 3522 11258 3628
rect 11292 3522 11495 3628
rect 11175 3515 11215 3522
rect 11258 3515 11495 3522
rect 11725 3628 11842 3635
rect 11885 3628 12045 3635
rect 11725 3522 11808 3628
rect 11842 3522 12045 3628
rect 11725 3515 11765 3522
rect 11808 3515 12045 3522
rect 12275 3628 12392 3635
rect 12435 3628 12595 3635
rect 12275 3522 12358 3628
rect 12392 3522 12595 3628
rect 12275 3515 12315 3522
rect 12358 3515 12595 3522
rect 12825 3628 12942 3635
rect 12985 3628 13145 3635
rect 12825 3522 12908 3628
rect 12942 3522 13145 3628
rect 12825 3515 12865 3522
rect 12908 3515 13145 3522
rect 13375 3628 13492 3635
rect 13535 3628 13695 3635
rect 13375 3522 13458 3628
rect 13492 3522 13695 3628
rect 13375 3515 13415 3522
rect 13458 3515 13695 3522
rect 13925 3628 14042 3635
rect 14085 3628 14245 3635
rect 13925 3522 14008 3628
rect 14042 3522 14245 3628
rect 13925 3515 13965 3522
rect 14008 3515 14245 3522
rect 14475 3628 14592 3635
rect 14635 3628 14795 3635
rect 14475 3522 14558 3628
rect 14592 3522 14795 3628
rect 14475 3515 14515 3522
rect 14558 3515 14795 3522
rect 15025 3628 15142 3635
rect 15185 3628 15345 3635
rect 15025 3522 15108 3628
rect 15142 3522 15345 3628
rect 15025 3515 15065 3522
rect 15108 3515 15345 3522
rect 15575 3628 15692 3635
rect 15735 3628 15895 3635
rect 15575 3522 15658 3628
rect 15692 3522 15895 3628
rect 15575 3515 15615 3522
rect 15658 3515 15895 3522
rect 16125 3628 16242 3635
rect 16285 3628 16445 3635
rect 16125 3522 16208 3628
rect 16242 3522 16445 3628
rect 16125 3515 16165 3522
rect 16208 3515 16445 3522
rect 16675 3628 16792 3635
rect 16835 3628 16995 3635
rect 16675 3522 16758 3628
rect 16792 3522 16995 3628
rect 16675 3515 16715 3522
rect 16758 3515 16995 3522
rect 17225 3628 17342 3635
rect 17385 3628 17545 3635
rect 17225 3522 17308 3628
rect 17342 3522 17545 3628
rect 17225 3515 17265 3522
rect 17308 3515 17545 3522
rect 17775 3628 17892 3635
rect 17935 3628 18095 3635
rect 17775 3522 17858 3628
rect 17892 3522 18095 3628
rect 17775 3515 17815 3522
rect 17858 3515 18095 3522
rect 18325 3628 18442 3635
rect 18485 3628 18645 3635
rect 18325 3522 18408 3628
rect 18442 3522 18645 3628
rect 18325 3515 18365 3522
rect 18408 3515 18645 3522
rect 18875 3628 18992 3635
rect 19035 3628 19195 3635
rect 18875 3522 18958 3628
rect 18992 3522 19195 3628
rect 18875 3515 18915 3522
rect 18958 3515 19195 3522
rect 765 3475 885 3515
rect 1315 3475 1435 3515
rect 1865 3475 1985 3515
rect 2415 3475 2535 3515
rect 2965 3475 3085 3515
rect 3515 3475 3635 3515
rect 4065 3475 4185 3515
rect 4615 3475 4735 3515
rect 5165 3475 5285 3515
rect 5715 3475 5835 3515
rect 6265 3475 6385 3515
rect 6815 3475 6935 3515
rect 7365 3475 7485 3515
rect 7915 3475 8035 3515
rect 8465 3475 8585 3515
rect 9015 3475 9135 3515
rect 9565 3475 9685 3515
rect 10115 3475 10235 3515
rect 10665 3475 10785 3515
rect 11215 3475 11335 3515
rect 11765 3475 11885 3515
rect 12315 3475 12435 3515
rect 12865 3475 12985 3515
rect 13415 3475 13535 3515
rect 13965 3475 14085 3515
rect 14515 3475 14635 3515
rect 15065 3475 15185 3515
rect 15615 3475 15735 3515
rect 16165 3475 16285 3515
rect 16715 3475 16835 3515
rect 17265 3475 17385 3515
rect 17815 3475 17935 3515
rect 18365 3475 18485 3515
rect 18915 3475 19035 3515
rect 19185 3354 19200 3371
rect 19202 3362 19204 3788
rect 19202 3348 19217 3354
rect 500 3275 507 3325
rect 500 2839 525 3240
rect 628 3222 885 3245
rect 1178 3222 1435 3245
rect 1728 3222 1985 3245
rect 2278 3222 2535 3245
rect 2828 3222 3085 3245
rect 3378 3222 3635 3245
rect 3928 3222 4185 3245
rect 4478 3222 4735 3245
rect 5028 3222 5285 3245
rect 5578 3222 5835 3245
rect 6128 3222 6385 3245
rect 6678 3222 6935 3245
rect 7228 3222 7485 3245
rect 7778 3222 8035 3245
rect 8328 3222 8585 3245
rect 8878 3222 9135 3245
rect 9428 3222 9685 3245
rect 9978 3222 10235 3245
rect 10528 3222 10785 3245
rect 11078 3222 11335 3245
rect 11628 3222 11885 3245
rect 12178 3222 12435 3245
rect 12728 3222 12985 3245
rect 13278 3222 13535 3245
rect 13828 3222 14085 3245
rect 14378 3222 14635 3245
rect 14928 3222 15185 3245
rect 15478 3222 15735 3245
rect 16028 3222 16285 3245
rect 16578 3222 16835 3245
rect 17128 3222 17385 3245
rect 17678 3222 17935 3245
rect 18228 3222 18485 3245
rect 18778 3222 19035 3245
rect 605 3085 609 3222
rect 784 3125 885 3222
rect 765 3085 885 3125
rect 1155 3085 1159 3222
rect 1334 3125 1435 3222
rect 1315 3085 1435 3125
rect 1705 3085 1709 3222
rect 1884 3125 1985 3222
rect 1865 3085 1985 3125
rect 2255 3085 2259 3222
rect 2434 3125 2535 3222
rect 2415 3085 2535 3125
rect 2805 3085 2809 3222
rect 2984 3125 3085 3222
rect 2965 3085 3085 3125
rect 3355 3085 3359 3222
rect 3534 3125 3635 3222
rect 3515 3085 3635 3125
rect 3905 3085 3909 3222
rect 4084 3125 4185 3222
rect 4065 3085 4185 3125
rect 4455 3085 4459 3222
rect 4634 3125 4735 3222
rect 4615 3085 4735 3125
rect 5005 3085 5009 3222
rect 5184 3125 5285 3222
rect 5165 3085 5285 3125
rect 5555 3085 5559 3222
rect 5734 3125 5835 3222
rect 5715 3085 5835 3125
rect 6105 3085 6109 3222
rect 6284 3125 6385 3222
rect 6265 3085 6385 3125
rect 6655 3085 6659 3222
rect 6834 3125 6935 3222
rect 6815 3085 6935 3125
rect 7205 3085 7209 3222
rect 7384 3125 7485 3222
rect 7365 3085 7485 3125
rect 7755 3085 7759 3222
rect 7934 3125 8035 3222
rect 7915 3085 8035 3125
rect 8305 3085 8309 3222
rect 8484 3125 8585 3222
rect 8465 3085 8585 3125
rect 8855 3085 8859 3222
rect 9034 3125 9135 3222
rect 9015 3085 9135 3125
rect 9405 3085 9409 3222
rect 9584 3125 9685 3222
rect 9565 3085 9685 3125
rect 9955 3085 9959 3222
rect 10134 3125 10235 3222
rect 10115 3085 10235 3125
rect 10505 3085 10509 3222
rect 10684 3125 10785 3222
rect 10665 3085 10785 3125
rect 11055 3085 11059 3222
rect 11234 3125 11335 3222
rect 11215 3085 11335 3125
rect 11605 3085 11609 3222
rect 11784 3125 11885 3222
rect 11765 3085 11885 3125
rect 12155 3085 12159 3222
rect 12334 3125 12435 3222
rect 12315 3085 12435 3125
rect 12705 3085 12709 3222
rect 12884 3125 12985 3222
rect 12865 3085 12985 3125
rect 13255 3085 13259 3222
rect 13434 3125 13535 3222
rect 13415 3085 13535 3125
rect 13805 3085 13809 3222
rect 13984 3125 14085 3222
rect 13965 3085 14085 3125
rect 14355 3085 14359 3222
rect 14534 3125 14635 3222
rect 14515 3085 14635 3125
rect 14905 3085 14909 3222
rect 15084 3125 15185 3222
rect 15065 3085 15185 3125
rect 15455 3085 15459 3222
rect 15634 3125 15735 3222
rect 15615 3085 15735 3125
rect 16005 3085 16009 3222
rect 16184 3125 16285 3222
rect 16165 3085 16285 3125
rect 16555 3085 16559 3222
rect 16734 3125 16835 3222
rect 16715 3085 16835 3125
rect 17105 3085 17109 3222
rect 17284 3125 17385 3222
rect 17265 3085 17385 3125
rect 17655 3085 17659 3222
rect 17834 3125 17935 3222
rect 17815 3085 17935 3125
rect 18205 3085 18209 3222
rect 18384 3125 18485 3222
rect 18365 3085 18485 3125
rect 18755 3085 18759 3222
rect 18934 3125 19035 3222
rect 18915 3085 19035 3125
rect 725 3078 842 3085
rect 885 3078 1045 3085
rect 725 2972 808 3078
rect 842 2972 1045 3078
rect 725 2965 765 2972
rect 808 2965 1045 2972
rect 1275 3078 1392 3085
rect 1435 3078 1595 3085
rect 1275 2972 1358 3078
rect 1392 2972 1595 3078
rect 1275 2965 1315 2972
rect 1358 2965 1595 2972
rect 1825 3078 1942 3085
rect 1985 3078 2145 3085
rect 1825 2972 1908 3078
rect 1942 2972 2145 3078
rect 1825 2965 1865 2972
rect 1908 2965 2145 2972
rect 2375 3078 2492 3085
rect 2535 3078 2695 3085
rect 2375 2972 2458 3078
rect 2492 2972 2695 3078
rect 2375 2965 2415 2972
rect 2458 2965 2695 2972
rect 2925 3078 3042 3085
rect 3085 3078 3245 3085
rect 2925 2972 3008 3078
rect 3042 2972 3245 3078
rect 2925 2965 2965 2972
rect 3008 2965 3245 2972
rect 3475 3078 3592 3085
rect 3635 3078 3795 3085
rect 3475 2972 3558 3078
rect 3592 2972 3795 3078
rect 3475 2965 3515 2972
rect 3558 2965 3795 2972
rect 4025 3078 4142 3085
rect 4185 3078 4345 3085
rect 4025 2972 4108 3078
rect 4142 2972 4345 3078
rect 4025 2965 4065 2972
rect 4108 2965 4345 2972
rect 4575 3078 4692 3085
rect 4735 3078 4895 3085
rect 4575 2972 4658 3078
rect 4692 2972 4895 3078
rect 4575 2965 4615 2972
rect 4658 2965 4895 2972
rect 5125 3078 5242 3085
rect 5285 3078 5445 3085
rect 5125 2972 5208 3078
rect 5242 2972 5445 3078
rect 5125 2965 5165 2972
rect 5208 2965 5445 2972
rect 5675 3078 5792 3085
rect 5835 3078 5995 3085
rect 5675 2972 5758 3078
rect 5792 2972 5995 3078
rect 5675 2965 5715 2972
rect 5758 2965 5995 2972
rect 6225 3078 6342 3085
rect 6385 3078 6545 3085
rect 6225 2972 6308 3078
rect 6342 2972 6545 3078
rect 6225 2965 6265 2972
rect 6308 2965 6545 2972
rect 6775 3078 6892 3085
rect 6935 3078 7095 3085
rect 6775 2972 6858 3078
rect 6892 2972 7095 3078
rect 6775 2965 6815 2972
rect 6858 2965 7095 2972
rect 7325 3078 7442 3085
rect 7485 3078 7645 3085
rect 7325 2972 7408 3078
rect 7442 2972 7645 3078
rect 7325 2965 7365 2972
rect 7408 2965 7645 2972
rect 7875 3078 7992 3085
rect 8035 3078 8195 3085
rect 7875 2972 7958 3078
rect 7992 2972 8195 3078
rect 7875 2965 7915 2972
rect 7958 2965 8195 2972
rect 8425 3078 8542 3085
rect 8585 3078 8745 3085
rect 8425 2972 8508 3078
rect 8542 2972 8745 3078
rect 8425 2965 8465 2972
rect 8508 2965 8745 2972
rect 8975 3078 9092 3085
rect 9135 3078 9295 3085
rect 8975 2972 9058 3078
rect 9092 2972 9295 3078
rect 8975 2965 9015 2972
rect 9058 2965 9295 2972
rect 9525 3078 9642 3085
rect 9685 3078 9845 3085
rect 9525 2972 9608 3078
rect 9642 2972 9845 3078
rect 9525 2965 9565 2972
rect 9608 2965 9845 2972
rect 10075 3078 10192 3085
rect 10235 3078 10395 3085
rect 10075 2972 10158 3078
rect 10192 2972 10395 3078
rect 10075 2965 10115 2972
rect 10158 2965 10395 2972
rect 10625 3078 10742 3085
rect 10785 3078 10945 3085
rect 10625 2972 10708 3078
rect 10742 2972 10945 3078
rect 10625 2965 10665 2972
rect 10708 2965 10945 2972
rect 11175 3078 11292 3085
rect 11335 3078 11495 3085
rect 11175 2972 11258 3078
rect 11292 2972 11495 3078
rect 11175 2965 11215 2972
rect 11258 2965 11495 2972
rect 11725 3078 11842 3085
rect 11885 3078 12045 3085
rect 11725 2972 11808 3078
rect 11842 2972 12045 3078
rect 11725 2965 11765 2972
rect 11808 2965 12045 2972
rect 12275 3078 12392 3085
rect 12435 3078 12595 3085
rect 12275 2972 12358 3078
rect 12392 2972 12595 3078
rect 12275 2965 12315 2972
rect 12358 2965 12595 2972
rect 12825 3078 12942 3085
rect 12985 3078 13145 3085
rect 12825 2972 12908 3078
rect 12942 2972 13145 3078
rect 12825 2965 12865 2972
rect 12908 2965 13145 2972
rect 13375 3078 13492 3085
rect 13535 3078 13695 3085
rect 13375 2972 13458 3078
rect 13492 2972 13695 3078
rect 13375 2965 13415 2972
rect 13458 2965 13695 2972
rect 13925 3078 14042 3085
rect 14085 3078 14245 3085
rect 13925 2972 14008 3078
rect 14042 2972 14245 3078
rect 13925 2965 13965 2972
rect 14008 2965 14245 2972
rect 14475 3078 14592 3085
rect 14635 3078 14795 3085
rect 14475 2972 14558 3078
rect 14592 2972 14795 3078
rect 14475 2965 14515 2972
rect 14558 2965 14795 2972
rect 15025 3078 15142 3085
rect 15185 3078 15345 3085
rect 15025 2972 15108 3078
rect 15142 2972 15345 3078
rect 15025 2965 15065 2972
rect 15108 2965 15345 2972
rect 15575 3078 15692 3085
rect 15735 3078 15895 3085
rect 15575 2972 15658 3078
rect 15692 2972 15895 3078
rect 15575 2965 15615 2972
rect 15658 2965 15895 2972
rect 16125 3078 16242 3085
rect 16285 3078 16445 3085
rect 16125 2972 16208 3078
rect 16242 2972 16445 3078
rect 16125 2965 16165 2972
rect 16208 2965 16445 2972
rect 16675 3078 16792 3085
rect 16835 3078 16995 3085
rect 16675 2972 16758 3078
rect 16792 2972 16995 3078
rect 16675 2965 16715 2972
rect 16758 2965 16995 2972
rect 17225 3078 17342 3085
rect 17385 3078 17545 3085
rect 17225 2972 17308 3078
rect 17342 2972 17545 3078
rect 17225 2965 17265 2972
rect 17308 2965 17545 2972
rect 17775 3078 17892 3085
rect 17935 3078 18095 3085
rect 17775 2972 17858 3078
rect 17892 2972 18095 3078
rect 17775 2965 17815 2972
rect 17858 2965 18095 2972
rect 18325 3078 18442 3085
rect 18485 3078 18645 3085
rect 18325 2972 18408 3078
rect 18442 2972 18645 3078
rect 18325 2965 18365 2972
rect 18408 2965 18645 2972
rect 18875 3078 18992 3085
rect 19035 3078 19195 3085
rect 18875 2972 18958 3078
rect 18992 2972 19195 3078
rect 18875 2965 18915 2972
rect 18958 2965 19195 2972
rect 765 2925 885 2965
rect 1315 2925 1435 2965
rect 1865 2925 1985 2965
rect 2415 2925 2535 2965
rect 2965 2925 3085 2965
rect 3515 2925 3635 2965
rect 4065 2925 4185 2965
rect 4615 2925 4735 2965
rect 5165 2925 5285 2965
rect 5715 2925 5835 2965
rect 6265 2925 6385 2965
rect 6815 2925 6935 2965
rect 7365 2925 7485 2965
rect 7915 2925 8035 2965
rect 8465 2925 8585 2965
rect 9015 2925 9135 2965
rect 9565 2925 9685 2965
rect 10115 2925 10235 2965
rect 10665 2925 10785 2965
rect 11215 2925 11335 2965
rect 11765 2925 11885 2965
rect 12315 2925 12435 2965
rect 12865 2925 12985 2965
rect 13415 2925 13535 2965
rect 13965 2925 14085 2965
rect 14515 2925 14635 2965
rect 15065 2925 15185 2965
rect 15615 2925 15735 2965
rect 16165 2925 16285 2965
rect 16715 2925 16835 2965
rect 17265 2925 17385 2965
rect 17815 2925 17935 2965
rect 18365 2925 18485 2965
rect 18915 2925 19035 2965
rect 19202 2812 19204 3238
rect 500 2725 507 2775
rect 19202 2696 19217 2702
rect 628 2672 885 2695
rect 1178 2672 1435 2695
rect 1728 2672 1985 2695
rect 2278 2672 2535 2695
rect 2828 2672 3085 2695
rect 3378 2672 3635 2695
rect 3928 2672 4185 2695
rect 4478 2672 4735 2695
rect 5028 2672 5285 2695
rect 5578 2672 5835 2695
rect 6128 2672 6385 2695
rect 6678 2672 6935 2695
rect 7228 2672 7485 2695
rect 7778 2672 8035 2695
rect 8328 2672 8585 2695
rect 8878 2672 9135 2695
rect 9428 2672 9685 2695
rect 9978 2672 10235 2695
rect 10528 2672 10785 2695
rect 11078 2672 11335 2695
rect 11628 2672 11885 2695
rect 12178 2672 12435 2695
rect 12728 2672 12985 2695
rect 13278 2672 13535 2695
rect 13828 2672 14085 2695
rect 14378 2672 14635 2695
rect 14928 2672 15185 2695
rect 15478 2672 15735 2695
rect 16028 2672 16285 2695
rect 16578 2672 16835 2695
rect 17128 2672 17385 2695
rect 17678 2672 17935 2695
rect 18228 2672 18485 2695
rect 18778 2672 19035 2695
rect 605 2535 609 2672
rect 784 2575 885 2672
rect 765 2535 885 2575
rect 1155 2535 1159 2672
rect 1334 2575 1435 2672
rect 1315 2535 1435 2575
rect 1705 2535 1709 2672
rect 1884 2575 1985 2672
rect 1865 2535 1985 2575
rect 2255 2535 2259 2672
rect 2434 2575 2535 2672
rect 2415 2535 2535 2575
rect 2805 2535 2809 2672
rect 2984 2575 3085 2672
rect 2965 2535 3085 2575
rect 3355 2535 3359 2672
rect 3534 2575 3635 2672
rect 3515 2535 3635 2575
rect 3905 2535 3909 2672
rect 4084 2575 4185 2672
rect 4065 2535 4185 2575
rect 4455 2535 4459 2672
rect 4634 2575 4735 2672
rect 4615 2535 4735 2575
rect 5005 2535 5009 2672
rect 5184 2575 5285 2672
rect 5165 2535 5285 2575
rect 5555 2535 5559 2672
rect 5734 2575 5835 2672
rect 5715 2535 5835 2575
rect 6105 2535 6109 2672
rect 6284 2575 6385 2672
rect 6265 2535 6385 2575
rect 6655 2535 6659 2672
rect 6834 2575 6935 2672
rect 6815 2535 6935 2575
rect 7205 2535 7209 2672
rect 7384 2575 7485 2672
rect 7365 2535 7485 2575
rect 7755 2535 7759 2672
rect 7934 2575 8035 2672
rect 7915 2535 8035 2575
rect 8305 2535 8309 2672
rect 8484 2575 8585 2672
rect 8465 2535 8585 2575
rect 8855 2535 8859 2672
rect 9034 2575 9135 2672
rect 9015 2535 9135 2575
rect 9405 2535 9409 2672
rect 9584 2575 9685 2672
rect 9565 2535 9685 2575
rect 9955 2535 9959 2672
rect 10134 2575 10235 2672
rect 10115 2535 10235 2575
rect 10505 2535 10509 2672
rect 10684 2575 10785 2672
rect 10665 2535 10785 2575
rect 11055 2535 11059 2672
rect 11234 2575 11335 2672
rect 11215 2535 11335 2575
rect 11605 2535 11609 2672
rect 11784 2575 11885 2672
rect 11765 2535 11885 2575
rect 12155 2535 12159 2672
rect 12334 2575 12435 2672
rect 12315 2535 12435 2575
rect 12705 2535 12709 2672
rect 12884 2575 12985 2672
rect 12865 2535 12985 2575
rect 13255 2535 13259 2672
rect 13434 2575 13535 2672
rect 13415 2535 13535 2575
rect 13805 2535 13809 2672
rect 13984 2575 14085 2672
rect 13965 2535 14085 2575
rect 14355 2535 14359 2672
rect 14534 2575 14635 2672
rect 14515 2535 14635 2575
rect 14905 2535 14909 2672
rect 15084 2575 15185 2672
rect 15065 2535 15185 2575
rect 15455 2535 15459 2672
rect 15634 2575 15735 2672
rect 15615 2535 15735 2575
rect 16005 2535 16009 2672
rect 16184 2575 16285 2672
rect 16165 2535 16285 2575
rect 16555 2535 16559 2672
rect 16734 2575 16835 2672
rect 16715 2535 16835 2575
rect 17105 2535 17109 2672
rect 17284 2575 17385 2672
rect 17265 2535 17385 2575
rect 17655 2535 17659 2672
rect 17834 2575 17935 2672
rect 17815 2535 17935 2575
rect 18205 2535 18209 2672
rect 18384 2575 18485 2672
rect 18365 2535 18485 2575
rect 18755 2535 18759 2672
rect 18934 2575 19035 2672
rect 18915 2535 19035 2575
rect 725 2528 842 2535
rect 885 2528 1045 2535
rect 725 2422 808 2528
rect 842 2422 1045 2528
rect 725 2415 765 2422
rect 808 2415 1045 2422
rect 1275 2528 1392 2535
rect 1435 2528 1595 2535
rect 1275 2422 1358 2528
rect 1392 2422 1595 2528
rect 1275 2415 1315 2422
rect 1358 2415 1595 2422
rect 1825 2528 1942 2535
rect 1985 2528 2145 2535
rect 1825 2422 1908 2528
rect 1942 2422 2145 2528
rect 1825 2415 1865 2422
rect 1908 2415 2145 2422
rect 2375 2528 2492 2535
rect 2535 2528 2695 2535
rect 2375 2422 2458 2528
rect 2492 2422 2695 2528
rect 2375 2415 2415 2422
rect 2458 2415 2695 2422
rect 2925 2528 3042 2535
rect 3085 2528 3245 2535
rect 2925 2422 3008 2528
rect 3042 2422 3245 2528
rect 2925 2415 2965 2422
rect 3008 2415 3245 2422
rect 3475 2528 3592 2535
rect 3635 2528 3795 2535
rect 3475 2422 3558 2528
rect 3592 2422 3795 2528
rect 3475 2415 3515 2422
rect 3558 2415 3795 2422
rect 4025 2528 4142 2535
rect 4185 2528 4345 2535
rect 4025 2422 4108 2528
rect 4142 2422 4345 2528
rect 4025 2415 4065 2422
rect 4108 2415 4345 2422
rect 4575 2528 4692 2535
rect 4735 2528 4895 2535
rect 4575 2422 4658 2528
rect 4692 2422 4895 2528
rect 4575 2415 4615 2422
rect 4658 2415 4895 2422
rect 5125 2528 5242 2535
rect 5285 2528 5445 2535
rect 5125 2422 5208 2528
rect 5242 2422 5445 2528
rect 5125 2415 5165 2422
rect 5208 2415 5445 2422
rect 5675 2528 5792 2535
rect 5835 2528 5995 2535
rect 5675 2422 5758 2528
rect 5792 2422 5995 2528
rect 5675 2415 5715 2422
rect 5758 2415 5995 2422
rect 6225 2528 6342 2535
rect 6385 2528 6545 2535
rect 6225 2422 6308 2528
rect 6342 2422 6545 2528
rect 6225 2415 6265 2422
rect 6308 2415 6545 2422
rect 6775 2528 6892 2535
rect 6935 2528 7095 2535
rect 6775 2422 6858 2528
rect 6892 2422 7095 2528
rect 6775 2415 6815 2422
rect 6858 2415 7095 2422
rect 7325 2528 7442 2535
rect 7485 2528 7645 2535
rect 7325 2422 7408 2528
rect 7442 2422 7645 2528
rect 7325 2415 7365 2422
rect 7408 2415 7645 2422
rect 7875 2528 7992 2535
rect 8035 2528 8195 2535
rect 7875 2422 7958 2528
rect 7992 2422 8195 2528
rect 7875 2415 7915 2422
rect 7958 2415 8195 2422
rect 8425 2528 8542 2535
rect 8585 2528 8745 2535
rect 8425 2422 8508 2528
rect 8542 2422 8745 2528
rect 8425 2415 8465 2422
rect 8508 2415 8745 2422
rect 8975 2528 9092 2535
rect 9135 2528 9295 2535
rect 8975 2422 9058 2528
rect 9092 2422 9295 2528
rect 8975 2415 9015 2422
rect 9058 2415 9295 2422
rect 9525 2528 9642 2535
rect 9685 2528 9845 2535
rect 9525 2422 9608 2528
rect 9642 2422 9845 2528
rect 9525 2415 9565 2422
rect 9608 2415 9845 2422
rect 10075 2528 10192 2535
rect 10235 2528 10395 2535
rect 10075 2422 10158 2528
rect 10192 2422 10395 2528
rect 10075 2415 10115 2422
rect 10158 2415 10395 2422
rect 10625 2528 10742 2535
rect 10785 2528 10945 2535
rect 10625 2422 10708 2528
rect 10742 2422 10945 2528
rect 10625 2415 10665 2422
rect 10708 2415 10945 2422
rect 11175 2528 11292 2535
rect 11335 2528 11495 2535
rect 11175 2422 11258 2528
rect 11292 2422 11495 2528
rect 11175 2415 11215 2422
rect 11258 2415 11495 2422
rect 11725 2528 11842 2535
rect 11885 2528 12045 2535
rect 11725 2422 11808 2528
rect 11842 2422 12045 2528
rect 11725 2415 11765 2422
rect 11808 2415 12045 2422
rect 12275 2528 12392 2535
rect 12435 2528 12595 2535
rect 12275 2422 12358 2528
rect 12392 2422 12595 2528
rect 12275 2415 12315 2422
rect 12358 2415 12595 2422
rect 12825 2528 12942 2535
rect 12985 2528 13145 2535
rect 12825 2422 12908 2528
rect 12942 2422 13145 2528
rect 12825 2415 12865 2422
rect 12908 2415 13145 2422
rect 13375 2528 13492 2535
rect 13535 2528 13695 2535
rect 13375 2422 13458 2528
rect 13492 2422 13695 2528
rect 13375 2415 13415 2422
rect 13458 2415 13695 2422
rect 13925 2528 14042 2535
rect 14085 2528 14245 2535
rect 13925 2422 14008 2528
rect 14042 2422 14245 2528
rect 13925 2415 13965 2422
rect 14008 2415 14245 2422
rect 14475 2528 14592 2535
rect 14635 2528 14795 2535
rect 14475 2422 14558 2528
rect 14592 2422 14795 2528
rect 14475 2415 14515 2422
rect 14558 2415 14795 2422
rect 15025 2528 15142 2535
rect 15185 2528 15345 2535
rect 15025 2422 15108 2528
rect 15142 2422 15345 2528
rect 15025 2415 15065 2422
rect 15108 2415 15345 2422
rect 15575 2528 15692 2535
rect 15735 2528 15895 2535
rect 15575 2422 15658 2528
rect 15692 2422 15895 2528
rect 15575 2415 15615 2422
rect 15658 2415 15895 2422
rect 16125 2528 16242 2535
rect 16285 2528 16445 2535
rect 16125 2422 16208 2528
rect 16242 2422 16445 2528
rect 16125 2415 16165 2422
rect 16208 2415 16445 2422
rect 16675 2528 16792 2535
rect 16835 2528 16995 2535
rect 16675 2422 16758 2528
rect 16792 2422 16995 2528
rect 16675 2415 16715 2422
rect 16758 2415 16995 2422
rect 17225 2528 17342 2535
rect 17385 2528 17545 2535
rect 17225 2422 17308 2528
rect 17342 2422 17545 2528
rect 17225 2415 17265 2422
rect 17308 2415 17545 2422
rect 17775 2528 17892 2535
rect 17935 2528 18095 2535
rect 17775 2422 17858 2528
rect 17892 2422 18095 2528
rect 17775 2415 17815 2422
rect 17858 2415 18095 2422
rect 18325 2528 18442 2535
rect 18485 2528 18645 2535
rect 18325 2422 18408 2528
rect 18442 2422 18645 2528
rect 18325 2415 18365 2422
rect 18408 2415 18645 2422
rect 18875 2528 18992 2535
rect 19035 2528 19195 2535
rect 18875 2422 18958 2528
rect 18992 2422 19195 2528
rect 18875 2415 18915 2422
rect 18958 2415 19195 2422
rect 765 2375 885 2415
rect 1315 2375 1435 2415
rect 1865 2375 1985 2415
rect 2415 2375 2535 2415
rect 2965 2375 3085 2415
rect 3515 2375 3635 2415
rect 4065 2375 4185 2415
rect 4615 2375 4735 2415
rect 5165 2375 5285 2415
rect 5715 2375 5835 2415
rect 6265 2375 6385 2415
rect 6815 2375 6935 2415
rect 7365 2375 7485 2415
rect 7915 2375 8035 2415
rect 8465 2375 8585 2415
rect 9015 2375 9135 2415
rect 9565 2375 9685 2415
rect 10115 2375 10235 2415
rect 10665 2375 10785 2415
rect 11215 2375 11335 2415
rect 11765 2375 11885 2415
rect 12315 2375 12435 2415
rect 12865 2375 12985 2415
rect 13415 2375 13535 2415
rect 13965 2375 14085 2415
rect 14515 2375 14635 2415
rect 15065 2375 15185 2415
rect 15615 2375 15735 2415
rect 16165 2375 16285 2415
rect 16715 2375 16835 2415
rect 17265 2375 17385 2415
rect 17815 2375 17935 2415
rect 18365 2375 18485 2415
rect 18915 2375 19035 2415
rect 19185 2254 19200 2271
rect 19202 2262 19204 2688
rect 19202 2248 19217 2254
rect 500 2175 507 2225
rect 500 1739 525 2140
rect 628 2122 885 2145
rect 1178 2122 1435 2145
rect 1728 2122 1985 2145
rect 2278 2122 2535 2145
rect 2828 2122 3085 2145
rect 3378 2122 3635 2145
rect 3928 2122 4185 2145
rect 4478 2122 4735 2145
rect 5028 2122 5285 2145
rect 5578 2122 5835 2145
rect 6128 2122 6385 2145
rect 6678 2122 6935 2145
rect 7228 2122 7485 2145
rect 7778 2122 8035 2145
rect 8328 2122 8585 2145
rect 8878 2122 9135 2145
rect 9428 2122 9685 2145
rect 9978 2122 10235 2145
rect 10528 2122 10785 2145
rect 11078 2122 11335 2145
rect 11628 2122 11885 2145
rect 12178 2122 12435 2145
rect 12728 2122 12985 2145
rect 13278 2122 13535 2145
rect 13828 2122 14085 2145
rect 14378 2122 14635 2145
rect 14928 2122 15185 2145
rect 15478 2122 15735 2145
rect 16028 2122 16285 2145
rect 16578 2122 16835 2145
rect 17128 2122 17385 2145
rect 17678 2122 17935 2145
rect 18228 2122 18485 2145
rect 18778 2122 19035 2145
rect 605 1985 609 2122
rect 784 2025 885 2122
rect 765 1985 885 2025
rect 1155 1985 1159 2122
rect 1334 2025 1435 2122
rect 1315 1985 1435 2025
rect 1705 1985 1709 2122
rect 1884 2025 1985 2122
rect 1865 1985 1985 2025
rect 2255 1985 2259 2122
rect 2434 2025 2535 2122
rect 2415 1985 2535 2025
rect 2805 1985 2809 2122
rect 2984 2025 3085 2122
rect 2965 1985 3085 2025
rect 3355 1985 3359 2122
rect 3534 2025 3635 2122
rect 3515 1985 3635 2025
rect 3905 1985 3909 2122
rect 4084 2025 4185 2122
rect 4065 1985 4185 2025
rect 4455 1985 4459 2122
rect 4634 2025 4735 2122
rect 4615 1985 4735 2025
rect 5005 1985 5009 2122
rect 5184 2025 5285 2122
rect 5165 1985 5285 2025
rect 5555 1985 5559 2122
rect 5734 2025 5835 2122
rect 5715 1985 5835 2025
rect 6105 1985 6109 2122
rect 6284 2025 6385 2122
rect 6265 1985 6385 2025
rect 6655 1985 6659 2122
rect 6834 2025 6935 2122
rect 6815 1985 6935 2025
rect 7205 1985 7209 2122
rect 7384 2025 7485 2122
rect 7365 1985 7485 2025
rect 7755 1985 7759 2122
rect 7934 2025 8035 2122
rect 7915 1985 8035 2025
rect 8305 1985 8309 2122
rect 8484 2025 8585 2122
rect 8465 1985 8585 2025
rect 8855 1985 8859 2122
rect 9034 2025 9135 2122
rect 9015 1985 9135 2025
rect 9405 1985 9409 2122
rect 9584 2025 9685 2122
rect 9565 1985 9685 2025
rect 9955 1985 9959 2122
rect 10134 2025 10235 2122
rect 10115 1985 10235 2025
rect 10505 1985 10509 2122
rect 10684 2025 10785 2122
rect 10665 1985 10785 2025
rect 11055 1985 11059 2122
rect 11234 2025 11335 2122
rect 11215 1985 11335 2025
rect 11605 1985 11609 2122
rect 11784 2025 11885 2122
rect 11765 1985 11885 2025
rect 12155 1985 12159 2122
rect 12334 2025 12435 2122
rect 12315 1985 12435 2025
rect 12705 1985 12709 2122
rect 12884 2025 12985 2122
rect 12865 1985 12985 2025
rect 13255 1985 13259 2122
rect 13434 2025 13535 2122
rect 13415 1985 13535 2025
rect 13805 1985 13809 2122
rect 13984 2025 14085 2122
rect 13965 1985 14085 2025
rect 14355 1985 14359 2122
rect 14534 2025 14635 2122
rect 14515 1985 14635 2025
rect 14905 1985 14909 2122
rect 15084 2025 15185 2122
rect 15065 1985 15185 2025
rect 15455 1985 15459 2122
rect 15634 2025 15735 2122
rect 15615 1985 15735 2025
rect 16005 1985 16009 2122
rect 16184 2025 16285 2122
rect 16165 1985 16285 2025
rect 16555 1985 16559 2122
rect 16734 2025 16835 2122
rect 16715 1985 16835 2025
rect 17105 1985 17109 2122
rect 17284 2025 17385 2122
rect 17265 1985 17385 2025
rect 17655 1985 17659 2122
rect 17834 2025 17935 2122
rect 17815 1985 17935 2025
rect 18205 1985 18209 2122
rect 18384 2025 18485 2122
rect 18365 1985 18485 2025
rect 18755 1985 18759 2122
rect 18934 2025 19035 2122
rect 18915 1985 19035 2025
rect 725 1978 842 1985
rect 885 1978 1045 1985
rect 725 1872 808 1978
rect 842 1872 1045 1978
rect 725 1865 765 1872
rect 808 1865 1045 1872
rect 1275 1978 1392 1985
rect 1435 1978 1595 1985
rect 1275 1872 1358 1978
rect 1392 1872 1595 1978
rect 1275 1865 1315 1872
rect 1358 1865 1595 1872
rect 1825 1978 1942 1985
rect 1985 1978 2145 1985
rect 1825 1872 1908 1978
rect 1942 1872 2145 1978
rect 1825 1865 1865 1872
rect 1908 1865 2145 1872
rect 2375 1978 2492 1985
rect 2535 1978 2695 1985
rect 2375 1872 2458 1978
rect 2492 1872 2695 1978
rect 2375 1865 2415 1872
rect 2458 1865 2695 1872
rect 2925 1978 3042 1985
rect 3085 1978 3245 1985
rect 2925 1872 3008 1978
rect 3042 1872 3245 1978
rect 2925 1865 2965 1872
rect 3008 1865 3245 1872
rect 3475 1978 3592 1985
rect 3635 1978 3795 1985
rect 3475 1872 3558 1978
rect 3592 1872 3795 1978
rect 3475 1865 3515 1872
rect 3558 1865 3795 1872
rect 4025 1978 4142 1985
rect 4185 1978 4345 1985
rect 4025 1872 4108 1978
rect 4142 1872 4345 1978
rect 4025 1865 4065 1872
rect 4108 1865 4345 1872
rect 4575 1978 4692 1985
rect 4735 1978 4895 1985
rect 4575 1872 4658 1978
rect 4692 1872 4895 1978
rect 4575 1865 4615 1872
rect 4658 1865 4895 1872
rect 5125 1978 5242 1985
rect 5285 1978 5445 1985
rect 5125 1872 5208 1978
rect 5242 1872 5445 1978
rect 5125 1865 5165 1872
rect 5208 1865 5445 1872
rect 5675 1978 5792 1985
rect 5835 1978 5995 1985
rect 5675 1872 5758 1978
rect 5792 1872 5995 1978
rect 5675 1865 5715 1872
rect 5758 1865 5995 1872
rect 6225 1978 6342 1985
rect 6385 1978 6545 1985
rect 6225 1872 6308 1978
rect 6342 1872 6545 1978
rect 6225 1865 6265 1872
rect 6308 1865 6545 1872
rect 6775 1978 6892 1985
rect 6935 1978 7095 1985
rect 6775 1872 6858 1978
rect 6892 1872 7095 1978
rect 6775 1865 6815 1872
rect 6858 1865 7095 1872
rect 7325 1978 7442 1985
rect 7485 1978 7645 1985
rect 7325 1872 7408 1978
rect 7442 1872 7645 1978
rect 7325 1865 7365 1872
rect 7408 1865 7645 1872
rect 7875 1978 7992 1985
rect 8035 1978 8195 1985
rect 7875 1872 7958 1978
rect 7992 1872 8195 1978
rect 7875 1865 7915 1872
rect 7958 1865 8195 1872
rect 8425 1978 8542 1985
rect 8585 1978 8745 1985
rect 8425 1872 8508 1978
rect 8542 1872 8745 1978
rect 8425 1865 8465 1872
rect 8508 1865 8745 1872
rect 8975 1978 9092 1985
rect 9135 1978 9295 1985
rect 8975 1872 9058 1978
rect 9092 1872 9295 1978
rect 8975 1865 9015 1872
rect 9058 1865 9295 1872
rect 9525 1978 9642 1985
rect 9685 1978 9845 1985
rect 9525 1872 9608 1978
rect 9642 1872 9845 1978
rect 9525 1865 9565 1872
rect 9608 1865 9845 1872
rect 10075 1978 10192 1985
rect 10235 1978 10395 1985
rect 10075 1872 10158 1978
rect 10192 1872 10395 1978
rect 10075 1865 10115 1872
rect 10158 1865 10395 1872
rect 10625 1978 10742 1985
rect 10785 1978 10945 1985
rect 10625 1872 10708 1978
rect 10742 1872 10945 1978
rect 10625 1865 10665 1872
rect 10708 1865 10945 1872
rect 11175 1978 11292 1985
rect 11335 1978 11495 1985
rect 11175 1872 11258 1978
rect 11292 1872 11495 1978
rect 11175 1865 11215 1872
rect 11258 1865 11495 1872
rect 11725 1978 11842 1985
rect 11885 1978 12045 1985
rect 11725 1872 11808 1978
rect 11842 1872 12045 1978
rect 11725 1865 11765 1872
rect 11808 1865 12045 1872
rect 12275 1978 12392 1985
rect 12435 1978 12595 1985
rect 12275 1872 12358 1978
rect 12392 1872 12595 1978
rect 12275 1865 12315 1872
rect 12358 1865 12595 1872
rect 12825 1978 12942 1985
rect 12985 1978 13145 1985
rect 12825 1872 12908 1978
rect 12942 1872 13145 1978
rect 12825 1865 12865 1872
rect 12908 1865 13145 1872
rect 13375 1978 13492 1985
rect 13535 1978 13695 1985
rect 13375 1872 13458 1978
rect 13492 1872 13695 1978
rect 13375 1865 13415 1872
rect 13458 1865 13695 1872
rect 13925 1978 14042 1985
rect 14085 1978 14245 1985
rect 13925 1872 14008 1978
rect 14042 1872 14245 1978
rect 13925 1865 13965 1872
rect 14008 1865 14245 1872
rect 14475 1978 14592 1985
rect 14635 1978 14795 1985
rect 14475 1872 14558 1978
rect 14592 1872 14795 1978
rect 14475 1865 14515 1872
rect 14558 1865 14795 1872
rect 15025 1978 15142 1985
rect 15185 1978 15345 1985
rect 15025 1872 15108 1978
rect 15142 1872 15345 1978
rect 15025 1865 15065 1872
rect 15108 1865 15345 1872
rect 15575 1978 15692 1985
rect 15735 1978 15895 1985
rect 15575 1872 15658 1978
rect 15692 1872 15895 1978
rect 15575 1865 15615 1872
rect 15658 1865 15895 1872
rect 16125 1978 16242 1985
rect 16285 1978 16445 1985
rect 16125 1872 16208 1978
rect 16242 1872 16445 1978
rect 16125 1865 16165 1872
rect 16208 1865 16445 1872
rect 16675 1978 16792 1985
rect 16835 1978 16995 1985
rect 16675 1872 16758 1978
rect 16792 1872 16995 1978
rect 16675 1865 16715 1872
rect 16758 1865 16995 1872
rect 17225 1978 17342 1985
rect 17385 1978 17545 1985
rect 17225 1872 17308 1978
rect 17342 1872 17545 1978
rect 17225 1865 17265 1872
rect 17308 1865 17545 1872
rect 17775 1978 17892 1985
rect 17935 1978 18095 1985
rect 17775 1872 17858 1978
rect 17892 1872 18095 1978
rect 17775 1865 17815 1872
rect 17858 1865 18095 1872
rect 18325 1978 18442 1985
rect 18485 1978 18645 1985
rect 18325 1872 18408 1978
rect 18442 1872 18645 1978
rect 18325 1865 18365 1872
rect 18408 1865 18645 1872
rect 18875 1978 18992 1985
rect 19035 1978 19195 1985
rect 18875 1872 18958 1978
rect 18992 1872 19195 1978
rect 18875 1865 18915 1872
rect 18958 1865 19195 1872
rect 765 1825 885 1865
rect 1315 1825 1435 1865
rect 1865 1825 1985 1865
rect 2415 1825 2535 1865
rect 2965 1825 3085 1865
rect 3515 1825 3635 1865
rect 4065 1825 4185 1865
rect 4615 1825 4735 1865
rect 5165 1825 5285 1865
rect 5715 1825 5835 1865
rect 6265 1825 6385 1865
rect 6815 1825 6935 1865
rect 7365 1825 7485 1865
rect 7915 1825 8035 1865
rect 8465 1825 8585 1865
rect 9015 1825 9135 1865
rect 9565 1825 9685 1865
rect 10115 1825 10235 1865
rect 10665 1825 10785 1865
rect 11215 1825 11335 1865
rect 11765 1825 11885 1865
rect 12315 1825 12435 1865
rect 12865 1825 12985 1865
rect 13415 1825 13535 1865
rect 13965 1825 14085 1865
rect 14515 1825 14635 1865
rect 15065 1825 15185 1865
rect 15615 1825 15735 1865
rect 16165 1825 16285 1865
rect 16715 1825 16835 1865
rect 17265 1825 17385 1865
rect 17815 1825 17935 1865
rect 18365 1825 18485 1865
rect 18915 1825 19035 1865
rect 19202 1712 19204 2138
rect 500 1625 507 1675
rect 19202 1596 19217 1602
rect 628 1572 885 1595
rect 1178 1572 1435 1595
rect 1728 1572 1985 1595
rect 2278 1572 2535 1595
rect 2828 1572 3085 1595
rect 3378 1572 3635 1595
rect 3928 1572 4185 1595
rect 4478 1572 4735 1595
rect 5028 1572 5285 1595
rect 5578 1572 5835 1595
rect 6128 1572 6385 1595
rect 6678 1572 6935 1595
rect 7228 1572 7485 1595
rect 7778 1572 8035 1595
rect 8328 1572 8585 1595
rect 8878 1572 9135 1595
rect 9428 1572 9685 1595
rect 9978 1572 10235 1595
rect 10528 1572 10785 1595
rect 11078 1572 11335 1595
rect 11628 1572 11885 1595
rect 12178 1572 12435 1595
rect 12728 1572 12985 1595
rect 13278 1572 13535 1595
rect 13828 1572 14085 1595
rect 14378 1572 14635 1595
rect 14928 1572 15185 1595
rect 15478 1572 15735 1595
rect 16028 1572 16285 1595
rect 16578 1572 16835 1595
rect 17128 1572 17385 1595
rect 17678 1572 17935 1595
rect 18228 1572 18485 1595
rect 18778 1572 19035 1595
rect 605 1435 609 1572
rect 784 1475 885 1572
rect 765 1435 885 1475
rect 1155 1435 1159 1572
rect 1334 1475 1435 1572
rect 1315 1435 1435 1475
rect 1705 1435 1709 1572
rect 1884 1475 1985 1572
rect 1865 1435 1985 1475
rect 2255 1435 2259 1572
rect 2434 1475 2535 1572
rect 2415 1435 2535 1475
rect 2805 1435 2809 1572
rect 2984 1475 3085 1572
rect 2965 1435 3085 1475
rect 3355 1435 3359 1572
rect 3534 1475 3635 1572
rect 3515 1435 3635 1475
rect 3905 1435 3909 1572
rect 4084 1475 4185 1572
rect 4065 1435 4185 1475
rect 4455 1435 4459 1572
rect 4634 1475 4735 1572
rect 4615 1435 4735 1475
rect 5005 1435 5009 1572
rect 5184 1475 5285 1572
rect 5165 1435 5285 1475
rect 5555 1435 5559 1572
rect 5734 1475 5835 1572
rect 5715 1435 5835 1475
rect 6105 1435 6109 1572
rect 6284 1475 6385 1572
rect 6265 1435 6385 1475
rect 6655 1435 6659 1572
rect 6834 1475 6935 1572
rect 6815 1435 6935 1475
rect 7205 1435 7209 1572
rect 7384 1475 7485 1572
rect 7365 1435 7485 1475
rect 7755 1435 7759 1572
rect 7934 1475 8035 1572
rect 7915 1435 8035 1475
rect 8305 1435 8309 1572
rect 8484 1475 8585 1572
rect 8465 1435 8585 1475
rect 8855 1435 8859 1572
rect 9034 1475 9135 1572
rect 9015 1435 9135 1475
rect 9405 1435 9409 1572
rect 9584 1475 9685 1572
rect 9565 1435 9685 1475
rect 9955 1435 9959 1572
rect 10134 1475 10235 1572
rect 10115 1435 10235 1475
rect 10505 1435 10509 1572
rect 10684 1475 10785 1572
rect 10665 1435 10785 1475
rect 11055 1435 11059 1572
rect 11234 1475 11335 1572
rect 11215 1435 11335 1475
rect 11605 1435 11609 1572
rect 11784 1475 11885 1572
rect 11765 1435 11885 1475
rect 12155 1435 12159 1572
rect 12334 1475 12435 1572
rect 12315 1435 12435 1475
rect 12705 1435 12709 1572
rect 12884 1475 12985 1572
rect 12865 1435 12985 1475
rect 13255 1435 13259 1572
rect 13434 1475 13535 1572
rect 13415 1435 13535 1475
rect 13805 1435 13809 1572
rect 13984 1475 14085 1572
rect 13965 1435 14085 1475
rect 14355 1435 14359 1572
rect 14534 1475 14635 1572
rect 14515 1435 14635 1475
rect 14905 1435 14909 1572
rect 15084 1475 15185 1572
rect 15065 1435 15185 1475
rect 15455 1435 15459 1572
rect 15634 1475 15735 1572
rect 15615 1435 15735 1475
rect 16005 1435 16009 1572
rect 16184 1475 16285 1572
rect 16165 1435 16285 1475
rect 16555 1435 16559 1572
rect 16734 1475 16835 1572
rect 16715 1435 16835 1475
rect 17105 1435 17109 1572
rect 17284 1475 17385 1572
rect 17265 1435 17385 1475
rect 17655 1435 17659 1572
rect 17834 1475 17935 1572
rect 17815 1435 17935 1475
rect 18205 1435 18209 1572
rect 18384 1475 18485 1572
rect 18365 1435 18485 1475
rect 18755 1435 18759 1572
rect 18934 1475 19035 1572
rect 18915 1435 19035 1475
rect 725 1428 842 1435
rect 885 1428 1045 1435
rect 725 1322 808 1428
rect 842 1322 1045 1428
rect 725 1315 765 1322
rect 808 1315 1045 1322
rect 1275 1428 1392 1435
rect 1435 1428 1595 1435
rect 1275 1322 1358 1428
rect 1392 1322 1595 1428
rect 1275 1315 1315 1322
rect 1358 1315 1595 1322
rect 1825 1428 1942 1435
rect 1985 1428 2145 1435
rect 1825 1322 1908 1428
rect 1942 1322 2145 1428
rect 1825 1315 1865 1322
rect 1908 1315 2145 1322
rect 2375 1428 2492 1435
rect 2535 1428 2695 1435
rect 2375 1322 2458 1428
rect 2492 1322 2695 1428
rect 2375 1315 2415 1322
rect 2458 1315 2695 1322
rect 2925 1428 3042 1435
rect 3085 1428 3245 1435
rect 2925 1322 3008 1428
rect 3042 1322 3245 1428
rect 2925 1315 2965 1322
rect 3008 1315 3245 1322
rect 3475 1428 3592 1435
rect 3635 1428 3795 1435
rect 3475 1322 3558 1428
rect 3592 1322 3795 1428
rect 3475 1315 3515 1322
rect 3558 1315 3795 1322
rect 4025 1428 4142 1435
rect 4185 1428 4345 1435
rect 4025 1322 4108 1428
rect 4142 1322 4345 1428
rect 4025 1315 4065 1322
rect 4108 1315 4345 1322
rect 4575 1428 4692 1435
rect 4735 1428 4895 1435
rect 4575 1322 4658 1428
rect 4692 1322 4895 1428
rect 4575 1315 4615 1322
rect 4658 1315 4895 1322
rect 5125 1428 5242 1435
rect 5285 1428 5445 1435
rect 5125 1322 5208 1428
rect 5242 1322 5445 1428
rect 5125 1315 5165 1322
rect 5208 1315 5445 1322
rect 5675 1428 5792 1435
rect 5835 1428 5995 1435
rect 5675 1322 5758 1428
rect 5792 1322 5995 1428
rect 5675 1315 5715 1322
rect 5758 1315 5995 1322
rect 6225 1428 6342 1435
rect 6385 1428 6545 1435
rect 6225 1322 6308 1428
rect 6342 1322 6545 1428
rect 6225 1315 6265 1322
rect 6308 1315 6545 1322
rect 6775 1428 6892 1435
rect 6935 1428 7095 1435
rect 6775 1322 6858 1428
rect 6892 1322 7095 1428
rect 6775 1315 6815 1322
rect 6858 1315 7095 1322
rect 7325 1428 7442 1435
rect 7485 1428 7645 1435
rect 7325 1322 7408 1428
rect 7442 1322 7645 1428
rect 7325 1315 7365 1322
rect 7408 1315 7645 1322
rect 7875 1428 7992 1435
rect 8035 1428 8195 1435
rect 7875 1322 7958 1428
rect 7992 1322 8195 1428
rect 7875 1315 7915 1322
rect 7958 1315 8195 1322
rect 8425 1428 8542 1435
rect 8585 1428 8745 1435
rect 8425 1322 8508 1428
rect 8542 1322 8745 1428
rect 8425 1315 8465 1322
rect 8508 1315 8745 1322
rect 8975 1428 9092 1435
rect 9135 1428 9295 1435
rect 8975 1322 9058 1428
rect 9092 1322 9295 1428
rect 8975 1315 9015 1322
rect 9058 1315 9295 1322
rect 9525 1428 9642 1435
rect 9685 1428 9845 1435
rect 9525 1322 9608 1428
rect 9642 1322 9845 1428
rect 9525 1315 9565 1322
rect 9608 1315 9845 1322
rect 10075 1428 10192 1435
rect 10235 1428 10395 1435
rect 10075 1322 10158 1428
rect 10192 1322 10395 1428
rect 10075 1315 10115 1322
rect 10158 1315 10395 1322
rect 10625 1428 10742 1435
rect 10785 1428 10945 1435
rect 10625 1322 10708 1428
rect 10742 1322 10945 1428
rect 10625 1315 10665 1322
rect 10708 1315 10945 1322
rect 11175 1428 11292 1435
rect 11335 1428 11495 1435
rect 11175 1322 11258 1428
rect 11292 1322 11495 1428
rect 11175 1315 11215 1322
rect 11258 1315 11495 1322
rect 11725 1428 11842 1435
rect 11885 1428 12045 1435
rect 11725 1322 11808 1428
rect 11842 1322 12045 1428
rect 11725 1315 11765 1322
rect 11808 1315 12045 1322
rect 12275 1428 12392 1435
rect 12435 1428 12595 1435
rect 12275 1322 12358 1428
rect 12392 1322 12595 1428
rect 12275 1315 12315 1322
rect 12358 1315 12595 1322
rect 12825 1428 12942 1435
rect 12985 1428 13145 1435
rect 12825 1322 12908 1428
rect 12942 1322 13145 1428
rect 12825 1315 12865 1322
rect 12908 1315 13145 1322
rect 13375 1428 13492 1435
rect 13535 1428 13695 1435
rect 13375 1322 13458 1428
rect 13492 1322 13695 1428
rect 13375 1315 13415 1322
rect 13458 1315 13695 1322
rect 13925 1428 14042 1435
rect 14085 1428 14245 1435
rect 13925 1322 14008 1428
rect 14042 1322 14245 1428
rect 13925 1315 13965 1322
rect 14008 1315 14245 1322
rect 14475 1428 14592 1435
rect 14635 1428 14795 1435
rect 14475 1322 14558 1428
rect 14592 1322 14795 1428
rect 14475 1315 14515 1322
rect 14558 1315 14795 1322
rect 15025 1428 15142 1435
rect 15185 1428 15345 1435
rect 15025 1322 15108 1428
rect 15142 1322 15345 1428
rect 15025 1315 15065 1322
rect 15108 1315 15345 1322
rect 15575 1428 15692 1435
rect 15735 1428 15895 1435
rect 15575 1322 15658 1428
rect 15692 1322 15895 1428
rect 15575 1315 15615 1322
rect 15658 1315 15895 1322
rect 16125 1428 16242 1435
rect 16285 1428 16445 1435
rect 16125 1322 16208 1428
rect 16242 1322 16445 1428
rect 16125 1315 16165 1322
rect 16208 1315 16445 1322
rect 16675 1428 16792 1435
rect 16835 1428 16995 1435
rect 16675 1322 16758 1428
rect 16792 1322 16995 1428
rect 16675 1315 16715 1322
rect 16758 1315 16995 1322
rect 17225 1428 17342 1435
rect 17385 1428 17545 1435
rect 17225 1322 17308 1428
rect 17342 1322 17545 1428
rect 17225 1315 17265 1322
rect 17308 1315 17545 1322
rect 17775 1428 17892 1435
rect 17935 1428 18095 1435
rect 17775 1322 17858 1428
rect 17892 1322 18095 1428
rect 17775 1315 17815 1322
rect 17858 1315 18095 1322
rect 18325 1428 18442 1435
rect 18485 1428 18645 1435
rect 18325 1322 18408 1428
rect 18442 1322 18645 1428
rect 18325 1315 18365 1322
rect 18408 1315 18645 1322
rect 18875 1428 18992 1435
rect 19035 1428 19195 1435
rect 18875 1322 18958 1428
rect 18992 1322 19195 1428
rect 18875 1315 18915 1322
rect 18958 1315 19195 1322
rect 765 1275 885 1315
rect 1315 1275 1435 1315
rect 1865 1275 1985 1315
rect 2415 1275 2535 1315
rect 2965 1275 3085 1315
rect 3515 1275 3635 1315
rect 4065 1275 4185 1315
rect 4615 1275 4735 1315
rect 5165 1275 5285 1315
rect 5715 1275 5835 1315
rect 6265 1275 6385 1315
rect 6815 1275 6935 1315
rect 7365 1275 7485 1315
rect 7915 1275 8035 1315
rect 8465 1275 8585 1315
rect 9015 1275 9135 1315
rect 9565 1275 9685 1315
rect 10115 1275 10235 1315
rect 10665 1275 10785 1315
rect 11215 1275 11335 1315
rect 11765 1275 11885 1315
rect 12315 1275 12435 1315
rect 12865 1275 12985 1315
rect 13415 1275 13535 1315
rect 13965 1275 14085 1315
rect 14515 1275 14635 1315
rect 15065 1275 15185 1315
rect 15615 1275 15735 1315
rect 16165 1275 16285 1315
rect 16715 1275 16835 1315
rect 17265 1275 17385 1315
rect 17815 1275 17935 1315
rect 18365 1275 18485 1315
rect 18915 1275 19035 1315
rect 19185 1154 19200 1171
rect 19202 1162 19204 1588
rect 19202 1148 19217 1154
rect 500 1075 507 1125
rect 500 639 525 1040
rect 628 1022 885 1045
rect 1178 1022 1435 1045
rect 1728 1022 1985 1045
rect 2278 1022 2535 1045
rect 2828 1022 3085 1045
rect 3378 1022 3635 1045
rect 3928 1022 4185 1045
rect 4478 1022 4735 1045
rect 5028 1022 5285 1045
rect 5578 1022 5835 1045
rect 6128 1022 6385 1045
rect 6678 1022 6935 1045
rect 7228 1022 7485 1045
rect 7778 1022 8035 1045
rect 8328 1022 8585 1045
rect 8878 1022 9135 1045
rect 9428 1022 9685 1045
rect 9978 1022 10235 1045
rect 10528 1022 10785 1045
rect 11078 1022 11335 1045
rect 11628 1022 11885 1045
rect 12178 1022 12435 1045
rect 12728 1022 12985 1045
rect 13278 1022 13535 1045
rect 13828 1022 14085 1045
rect 14378 1022 14635 1045
rect 14928 1022 15185 1045
rect 15478 1022 15735 1045
rect 16028 1022 16285 1045
rect 16578 1022 16835 1045
rect 17128 1022 17385 1045
rect 17678 1022 17935 1045
rect 18228 1022 18485 1045
rect 18778 1022 19035 1045
rect 605 885 609 1022
rect 784 925 885 1022
rect 765 885 885 925
rect 1155 885 1159 1022
rect 1334 925 1435 1022
rect 1315 885 1435 925
rect 1705 885 1709 1022
rect 1884 925 1985 1022
rect 1865 885 1985 925
rect 2255 885 2259 1022
rect 2434 925 2535 1022
rect 2415 885 2535 925
rect 2805 885 2809 1022
rect 2984 925 3085 1022
rect 2965 885 3085 925
rect 3355 885 3359 1022
rect 3534 925 3635 1022
rect 3515 885 3635 925
rect 3905 885 3909 1022
rect 4084 925 4185 1022
rect 4065 885 4185 925
rect 4455 885 4459 1022
rect 4634 925 4735 1022
rect 4615 885 4735 925
rect 5005 885 5009 1022
rect 5184 925 5285 1022
rect 5165 885 5285 925
rect 5555 885 5559 1022
rect 5734 925 5835 1022
rect 5715 885 5835 925
rect 6105 885 6109 1022
rect 6284 925 6385 1022
rect 6265 885 6385 925
rect 6655 885 6659 1022
rect 6834 925 6935 1022
rect 6815 885 6935 925
rect 7205 885 7209 1022
rect 7384 925 7485 1022
rect 7365 885 7485 925
rect 7755 885 7759 1022
rect 7934 925 8035 1022
rect 7915 885 8035 925
rect 8305 885 8309 1022
rect 8484 925 8585 1022
rect 8465 885 8585 925
rect 8855 885 8859 1022
rect 9034 925 9135 1022
rect 9015 885 9135 925
rect 9405 885 9409 1022
rect 9584 925 9685 1022
rect 9565 885 9685 925
rect 9955 885 9959 1022
rect 10134 925 10235 1022
rect 10115 885 10235 925
rect 10505 885 10509 1022
rect 10684 925 10785 1022
rect 10665 885 10785 925
rect 11055 885 11059 1022
rect 11234 925 11335 1022
rect 11215 885 11335 925
rect 11605 885 11609 1022
rect 11784 925 11885 1022
rect 11765 885 11885 925
rect 12155 885 12159 1022
rect 12334 925 12435 1022
rect 12315 885 12435 925
rect 12705 885 12709 1022
rect 12884 925 12985 1022
rect 12865 885 12985 925
rect 13255 885 13259 1022
rect 13434 925 13535 1022
rect 13415 885 13535 925
rect 13805 885 13809 1022
rect 13984 925 14085 1022
rect 13965 885 14085 925
rect 14355 885 14359 1022
rect 14534 925 14635 1022
rect 14515 885 14635 925
rect 14905 885 14909 1022
rect 15084 925 15185 1022
rect 15065 885 15185 925
rect 15455 885 15459 1022
rect 15634 925 15735 1022
rect 15615 885 15735 925
rect 16005 885 16009 1022
rect 16184 925 16285 1022
rect 16165 885 16285 925
rect 16555 885 16559 1022
rect 16734 925 16835 1022
rect 16715 885 16835 925
rect 17105 885 17109 1022
rect 17284 925 17385 1022
rect 17265 885 17385 925
rect 17655 885 17659 1022
rect 17834 925 17935 1022
rect 17815 885 17935 925
rect 18205 885 18209 1022
rect 18384 925 18485 1022
rect 18365 885 18485 925
rect 18755 885 18759 1022
rect 18934 925 19035 1022
rect 18915 885 19035 925
rect 725 878 842 885
rect 885 878 1045 885
rect 725 772 808 878
rect 842 772 1045 878
rect 725 765 765 772
rect 808 765 1045 772
rect 1275 878 1392 885
rect 1435 878 1595 885
rect 1275 772 1358 878
rect 1392 772 1595 878
rect 1275 765 1315 772
rect 1358 765 1595 772
rect 1825 878 1942 885
rect 1985 878 2145 885
rect 1825 772 1908 878
rect 1942 772 2145 878
rect 1825 765 1865 772
rect 1908 765 2145 772
rect 2375 878 2492 885
rect 2535 878 2695 885
rect 2375 772 2458 878
rect 2492 772 2695 878
rect 2375 765 2415 772
rect 2458 765 2695 772
rect 2925 878 3042 885
rect 3085 878 3245 885
rect 2925 772 3008 878
rect 3042 772 3245 878
rect 2925 765 2965 772
rect 3008 765 3245 772
rect 3475 878 3592 885
rect 3635 878 3795 885
rect 3475 772 3558 878
rect 3592 772 3795 878
rect 3475 765 3515 772
rect 3558 765 3795 772
rect 4025 878 4142 885
rect 4185 878 4345 885
rect 4025 772 4108 878
rect 4142 772 4345 878
rect 4025 765 4065 772
rect 4108 765 4345 772
rect 4575 878 4692 885
rect 4735 878 4895 885
rect 4575 772 4658 878
rect 4692 772 4895 878
rect 4575 765 4615 772
rect 4658 765 4895 772
rect 5125 878 5242 885
rect 5285 878 5445 885
rect 5125 772 5208 878
rect 5242 772 5445 878
rect 5125 765 5165 772
rect 5208 765 5445 772
rect 5675 878 5792 885
rect 5835 878 5995 885
rect 5675 772 5758 878
rect 5792 772 5995 878
rect 5675 765 5715 772
rect 5758 765 5995 772
rect 6225 878 6342 885
rect 6385 878 6545 885
rect 6225 772 6308 878
rect 6342 772 6545 878
rect 6225 765 6265 772
rect 6308 765 6545 772
rect 6775 878 6892 885
rect 6935 878 7095 885
rect 6775 772 6858 878
rect 6892 772 7095 878
rect 6775 765 6815 772
rect 6858 765 7095 772
rect 7325 878 7442 885
rect 7485 878 7645 885
rect 7325 772 7408 878
rect 7442 772 7645 878
rect 7325 765 7365 772
rect 7408 765 7645 772
rect 7875 878 7992 885
rect 8035 878 8195 885
rect 7875 772 7958 878
rect 7992 772 8195 878
rect 7875 765 7915 772
rect 7958 765 8195 772
rect 8425 878 8542 885
rect 8585 878 8745 885
rect 8425 772 8508 878
rect 8542 772 8745 878
rect 8425 765 8465 772
rect 8508 765 8745 772
rect 8975 878 9092 885
rect 9135 878 9295 885
rect 8975 772 9058 878
rect 9092 772 9295 878
rect 8975 765 9015 772
rect 9058 765 9295 772
rect 9525 878 9642 885
rect 9685 878 9845 885
rect 9525 772 9608 878
rect 9642 772 9845 878
rect 9525 765 9565 772
rect 9608 765 9845 772
rect 10075 878 10192 885
rect 10235 878 10395 885
rect 10075 772 10158 878
rect 10192 772 10395 878
rect 10075 765 10115 772
rect 10158 765 10395 772
rect 10625 878 10742 885
rect 10785 878 10945 885
rect 10625 772 10708 878
rect 10742 772 10945 878
rect 10625 765 10665 772
rect 10708 765 10945 772
rect 11175 878 11292 885
rect 11335 878 11495 885
rect 11175 772 11258 878
rect 11292 772 11495 878
rect 11175 765 11215 772
rect 11258 765 11495 772
rect 11725 878 11842 885
rect 11885 878 12045 885
rect 11725 772 11808 878
rect 11842 772 12045 878
rect 11725 765 11765 772
rect 11808 765 12045 772
rect 12275 878 12392 885
rect 12435 878 12595 885
rect 12275 772 12358 878
rect 12392 772 12595 878
rect 12275 765 12315 772
rect 12358 765 12595 772
rect 12825 878 12942 885
rect 12985 878 13145 885
rect 12825 772 12908 878
rect 12942 772 13145 878
rect 12825 765 12865 772
rect 12908 765 13145 772
rect 13375 878 13492 885
rect 13535 878 13695 885
rect 13375 772 13458 878
rect 13492 772 13695 878
rect 13375 765 13415 772
rect 13458 765 13695 772
rect 13925 878 14042 885
rect 14085 878 14245 885
rect 13925 772 14008 878
rect 14042 772 14245 878
rect 13925 765 13965 772
rect 14008 765 14245 772
rect 14475 878 14592 885
rect 14635 878 14795 885
rect 14475 772 14558 878
rect 14592 772 14795 878
rect 14475 765 14515 772
rect 14558 765 14795 772
rect 15025 878 15142 885
rect 15185 878 15345 885
rect 15025 772 15108 878
rect 15142 772 15345 878
rect 15025 765 15065 772
rect 15108 765 15345 772
rect 15575 878 15692 885
rect 15735 878 15895 885
rect 15575 772 15658 878
rect 15692 772 15895 878
rect 15575 765 15615 772
rect 15658 765 15895 772
rect 16125 878 16242 885
rect 16285 878 16445 885
rect 16125 772 16208 878
rect 16242 772 16445 878
rect 16125 765 16165 772
rect 16208 765 16445 772
rect 16675 878 16792 885
rect 16835 878 16995 885
rect 16675 772 16758 878
rect 16792 772 16995 878
rect 16675 765 16715 772
rect 16758 765 16995 772
rect 17225 878 17342 885
rect 17385 878 17545 885
rect 17225 772 17308 878
rect 17342 772 17545 878
rect 17225 765 17265 772
rect 17308 765 17545 772
rect 17775 878 17892 885
rect 17935 878 18095 885
rect 17775 772 17858 878
rect 17892 772 18095 878
rect 17775 765 17815 772
rect 17858 765 18095 772
rect 18325 878 18442 885
rect 18485 878 18645 885
rect 18325 772 18408 878
rect 18442 772 18645 878
rect 18325 765 18365 772
rect 18408 765 18645 772
rect 18875 878 18992 885
rect 19035 878 19195 885
rect 18875 772 18958 878
rect 18992 772 19195 878
rect 18875 765 18915 772
rect 18958 765 19195 772
rect 765 725 885 765
rect 1315 725 1435 765
rect 1865 725 1985 765
rect 2415 725 2535 765
rect 2965 725 3085 765
rect 3515 725 3635 765
rect 4065 725 4185 765
rect 4615 725 4735 765
rect 5165 725 5285 765
rect 5715 725 5835 765
rect 6265 725 6385 765
rect 6815 725 6935 765
rect 7365 725 7485 765
rect 7915 725 8035 765
rect 8465 725 8585 765
rect 9015 725 9135 765
rect 9565 725 9685 765
rect 10115 725 10235 765
rect 10665 725 10785 765
rect 11215 725 11335 765
rect 11765 725 11885 765
rect 12315 725 12435 765
rect 12865 725 12985 765
rect 13415 725 13535 765
rect 13965 725 14085 765
rect 14515 725 14635 765
rect 15065 725 15185 765
rect 15615 725 15735 765
rect 16165 725 16285 765
rect 16715 725 16835 765
rect 17265 725 17385 765
rect 17815 725 17935 765
rect 18365 725 18485 765
rect 18915 725 19035 765
rect 19202 612 19204 1038
rect 500 525 507 575
rect 525 500 575 507
rect 610 500 1040 525
rect 1075 500 1125 507
rect 1625 500 1675 507
rect 1710 500 2140 525
rect 2175 500 2225 507
rect 2725 500 2775 507
rect 2810 500 3240 525
rect 3275 500 3325 507
rect 3825 500 3875 507
rect 3910 500 4340 525
rect 4375 500 4425 507
rect 4925 500 4975 507
rect 5010 500 5440 525
rect 5475 500 5525 507
rect 6025 500 6075 507
rect 6110 500 6540 525
rect 6575 500 6625 507
rect 7125 500 7175 507
rect 7210 500 7640 525
rect 7675 500 7725 507
rect 8225 500 8275 507
rect 8310 500 8740 525
rect 8775 500 8825 507
rect 9325 500 9375 507
rect 9410 500 9840 525
rect 9875 500 9925 507
rect 10425 500 10475 507
rect 10510 500 10940 525
rect 10975 500 11025 507
rect 11525 500 11575 507
rect 11610 500 12040 525
rect 12075 500 12125 507
rect 12625 500 12675 507
rect 12710 500 13140 525
rect 13175 500 13225 507
rect 13725 500 13775 507
rect 13810 500 14240 525
rect 14275 500 14325 507
rect 14825 500 14875 507
rect 14910 500 15340 525
rect 15375 500 15425 507
rect 15925 500 15975 507
rect 16010 500 16440 525
rect 16475 500 16525 507
rect 17025 500 17075 507
rect 17110 500 17540 525
rect 17575 500 17625 507
rect 18125 500 18175 507
rect 18210 500 18640 525
rect 18675 500 18725 507
rect 19202 500 19217 502
<< dnwell >>
rect -2950 19200 22750 22750
rect -2950 500 500 19200
rect 19200 500 22750 19200
rect -2950 -2950 22750 500
<< nwell >>
rect -5400 20400 25200 25200
rect -5400 -600 -600 20400
rect 20400 -600 25200 20400
rect -5400 -5400 25200 -600
<< pwell >>
rect -600 19200 20400 20400
rect -600 500 500 19200
rect 19200 500 20400 19200
rect -600 -600 20400 500
<< mvnmos >>
rect 525 19306 575 19744
rect 1075 19306 1125 19744
rect 1625 19306 1675 19744
rect 2175 19306 2225 19744
rect 2725 19306 2775 19744
rect 3275 19306 3325 19744
rect 3825 19306 3875 19744
rect 4375 19306 4425 19744
rect 4925 19306 4975 19744
rect 5475 19306 5525 19744
rect 6025 19306 6075 19744
rect 6575 19306 6625 19744
rect 7125 19306 7175 19744
rect 7675 19306 7725 19744
rect 8225 19306 8275 19744
rect 8775 19306 8825 19744
rect 9325 19306 9375 19744
rect 9875 19306 9925 19744
rect 10425 19306 10475 19744
rect 10975 19306 11025 19744
rect 11525 19306 11575 19744
rect 12075 19306 12125 19744
rect 12625 19306 12675 19744
rect 13175 19306 13225 19744
rect 13725 19306 13775 19744
rect 14275 19306 14325 19744
rect 14825 19306 14875 19744
rect 15375 19306 15425 19744
rect 15925 19306 15975 19744
rect 16475 19306 16525 19744
rect 17025 19306 17075 19744
rect 17575 19306 17625 19744
rect 18125 19306 18175 19744
rect 18675 19306 18725 19744
rect 19225 19306 19275 19744
rect 56 19225 494 19275
rect 606 19225 1044 19275
rect 1156 19225 1594 19275
rect 1706 19225 2144 19275
rect 2256 19225 2694 19275
rect 2806 19225 3244 19275
rect 3356 19225 3794 19275
rect 3906 19225 4344 19275
rect 4456 19225 4894 19275
rect 5006 19225 5444 19275
rect 5556 19225 5994 19275
rect 6106 19225 6544 19275
rect 6656 19225 7094 19275
rect 7206 19225 7644 19275
rect 7756 19225 8194 19275
rect 8306 19225 8744 19275
rect 8856 19225 9294 19275
rect 9406 19225 9844 19275
rect 9956 19225 10394 19275
rect 10506 19225 10944 19275
rect 11056 19225 11494 19275
rect 11606 19225 12044 19275
rect 12156 19225 12594 19275
rect 12706 19225 13144 19275
rect 13256 19225 13694 19275
rect 13806 19225 14244 19275
rect 14356 19225 14794 19275
rect 14906 19225 15344 19275
rect 15456 19225 15894 19275
rect 16006 19225 16444 19275
rect 16556 19225 16994 19275
rect 17106 19225 17544 19275
rect 17656 19225 18094 19275
rect 18206 19225 18644 19275
rect 18756 19225 19194 19275
rect 19306 19225 19744 19275
rect 19225 18756 19275 19194
rect 56 18675 494 18725
rect 19306 18675 19744 18725
rect 19225 18206 19275 18644
rect 56 18125 494 18175
rect 19306 18125 19744 18175
rect 19225 17656 19275 18094
rect 56 17575 494 17625
rect 19306 17575 19744 17625
rect 19225 17106 19275 17544
rect 56 17025 494 17075
rect 19306 17025 19744 17075
rect 19225 16556 19275 16994
rect 56 16475 494 16525
rect 19306 16475 19744 16525
rect 19225 16006 19275 16444
rect 56 15925 494 15975
rect 19306 15925 19744 15975
rect 19225 15456 19275 15894
rect 56 15375 494 15425
rect 19306 15375 19744 15425
rect 19225 14906 19275 15344
rect 56 14825 494 14875
rect 19306 14825 19744 14875
rect 19225 14356 19275 14794
rect 56 14275 494 14325
rect 19306 14275 19744 14325
rect 19225 13806 19275 14244
rect 56 13725 494 13775
rect 19306 13725 19744 13775
rect 19225 13256 19275 13694
rect 56 13175 494 13225
rect 19306 13175 19744 13225
rect 19225 12706 19275 13144
rect 56 12625 494 12675
rect 19306 12625 19744 12675
rect 19225 12156 19275 12594
rect 56 12075 494 12125
rect 19306 12075 19744 12125
rect 19225 11606 19275 12044
rect 56 11525 494 11575
rect 19306 11525 19744 11575
rect 19225 11056 19275 11494
rect 56 10975 494 11025
rect 19306 10975 19744 11025
rect 19225 10506 19275 10944
rect 56 10425 494 10475
rect 19306 10425 19744 10475
rect 19225 9956 19275 10394
rect 56 9875 494 9925
rect 19306 9875 19744 9925
rect 19225 9406 19275 9844
rect 56 9325 494 9375
rect 19306 9325 19744 9375
rect 19225 8856 19275 9294
rect 56 8775 494 8825
rect 19306 8775 19744 8825
rect 19225 8306 19275 8744
rect 56 8225 494 8275
rect 19306 8225 19744 8275
rect 19225 7756 19275 8194
rect 56 7675 494 7725
rect 19306 7675 19744 7725
rect 19225 7206 19275 7644
rect 56 7125 494 7175
rect 19306 7125 19744 7175
rect 19225 6656 19275 7094
rect 56 6575 494 6625
rect 19306 6575 19744 6625
rect 19225 6106 19275 6544
rect 56 6025 494 6075
rect 19306 6025 19744 6075
rect 19225 5556 19275 5994
rect 56 5475 494 5525
rect 19306 5475 19744 5525
rect 19225 5006 19275 5444
rect 56 4925 494 4975
rect 19306 4925 19744 4975
rect 19225 4456 19275 4894
rect 56 4375 494 4425
rect 19306 4375 19744 4425
rect 19225 3906 19275 4344
rect 56 3825 494 3875
rect 19306 3825 19744 3875
rect 19225 3356 19275 3794
rect 56 3275 494 3325
rect 19306 3275 19744 3325
rect 19225 2806 19275 3244
rect 56 2725 494 2775
rect 19306 2725 19744 2775
rect 19225 2256 19275 2694
rect 56 2175 494 2225
rect 19306 2175 19744 2225
rect 19225 1706 19275 2144
rect 56 1625 494 1675
rect 19306 1625 19744 1675
rect 19225 1156 19275 1594
rect 56 1075 494 1125
rect 19306 1075 19744 1125
rect 19225 606 19275 1044
rect 56 525 494 575
rect 19306 525 19744 575
rect 525 56 575 494
rect 1075 56 1125 494
rect 1625 56 1675 494
rect 2175 56 2225 494
rect 2725 56 2775 494
rect 3275 56 3325 494
rect 3825 56 3875 494
rect 4375 56 4425 494
rect 4925 56 4975 494
rect 5475 56 5525 494
rect 6025 56 6075 494
rect 6575 56 6625 494
rect 7125 56 7175 494
rect 7675 56 7725 494
rect 8225 56 8275 494
rect 8775 56 8825 494
rect 9325 56 9375 494
rect 9875 56 9925 494
rect 10425 56 10475 494
rect 10975 56 11025 494
rect 11525 56 11575 494
rect 12075 56 12125 494
rect 12625 56 12675 494
rect 13175 56 13225 494
rect 13725 56 13775 494
rect 14275 56 14325 494
rect 14825 56 14875 494
rect 15375 56 15425 494
rect 15925 56 15975 494
rect 16475 56 16525 494
rect 17025 56 17075 494
rect 17575 56 17625 494
rect 18125 56 18175 494
rect 18675 56 18725 494
rect 19225 56 19275 494
<< mvndiff >>
rect 604 19744 1046 19746
rect 1704 19744 2146 19746
rect 2804 19744 3246 19746
rect 3904 19744 4346 19746
rect 5004 19744 5446 19746
rect 6104 19744 6546 19746
rect 7204 19744 7646 19746
rect 8304 19744 8746 19746
rect 9404 19744 9846 19746
rect 10504 19744 10946 19746
rect 11604 19744 12046 19746
rect 12704 19744 13146 19746
rect 13804 19744 14246 19746
rect 14904 19744 15346 19746
rect 16004 19744 16446 19746
rect 17104 19744 17546 19746
rect 18204 19744 18646 19746
rect 19304 19744 19746 19746
rect 496 19738 525 19744
rect 496 19339 502 19738
rect 461 19312 502 19339
rect 519 19312 525 19738
rect 461 19306 525 19312
rect 575 19738 1075 19744
rect 575 19312 581 19738
rect 598 19690 1052 19738
rect 598 19360 660 19690
rect 990 19360 1052 19690
rect 598 19312 1052 19360
rect 1069 19312 1075 19738
rect 575 19306 1075 19312
rect 1125 19738 1154 19744
rect 1125 19312 1131 19738
rect 1148 19339 1154 19738
rect 1596 19738 1625 19744
rect 1596 19339 1602 19738
rect 1148 19312 1189 19339
rect 1125 19306 1189 19312
rect 461 19304 494 19306
rect 56 19298 494 19304
rect 56 19281 62 19298
rect 488 19281 494 19298
rect 56 19275 494 19281
rect 604 19304 1046 19306
rect 606 19298 1044 19304
rect 606 19281 612 19298
rect 1038 19281 1044 19298
rect 606 19275 1044 19281
rect 1156 19304 1189 19306
rect 1561 19312 1602 19339
rect 1619 19312 1625 19738
rect 1561 19306 1625 19312
rect 1675 19738 2175 19744
rect 1675 19312 1681 19738
rect 1698 19690 2152 19738
rect 1698 19360 1760 19690
rect 2090 19360 2152 19690
rect 1698 19312 2152 19360
rect 2169 19312 2175 19738
rect 1675 19306 2175 19312
rect 2225 19738 2254 19744
rect 2225 19312 2231 19738
rect 2248 19339 2254 19738
rect 2696 19738 2725 19744
rect 2696 19339 2702 19738
rect 2248 19312 2289 19339
rect 2225 19306 2289 19312
rect 1561 19304 1594 19306
rect 1156 19298 1594 19304
rect 1156 19281 1162 19298
rect 1588 19281 1594 19298
rect 1156 19275 1594 19281
rect 1704 19304 2146 19306
rect 1706 19298 2144 19304
rect 1706 19281 1712 19298
rect 2138 19281 2144 19298
rect 1706 19275 2144 19281
rect 2256 19304 2289 19306
rect 2661 19312 2702 19339
rect 2719 19312 2725 19738
rect 2661 19306 2725 19312
rect 2775 19738 3275 19744
rect 2775 19312 2781 19738
rect 2798 19690 3252 19738
rect 2798 19360 2860 19690
rect 3190 19360 3252 19690
rect 2798 19312 3252 19360
rect 3269 19312 3275 19738
rect 2775 19306 3275 19312
rect 3325 19738 3354 19744
rect 3325 19312 3331 19738
rect 3348 19339 3354 19738
rect 3796 19738 3825 19744
rect 3796 19339 3802 19738
rect 3348 19312 3389 19339
rect 3325 19306 3389 19312
rect 2661 19304 2694 19306
rect 2256 19298 2694 19304
rect 2256 19281 2262 19298
rect 2688 19281 2694 19298
rect 2256 19275 2694 19281
rect 2804 19304 3246 19306
rect 2806 19298 3244 19304
rect 2806 19281 2812 19298
rect 3238 19281 3244 19298
rect 2806 19275 3244 19281
rect 3356 19304 3389 19306
rect 3761 19312 3802 19339
rect 3819 19312 3825 19738
rect 3761 19306 3825 19312
rect 3875 19738 4375 19744
rect 3875 19312 3881 19738
rect 3898 19690 4352 19738
rect 3898 19360 3960 19690
rect 4290 19360 4352 19690
rect 3898 19312 4352 19360
rect 4369 19312 4375 19738
rect 3875 19306 4375 19312
rect 4425 19738 4454 19744
rect 4425 19312 4431 19738
rect 4448 19339 4454 19738
rect 4896 19738 4925 19744
rect 4896 19339 4902 19738
rect 4448 19312 4489 19339
rect 4425 19306 4489 19312
rect 3761 19304 3794 19306
rect 3356 19298 3794 19304
rect 3356 19281 3362 19298
rect 3788 19281 3794 19298
rect 3356 19275 3794 19281
rect 3904 19304 4346 19306
rect 3906 19298 4344 19304
rect 3906 19281 3912 19298
rect 4338 19281 4344 19298
rect 3906 19275 4344 19281
rect 4456 19304 4489 19306
rect 4861 19312 4902 19339
rect 4919 19312 4925 19738
rect 4861 19306 4925 19312
rect 4975 19738 5475 19744
rect 4975 19312 4981 19738
rect 4998 19690 5452 19738
rect 4998 19360 5060 19690
rect 5390 19360 5452 19690
rect 4998 19312 5452 19360
rect 5469 19312 5475 19738
rect 4975 19306 5475 19312
rect 5525 19738 5554 19744
rect 5525 19312 5531 19738
rect 5548 19339 5554 19738
rect 5996 19738 6025 19744
rect 5996 19339 6002 19738
rect 5548 19312 5589 19339
rect 5525 19306 5589 19312
rect 4861 19304 4894 19306
rect 4456 19298 4894 19304
rect 4456 19281 4462 19298
rect 4888 19281 4894 19298
rect 4456 19275 4894 19281
rect 5004 19304 5446 19306
rect 5006 19298 5444 19304
rect 5006 19281 5012 19298
rect 5438 19281 5444 19298
rect 5006 19275 5444 19281
rect 5556 19304 5589 19306
rect 5961 19312 6002 19339
rect 6019 19312 6025 19738
rect 5961 19306 6025 19312
rect 6075 19738 6575 19744
rect 6075 19312 6081 19738
rect 6098 19690 6552 19738
rect 6098 19360 6160 19690
rect 6490 19360 6552 19690
rect 6098 19312 6552 19360
rect 6569 19312 6575 19738
rect 6075 19306 6575 19312
rect 6625 19738 6654 19744
rect 6625 19312 6631 19738
rect 6648 19339 6654 19738
rect 7096 19738 7125 19744
rect 7096 19339 7102 19738
rect 6648 19312 6689 19339
rect 6625 19306 6689 19312
rect 5961 19304 5994 19306
rect 5556 19298 5994 19304
rect 5556 19281 5562 19298
rect 5988 19281 5994 19298
rect 5556 19275 5994 19281
rect 6104 19304 6546 19306
rect 6106 19298 6544 19304
rect 6106 19281 6112 19298
rect 6538 19281 6544 19298
rect 6106 19275 6544 19281
rect 6656 19304 6689 19306
rect 7061 19312 7102 19339
rect 7119 19312 7125 19738
rect 7061 19306 7125 19312
rect 7175 19738 7675 19744
rect 7175 19312 7181 19738
rect 7198 19690 7652 19738
rect 7198 19360 7260 19690
rect 7590 19360 7652 19690
rect 7198 19312 7652 19360
rect 7669 19312 7675 19738
rect 7175 19306 7675 19312
rect 7725 19738 7754 19744
rect 7725 19312 7731 19738
rect 7748 19339 7754 19738
rect 8196 19738 8225 19744
rect 8196 19339 8202 19738
rect 7748 19312 7789 19339
rect 7725 19306 7789 19312
rect 7061 19304 7094 19306
rect 6656 19298 7094 19304
rect 6656 19281 6662 19298
rect 7088 19281 7094 19298
rect 6656 19275 7094 19281
rect 7204 19304 7646 19306
rect 7206 19298 7644 19304
rect 7206 19281 7212 19298
rect 7638 19281 7644 19298
rect 7206 19275 7644 19281
rect 7756 19304 7789 19306
rect 8161 19312 8202 19339
rect 8219 19312 8225 19738
rect 8161 19306 8225 19312
rect 8275 19738 8775 19744
rect 8275 19312 8281 19738
rect 8298 19690 8752 19738
rect 8298 19360 8360 19690
rect 8690 19360 8752 19690
rect 8298 19312 8752 19360
rect 8769 19312 8775 19738
rect 8275 19306 8775 19312
rect 8825 19738 8854 19744
rect 8825 19312 8831 19738
rect 8848 19339 8854 19738
rect 9296 19738 9325 19744
rect 9296 19339 9302 19738
rect 8848 19312 8889 19339
rect 8825 19306 8889 19312
rect 8161 19304 8194 19306
rect 7756 19298 8194 19304
rect 7756 19281 7762 19298
rect 8188 19281 8194 19298
rect 7756 19275 8194 19281
rect 8304 19304 8746 19306
rect 8306 19298 8744 19304
rect 8306 19281 8312 19298
rect 8738 19281 8744 19298
rect 8306 19275 8744 19281
rect 8856 19304 8889 19306
rect 9261 19312 9302 19339
rect 9319 19312 9325 19738
rect 9261 19306 9325 19312
rect 9375 19738 9875 19744
rect 9375 19312 9381 19738
rect 9398 19690 9852 19738
rect 9398 19360 9460 19690
rect 9790 19360 9852 19690
rect 9398 19312 9852 19360
rect 9869 19312 9875 19738
rect 9375 19306 9875 19312
rect 9925 19738 9954 19744
rect 9925 19312 9931 19738
rect 9948 19339 9954 19738
rect 10396 19738 10425 19744
rect 10396 19339 10402 19738
rect 9948 19312 9989 19339
rect 9925 19306 9989 19312
rect 9261 19304 9294 19306
rect 8856 19298 9294 19304
rect 8856 19281 8862 19298
rect 9288 19281 9294 19298
rect 8856 19275 9294 19281
rect 9404 19304 9846 19306
rect 9406 19298 9844 19304
rect 9406 19281 9412 19298
rect 9838 19281 9844 19298
rect 9406 19275 9844 19281
rect 9956 19304 9989 19306
rect 10361 19312 10402 19339
rect 10419 19312 10425 19738
rect 10361 19306 10425 19312
rect 10475 19738 10975 19744
rect 10475 19312 10481 19738
rect 10498 19690 10952 19738
rect 10498 19360 10560 19690
rect 10890 19360 10952 19690
rect 10498 19312 10952 19360
rect 10969 19312 10975 19738
rect 10475 19306 10975 19312
rect 11025 19738 11054 19744
rect 11025 19312 11031 19738
rect 11048 19339 11054 19738
rect 11496 19738 11525 19744
rect 11496 19339 11502 19738
rect 11048 19312 11089 19339
rect 11025 19306 11089 19312
rect 10361 19304 10394 19306
rect 9956 19298 10394 19304
rect 9956 19281 9962 19298
rect 10388 19281 10394 19298
rect 9956 19275 10394 19281
rect 10504 19304 10946 19306
rect 10506 19298 10944 19304
rect 10506 19281 10512 19298
rect 10938 19281 10944 19298
rect 10506 19275 10944 19281
rect 11056 19304 11089 19306
rect 11461 19312 11502 19339
rect 11519 19312 11525 19738
rect 11461 19306 11525 19312
rect 11575 19738 12075 19744
rect 11575 19312 11581 19738
rect 11598 19690 12052 19738
rect 11598 19360 11660 19690
rect 11990 19360 12052 19690
rect 11598 19312 12052 19360
rect 12069 19312 12075 19738
rect 11575 19306 12075 19312
rect 12125 19738 12154 19744
rect 12125 19312 12131 19738
rect 12148 19339 12154 19738
rect 12596 19738 12625 19744
rect 12596 19339 12602 19738
rect 12148 19312 12189 19339
rect 12125 19306 12189 19312
rect 11461 19304 11494 19306
rect 11056 19298 11494 19304
rect 11056 19281 11062 19298
rect 11488 19281 11494 19298
rect 11056 19275 11494 19281
rect 11604 19304 12046 19306
rect 11606 19298 12044 19304
rect 11606 19281 11612 19298
rect 12038 19281 12044 19298
rect 11606 19275 12044 19281
rect 12156 19304 12189 19306
rect 12561 19312 12602 19339
rect 12619 19312 12625 19738
rect 12561 19306 12625 19312
rect 12675 19738 13175 19744
rect 12675 19312 12681 19738
rect 12698 19690 13152 19738
rect 12698 19360 12760 19690
rect 13090 19360 13152 19690
rect 12698 19312 13152 19360
rect 13169 19312 13175 19738
rect 12675 19306 13175 19312
rect 13225 19738 13254 19744
rect 13225 19312 13231 19738
rect 13248 19339 13254 19738
rect 13696 19738 13725 19744
rect 13696 19339 13702 19738
rect 13248 19312 13289 19339
rect 13225 19306 13289 19312
rect 12561 19304 12594 19306
rect 12156 19298 12594 19304
rect 12156 19281 12162 19298
rect 12588 19281 12594 19298
rect 12156 19275 12594 19281
rect 12704 19304 13146 19306
rect 12706 19298 13144 19304
rect 12706 19281 12712 19298
rect 13138 19281 13144 19298
rect 12706 19275 13144 19281
rect 13256 19304 13289 19306
rect 13661 19312 13702 19339
rect 13719 19312 13725 19738
rect 13661 19306 13725 19312
rect 13775 19738 14275 19744
rect 13775 19312 13781 19738
rect 13798 19690 14252 19738
rect 13798 19360 13860 19690
rect 14190 19360 14252 19690
rect 13798 19312 14252 19360
rect 14269 19312 14275 19738
rect 13775 19306 14275 19312
rect 14325 19738 14354 19744
rect 14325 19312 14331 19738
rect 14348 19339 14354 19738
rect 14796 19738 14825 19744
rect 14796 19339 14802 19738
rect 14348 19312 14389 19339
rect 14325 19306 14389 19312
rect 13661 19304 13694 19306
rect 13256 19298 13694 19304
rect 13256 19281 13262 19298
rect 13688 19281 13694 19298
rect 13256 19275 13694 19281
rect 13804 19304 14246 19306
rect 13806 19298 14244 19304
rect 13806 19281 13812 19298
rect 14238 19281 14244 19298
rect 13806 19275 14244 19281
rect 14356 19304 14389 19306
rect 14761 19312 14802 19339
rect 14819 19312 14825 19738
rect 14761 19306 14825 19312
rect 14875 19738 15375 19744
rect 14875 19312 14881 19738
rect 14898 19690 15352 19738
rect 14898 19360 14960 19690
rect 15290 19360 15352 19690
rect 14898 19312 15352 19360
rect 15369 19312 15375 19738
rect 14875 19306 15375 19312
rect 15425 19738 15454 19744
rect 15425 19312 15431 19738
rect 15448 19339 15454 19738
rect 15896 19738 15925 19744
rect 15896 19339 15902 19738
rect 15448 19312 15489 19339
rect 15425 19306 15489 19312
rect 14761 19304 14794 19306
rect 14356 19298 14794 19304
rect 14356 19281 14362 19298
rect 14788 19281 14794 19298
rect 14356 19275 14794 19281
rect 14904 19304 15346 19306
rect 14906 19298 15344 19304
rect 14906 19281 14912 19298
rect 15338 19281 15344 19298
rect 14906 19275 15344 19281
rect 15456 19304 15489 19306
rect 15861 19312 15902 19339
rect 15919 19312 15925 19738
rect 15861 19306 15925 19312
rect 15975 19738 16475 19744
rect 15975 19312 15981 19738
rect 15998 19690 16452 19738
rect 15998 19360 16060 19690
rect 16390 19360 16452 19690
rect 15998 19312 16452 19360
rect 16469 19312 16475 19738
rect 15975 19306 16475 19312
rect 16525 19738 16554 19744
rect 16525 19312 16531 19738
rect 16548 19339 16554 19738
rect 16996 19738 17025 19744
rect 16996 19339 17002 19738
rect 16548 19312 16589 19339
rect 16525 19306 16589 19312
rect 15861 19304 15894 19306
rect 15456 19298 15894 19304
rect 15456 19281 15462 19298
rect 15888 19281 15894 19298
rect 15456 19275 15894 19281
rect 16004 19304 16446 19306
rect 16006 19298 16444 19304
rect 16006 19281 16012 19298
rect 16438 19281 16444 19298
rect 16006 19275 16444 19281
rect 16556 19304 16589 19306
rect 16961 19312 17002 19339
rect 17019 19312 17025 19738
rect 16961 19306 17025 19312
rect 17075 19738 17575 19744
rect 17075 19312 17081 19738
rect 17098 19690 17552 19738
rect 17098 19360 17160 19690
rect 17490 19360 17552 19690
rect 17098 19312 17552 19360
rect 17569 19312 17575 19738
rect 17075 19306 17575 19312
rect 17625 19738 17654 19744
rect 17625 19312 17631 19738
rect 17648 19339 17654 19738
rect 18096 19738 18125 19744
rect 18096 19339 18102 19738
rect 17648 19312 17689 19339
rect 17625 19306 17689 19312
rect 16961 19304 16994 19306
rect 16556 19298 16994 19304
rect 16556 19281 16562 19298
rect 16988 19281 16994 19298
rect 16556 19275 16994 19281
rect 17104 19304 17546 19306
rect 17106 19298 17544 19304
rect 17106 19281 17112 19298
rect 17538 19281 17544 19298
rect 17106 19275 17544 19281
rect 17656 19304 17689 19306
rect 18061 19312 18102 19339
rect 18119 19312 18125 19738
rect 18061 19306 18125 19312
rect 18175 19738 18675 19744
rect 18175 19312 18181 19738
rect 18198 19690 18652 19738
rect 18198 19360 18260 19690
rect 18590 19360 18652 19690
rect 18198 19312 18652 19360
rect 18669 19312 18675 19738
rect 18175 19306 18675 19312
rect 18725 19738 18754 19744
rect 18725 19312 18731 19738
rect 18748 19339 18754 19738
rect 19196 19738 19225 19744
rect 19196 19339 19202 19738
rect 18748 19312 18789 19339
rect 18725 19306 18789 19312
rect 18061 19304 18094 19306
rect 17656 19298 18094 19304
rect 17656 19281 17662 19298
rect 18088 19281 18094 19298
rect 17656 19275 18094 19281
rect 18204 19304 18646 19306
rect 18206 19298 18644 19304
rect 18206 19281 18212 19298
rect 18638 19281 18644 19298
rect 18206 19275 18644 19281
rect 18756 19304 18789 19306
rect 19161 19312 19202 19339
rect 19219 19312 19225 19738
rect 19161 19306 19225 19312
rect 19275 19738 19746 19744
rect 19275 19312 19281 19738
rect 19298 19690 19746 19738
rect 19298 19360 19360 19690
rect 19690 19360 19746 19690
rect 19298 19312 19746 19360
rect 19275 19306 19746 19312
rect 19161 19304 19194 19306
rect 18756 19298 19194 19304
rect 18756 19281 18762 19298
rect 19188 19281 19194 19298
rect 18756 19275 19194 19281
rect 19304 19304 19746 19306
rect 19306 19298 19744 19304
rect 19306 19281 19312 19298
rect 19738 19281 19744 19298
rect 19306 19275 19744 19281
rect 56 19219 494 19225
rect 56 19202 62 19219
rect 488 19202 494 19219
rect 56 19196 494 19202
rect 606 19219 1044 19225
rect 606 19202 612 19219
rect 1038 19202 1044 19219
rect 606 19200 1044 19202
rect 1156 19219 1594 19225
rect 1156 19202 1162 19219
rect 1588 19202 1594 19219
rect 1156 19200 1594 19202
rect 1706 19219 2144 19225
rect 1706 19202 1712 19219
rect 2138 19202 2144 19219
rect 1706 19200 2144 19202
rect 2256 19219 2694 19225
rect 2256 19202 2262 19219
rect 2688 19202 2694 19219
rect 2256 19200 2694 19202
rect 2806 19219 3244 19225
rect 2806 19202 2812 19219
rect 3238 19202 3244 19219
rect 2806 19200 3244 19202
rect 3356 19219 3794 19225
rect 3356 19202 3362 19219
rect 3788 19202 3794 19219
rect 3356 19200 3794 19202
rect 3906 19219 4344 19225
rect 3906 19202 3912 19219
rect 4338 19202 4344 19219
rect 3906 19200 4344 19202
rect 4456 19219 4894 19225
rect 4456 19202 4462 19219
rect 4888 19202 4894 19219
rect 4456 19200 4894 19202
rect 5006 19219 5444 19225
rect 5006 19202 5012 19219
rect 5438 19202 5444 19219
rect 5006 19200 5444 19202
rect 5556 19219 5994 19225
rect 5556 19202 5562 19219
rect 5988 19202 5994 19219
rect 5556 19200 5994 19202
rect 6106 19219 6544 19225
rect 6106 19202 6112 19219
rect 6538 19202 6544 19219
rect 6106 19200 6544 19202
rect 6656 19219 7094 19225
rect 6656 19202 6662 19219
rect 7088 19202 7094 19219
rect 6656 19200 7094 19202
rect 7206 19219 7644 19225
rect 7206 19202 7212 19219
rect 7638 19202 7644 19219
rect 7206 19200 7644 19202
rect 7756 19219 8194 19225
rect 7756 19202 7762 19219
rect 8188 19202 8194 19219
rect 7756 19200 8194 19202
rect 8306 19219 8744 19225
rect 8306 19202 8312 19219
rect 8738 19202 8744 19219
rect 8306 19200 8744 19202
rect 8856 19219 9294 19225
rect 8856 19202 8862 19219
rect 9288 19202 9294 19219
rect 8856 19200 9294 19202
rect 9406 19219 9844 19225
rect 9406 19202 9412 19219
rect 9838 19202 9844 19219
rect 9406 19200 9844 19202
rect 9956 19219 10394 19225
rect 9956 19202 9962 19219
rect 10388 19202 10394 19219
rect 9956 19200 10394 19202
rect 10506 19219 10944 19225
rect 10506 19202 10512 19219
rect 10938 19202 10944 19219
rect 10506 19200 10944 19202
rect 11056 19219 11494 19225
rect 11056 19202 11062 19219
rect 11488 19202 11494 19219
rect 11056 19200 11494 19202
rect 11606 19219 12044 19225
rect 11606 19202 11612 19219
rect 12038 19202 12044 19219
rect 11606 19200 12044 19202
rect 12156 19219 12594 19225
rect 12156 19202 12162 19219
rect 12588 19202 12594 19219
rect 12156 19200 12594 19202
rect 12706 19219 13144 19225
rect 12706 19202 12712 19219
rect 13138 19202 13144 19219
rect 12706 19200 13144 19202
rect 13256 19219 13694 19225
rect 13256 19202 13262 19219
rect 13688 19202 13694 19219
rect 13256 19200 13694 19202
rect 13806 19219 14244 19225
rect 13806 19202 13812 19219
rect 14238 19202 14244 19219
rect 13806 19200 14244 19202
rect 14356 19219 14794 19225
rect 14356 19202 14362 19219
rect 14788 19202 14794 19219
rect 14356 19200 14794 19202
rect 14906 19219 15344 19225
rect 14906 19202 14912 19219
rect 15338 19202 15344 19219
rect 14906 19200 15344 19202
rect 15456 19219 15894 19225
rect 15456 19202 15462 19219
rect 15888 19202 15894 19219
rect 15456 19200 15894 19202
rect 16006 19219 16444 19225
rect 16006 19202 16012 19219
rect 16438 19202 16444 19219
rect 16006 19200 16444 19202
rect 16556 19219 16994 19225
rect 16556 19202 16562 19219
rect 16988 19202 16994 19219
rect 16556 19200 16994 19202
rect 17106 19219 17544 19225
rect 17106 19202 17112 19219
rect 17538 19202 17544 19219
rect 17106 19200 17544 19202
rect 17656 19219 18094 19225
rect 17656 19202 17662 19219
rect 18088 19202 18094 19219
rect 17656 19200 18094 19202
rect 18206 19219 18644 19225
rect 18206 19202 18212 19219
rect 18638 19202 18644 19219
rect 18206 19200 18644 19202
rect 18756 19219 19194 19225
rect 18756 19202 18762 19219
rect 19188 19202 19194 19219
rect 18756 19200 19194 19202
rect 54 19194 496 19196
rect 19306 19219 19744 19225
rect 19306 19202 19312 19219
rect 19738 19202 19744 19219
rect 19306 19196 19744 19202
rect 19306 19194 19339 19196
rect 54 19140 500 19194
rect 54 18810 110 19140
rect 440 18810 500 19140
rect 54 18756 500 18810
rect 19200 19188 19225 19194
rect 19200 18762 19202 19188
rect 19219 18762 19225 19188
rect 19200 18756 19225 18762
rect 19275 19188 19339 19194
rect 19275 18762 19281 19188
rect 19298 19161 19339 19188
rect 19298 18789 19304 19161
rect 19298 18762 19339 18789
rect 19275 18756 19339 18762
rect 54 18754 496 18756
rect 56 18748 494 18754
rect 56 18731 62 18748
rect 488 18731 494 18748
rect 56 18725 494 18731
rect 19306 18754 19339 18756
rect 19306 18748 19744 18754
rect 19306 18731 19312 18748
rect 19738 18731 19744 18748
rect 19306 18725 19744 18731
rect 56 18669 494 18675
rect 56 18652 62 18669
rect 488 18652 494 18669
rect 56 18646 494 18652
rect 461 18644 494 18646
rect 19306 18669 19744 18675
rect 19306 18652 19312 18669
rect 19738 18652 19744 18669
rect 19306 18646 19744 18652
rect 19304 18644 19746 18646
rect 461 18611 500 18644
rect 496 18239 500 18611
rect 461 18206 500 18239
rect 19200 18638 19225 18644
rect 19200 18212 19202 18638
rect 19219 18212 19225 18638
rect 19200 18206 19225 18212
rect 19275 18638 19746 18644
rect 19275 18212 19281 18638
rect 19298 18590 19746 18638
rect 19298 18260 19360 18590
rect 19690 18260 19746 18590
rect 19298 18212 19746 18260
rect 19275 18206 19746 18212
rect 461 18204 494 18206
rect 56 18198 494 18204
rect 56 18181 62 18198
rect 488 18181 494 18198
rect 56 18175 494 18181
rect 19304 18204 19746 18206
rect 19306 18198 19744 18204
rect 19306 18181 19312 18198
rect 19738 18181 19744 18198
rect 19306 18175 19744 18181
rect 56 18119 494 18125
rect 56 18102 62 18119
rect 488 18102 494 18119
rect 56 18096 494 18102
rect 54 18094 496 18096
rect 19306 18119 19744 18125
rect 19306 18102 19312 18119
rect 19738 18102 19744 18119
rect 19306 18096 19744 18102
rect 19306 18094 19339 18096
rect 54 18040 500 18094
rect 54 17710 110 18040
rect 440 17710 500 18040
rect 54 17656 500 17710
rect 19200 18088 19225 18094
rect 19200 17662 19202 18088
rect 19219 17662 19225 18088
rect 19200 17656 19225 17662
rect 19275 18088 19339 18094
rect 19275 17662 19281 18088
rect 19298 18061 19339 18088
rect 19298 17689 19304 18061
rect 19298 17662 19339 17689
rect 19275 17656 19339 17662
rect 54 17654 496 17656
rect 56 17648 494 17654
rect 56 17631 62 17648
rect 488 17631 494 17648
rect 56 17625 494 17631
rect 19306 17654 19339 17656
rect 19306 17648 19744 17654
rect 19306 17631 19312 17648
rect 19738 17631 19744 17648
rect 19306 17625 19744 17631
rect 56 17569 494 17575
rect 56 17552 62 17569
rect 488 17552 494 17569
rect 56 17546 494 17552
rect 461 17544 494 17546
rect 19306 17569 19744 17575
rect 19306 17552 19312 17569
rect 19738 17552 19744 17569
rect 19306 17546 19744 17552
rect 19304 17544 19746 17546
rect 461 17511 500 17544
rect 496 17139 500 17511
rect 461 17106 500 17139
rect 19200 17538 19225 17544
rect 19200 17112 19202 17538
rect 19219 17112 19225 17538
rect 19200 17106 19225 17112
rect 19275 17538 19746 17544
rect 19275 17112 19281 17538
rect 19298 17490 19746 17538
rect 19298 17160 19360 17490
rect 19690 17160 19746 17490
rect 19298 17112 19746 17160
rect 19275 17106 19746 17112
rect 461 17104 494 17106
rect 56 17098 494 17104
rect 56 17081 62 17098
rect 488 17081 494 17098
rect 56 17075 494 17081
rect 19304 17104 19746 17106
rect 19306 17098 19744 17104
rect 19306 17081 19312 17098
rect 19738 17081 19744 17098
rect 19306 17075 19744 17081
rect 56 17019 494 17025
rect 56 17002 62 17019
rect 488 17002 494 17019
rect 56 16996 494 17002
rect 54 16994 496 16996
rect 19306 17019 19744 17025
rect 19306 17002 19312 17019
rect 19738 17002 19744 17019
rect 19306 16996 19744 17002
rect 19306 16994 19339 16996
rect 54 16940 500 16994
rect 54 16610 110 16940
rect 440 16610 500 16940
rect 54 16556 500 16610
rect 19200 16988 19225 16994
rect 19200 16562 19202 16988
rect 19219 16562 19225 16988
rect 19200 16556 19225 16562
rect 19275 16988 19339 16994
rect 19275 16562 19281 16988
rect 19298 16961 19339 16988
rect 19298 16589 19304 16961
rect 19298 16562 19339 16589
rect 19275 16556 19339 16562
rect 54 16554 496 16556
rect 56 16548 494 16554
rect 56 16531 62 16548
rect 488 16531 494 16548
rect 56 16525 494 16531
rect 19306 16554 19339 16556
rect 19306 16548 19744 16554
rect 19306 16531 19312 16548
rect 19738 16531 19744 16548
rect 19306 16525 19744 16531
rect 56 16469 494 16475
rect 56 16452 62 16469
rect 488 16452 494 16469
rect 56 16446 494 16452
rect 461 16444 494 16446
rect 19306 16469 19744 16475
rect 19306 16452 19312 16469
rect 19738 16452 19744 16469
rect 19306 16446 19744 16452
rect 19304 16444 19746 16446
rect 461 16411 500 16444
rect 496 16039 500 16411
rect 461 16006 500 16039
rect 19200 16438 19225 16444
rect 19200 16012 19202 16438
rect 19219 16012 19225 16438
rect 19200 16006 19225 16012
rect 19275 16438 19746 16444
rect 19275 16012 19281 16438
rect 19298 16390 19746 16438
rect 19298 16060 19360 16390
rect 19690 16060 19746 16390
rect 19298 16012 19746 16060
rect 19275 16006 19746 16012
rect 461 16004 494 16006
rect 56 15998 494 16004
rect 56 15981 62 15998
rect 488 15981 494 15998
rect 56 15975 494 15981
rect 19304 16004 19746 16006
rect 19306 15998 19744 16004
rect 19306 15981 19312 15998
rect 19738 15981 19744 15998
rect 19306 15975 19744 15981
rect 56 15919 494 15925
rect 56 15902 62 15919
rect 488 15902 494 15919
rect 56 15896 494 15902
rect 54 15894 496 15896
rect 19306 15919 19744 15925
rect 19306 15902 19312 15919
rect 19738 15902 19744 15919
rect 19306 15896 19744 15902
rect 19306 15894 19339 15896
rect 54 15840 500 15894
rect 54 15510 110 15840
rect 440 15510 500 15840
rect 54 15456 500 15510
rect 19200 15888 19225 15894
rect 19200 15462 19202 15888
rect 19219 15462 19225 15888
rect 19200 15456 19225 15462
rect 19275 15888 19339 15894
rect 19275 15462 19281 15888
rect 19298 15861 19339 15888
rect 19298 15489 19304 15861
rect 19298 15462 19339 15489
rect 19275 15456 19339 15462
rect 54 15454 496 15456
rect 56 15448 494 15454
rect 56 15431 62 15448
rect 488 15431 494 15448
rect 56 15425 494 15431
rect 19306 15454 19339 15456
rect 19306 15448 19744 15454
rect 19306 15431 19312 15448
rect 19738 15431 19744 15448
rect 19306 15425 19744 15431
rect 56 15369 494 15375
rect 56 15352 62 15369
rect 488 15352 494 15369
rect 56 15346 494 15352
rect 461 15344 494 15346
rect 19306 15369 19744 15375
rect 19306 15352 19312 15369
rect 19738 15352 19744 15369
rect 19306 15346 19744 15352
rect 19304 15344 19746 15346
rect 461 15311 500 15344
rect 496 14939 500 15311
rect 461 14906 500 14939
rect 19200 15338 19225 15344
rect 19200 14912 19202 15338
rect 19219 14912 19225 15338
rect 19200 14906 19225 14912
rect 19275 15338 19746 15344
rect 19275 14912 19281 15338
rect 19298 15290 19746 15338
rect 19298 14960 19360 15290
rect 19690 14960 19746 15290
rect 19298 14912 19746 14960
rect 19275 14906 19746 14912
rect 461 14904 494 14906
rect 56 14898 494 14904
rect 56 14881 62 14898
rect 488 14881 494 14898
rect 56 14875 494 14881
rect 19304 14904 19746 14906
rect 19306 14898 19744 14904
rect 19306 14881 19312 14898
rect 19738 14881 19744 14898
rect 19306 14875 19744 14881
rect 56 14819 494 14825
rect 56 14802 62 14819
rect 488 14802 494 14819
rect 56 14796 494 14802
rect 54 14794 496 14796
rect 19306 14819 19744 14825
rect 19306 14802 19312 14819
rect 19738 14802 19744 14819
rect 19306 14796 19744 14802
rect 19306 14794 19339 14796
rect 54 14740 500 14794
rect 54 14410 110 14740
rect 440 14410 500 14740
rect 54 14356 500 14410
rect 19200 14788 19225 14794
rect 19200 14362 19202 14788
rect 19219 14362 19225 14788
rect 19200 14356 19225 14362
rect 19275 14788 19339 14794
rect 19275 14362 19281 14788
rect 19298 14761 19339 14788
rect 19298 14389 19304 14761
rect 19298 14362 19339 14389
rect 19275 14356 19339 14362
rect 54 14354 496 14356
rect 56 14348 494 14354
rect 56 14331 62 14348
rect 488 14331 494 14348
rect 56 14325 494 14331
rect 19306 14354 19339 14356
rect 19306 14348 19744 14354
rect 19306 14331 19312 14348
rect 19738 14331 19744 14348
rect 19306 14325 19744 14331
rect 56 14269 494 14275
rect 56 14252 62 14269
rect 488 14252 494 14269
rect 56 14246 494 14252
rect 461 14244 494 14246
rect 19306 14269 19744 14275
rect 19306 14252 19312 14269
rect 19738 14252 19744 14269
rect 19306 14246 19744 14252
rect 19304 14244 19746 14246
rect 461 14211 500 14244
rect 496 13839 500 14211
rect 461 13806 500 13839
rect 19200 14238 19225 14244
rect 19200 13812 19202 14238
rect 19219 13812 19225 14238
rect 19200 13806 19225 13812
rect 19275 14238 19746 14244
rect 19275 13812 19281 14238
rect 19298 14190 19746 14238
rect 19298 13860 19360 14190
rect 19690 13860 19746 14190
rect 19298 13812 19746 13860
rect 19275 13806 19746 13812
rect 461 13804 494 13806
rect 56 13798 494 13804
rect 56 13781 62 13798
rect 488 13781 494 13798
rect 56 13775 494 13781
rect 19304 13804 19746 13806
rect 19306 13798 19744 13804
rect 19306 13781 19312 13798
rect 19738 13781 19744 13798
rect 19306 13775 19744 13781
rect 56 13719 494 13725
rect 56 13702 62 13719
rect 488 13702 494 13719
rect 56 13696 494 13702
rect 54 13694 496 13696
rect 19306 13719 19744 13725
rect 19306 13702 19312 13719
rect 19738 13702 19744 13719
rect 19306 13696 19744 13702
rect 19306 13694 19339 13696
rect 54 13640 500 13694
rect 54 13310 110 13640
rect 440 13310 500 13640
rect 54 13256 500 13310
rect 19200 13688 19225 13694
rect 19200 13262 19202 13688
rect 19219 13262 19225 13688
rect 19200 13256 19225 13262
rect 19275 13688 19339 13694
rect 19275 13262 19281 13688
rect 19298 13661 19339 13688
rect 19298 13289 19304 13661
rect 19298 13262 19339 13289
rect 19275 13256 19339 13262
rect 54 13254 496 13256
rect 56 13248 494 13254
rect 56 13231 62 13248
rect 488 13231 494 13248
rect 56 13225 494 13231
rect 19306 13254 19339 13256
rect 19306 13248 19744 13254
rect 19306 13231 19312 13248
rect 19738 13231 19744 13248
rect 19306 13225 19744 13231
rect 56 13169 494 13175
rect 56 13152 62 13169
rect 488 13152 494 13169
rect 56 13146 494 13152
rect 461 13144 494 13146
rect 19306 13169 19744 13175
rect 19306 13152 19312 13169
rect 19738 13152 19744 13169
rect 19306 13146 19744 13152
rect 19304 13144 19746 13146
rect 461 13111 500 13144
rect 496 12739 500 13111
rect 461 12706 500 12739
rect 19200 13138 19225 13144
rect 19200 12712 19202 13138
rect 19219 12712 19225 13138
rect 19200 12706 19225 12712
rect 19275 13138 19746 13144
rect 19275 12712 19281 13138
rect 19298 13090 19746 13138
rect 19298 12760 19360 13090
rect 19690 12760 19746 13090
rect 19298 12712 19746 12760
rect 19275 12706 19746 12712
rect 461 12704 494 12706
rect 56 12698 494 12704
rect 56 12681 62 12698
rect 488 12681 494 12698
rect 56 12675 494 12681
rect 19304 12704 19746 12706
rect 19306 12698 19744 12704
rect 19306 12681 19312 12698
rect 19738 12681 19744 12698
rect 19306 12675 19744 12681
rect 56 12619 494 12625
rect 56 12602 62 12619
rect 488 12602 494 12619
rect 56 12596 494 12602
rect 54 12594 496 12596
rect 19306 12619 19744 12625
rect 19306 12602 19312 12619
rect 19738 12602 19744 12619
rect 19306 12596 19744 12602
rect 19306 12594 19339 12596
rect 54 12540 500 12594
rect 54 12210 110 12540
rect 440 12210 500 12540
rect 54 12156 500 12210
rect 19200 12588 19225 12594
rect 19200 12162 19202 12588
rect 19219 12162 19225 12588
rect 19200 12156 19225 12162
rect 19275 12588 19339 12594
rect 19275 12162 19281 12588
rect 19298 12561 19339 12588
rect 19298 12189 19304 12561
rect 19298 12162 19339 12189
rect 19275 12156 19339 12162
rect 54 12154 496 12156
rect 56 12148 494 12154
rect 56 12131 62 12148
rect 488 12131 494 12148
rect 56 12125 494 12131
rect 19306 12154 19339 12156
rect 19306 12148 19744 12154
rect 19306 12131 19312 12148
rect 19738 12131 19744 12148
rect 19306 12125 19744 12131
rect 56 12069 494 12075
rect 56 12052 62 12069
rect 488 12052 494 12069
rect 56 12046 494 12052
rect 461 12044 494 12046
rect 19306 12069 19744 12075
rect 19306 12052 19312 12069
rect 19738 12052 19744 12069
rect 19306 12046 19744 12052
rect 19304 12044 19746 12046
rect 461 12011 500 12044
rect 496 11639 500 12011
rect 461 11606 500 11639
rect 19200 12038 19225 12044
rect 19200 11612 19202 12038
rect 19219 11612 19225 12038
rect 19200 11606 19225 11612
rect 19275 12038 19746 12044
rect 19275 11612 19281 12038
rect 19298 11990 19746 12038
rect 19298 11660 19360 11990
rect 19690 11660 19746 11990
rect 19298 11612 19746 11660
rect 19275 11606 19746 11612
rect 461 11604 494 11606
rect 56 11598 494 11604
rect 56 11581 62 11598
rect 488 11581 494 11598
rect 56 11575 494 11581
rect 19304 11604 19746 11606
rect 19306 11598 19744 11604
rect 19306 11581 19312 11598
rect 19738 11581 19744 11598
rect 19306 11575 19744 11581
rect 56 11519 494 11525
rect 56 11502 62 11519
rect 488 11502 494 11519
rect 56 11496 494 11502
rect 54 11494 496 11496
rect 19306 11519 19744 11525
rect 19306 11502 19312 11519
rect 19738 11502 19744 11519
rect 19306 11496 19744 11502
rect 19306 11494 19339 11496
rect 54 11440 500 11494
rect 54 11110 110 11440
rect 440 11110 500 11440
rect 54 11056 500 11110
rect 19200 11488 19225 11494
rect 19200 11062 19202 11488
rect 19219 11062 19225 11488
rect 19200 11056 19225 11062
rect 19275 11488 19339 11494
rect 19275 11062 19281 11488
rect 19298 11461 19339 11488
rect 19298 11089 19304 11461
rect 19298 11062 19339 11089
rect 19275 11056 19339 11062
rect 54 11054 496 11056
rect 56 11048 494 11054
rect 56 11031 62 11048
rect 488 11031 494 11048
rect 56 11025 494 11031
rect 19306 11054 19339 11056
rect 19306 11048 19744 11054
rect 19306 11031 19312 11048
rect 19738 11031 19744 11048
rect 19306 11025 19744 11031
rect 56 10969 494 10975
rect 56 10952 62 10969
rect 488 10952 494 10969
rect 56 10946 494 10952
rect 461 10944 494 10946
rect 19306 10969 19744 10975
rect 19306 10952 19312 10969
rect 19738 10952 19744 10969
rect 19306 10946 19744 10952
rect 19304 10944 19746 10946
rect 461 10911 500 10944
rect 496 10539 500 10911
rect 461 10506 500 10539
rect 19200 10938 19225 10944
rect 19200 10512 19202 10938
rect 19219 10512 19225 10938
rect 19200 10506 19225 10512
rect 19275 10938 19746 10944
rect 19275 10512 19281 10938
rect 19298 10890 19746 10938
rect 19298 10560 19360 10890
rect 19690 10560 19746 10890
rect 19298 10512 19746 10560
rect 19275 10506 19746 10512
rect 461 10504 494 10506
rect 56 10498 494 10504
rect 56 10481 62 10498
rect 488 10481 494 10498
rect 56 10475 494 10481
rect 19304 10504 19746 10506
rect 19306 10498 19744 10504
rect 19306 10481 19312 10498
rect 19738 10481 19744 10498
rect 19306 10475 19744 10481
rect 56 10419 494 10425
rect 56 10402 62 10419
rect 488 10402 494 10419
rect 56 10396 494 10402
rect 54 10394 496 10396
rect 19306 10419 19744 10425
rect 19306 10402 19312 10419
rect 19738 10402 19744 10419
rect 19306 10396 19744 10402
rect 19306 10394 19339 10396
rect 54 10340 500 10394
rect 54 10010 110 10340
rect 440 10010 500 10340
rect 54 9956 500 10010
rect 19200 10388 19225 10394
rect 19200 9962 19202 10388
rect 19219 9962 19225 10388
rect 19200 9956 19225 9962
rect 19275 10388 19339 10394
rect 19275 9962 19281 10388
rect 19298 10361 19339 10388
rect 19298 9989 19304 10361
rect 19298 9962 19339 9989
rect 19275 9956 19339 9962
rect 54 9954 496 9956
rect 56 9948 494 9954
rect 56 9931 62 9948
rect 488 9931 494 9948
rect 56 9925 494 9931
rect 19306 9954 19339 9956
rect 19306 9948 19744 9954
rect 19306 9931 19312 9948
rect 19738 9931 19744 9948
rect 19306 9925 19744 9931
rect 56 9869 494 9875
rect 56 9852 62 9869
rect 488 9852 494 9869
rect 56 9846 494 9852
rect 461 9844 494 9846
rect 19306 9869 19744 9875
rect 19306 9852 19312 9869
rect 19738 9852 19744 9869
rect 19306 9846 19744 9852
rect 19304 9844 19746 9846
rect 461 9811 500 9844
rect 496 9439 500 9811
rect 461 9406 500 9439
rect 19200 9838 19225 9844
rect 19200 9412 19202 9838
rect 19219 9412 19225 9838
rect 19200 9406 19225 9412
rect 19275 9838 19746 9844
rect 19275 9412 19281 9838
rect 19298 9790 19746 9838
rect 19298 9460 19360 9790
rect 19690 9460 19746 9790
rect 19298 9412 19746 9460
rect 19275 9406 19746 9412
rect 461 9404 494 9406
rect 56 9398 494 9404
rect 56 9381 62 9398
rect 488 9381 494 9398
rect 56 9375 494 9381
rect 19304 9404 19746 9406
rect 19306 9398 19744 9404
rect 19306 9381 19312 9398
rect 19738 9381 19744 9398
rect 19306 9375 19744 9381
rect 56 9319 494 9325
rect 56 9302 62 9319
rect 488 9302 494 9319
rect 56 9296 494 9302
rect 54 9294 496 9296
rect 19306 9319 19744 9325
rect 19306 9302 19312 9319
rect 19738 9302 19744 9319
rect 19306 9296 19744 9302
rect 19306 9294 19339 9296
rect 54 9240 500 9294
rect 54 8910 110 9240
rect 440 8910 500 9240
rect 54 8856 500 8910
rect 19200 9288 19225 9294
rect 19200 8862 19202 9288
rect 19219 8862 19225 9288
rect 19200 8856 19225 8862
rect 19275 9288 19339 9294
rect 19275 8862 19281 9288
rect 19298 9261 19339 9288
rect 19298 8889 19304 9261
rect 19298 8862 19339 8889
rect 19275 8856 19339 8862
rect 54 8854 496 8856
rect 56 8848 494 8854
rect 56 8831 62 8848
rect 488 8831 494 8848
rect 56 8825 494 8831
rect 19306 8854 19339 8856
rect 19306 8848 19744 8854
rect 19306 8831 19312 8848
rect 19738 8831 19744 8848
rect 19306 8825 19744 8831
rect 56 8769 494 8775
rect 56 8752 62 8769
rect 488 8752 494 8769
rect 56 8746 494 8752
rect 461 8744 494 8746
rect 19306 8769 19744 8775
rect 19306 8752 19312 8769
rect 19738 8752 19744 8769
rect 19306 8746 19744 8752
rect 19304 8744 19746 8746
rect 461 8711 500 8744
rect 496 8339 500 8711
rect 461 8306 500 8339
rect 19200 8738 19225 8744
rect 19200 8312 19202 8738
rect 19219 8312 19225 8738
rect 19200 8306 19225 8312
rect 19275 8738 19746 8744
rect 19275 8312 19281 8738
rect 19298 8690 19746 8738
rect 19298 8360 19360 8690
rect 19690 8360 19746 8690
rect 19298 8312 19746 8360
rect 19275 8306 19746 8312
rect 461 8304 494 8306
rect 56 8298 494 8304
rect 56 8281 62 8298
rect 488 8281 494 8298
rect 56 8275 494 8281
rect 19304 8304 19746 8306
rect 19306 8298 19744 8304
rect 19306 8281 19312 8298
rect 19738 8281 19744 8298
rect 19306 8275 19744 8281
rect 56 8219 494 8225
rect 56 8202 62 8219
rect 488 8202 494 8219
rect 56 8196 494 8202
rect 54 8194 496 8196
rect 19306 8219 19744 8225
rect 19306 8202 19312 8219
rect 19738 8202 19744 8219
rect 19306 8196 19744 8202
rect 19306 8194 19339 8196
rect 54 8140 500 8194
rect 54 7810 110 8140
rect 440 7810 500 8140
rect 54 7756 500 7810
rect 19200 8188 19225 8194
rect 19200 7762 19202 8188
rect 19219 7762 19225 8188
rect 19200 7756 19225 7762
rect 19275 8188 19339 8194
rect 19275 7762 19281 8188
rect 19298 8161 19339 8188
rect 19298 7789 19304 8161
rect 19298 7762 19339 7789
rect 19275 7756 19339 7762
rect 54 7754 496 7756
rect 56 7748 494 7754
rect 56 7731 62 7748
rect 488 7731 494 7748
rect 56 7725 494 7731
rect 19306 7754 19339 7756
rect 19306 7748 19744 7754
rect 19306 7731 19312 7748
rect 19738 7731 19744 7748
rect 19306 7725 19744 7731
rect 56 7669 494 7675
rect 56 7652 62 7669
rect 488 7652 494 7669
rect 56 7646 494 7652
rect 461 7644 494 7646
rect 19306 7669 19744 7675
rect 19306 7652 19312 7669
rect 19738 7652 19744 7669
rect 19306 7646 19744 7652
rect 19304 7644 19746 7646
rect 461 7611 500 7644
rect 496 7239 500 7611
rect 461 7206 500 7239
rect 19200 7638 19225 7644
rect 19200 7212 19202 7638
rect 19219 7212 19225 7638
rect 19200 7206 19225 7212
rect 19275 7638 19746 7644
rect 19275 7212 19281 7638
rect 19298 7590 19746 7638
rect 19298 7260 19360 7590
rect 19690 7260 19746 7590
rect 19298 7212 19746 7260
rect 19275 7206 19746 7212
rect 461 7204 494 7206
rect 56 7198 494 7204
rect 56 7181 62 7198
rect 488 7181 494 7198
rect 56 7175 494 7181
rect 19304 7204 19746 7206
rect 19306 7198 19744 7204
rect 19306 7181 19312 7198
rect 19738 7181 19744 7198
rect 19306 7175 19744 7181
rect 56 7119 494 7125
rect 56 7102 62 7119
rect 488 7102 494 7119
rect 56 7096 494 7102
rect 54 7094 496 7096
rect 19306 7119 19744 7125
rect 19306 7102 19312 7119
rect 19738 7102 19744 7119
rect 19306 7096 19744 7102
rect 19306 7094 19339 7096
rect 54 7040 500 7094
rect 54 6710 110 7040
rect 440 6710 500 7040
rect 54 6656 500 6710
rect 19200 7088 19225 7094
rect 19200 6662 19202 7088
rect 19219 6662 19225 7088
rect 19200 6656 19225 6662
rect 19275 7088 19339 7094
rect 19275 6662 19281 7088
rect 19298 7061 19339 7088
rect 19298 6689 19304 7061
rect 19298 6662 19339 6689
rect 19275 6656 19339 6662
rect 54 6654 496 6656
rect 56 6648 494 6654
rect 56 6631 62 6648
rect 488 6631 494 6648
rect 56 6625 494 6631
rect 19306 6654 19339 6656
rect 19306 6648 19744 6654
rect 19306 6631 19312 6648
rect 19738 6631 19744 6648
rect 19306 6625 19744 6631
rect 56 6569 494 6575
rect 56 6552 62 6569
rect 488 6552 494 6569
rect 56 6546 494 6552
rect 461 6544 494 6546
rect 19306 6569 19744 6575
rect 19306 6552 19312 6569
rect 19738 6552 19744 6569
rect 19306 6546 19744 6552
rect 19304 6544 19746 6546
rect 461 6511 500 6544
rect 496 6139 500 6511
rect 461 6106 500 6139
rect 19200 6538 19225 6544
rect 19200 6112 19202 6538
rect 19219 6112 19225 6538
rect 19200 6106 19225 6112
rect 19275 6538 19746 6544
rect 19275 6112 19281 6538
rect 19298 6490 19746 6538
rect 19298 6160 19360 6490
rect 19690 6160 19746 6490
rect 19298 6112 19746 6160
rect 19275 6106 19746 6112
rect 461 6104 494 6106
rect 56 6098 494 6104
rect 56 6081 62 6098
rect 488 6081 494 6098
rect 56 6075 494 6081
rect 19304 6104 19746 6106
rect 19306 6098 19744 6104
rect 19306 6081 19312 6098
rect 19738 6081 19744 6098
rect 19306 6075 19744 6081
rect 56 6019 494 6025
rect 56 6002 62 6019
rect 488 6002 494 6019
rect 56 5996 494 6002
rect 54 5994 496 5996
rect 19306 6019 19744 6025
rect 19306 6002 19312 6019
rect 19738 6002 19744 6019
rect 19306 5996 19744 6002
rect 19306 5994 19339 5996
rect 54 5940 500 5994
rect 54 5610 110 5940
rect 440 5610 500 5940
rect 54 5556 500 5610
rect 19200 5988 19225 5994
rect 19200 5562 19202 5988
rect 19219 5562 19225 5988
rect 19200 5556 19225 5562
rect 19275 5988 19339 5994
rect 19275 5562 19281 5988
rect 19298 5961 19339 5988
rect 19298 5589 19304 5961
rect 19298 5562 19339 5589
rect 19275 5556 19339 5562
rect 54 5554 496 5556
rect 56 5548 494 5554
rect 56 5531 62 5548
rect 488 5531 494 5548
rect 56 5525 494 5531
rect 19306 5554 19339 5556
rect 19306 5548 19744 5554
rect 19306 5531 19312 5548
rect 19738 5531 19744 5548
rect 19306 5525 19744 5531
rect 56 5469 494 5475
rect 56 5452 62 5469
rect 488 5452 494 5469
rect 56 5446 494 5452
rect 461 5444 494 5446
rect 19306 5469 19744 5475
rect 19306 5452 19312 5469
rect 19738 5452 19744 5469
rect 19306 5446 19744 5452
rect 19304 5444 19746 5446
rect 461 5411 500 5444
rect 496 5039 500 5411
rect 461 5006 500 5039
rect 19200 5438 19225 5444
rect 19200 5012 19202 5438
rect 19219 5012 19225 5438
rect 19200 5006 19225 5012
rect 19275 5438 19746 5444
rect 19275 5012 19281 5438
rect 19298 5390 19746 5438
rect 19298 5060 19360 5390
rect 19690 5060 19746 5390
rect 19298 5012 19746 5060
rect 19275 5006 19746 5012
rect 461 5004 494 5006
rect 56 4998 494 5004
rect 56 4981 62 4998
rect 488 4981 494 4998
rect 56 4975 494 4981
rect 19304 5004 19746 5006
rect 19306 4998 19744 5004
rect 19306 4981 19312 4998
rect 19738 4981 19744 4998
rect 19306 4975 19744 4981
rect 56 4919 494 4925
rect 56 4902 62 4919
rect 488 4902 494 4919
rect 56 4896 494 4902
rect 54 4894 496 4896
rect 19306 4919 19744 4925
rect 19306 4902 19312 4919
rect 19738 4902 19744 4919
rect 19306 4896 19744 4902
rect 19306 4894 19339 4896
rect 54 4840 500 4894
rect 54 4510 110 4840
rect 440 4510 500 4840
rect 54 4456 500 4510
rect 19200 4888 19225 4894
rect 19200 4462 19202 4888
rect 19219 4462 19225 4888
rect 19200 4456 19225 4462
rect 19275 4888 19339 4894
rect 19275 4462 19281 4888
rect 19298 4861 19339 4888
rect 19298 4489 19304 4861
rect 19298 4462 19339 4489
rect 19275 4456 19339 4462
rect 54 4454 496 4456
rect 56 4448 494 4454
rect 56 4431 62 4448
rect 488 4431 494 4448
rect 56 4425 494 4431
rect 19306 4454 19339 4456
rect 19306 4448 19744 4454
rect 19306 4431 19312 4448
rect 19738 4431 19744 4448
rect 19306 4425 19744 4431
rect 56 4369 494 4375
rect 56 4352 62 4369
rect 488 4352 494 4369
rect 56 4346 494 4352
rect 461 4344 494 4346
rect 19306 4369 19744 4375
rect 19306 4352 19312 4369
rect 19738 4352 19744 4369
rect 19306 4346 19744 4352
rect 19304 4344 19746 4346
rect 461 4311 500 4344
rect 496 3939 500 4311
rect 461 3906 500 3939
rect 19200 4338 19225 4344
rect 19200 3912 19202 4338
rect 19219 3912 19225 4338
rect 19200 3906 19225 3912
rect 19275 4338 19746 4344
rect 19275 3912 19281 4338
rect 19298 4290 19746 4338
rect 19298 3960 19360 4290
rect 19690 3960 19746 4290
rect 19298 3912 19746 3960
rect 19275 3906 19746 3912
rect 461 3904 494 3906
rect 56 3898 494 3904
rect 56 3881 62 3898
rect 488 3881 494 3898
rect 56 3875 494 3881
rect 19304 3904 19746 3906
rect 19306 3898 19744 3904
rect 19306 3881 19312 3898
rect 19738 3881 19744 3898
rect 19306 3875 19744 3881
rect 56 3819 494 3825
rect 56 3802 62 3819
rect 488 3802 494 3819
rect 56 3796 494 3802
rect 54 3794 496 3796
rect 19306 3819 19744 3825
rect 19306 3802 19312 3819
rect 19738 3802 19744 3819
rect 19306 3796 19744 3802
rect 19306 3794 19339 3796
rect 54 3740 500 3794
rect 54 3410 110 3740
rect 440 3410 500 3740
rect 54 3356 500 3410
rect 19200 3788 19225 3794
rect 19200 3362 19202 3788
rect 19219 3362 19225 3788
rect 19200 3356 19225 3362
rect 19275 3788 19339 3794
rect 19275 3362 19281 3788
rect 19298 3761 19339 3788
rect 19298 3389 19304 3761
rect 19298 3362 19339 3389
rect 19275 3356 19339 3362
rect 54 3354 496 3356
rect 56 3348 494 3354
rect 56 3331 62 3348
rect 488 3331 494 3348
rect 56 3325 494 3331
rect 19306 3354 19339 3356
rect 19306 3348 19744 3354
rect 19306 3331 19312 3348
rect 19738 3331 19744 3348
rect 19306 3325 19744 3331
rect 56 3269 494 3275
rect 56 3252 62 3269
rect 488 3252 494 3269
rect 56 3246 494 3252
rect 461 3244 494 3246
rect 19306 3269 19744 3275
rect 19306 3252 19312 3269
rect 19738 3252 19744 3269
rect 19306 3246 19744 3252
rect 19304 3244 19746 3246
rect 461 3211 500 3244
rect 496 2839 500 3211
rect 461 2806 500 2839
rect 19200 3238 19225 3244
rect 19200 2812 19202 3238
rect 19219 2812 19225 3238
rect 19200 2806 19225 2812
rect 19275 3238 19746 3244
rect 19275 2812 19281 3238
rect 19298 3190 19746 3238
rect 19298 2860 19360 3190
rect 19690 2860 19746 3190
rect 19298 2812 19746 2860
rect 19275 2806 19746 2812
rect 461 2804 494 2806
rect 56 2798 494 2804
rect 56 2781 62 2798
rect 488 2781 494 2798
rect 56 2775 494 2781
rect 19304 2804 19746 2806
rect 19306 2798 19744 2804
rect 19306 2781 19312 2798
rect 19738 2781 19744 2798
rect 19306 2775 19744 2781
rect 56 2719 494 2725
rect 56 2702 62 2719
rect 488 2702 494 2719
rect 56 2696 494 2702
rect 54 2694 496 2696
rect 19306 2719 19744 2725
rect 19306 2702 19312 2719
rect 19738 2702 19744 2719
rect 19306 2696 19744 2702
rect 19306 2694 19339 2696
rect 54 2640 500 2694
rect 54 2310 110 2640
rect 440 2310 500 2640
rect 54 2256 500 2310
rect 19200 2688 19225 2694
rect 19200 2262 19202 2688
rect 19219 2262 19225 2688
rect 19200 2256 19225 2262
rect 19275 2688 19339 2694
rect 19275 2262 19281 2688
rect 19298 2661 19339 2688
rect 19298 2289 19304 2661
rect 19298 2262 19339 2289
rect 19275 2256 19339 2262
rect 54 2254 496 2256
rect 56 2248 494 2254
rect 56 2231 62 2248
rect 488 2231 494 2248
rect 56 2225 494 2231
rect 19306 2254 19339 2256
rect 19306 2248 19744 2254
rect 19306 2231 19312 2248
rect 19738 2231 19744 2248
rect 19306 2225 19744 2231
rect 56 2169 494 2175
rect 56 2152 62 2169
rect 488 2152 494 2169
rect 56 2146 494 2152
rect 461 2144 494 2146
rect 19306 2169 19744 2175
rect 19306 2152 19312 2169
rect 19738 2152 19744 2169
rect 19306 2146 19744 2152
rect 19304 2144 19746 2146
rect 461 2111 500 2144
rect 496 1739 500 2111
rect 461 1706 500 1739
rect 19200 2138 19225 2144
rect 19200 1712 19202 2138
rect 19219 1712 19225 2138
rect 19200 1706 19225 1712
rect 19275 2138 19746 2144
rect 19275 1712 19281 2138
rect 19298 2090 19746 2138
rect 19298 1760 19360 2090
rect 19690 1760 19746 2090
rect 19298 1712 19746 1760
rect 19275 1706 19746 1712
rect 461 1704 494 1706
rect 56 1698 494 1704
rect 56 1681 62 1698
rect 488 1681 494 1698
rect 56 1675 494 1681
rect 19304 1704 19746 1706
rect 19306 1698 19744 1704
rect 19306 1681 19312 1698
rect 19738 1681 19744 1698
rect 19306 1675 19744 1681
rect 56 1619 494 1625
rect 56 1602 62 1619
rect 488 1602 494 1619
rect 56 1596 494 1602
rect 54 1594 496 1596
rect 19306 1619 19744 1625
rect 19306 1602 19312 1619
rect 19738 1602 19744 1619
rect 19306 1596 19744 1602
rect 19306 1594 19339 1596
rect 54 1540 500 1594
rect 54 1210 110 1540
rect 440 1210 500 1540
rect 54 1156 500 1210
rect 19200 1588 19225 1594
rect 19200 1162 19202 1588
rect 19219 1162 19225 1588
rect 19200 1156 19225 1162
rect 19275 1588 19339 1594
rect 19275 1162 19281 1588
rect 19298 1561 19339 1588
rect 19298 1189 19304 1561
rect 19298 1162 19339 1189
rect 19275 1156 19339 1162
rect 54 1154 496 1156
rect 56 1148 494 1154
rect 56 1131 62 1148
rect 488 1131 494 1148
rect 56 1125 494 1131
rect 19306 1154 19339 1156
rect 19306 1148 19744 1154
rect 19306 1131 19312 1148
rect 19738 1131 19744 1148
rect 19306 1125 19744 1131
rect 56 1069 494 1075
rect 56 1052 62 1069
rect 488 1052 494 1069
rect 56 1046 494 1052
rect 461 1044 494 1046
rect 19306 1069 19744 1075
rect 19306 1052 19312 1069
rect 19738 1052 19744 1069
rect 19306 1046 19744 1052
rect 19304 1044 19746 1046
rect 461 1011 500 1044
rect 496 639 500 1011
rect 461 606 500 639
rect 19200 1038 19225 1044
rect 19200 612 19202 1038
rect 19219 612 19225 1038
rect 19200 606 19225 612
rect 19275 1038 19746 1044
rect 19275 612 19281 1038
rect 19298 990 19746 1038
rect 19298 660 19360 990
rect 19690 660 19746 990
rect 19298 612 19746 660
rect 19275 606 19746 612
rect 461 604 494 606
rect 56 598 494 604
rect 56 581 62 598
rect 488 581 494 598
rect 56 575 494 581
rect 19304 604 19746 606
rect 19306 598 19744 604
rect 19306 581 19312 598
rect 19738 581 19744 598
rect 19306 575 19744 581
rect 56 519 494 525
rect 56 502 62 519
rect 488 502 494 519
rect 56 496 494 502
rect 54 494 496 496
rect 606 496 1044 500
rect 606 494 639 496
rect 54 488 525 494
rect 54 440 502 488
rect 54 110 110 440
rect 440 110 502 440
rect 54 62 502 110
rect 519 62 525 488
rect 54 56 525 62
rect 575 488 639 494
rect 575 62 581 488
rect 598 461 639 488
rect 1011 494 1044 496
rect 1156 496 1594 500
rect 1154 494 1596 496
rect 1706 496 2144 500
rect 1706 494 1739 496
rect 1011 488 1075 494
rect 1011 461 1052 488
rect 598 62 604 461
rect 575 56 604 62
rect 1046 62 1052 461
rect 1069 62 1075 488
rect 1046 56 1075 62
rect 1125 488 1625 494
rect 1125 62 1131 488
rect 1148 440 1602 488
rect 1148 110 1210 440
rect 1540 110 1602 440
rect 1148 62 1602 110
rect 1619 62 1625 488
rect 1125 56 1625 62
rect 1675 488 1739 494
rect 1675 62 1681 488
rect 1698 461 1739 488
rect 2111 494 2144 496
rect 2256 496 2694 500
rect 2254 494 2696 496
rect 2806 496 3244 500
rect 2806 494 2839 496
rect 2111 488 2175 494
rect 2111 461 2152 488
rect 1698 62 1704 461
rect 1675 56 1704 62
rect 2146 62 2152 461
rect 2169 62 2175 488
rect 2146 56 2175 62
rect 2225 488 2725 494
rect 2225 62 2231 488
rect 2248 440 2702 488
rect 2248 110 2310 440
rect 2640 110 2702 440
rect 2248 62 2702 110
rect 2719 62 2725 488
rect 2225 56 2725 62
rect 2775 488 2839 494
rect 2775 62 2781 488
rect 2798 461 2839 488
rect 3211 494 3244 496
rect 3356 496 3794 500
rect 3354 494 3796 496
rect 3906 496 4344 500
rect 3906 494 3939 496
rect 3211 488 3275 494
rect 3211 461 3252 488
rect 2798 62 2804 461
rect 2775 56 2804 62
rect 3246 62 3252 461
rect 3269 62 3275 488
rect 3246 56 3275 62
rect 3325 488 3825 494
rect 3325 62 3331 488
rect 3348 440 3802 488
rect 3348 110 3410 440
rect 3740 110 3802 440
rect 3348 62 3802 110
rect 3819 62 3825 488
rect 3325 56 3825 62
rect 3875 488 3939 494
rect 3875 62 3881 488
rect 3898 461 3939 488
rect 4311 494 4344 496
rect 4456 496 4894 500
rect 4454 494 4896 496
rect 5006 496 5444 500
rect 5006 494 5039 496
rect 4311 488 4375 494
rect 4311 461 4352 488
rect 3898 62 3904 461
rect 3875 56 3904 62
rect 4346 62 4352 461
rect 4369 62 4375 488
rect 4346 56 4375 62
rect 4425 488 4925 494
rect 4425 62 4431 488
rect 4448 440 4902 488
rect 4448 110 4510 440
rect 4840 110 4902 440
rect 4448 62 4902 110
rect 4919 62 4925 488
rect 4425 56 4925 62
rect 4975 488 5039 494
rect 4975 62 4981 488
rect 4998 461 5039 488
rect 5411 494 5444 496
rect 5556 496 5994 500
rect 5554 494 5996 496
rect 6106 496 6544 500
rect 6106 494 6139 496
rect 5411 488 5475 494
rect 5411 461 5452 488
rect 4998 62 5004 461
rect 4975 56 5004 62
rect 5446 62 5452 461
rect 5469 62 5475 488
rect 5446 56 5475 62
rect 5525 488 6025 494
rect 5525 62 5531 488
rect 5548 440 6002 488
rect 5548 110 5610 440
rect 5940 110 6002 440
rect 5548 62 6002 110
rect 6019 62 6025 488
rect 5525 56 6025 62
rect 6075 488 6139 494
rect 6075 62 6081 488
rect 6098 461 6139 488
rect 6511 494 6544 496
rect 6656 496 7094 500
rect 6654 494 7096 496
rect 7206 496 7644 500
rect 7206 494 7239 496
rect 6511 488 6575 494
rect 6511 461 6552 488
rect 6098 62 6104 461
rect 6075 56 6104 62
rect 6546 62 6552 461
rect 6569 62 6575 488
rect 6546 56 6575 62
rect 6625 488 7125 494
rect 6625 62 6631 488
rect 6648 440 7102 488
rect 6648 110 6710 440
rect 7040 110 7102 440
rect 6648 62 7102 110
rect 7119 62 7125 488
rect 6625 56 7125 62
rect 7175 488 7239 494
rect 7175 62 7181 488
rect 7198 461 7239 488
rect 7611 494 7644 496
rect 7756 496 8194 500
rect 7754 494 8196 496
rect 8306 496 8744 500
rect 8306 494 8339 496
rect 7611 488 7675 494
rect 7611 461 7652 488
rect 7198 62 7204 461
rect 7175 56 7204 62
rect 7646 62 7652 461
rect 7669 62 7675 488
rect 7646 56 7675 62
rect 7725 488 8225 494
rect 7725 62 7731 488
rect 7748 440 8202 488
rect 7748 110 7810 440
rect 8140 110 8202 440
rect 7748 62 8202 110
rect 8219 62 8225 488
rect 7725 56 8225 62
rect 8275 488 8339 494
rect 8275 62 8281 488
rect 8298 461 8339 488
rect 8711 494 8744 496
rect 8856 496 9294 500
rect 8854 494 9296 496
rect 9406 496 9844 500
rect 9406 494 9439 496
rect 8711 488 8775 494
rect 8711 461 8752 488
rect 8298 62 8304 461
rect 8275 56 8304 62
rect 8746 62 8752 461
rect 8769 62 8775 488
rect 8746 56 8775 62
rect 8825 488 9325 494
rect 8825 62 8831 488
rect 8848 440 9302 488
rect 8848 110 8910 440
rect 9240 110 9302 440
rect 8848 62 9302 110
rect 9319 62 9325 488
rect 8825 56 9325 62
rect 9375 488 9439 494
rect 9375 62 9381 488
rect 9398 461 9439 488
rect 9811 494 9844 496
rect 9956 496 10394 500
rect 9954 494 10396 496
rect 10506 496 10944 500
rect 10506 494 10539 496
rect 9811 488 9875 494
rect 9811 461 9852 488
rect 9398 62 9404 461
rect 9375 56 9404 62
rect 9846 62 9852 461
rect 9869 62 9875 488
rect 9846 56 9875 62
rect 9925 488 10425 494
rect 9925 62 9931 488
rect 9948 440 10402 488
rect 9948 110 10010 440
rect 10340 110 10402 440
rect 9948 62 10402 110
rect 10419 62 10425 488
rect 9925 56 10425 62
rect 10475 488 10539 494
rect 10475 62 10481 488
rect 10498 461 10539 488
rect 10911 494 10944 496
rect 11056 496 11494 500
rect 11054 494 11496 496
rect 11606 496 12044 500
rect 11606 494 11639 496
rect 10911 488 10975 494
rect 10911 461 10952 488
rect 10498 62 10504 461
rect 10475 56 10504 62
rect 10946 62 10952 461
rect 10969 62 10975 488
rect 10946 56 10975 62
rect 11025 488 11525 494
rect 11025 62 11031 488
rect 11048 440 11502 488
rect 11048 110 11110 440
rect 11440 110 11502 440
rect 11048 62 11502 110
rect 11519 62 11525 488
rect 11025 56 11525 62
rect 11575 488 11639 494
rect 11575 62 11581 488
rect 11598 461 11639 488
rect 12011 494 12044 496
rect 12156 496 12594 500
rect 12154 494 12596 496
rect 12706 496 13144 500
rect 12706 494 12739 496
rect 12011 488 12075 494
rect 12011 461 12052 488
rect 11598 62 11604 461
rect 11575 56 11604 62
rect 12046 62 12052 461
rect 12069 62 12075 488
rect 12046 56 12075 62
rect 12125 488 12625 494
rect 12125 62 12131 488
rect 12148 440 12602 488
rect 12148 110 12210 440
rect 12540 110 12602 440
rect 12148 62 12602 110
rect 12619 62 12625 488
rect 12125 56 12625 62
rect 12675 488 12739 494
rect 12675 62 12681 488
rect 12698 461 12739 488
rect 13111 494 13144 496
rect 13256 496 13694 500
rect 13254 494 13696 496
rect 13806 496 14244 500
rect 13806 494 13839 496
rect 13111 488 13175 494
rect 13111 461 13152 488
rect 12698 62 12704 461
rect 12675 56 12704 62
rect 13146 62 13152 461
rect 13169 62 13175 488
rect 13146 56 13175 62
rect 13225 488 13725 494
rect 13225 62 13231 488
rect 13248 440 13702 488
rect 13248 110 13310 440
rect 13640 110 13702 440
rect 13248 62 13702 110
rect 13719 62 13725 488
rect 13225 56 13725 62
rect 13775 488 13839 494
rect 13775 62 13781 488
rect 13798 461 13839 488
rect 14211 494 14244 496
rect 14356 496 14794 500
rect 14354 494 14796 496
rect 14906 496 15344 500
rect 14906 494 14939 496
rect 14211 488 14275 494
rect 14211 461 14252 488
rect 13798 62 13804 461
rect 13775 56 13804 62
rect 14246 62 14252 461
rect 14269 62 14275 488
rect 14246 56 14275 62
rect 14325 488 14825 494
rect 14325 62 14331 488
rect 14348 440 14802 488
rect 14348 110 14410 440
rect 14740 110 14802 440
rect 14348 62 14802 110
rect 14819 62 14825 488
rect 14325 56 14825 62
rect 14875 488 14939 494
rect 14875 62 14881 488
rect 14898 461 14939 488
rect 15311 494 15344 496
rect 15456 496 15894 500
rect 15454 494 15896 496
rect 16006 496 16444 500
rect 16006 494 16039 496
rect 15311 488 15375 494
rect 15311 461 15352 488
rect 14898 62 14904 461
rect 14875 56 14904 62
rect 15346 62 15352 461
rect 15369 62 15375 488
rect 15346 56 15375 62
rect 15425 488 15925 494
rect 15425 62 15431 488
rect 15448 440 15902 488
rect 15448 110 15510 440
rect 15840 110 15902 440
rect 15448 62 15902 110
rect 15919 62 15925 488
rect 15425 56 15925 62
rect 15975 488 16039 494
rect 15975 62 15981 488
rect 15998 461 16039 488
rect 16411 494 16444 496
rect 16556 496 16994 500
rect 16554 494 16996 496
rect 17106 496 17544 500
rect 17106 494 17139 496
rect 16411 488 16475 494
rect 16411 461 16452 488
rect 15998 62 16004 461
rect 15975 56 16004 62
rect 16446 62 16452 461
rect 16469 62 16475 488
rect 16446 56 16475 62
rect 16525 488 17025 494
rect 16525 62 16531 488
rect 16548 440 17002 488
rect 16548 110 16610 440
rect 16940 110 17002 440
rect 16548 62 17002 110
rect 17019 62 17025 488
rect 16525 56 17025 62
rect 17075 488 17139 494
rect 17075 62 17081 488
rect 17098 461 17139 488
rect 17511 494 17544 496
rect 17656 496 18094 500
rect 17654 494 18096 496
rect 18206 496 18644 500
rect 18206 494 18239 496
rect 17511 488 17575 494
rect 17511 461 17552 488
rect 17098 62 17104 461
rect 17075 56 17104 62
rect 17546 62 17552 461
rect 17569 62 17575 488
rect 17546 56 17575 62
rect 17625 488 18125 494
rect 17625 62 17631 488
rect 17648 440 18102 488
rect 17648 110 17710 440
rect 18040 110 18102 440
rect 17648 62 18102 110
rect 18119 62 18125 488
rect 17625 56 18125 62
rect 18175 488 18239 494
rect 18175 62 18181 488
rect 18198 461 18239 488
rect 18611 494 18644 496
rect 18756 496 19194 500
rect 18754 494 19196 496
rect 19306 519 19744 525
rect 19306 502 19312 519
rect 19738 502 19744 519
rect 19306 496 19744 502
rect 19306 494 19339 496
rect 18611 488 18675 494
rect 18611 461 18652 488
rect 18198 62 18204 461
rect 18175 56 18204 62
rect 18646 62 18652 461
rect 18669 62 18675 488
rect 18646 56 18675 62
rect 18725 488 19225 494
rect 18725 62 18731 488
rect 18748 440 19202 488
rect 18748 110 18810 440
rect 19140 110 19202 440
rect 18748 62 19202 110
rect 19219 62 19225 488
rect 18725 56 19225 62
rect 19275 488 19339 494
rect 19275 62 19281 488
rect 19298 461 19339 488
rect 19298 62 19304 461
rect 19275 56 19304 62
rect 54 54 496 56
rect 1154 54 1596 56
rect 2254 54 2696 56
rect 3354 54 3796 56
rect 4454 54 4896 56
rect 5554 54 5996 56
rect 6654 54 7096 56
rect 7754 54 8196 56
rect 8854 54 9296 56
rect 9954 54 10396 56
rect 11054 54 11496 56
rect 12154 54 12596 56
rect 13254 54 13696 56
rect 14354 54 14796 56
rect 15454 54 15896 56
rect 16554 54 16996 56
rect 17654 54 18096 56
rect 18754 54 19196 56
<< mvndiffc >>
rect 502 19312 519 19738
rect 581 19312 598 19738
rect 1052 19312 1069 19738
rect 1131 19312 1148 19738
rect 62 19281 488 19298
rect 612 19281 1038 19298
rect 1602 19312 1619 19738
rect 1681 19312 1698 19738
rect 2152 19312 2169 19738
rect 2231 19312 2248 19738
rect 1162 19281 1588 19298
rect 1712 19281 2138 19298
rect 2702 19312 2719 19738
rect 2781 19312 2798 19738
rect 3252 19312 3269 19738
rect 3331 19312 3348 19738
rect 2262 19281 2688 19298
rect 2812 19281 3238 19298
rect 3802 19312 3819 19738
rect 3881 19312 3898 19738
rect 4352 19312 4369 19738
rect 4431 19312 4448 19738
rect 3362 19281 3788 19298
rect 3912 19281 4338 19298
rect 4902 19312 4919 19738
rect 4981 19312 4998 19738
rect 5452 19312 5469 19738
rect 5531 19312 5548 19738
rect 4462 19281 4888 19298
rect 5012 19281 5438 19298
rect 6002 19312 6019 19738
rect 6081 19312 6098 19738
rect 6552 19312 6569 19738
rect 6631 19312 6648 19738
rect 5562 19281 5988 19298
rect 6112 19281 6538 19298
rect 7102 19312 7119 19738
rect 7181 19312 7198 19738
rect 7652 19312 7669 19738
rect 7731 19312 7748 19738
rect 6662 19281 7088 19298
rect 7212 19281 7638 19298
rect 8202 19312 8219 19738
rect 8281 19312 8298 19738
rect 8752 19312 8769 19738
rect 8831 19312 8848 19738
rect 7762 19281 8188 19298
rect 8312 19281 8738 19298
rect 9302 19312 9319 19738
rect 9381 19312 9398 19738
rect 9852 19312 9869 19738
rect 9931 19312 9948 19738
rect 8862 19281 9288 19298
rect 9412 19281 9838 19298
rect 10402 19312 10419 19738
rect 10481 19312 10498 19738
rect 10952 19312 10969 19738
rect 11031 19312 11048 19738
rect 9962 19281 10388 19298
rect 10512 19281 10938 19298
rect 11502 19312 11519 19738
rect 11581 19312 11598 19738
rect 12052 19312 12069 19738
rect 12131 19312 12148 19738
rect 11062 19281 11488 19298
rect 11612 19281 12038 19298
rect 12602 19312 12619 19738
rect 12681 19312 12698 19738
rect 13152 19312 13169 19738
rect 13231 19312 13248 19738
rect 12162 19281 12588 19298
rect 12712 19281 13138 19298
rect 13702 19312 13719 19738
rect 13781 19312 13798 19738
rect 14252 19312 14269 19738
rect 14331 19312 14348 19738
rect 13262 19281 13688 19298
rect 13812 19281 14238 19298
rect 14802 19312 14819 19738
rect 14881 19312 14898 19738
rect 15352 19312 15369 19738
rect 15431 19312 15448 19738
rect 14362 19281 14788 19298
rect 14912 19281 15338 19298
rect 15902 19312 15919 19738
rect 15981 19312 15998 19738
rect 16452 19312 16469 19738
rect 16531 19312 16548 19738
rect 15462 19281 15888 19298
rect 16012 19281 16438 19298
rect 17002 19312 17019 19738
rect 17081 19312 17098 19738
rect 17552 19312 17569 19738
rect 17631 19312 17648 19738
rect 16562 19281 16988 19298
rect 17112 19281 17538 19298
rect 18102 19312 18119 19738
rect 18181 19312 18198 19738
rect 18652 19312 18669 19738
rect 18731 19312 18748 19738
rect 17662 19281 18088 19298
rect 18212 19281 18638 19298
rect 19202 19312 19219 19738
rect 19281 19312 19298 19738
rect 18762 19281 19188 19298
rect 19312 19281 19738 19298
rect 62 19202 488 19219
rect 612 19202 1038 19219
rect 1162 19202 1588 19219
rect 1712 19202 2138 19219
rect 2262 19202 2688 19219
rect 2812 19202 3238 19219
rect 3362 19202 3788 19219
rect 3912 19202 4338 19219
rect 4462 19202 4888 19219
rect 5012 19202 5438 19219
rect 5562 19202 5988 19219
rect 6112 19202 6538 19219
rect 6662 19202 7088 19219
rect 7212 19202 7638 19219
rect 7762 19202 8188 19219
rect 8312 19202 8738 19219
rect 8862 19202 9288 19219
rect 9412 19202 9838 19219
rect 9962 19202 10388 19219
rect 10512 19202 10938 19219
rect 11062 19202 11488 19219
rect 11612 19202 12038 19219
rect 12162 19202 12588 19219
rect 12712 19202 13138 19219
rect 13262 19202 13688 19219
rect 13812 19202 14238 19219
rect 14362 19202 14788 19219
rect 14912 19202 15338 19219
rect 15462 19202 15888 19219
rect 16012 19202 16438 19219
rect 16562 19202 16988 19219
rect 17112 19202 17538 19219
rect 17662 19202 18088 19219
rect 18212 19202 18638 19219
rect 18762 19202 19188 19219
rect 19312 19202 19738 19219
rect 19202 18762 19219 19188
rect 19281 18762 19298 19188
rect 62 18731 488 18748
rect 19312 18731 19738 18748
rect 62 18652 488 18669
rect 19312 18652 19738 18669
rect 19202 18212 19219 18638
rect 19281 18212 19298 18638
rect 62 18181 488 18198
rect 19312 18181 19738 18198
rect 62 18102 488 18119
rect 19312 18102 19738 18119
rect 19202 17662 19219 18088
rect 19281 17662 19298 18088
rect 62 17631 488 17648
rect 19312 17631 19738 17648
rect 62 17552 488 17569
rect 19312 17552 19738 17569
rect 19202 17112 19219 17538
rect 19281 17112 19298 17538
rect 62 17081 488 17098
rect 19312 17081 19738 17098
rect 62 17002 488 17019
rect 19312 17002 19738 17019
rect 19202 16562 19219 16988
rect 19281 16562 19298 16988
rect 62 16531 488 16548
rect 19312 16531 19738 16548
rect 62 16452 488 16469
rect 19312 16452 19738 16469
rect 19202 16012 19219 16438
rect 19281 16012 19298 16438
rect 62 15981 488 15998
rect 19312 15981 19738 15998
rect 62 15902 488 15919
rect 19312 15902 19738 15919
rect 19202 15462 19219 15888
rect 19281 15462 19298 15888
rect 62 15431 488 15448
rect 19312 15431 19738 15448
rect 62 15352 488 15369
rect 19312 15352 19738 15369
rect 19202 14912 19219 15338
rect 19281 14912 19298 15338
rect 62 14881 488 14898
rect 19312 14881 19738 14898
rect 62 14802 488 14819
rect 19312 14802 19738 14819
rect 19202 14362 19219 14788
rect 19281 14362 19298 14788
rect 62 14331 488 14348
rect 19312 14331 19738 14348
rect 62 14252 488 14269
rect 19312 14252 19738 14269
rect 19202 13812 19219 14238
rect 19281 13812 19298 14238
rect 62 13781 488 13798
rect 19312 13781 19738 13798
rect 62 13702 488 13719
rect 19312 13702 19738 13719
rect 19202 13262 19219 13688
rect 19281 13262 19298 13688
rect 62 13231 488 13248
rect 19312 13231 19738 13248
rect 62 13152 488 13169
rect 19312 13152 19738 13169
rect 19202 12712 19219 13138
rect 19281 12712 19298 13138
rect 62 12681 488 12698
rect 19312 12681 19738 12698
rect 62 12602 488 12619
rect 19312 12602 19738 12619
rect 19202 12162 19219 12588
rect 19281 12162 19298 12588
rect 62 12131 488 12148
rect 19312 12131 19738 12148
rect 62 12052 488 12069
rect 19312 12052 19738 12069
rect 19202 11612 19219 12038
rect 19281 11612 19298 12038
rect 62 11581 488 11598
rect 19312 11581 19738 11598
rect 62 11502 488 11519
rect 19312 11502 19738 11519
rect 19202 11062 19219 11488
rect 19281 11062 19298 11488
rect 62 11031 488 11048
rect 19312 11031 19738 11048
rect 62 10952 488 10969
rect 19312 10952 19738 10969
rect 19202 10512 19219 10938
rect 19281 10512 19298 10938
rect 62 10481 488 10498
rect 19312 10481 19738 10498
rect 62 10402 488 10419
rect 19312 10402 19738 10419
rect 19202 9962 19219 10388
rect 19281 9962 19298 10388
rect 62 9931 488 9948
rect 19312 9931 19738 9948
rect 62 9852 488 9869
rect 19312 9852 19738 9869
rect 19202 9412 19219 9838
rect 19281 9412 19298 9838
rect 62 9381 488 9398
rect 19312 9381 19738 9398
rect 62 9302 488 9319
rect 19312 9302 19738 9319
rect 19202 8862 19219 9288
rect 19281 8862 19298 9288
rect 62 8831 488 8848
rect 19312 8831 19738 8848
rect 62 8752 488 8769
rect 19312 8752 19738 8769
rect 19202 8312 19219 8738
rect 19281 8312 19298 8738
rect 62 8281 488 8298
rect 19312 8281 19738 8298
rect 62 8202 488 8219
rect 19312 8202 19738 8219
rect 19202 7762 19219 8188
rect 19281 7762 19298 8188
rect 62 7731 488 7748
rect 19312 7731 19738 7748
rect 62 7652 488 7669
rect 19312 7652 19738 7669
rect 19202 7212 19219 7638
rect 19281 7212 19298 7638
rect 62 7181 488 7198
rect 19312 7181 19738 7198
rect 62 7102 488 7119
rect 19312 7102 19738 7119
rect 19202 6662 19219 7088
rect 19281 6662 19298 7088
rect 62 6631 488 6648
rect 19312 6631 19738 6648
rect 62 6552 488 6569
rect 19312 6552 19738 6569
rect 19202 6112 19219 6538
rect 19281 6112 19298 6538
rect 62 6081 488 6098
rect 19312 6081 19738 6098
rect 62 6002 488 6019
rect 19312 6002 19738 6019
rect 19202 5562 19219 5988
rect 19281 5562 19298 5988
rect 62 5531 488 5548
rect 19312 5531 19738 5548
rect 62 5452 488 5469
rect 19312 5452 19738 5469
rect 19202 5012 19219 5438
rect 19281 5012 19298 5438
rect 62 4981 488 4998
rect 19312 4981 19738 4998
rect 62 4902 488 4919
rect 19312 4902 19738 4919
rect 19202 4462 19219 4888
rect 19281 4462 19298 4888
rect 62 4431 488 4448
rect 19312 4431 19738 4448
rect 62 4352 488 4369
rect 19312 4352 19738 4369
rect 19202 3912 19219 4338
rect 19281 3912 19298 4338
rect 62 3881 488 3898
rect 19312 3881 19738 3898
rect 62 3802 488 3819
rect 19312 3802 19738 3819
rect 19202 3362 19219 3788
rect 19281 3362 19298 3788
rect 62 3331 488 3348
rect 19312 3331 19738 3348
rect 62 3252 488 3269
rect 19312 3252 19738 3269
rect 19202 2812 19219 3238
rect 19281 2812 19298 3238
rect 62 2781 488 2798
rect 19312 2781 19738 2798
rect 62 2702 488 2719
rect 19312 2702 19738 2719
rect 19202 2262 19219 2688
rect 19281 2262 19298 2688
rect 62 2231 488 2248
rect 19312 2231 19738 2248
rect 62 2152 488 2169
rect 19312 2152 19738 2169
rect 19202 1712 19219 2138
rect 19281 1712 19298 2138
rect 62 1681 488 1698
rect 19312 1681 19738 1698
rect 62 1602 488 1619
rect 19312 1602 19738 1619
rect 19202 1162 19219 1588
rect 19281 1162 19298 1588
rect 62 1131 488 1148
rect 19312 1131 19738 1148
rect 62 1052 488 1069
rect 19312 1052 19738 1069
rect 19202 612 19219 1038
rect 19281 612 19298 1038
rect 62 581 488 598
rect 19312 581 19738 598
rect 62 502 488 519
rect 502 62 519 488
rect 581 62 598 488
rect 1052 62 1069 488
rect 1131 62 1148 488
rect 1602 62 1619 488
rect 1681 62 1698 488
rect 2152 62 2169 488
rect 2231 62 2248 488
rect 2702 62 2719 488
rect 2781 62 2798 488
rect 3252 62 3269 488
rect 3331 62 3348 488
rect 3802 62 3819 488
rect 3881 62 3898 488
rect 4352 62 4369 488
rect 4431 62 4448 488
rect 4902 62 4919 488
rect 4981 62 4998 488
rect 5452 62 5469 488
rect 5531 62 5548 488
rect 6002 62 6019 488
rect 6081 62 6098 488
rect 6552 62 6569 488
rect 6631 62 6648 488
rect 7102 62 7119 488
rect 7181 62 7198 488
rect 7652 62 7669 488
rect 7731 62 7748 488
rect 8202 62 8219 488
rect 8281 62 8298 488
rect 8752 62 8769 488
rect 8831 62 8848 488
rect 9302 62 9319 488
rect 9381 62 9398 488
rect 9852 62 9869 488
rect 9931 62 9948 488
rect 10402 62 10419 488
rect 10481 62 10498 488
rect 10952 62 10969 488
rect 11031 62 11048 488
rect 11502 62 11519 488
rect 11581 62 11598 488
rect 12052 62 12069 488
rect 12131 62 12148 488
rect 12602 62 12619 488
rect 12681 62 12698 488
rect 13152 62 13169 488
rect 13231 62 13248 488
rect 13702 62 13719 488
rect 13781 62 13798 488
rect 14252 62 14269 488
rect 14331 62 14348 488
rect 14802 62 14819 488
rect 14881 62 14898 488
rect 15352 62 15369 488
rect 15431 62 15448 488
rect 15902 62 15919 488
rect 15981 62 15998 488
rect 16452 62 16469 488
rect 16531 62 16548 488
rect 17002 62 17019 488
rect 17081 62 17098 488
rect 17552 62 17569 488
rect 17631 62 17648 488
rect 18102 62 18119 488
rect 18181 62 18198 488
rect 19312 502 19738 519
rect 18652 62 18669 488
rect 18731 62 18748 488
rect 19202 62 19219 488
rect 19281 62 19298 488
<< mvpsubdiff >>
rect -500 20288 20300 20300
rect -500 -488 -488 20288
rect -212 20000 20012 20012
rect -212 -200 -200 20000
rect 660 19678 990 19690
rect 660 19372 672 19678
rect 978 19372 990 19678
rect 660 19360 990 19372
rect 1760 19678 2090 19690
rect 1760 19372 1772 19678
rect 2078 19372 2090 19678
rect 1760 19360 2090 19372
rect 2860 19678 3190 19690
rect 2860 19372 2872 19678
rect 3178 19372 3190 19678
rect 2860 19360 3190 19372
rect 3960 19678 4290 19690
rect 3960 19372 3972 19678
rect 4278 19372 4290 19678
rect 3960 19360 4290 19372
rect 5060 19678 5390 19690
rect 5060 19372 5072 19678
rect 5378 19372 5390 19678
rect 5060 19360 5390 19372
rect 6160 19678 6490 19690
rect 6160 19372 6172 19678
rect 6478 19372 6490 19678
rect 6160 19360 6490 19372
rect 7260 19678 7590 19690
rect 7260 19372 7272 19678
rect 7578 19372 7590 19678
rect 7260 19360 7590 19372
rect 8360 19678 8690 19690
rect 8360 19372 8372 19678
rect 8678 19372 8690 19678
rect 8360 19360 8690 19372
rect 9460 19678 9790 19690
rect 9460 19372 9472 19678
rect 9778 19372 9790 19678
rect 9460 19360 9790 19372
rect 10560 19678 10890 19690
rect 10560 19372 10572 19678
rect 10878 19372 10890 19678
rect 10560 19360 10890 19372
rect 11660 19678 11990 19690
rect 11660 19372 11672 19678
rect 11978 19372 11990 19678
rect 11660 19360 11990 19372
rect 12760 19678 13090 19690
rect 12760 19372 12772 19678
rect 13078 19372 13090 19678
rect 12760 19360 13090 19372
rect 13860 19678 14190 19690
rect 13860 19372 13872 19678
rect 14178 19372 14190 19678
rect 13860 19360 14190 19372
rect 14960 19678 15290 19690
rect 14960 19372 14972 19678
rect 15278 19372 15290 19678
rect 14960 19360 15290 19372
rect 16060 19678 16390 19690
rect 16060 19372 16072 19678
rect 16378 19372 16390 19678
rect 16060 19360 16390 19372
rect 17160 19678 17490 19690
rect 17160 19372 17172 19678
rect 17478 19372 17490 19678
rect 17160 19360 17490 19372
rect 18260 19678 18590 19690
rect 18260 19372 18272 19678
rect 18578 19372 18590 19678
rect 18260 19360 18590 19372
rect 19360 19678 19690 19690
rect 19360 19372 19372 19678
rect 19678 19372 19690 19678
rect 19360 19360 19690 19372
rect 110 19128 440 19140
rect 110 18822 122 19128
rect 428 18822 440 19128
rect 110 18810 440 18822
rect 19360 18578 19690 18590
rect 19360 18272 19372 18578
rect 19678 18272 19690 18578
rect 19360 18260 19690 18272
rect 110 18028 440 18040
rect 110 17722 122 18028
rect 428 17722 440 18028
rect 110 17710 440 17722
rect 19360 17478 19690 17490
rect 19360 17172 19372 17478
rect 19678 17172 19690 17478
rect 19360 17160 19690 17172
rect 110 16928 440 16940
rect 110 16622 122 16928
rect 428 16622 440 16928
rect 110 16610 440 16622
rect 19360 16378 19690 16390
rect 19360 16072 19372 16378
rect 19678 16072 19690 16378
rect 19360 16060 19690 16072
rect 110 15828 440 15840
rect 110 15522 122 15828
rect 428 15522 440 15828
rect 110 15510 440 15522
rect 19360 15278 19690 15290
rect 19360 14972 19372 15278
rect 19678 14972 19690 15278
rect 19360 14960 19690 14972
rect 110 14728 440 14740
rect 110 14422 122 14728
rect 428 14422 440 14728
rect 110 14410 440 14422
rect 19360 14178 19690 14190
rect 19360 13872 19372 14178
rect 19678 13872 19690 14178
rect 19360 13860 19690 13872
rect 110 13628 440 13640
rect 110 13322 122 13628
rect 428 13322 440 13628
rect 110 13310 440 13322
rect 19360 13078 19690 13090
rect 19360 12772 19372 13078
rect 19678 12772 19690 13078
rect 19360 12760 19690 12772
rect 110 12528 440 12540
rect 110 12222 122 12528
rect 428 12222 440 12528
rect 110 12210 440 12222
rect 19360 11978 19690 11990
rect 19360 11672 19372 11978
rect 19678 11672 19690 11978
rect 19360 11660 19690 11672
rect 110 11428 440 11440
rect 110 11122 122 11428
rect 428 11122 440 11428
rect 110 11110 440 11122
rect 19360 10878 19690 10890
rect 19360 10572 19372 10878
rect 19678 10572 19690 10878
rect 19360 10560 19690 10572
rect 110 10328 440 10340
rect 110 10022 122 10328
rect 428 10022 440 10328
rect 110 10010 440 10022
rect 19360 9778 19690 9790
rect 19360 9472 19372 9778
rect 19678 9472 19690 9778
rect 19360 9460 19690 9472
rect 110 9228 440 9240
rect 110 8922 122 9228
rect 428 8922 440 9228
rect 110 8910 440 8922
rect 19360 8678 19690 8690
rect 19360 8372 19372 8678
rect 19678 8372 19690 8678
rect 19360 8360 19690 8372
rect 110 8128 440 8140
rect 110 7822 122 8128
rect 428 7822 440 8128
rect 110 7810 440 7822
rect 19360 7578 19690 7590
rect 19360 7272 19372 7578
rect 19678 7272 19690 7578
rect 19360 7260 19690 7272
rect 110 7028 440 7040
rect 110 6722 122 7028
rect 428 6722 440 7028
rect 110 6710 440 6722
rect 19360 6478 19690 6490
rect 19360 6172 19372 6478
rect 19678 6172 19690 6478
rect 19360 6160 19690 6172
rect 110 5928 440 5940
rect 110 5622 122 5928
rect 428 5622 440 5928
rect 110 5610 440 5622
rect 19360 5378 19690 5390
rect 19360 5072 19372 5378
rect 19678 5072 19690 5378
rect 19360 5060 19690 5072
rect 110 4828 440 4840
rect 110 4522 122 4828
rect 428 4522 440 4828
rect 110 4510 440 4522
rect 19360 4278 19690 4290
rect 19360 3972 19372 4278
rect 19678 3972 19690 4278
rect 19360 3960 19690 3972
rect 110 3728 440 3740
rect 110 3422 122 3728
rect 428 3422 440 3728
rect 110 3410 440 3422
rect 19360 3178 19690 3190
rect 19360 2872 19372 3178
rect 19678 2872 19690 3178
rect 19360 2860 19690 2872
rect 110 2628 440 2640
rect 110 2322 122 2628
rect 428 2322 440 2628
rect 110 2310 440 2322
rect 19360 2078 19690 2090
rect 19360 1772 19372 2078
rect 19678 1772 19690 2078
rect 19360 1760 19690 1772
rect 110 1528 440 1540
rect 110 1222 122 1528
rect 428 1222 440 1528
rect 110 1210 440 1222
rect 19360 978 19690 990
rect 19360 672 19372 978
rect 19678 672 19690 978
rect 19360 660 19690 672
rect 110 428 440 440
rect 110 122 122 428
rect 428 122 440 428
rect 110 110 440 122
rect 1210 428 1540 440
rect 1210 122 1222 428
rect 1528 122 1540 428
rect 1210 110 1540 122
rect 2310 428 2640 440
rect 2310 122 2322 428
rect 2628 122 2640 428
rect 2310 110 2640 122
rect 3410 428 3740 440
rect 3410 122 3422 428
rect 3728 122 3740 428
rect 3410 110 3740 122
rect 4510 428 4840 440
rect 4510 122 4522 428
rect 4828 122 4840 428
rect 4510 110 4840 122
rect 5610 428 5940 440
rect 5610 122 5622 428
rect 5928 122 5940 428
rect 5610 110 5940 122
rect 6710 428 7040 440
rect 6710 122 6722 428
rect 7028 122 7040 428
rect 6710 110 7040 122
rect 7810 428 8140 440
rect 7810 122 7822 428
rect 8128 122 8140 428
rect 7810 110 8140 122
rect 8910 428 9240 440
rect 8910 122 8922 428
rect 9228 122 9240 428
rect 8910 110 9240 122
rect 10010 428 10340 440
rect 10010 122 10022 428
rect 10328 122 10340 428
rect 10010 110 10340 122
rect 11110 428 11440 440
rect 11110 122 11122 428
rect 11428 122 11440 428
rect 11110 110 11440 122
rect 12210 428 12540 440
rect 12210 122 12222 428
rect 12528 122 12540 428
rect 12210 110 12540 122
rect 13310 428 13640 440
rect 13310 122 13322 428
rect 13628 122 13640 428
rect 13310 110 13640 122
rect 14410 428 14740 440
rect 14410 122 14422 428
rect 14728 122 14740 428
rect 14410 110 14740 122
rect 15510 428 15840 440
rect 15510 122 15522 428
rect 15828 122 15840 428
rect 15510 110 15840 122
rect 16610 428 16940 440
rect 16610 122 16622 428
rect 16928 122 16940 428
rect 16610 110 16940 122
rect 17710 428 18040 440
rect 17710 122 17722 428
rect 18028 122 18040 428
rect 17710 110 18040 122
rect 18810 428 19140 440
rect 18810 122 18822 428
rect 19128 122 19140 428
rect 18810 110 19140 122
rect 20000 -200 20012 20000
rect -212 -212 20012 -200
rect 20288 -488 20300 20288
rect -500 -500 20300 -488
<< mvnsubdiff >>
rect -5000 24788 24800 24800
rect -5000 -4988 -4988 24788
rect -1012 20800 20812 20812
rect -1012 -1000 -1000 20800
rect 20800 -1000 20812 20800
rect -1012 -1012 20812 -1000
rect 24788 -4988 24800 24788
rect -5000 -5000 24800 -4988
<< mvpsubdiffcont >>
rect -488 20012 20288 20288
rect -488 -212 -212 20012
rect 672 19372 978 19678
rect 1772 19372 2078 19678
rect 2872 19372 3178 19678
rect 3972 19372 4278 19678
rect 5072 19372 5378 19678
rect 6172 19372 6478 19678
rect 7272 19372 7578 19678
rect 8372 19372 8678 19678
rect 9472 19372 9778 19678
rect 10572 19372 10878 19678
rect 11672 19372 11978 19678
rect 12772 19372 13078 19678
rect 13872 19372 14178 19678
rect 14972 19372 15278 19678
rect 16072 19372 16378 19678
rect 17172 19372 17478 19678
rect 18272 19372 18578 19678
rect 19372 19372 19678 19678
rect 122 18822 428 19128
rect 19372 18272 19678 18578
rect 122 17722 428 18028
rect 19372 17172 19678 17478
rect 122 16622 428 16928
rect 19372 16072 19678 16378
rect 122 15522 428 15828
rect 19372 14972 19678 15278
rect 122 14422 428 14728
rect 19372 13872 19678 14178
rect 122 13322 428 13628
rect 19372 12772 19678 13078
rect 122 12222 428 12528
rect 19372 11672 19678 11978
rect 122 11122 428 11428
rect 19372 10572 19678 10878
rect 122 10022 428 10328
rect 19372 9472 19678 9778
rect 122 8922 428 9228
rect 19372 8372 19678 8678
rect 122 7822 428 8128
rect 19372 7272 19678 7578
rect 122 6722 428 7028
rect 19372 6172 19678 6478
rect 122 5622 428 5928
rect 19372 5072 19678 5378
rect 122 4522 428 4828
rect 19372 3972 19678 4278
rect 122 3422 428 3728
rect 19372 2872 19678 3178
rect 122 2322 428 2628
rect 19372 1772 19678 2078
rect 122 1222 428 1528
rect 19372 672 19678 978
rect 122 122 428 428
rect 1222 122 1528 428
rect 2322 122 2628 428
rect 3422 122 3728 428
rect 4522 122 4828 428
rect 5622 122 5928 428
rect 6722 122 7028 428
rect 7822 122 8128 428
rect 8922 122 9228 428
rect 10022 122 10328 428
rect 11122 122 11428 428
rect 12222 122 12528 428
rect 13322 122 13628 428
rect 14422 122 14728 428
rect 15522 122 15828 428
rect 16622 122 16928 428
rect 17722 122 18028 428
rect 18822 122 19128 428
rect 20012 -212 20288 20012
rect -488 -488 20288 -212
<< mvnsubdiffcont >>
rect -4988 20812 24788 24788
rect -4988 -1012 -1012 20812
rect 20812 -1012 24788 20812
rect -4988 -4988 24788 -1012
<< poly >>
rect -25 19817 19825 19825
rect -25 19783 -17 19817
rect 17 19783 533 19817
rect 567 19783 1083 19817
rect 1117 19783 1633 19817
rect 1667 19783 2183 19817
rect 2217 19783 2733 19817
rect 2767 19783 3283 19817
rect 3317 19783 3833 19817
rect 3867 19783 4383 19817
rect 4417 19783 4933 19817
rect 4967 19783 5483 19817
rect 5517 19783 6033 19817
rect 6067 19783 6583 19817
rect 6617 19783 7133 19817
rect 7167 19783 7683 19817
rect 7717 19783 8233 19817
rect 8267 19783 8783 19817
rect 8817 19783 9333 19817
rect 9367 19783 9883 19817
rect 9917 19783 10433 19817
rect 10467 19783 10983 19817
rect 11017 19783 11533 19817
rect 11567 19783 12083 19817
rect 12117 19783 12633 19817
rect 12667 19783 13183 19817
rect 13217 19783 13733 19817
rect 13767 19783 14283 19817
rect 14317 19783 14833 19817
rect 14867 19783 15383 19817
rect 15417 19783 15933 19817
rect 15967 19783 16483 19817
rect 16517 19783 17033 19817
rect 17067 19783 17583 19817
rect 17617 19783 18133 19817
rect 18167 19783 18683 19817
rect 18717 19783 19233 19817
rect 19267 19783 19783 19817
rect 19817 19783 19825 19817
rect -25 19775 19825 19783
rect -25 19275 25 19775
rect 525 19744 575 19775
rect 1075 19744 1125 19775
rect 1625 19744 1675 19775
rect 2175 19744 2225 19775
rect 2725 19744 2775 19775
rect 3275 19744 3325 19775
rect 3825 19744 3875 19775
rect 4375 19744 4425 19775
rect 4925 19744 4975 19775
rect 5475 19744 5525 19775
rect 6025 19744 6075 19775
rect 6575 19744 6625 19775
rect 7125 19744 7175 19775
rect 7675 19744 7725 19775
rect 8225 19744 8275 19775
rect 8775 19744 8825 19775
rect 9325 19744 9375 19775
rect 9875 19744 9925 19775
rect 10425 19744 10475 19775
rect 10975 19744 11025 19775
rect 11525 19744 11575 19775
rect 12075 19744 12125 19775
rect 12625 19744 12675 19775
rect 13175 19744 13225 19775
rect 13725 19744 13775 19775
rect 14275 19744 14325 19775
rect 14825 19744 14875 19775
rect 15375 19744 15425 19775
rect 15925 19744 15975 19775
rect 16475 19744 16525 19775
rect 17025 19744 17075 19775
rect 17575 19744 17625 19775
rect 18125 19744 18175 19775
rect 18675 19744 18725 19775
rect 19225 19744 19275 19775
rect 525 19275 575 19306
rect 1075 19275 1125 19306
rect 1625 19275 1675 19306
rect 2175 19275 2225 19306
rect 2725 19275 2775 19306
rect 3275 19275 3325 19306
rect 3825 19275 3875 19306
rect 4375 19275 4425 19306
rect 4925 19275 4975 19306
rect 5475 19275 5525 19306
rect 6025 19275 6075 19306
rect 6575 19275 6625 19306
rect 7125 19275 7175 19306
rect 7675 19275 7725 19306
rect 8225 19275 8275 19306
rect 8775 19275 8825 19306
rect 9325 19275 9375 19306
rect 9875 19275 9925 19306
rect 10425 19275 10475 19306
rect 10975 19275 11025 19306
rect 11525 19275 11575 19306
rect 12075 19275 12125 19306
rect 12625 19275 12675 19306
rect 13175 19275 13225 19306
rect 13725 19275 13775 19306
rect 14275 19275 14325 19306
rect 14825 19275 14875 19306
rect 15375 19275 15425 19306
rect 15925 19275 15975 19306
rect 16475 19275 16525 19306
rect 17025 19275 17075 19306
rect 17575 19275 17625 19306
rect 18125 19275 18175 19306
rect 18675 19275 18725 19306
rect 19225 19275 19275 19306
rect 19775 19275 19825 19775
rect -25 19267 56 19275
rect -25 19233 -17 19267
rect 17 19233 56 19267
rect -25 19225 56 19233
rect 494 19267 606 19275
rect 494 19233 533 19267
rect 567 19233 606 19267
rect 494 19225 606 19233
rect 1044 19267 1156 19275
rect 1044 19233 1083 19267
rect 1117 19233 1156 19267
rect 1044 19225 1156 19233
rect 1594 19267 1706 19275
rect 1594 19233 1633 19267
rect 1667 19233 1706 19267
rect 1594 19225 1706 19233
rect 2144 19267 2256 19275
rect 2144 19233 2183 19267
rect 2217 19233 2256 19267
rect 2144 19225 2256 19233
rect 2694 19267 2806 19275
rect 2694 19233 2733 19267
rect 2767 19233 2806 19267
rect 2694 19225 2806 19233
rect 3244 19267 3356 19275
rect 3244 19233 3283 19267
rect 3317 19233 3356 19267
rect 3244 19225 3356 19233
rect 3794 19267 3906 19275
rect 3794 19233 3833 19267
rect 3867 19233 3906 19267
rect 3794 19225 3906 19233
rect 4344 19267 4456 19275
rect 4344 19233 4383 19267
rect 4417 19233 4456 19267
rect 4344 19225 4456 19233
rect 4894 19267 5006 19275
rect 4894 19233 4933 19267
rect 4967 19233 5006 19267
rect 4894 19225 5006 19233
rect 5444 19267 5556 19275
rect 5444 19233 5483 19267
rect 5517 19233 5556 19267
rect 5444 19225 5556 19233
rect 5994 19267 6106 19275
rect 5994 19233 6033 19267
rect 6067 19233 6106 19267
rect 5994 19225 6106 19233
rect 6544 19267 6656 19275
rect 6544 19233 6583 19267
rect 6617 19233 6656 19267
rect 6544 19225 6656 19233
rect 7094 19267 7206 19275
rect 7094 19233 7133 19267
rect 7167 19233 7206 19267
rect 7094 19225 7206 19233
rect 7644 19267 7756 19275
rect 7644 19233 7683 19267
rect 7717 19233 7756 19267
rect 7644 19225 7756 19233
rect 8194 19267 8306 19275
rect 8194 19233 8233 19267
rect 8267 19233 8306 19267
rect 8194 19225 8306 19233
rect 8744 19267 8856 19275
rect 8744 19233 8783 19267
rect 8817 19233 8856 19267
rect 8744 19225 8856 19233
rect 9294 19267 9406 19275
rect 9294 19233 9333 19267
rect 9367 19233 9406 19267
rect 9294 19225 9406 19233
rect 9844 19267 9956 19275
rect 9844 19233 9883 19267
rect 9917 19233 9956 19267
rect 9844 19225 9956 19233
rect 10394 19267 10506 19275
rect 10394 19233 10433 19267
rect 10467 19233 10506 19267
rect 10394 19225 10506 19233
rect 10944 19267 11056 19275
rect 10944 19233 10983 19267
rect 11017 19233 11056 19267
rect 10944 19225 11056 19233
rect 11494 19267 11606 19275
rect 11494 19233 11533 19267
rect 11567 19233 11606 19267
rect 11494 19225 11606 19233
rect 12044 19267 12156 19275
rect 12044 19233 12083 19267
rect 12117 19233 12156 19267
rect 12044 19225 12156 19233
rect 12594 19267 12706 19275
rect 12594 19233 12633 19267
rect 12667 19233 12706 19267
rect 12594 19225 12706 19233
rect 13144 19267 13256 19275
rect 13144 19233 13183 19267
rect 13217 19233 13256 19267
rect 13144 19225 13256 19233
rect 13694 19267 13806 19275
rect 13694 19233 13733 19267
rect 13767 19233 13806 19267
rect 13694 19225 13806 19233
rect 14244 19267 14356 19275
rect 14244 19233 14283 19267
rect 14317 19233 14356 19267
rect 14244 19225 14356 19233
rect 14794 19267 14906 19275
rect 14794 19233 14833 19267
rect 14867 19233 14906 19267
rect 14794 19225 14906 19233
rect 15344 19267 15456 19275
rect 15344 19233 15383 19267
rect 15417 19233 15456 19267
rect 15344 19225 15456 19233
rect 15894 19267 16006 19275
rect 15894 19233 15933 19267
rect 15967 19233 16006 19267
rect 15894 19225 16006 19233
rect 16444 19267 16556 19275
rect 16444 19233 16483 19267
rect 16517 19233 16556 19267
rect 16444 19225 16556 19233
rect 16994 19267 17106 19275
rect 16994 19233 17033 19267
rect 17067 19233 17106 19267
rect 16994 19225 17106 19233
rect 17544 19267 17656 19275
rect 17544 19233 17583 19267
rect 17617 19233 17656 19267
rect 17544 19225 17656 19233
rect 18094 19267 18206 19275
rect 18094 19233 18133 19267
rect 18167 19233 18206 19267
rect 18094 19225 18206 19233
rect 18644 19267 18756 19275
rect 18644 19233 18683 19267
rect 18717 19233 18756 19267
rect 18644 19225 18756 19233
rect 19194 19267 19306 19275
rect 19194 19233 19233 19267
rect 19267 19233 19306 19267
rect 19194 19225 19306 19233
rect 19744 19267 19825 19275
rect 19744 19233 19783 19267
rect 19817 19233 19825 19267
rect 19744 19225 19825 19233
rect -25 18725 25 19225
rect 525 19200 575 19225
rect 1075 19200 1125 19225
rect 1625 19200 1675 19225
rect 2175 19200 2225 19225
rect 2725 19200 2775 19225
rect 3275 19200 3325 19225
rect 3825 19200 3875 19225
rect 4375 19200 4425 19225
rect 4925 19200 4975 19225
rect 5475 19200 5525 19225
rect 6025 19200 6075 19225
rect 6575 19200 6625 19225
rect 7125 19200 7175 19225
rect 7675 19200 7725 19225
rect 8225 19200 8275 19225
rect 8775 19200 8825 19225
rect 9325 19200 9375 19225
rect 9875 19200 9925 19225
rect 10425 19200 10475 19225
rect 10975 19200 11025 19225
rect 11525 19200 11575 19225
rect 12075 19200 12125 19225
rect 12625 19200 12675 19225
rect 13175 19200 13225 19225
rect 13725 19200 13775 19225
rect 14275 19200 14325 19225
rect 14825 19200 14875 19225
rect 15375 19200 15425 19225
rect 15925 19200 15975 19225
rect 16475 19200 16525 19225
rect 17025 19200 17075 19225
rect 17575 19200 17625 19225
rect 18125 19200 18175 19225
rect 18675 19200 18725 19225
rect 19225 19194 19275 19225
rect 19225 18725 19275 18756
rect 19775 18725 19825 19225
rect -25 18717 56 18725
rect -25 18683 -17 18717
rect 17 18683 56 18717
rect -25 18675 56 18683
rect 494 18675 500 18725
rect 19200 18717 19306 18725
rect 19200 18683 19233 18717
rect 19267 18683 19306 18717
rect 19200 18675 19306 18683
rect 19744 18717 19825 18725
rect 19744 18683 19783 18717
rect 19817 18683 19825 18717
rect 19744 18675 19825 18683
rect -25 18175 25 18675
rect 19225 18644 19275 18675
rect 19225 18175 19275 18206
rect 19775 18175 19825 18675
rect -25 18167 56 18175
rect -25 18133 -17 18167
rect 17 18133 56 18167
rect -25 18125 56 18133
rect 494 18125 500 18175
rect 19200 18167 19306 18175
rect 19200 18133 19233 18167
rect 19267 18133 19306 18167
rect 19200 18125 19306 18133
rect 19744 18167 19825 18175
rect 19744 18133 19783 18167
rect 19817 18133 19825 18167
rect 19744 18125 19825 18133
rect -25 17625 25 18125
rect 19225 18094 19275 18125
rect 19225 17625 19275 17656
rect 19775 17625 19825 18125
rect -25 17617 56 17625
rect -25 17583 -17 17617
rect 17 17583 56 17617
rect -25 17575 56 17583
rect 494 17575 500 17625
rect 19200 17617 19306 17625
rect 19200 17583 19233 17617
rect 19267 17583 19306 17617
rect 19200 17575 19306 17583
rect 19744 17617 19825 17625
rect 19744 17583 19783 17617
rect 19817 17583 19825 17617
rect 19744 17575 19825 17583
rect -25 17075 25 17575
rect 19225 17544 19275 17575
rect 19225 17075 19275 17106
rect 19775 17075 19825 17575
rect -25 17067 56 17075
rect -25 17033 -17 17067
rect 17 17033 56 17067
rect -25 17025 56 17033
rect 494 17025 500 17075
rect 19200 17067 19306 17075
rect 19200 17033 19233 17067
rect 19267 17033 19306 17067
rect 19200 17025 19306 17033
rect 19744 17067 19825 17075
rect 19744 17033 19783 17067
rect 19817 17033 19825 17067
rect 19744 17025 19825 17033
rect -25 16525 25 17025
rect 19225 16994 19275 17025
rect 19225 16525 19275 16556
rect 19775 16525 19825 17025
rect -25 16517 56 16525
rect -25 16483 -17 16517
rect 17 16483 56 16517
rect -25 16475 56 16483
rect 494 16475 500 16525
rect 19200 16517 19306 16525
rect 19200 16483 19233 16517
rect 19267 16483 19306 16517
rect 19200 16475 19306 16483
rect 19744 16517 19825 16525
rect 19744 16483 19783 16517
rect 19817 16483 19825 16517
rect 19744 16475 19825 16483
rect -25 15975 25 16475
rect 19225 16444 19275 16475
rect 19225 15975 19275 16006
rect 19775 15975 19825 16475
rect -25 15967 56 15975
rect -25 15933 -17 15967
rect 17 15933 56 15967
rect -25 15925 56 15933
rect 494 15925 500 15975
rect 19200 15967 19306 15975
rect 19200 15933 19233 15967
rect 19267 15933 19306 15967
rect 19200 15925 19306 15933
rect 19744 15967 19825 15975
rect 19744 15933 19783 15967
rect 19817 15933 19825 15967
rect 19744 15925 19825 15933
rect -25 15425 25 15925
rect 19225 15894 19275 15925
rect 19225 15425 19275 15456
rect 19775 15425 19825 15925
rect -25 15417 56 15425
rect -25 15383 -17 15417
rect 17 15383 56 15417
rect -25 15375 56 15383
rect 494 15375 500 15425
rect 19200 15417 19306 15425
rect 19200 15383 19233 15417
rect 19267 15383 19306 15417
rect 19200 15375 19306 15383
rect 19744 15417 19825 15425
rect 19744 15383 19783 15417
rect 19817 15383 19825 15417
rect 19744 15375 19825 15383
rect -25 14875 25 15375
rect 19225 15344 19275 15375
rect 19225 14875 19275 14906
rect 19775 14875 19825 15375
rect -25 14867 56 14875
rect -25 14833 -17 14867
rect 17 14833 56 14867
rect -25 14825 56 14833
rect 494 14825 500 14875
rect 19200 14867 19306 14875
rect 19200 14833 19233 14867
rect 19267 14833 19306 14867
rect 19200 14825 19306 14833
rect 19744 14867 19825 14875
rect 19744 14833 19783 14867
rect 19817 14833 19825 14867
rect 19744 14825 19825 14833
rect -25 14325 25 14825
rect 19225 14794 19275 14825
rect 19225 14325 19275 14356
rect 19775 14325 19825 14825
rect -25 14317 56 14325
rect -25 14283 -17 14317
rect 17 14283 56 14317
rect -25 14275 56 14283
rect 494 14275 500 14325
rect 19200 14317 19306 14325
rect 19200 14283 19233 14317
rect 19267 14283 19306 14317
rect 19200 14275 19306 14283
rect 19744 14317 19825 14325
rect 19744 14283 19783 14317
rect 19817 14283 19825 14317
rect 19744 14275 19825 14283
rect -25 13775 25 14275
rect 19225 14244 19275 14275
rect 19225 13775 19275 13806
rect 19775 13775 19825 14275
rect -25 13767 56 13775
rect -25 13733 -17 13767
rect 17 13733 56 13767
rect -25 13725 56 13733
rect 494 13725 500 13775
rect 19200 13767 19306 13775
rect 19200 13733 19233 13767
rect 19267 13733 19306 13767
rect 19200 13725 19306 13733
rect 19744 13767 19825 13775
rect 19744 13733 19783 13767
rect 19817 13733 19825 13767
rect 19744 13725 19825 13733
rect -25 13225 25 13725
rect 19225 13694 19275 13725
rect 19225 13225 19275 13256
rect 19775 13225 19825 13725
rect -25 13217 56 13225
rect -25 13183 -17 13217
rect 17 13183 56 13217
rect -25 13175 56 13183
rect 494 13175 500 13225
rect 19200 13217 19306 13225
rect 19200 13183 19233 13217
rect 19267 13183 19306 13217
rect 19200 13175 19306 13183
rect 19744 13217 19825 13225
rect 19744 13183 19783 13217
rect 19817 13183 19825 13217
rect 19744 13175 19825 13183
rect -25 12675 25 13175
rect 19225 13144 19275 13175
rect 19225 12675 19275 12706
rect 19775 12675 19825 13175
rect -25 12667 56 12675
rect -25 12633 -17 12667
rect 17 12633 56 12667
rect -25 12625 56 12633
rect 494 12625 500 12675
rect 19200 12667 19306 12675
rect 19200 12633 19233 12667
rect 19267 12633 19306 12667
rect 19200 12625 19306 12633
rect 19744 12667 19825 12675
rect 19744 12633 19783 12667
rect 19817 12633 19825 12667
rect 19744 12625 19825 12633
rect -25 12125 25 12625
rect 19225 12594 19275 12625
rect 19225 12125 19275 12156
rect 19775 12125 19825 12625
rect -25 12117 56 12125
rect -25 12083 -17 12117
rect 17 12083 56 12117
rect -25 12075 56 12083
rect 494 12075 500 12125
rect 19200 12117 19306 12125
rect 19200 12083 19233 12117
rect 19267 12083 19306 12117
rect 19200 12075 19306 12083
rect 19744 12117 19825 12125
rect 19744 12083 19783 12117
rect 19817 12083 19825 12117
rect 19744 12075 19825 12083
rect -25 11575 25 12075
rect 19225 12044 19275 12075
rect 19225 11575 19275 11606
rect 19775 11575 19825 12075
rect -25 11567 56 11575
rect -25 11533 -17 11567
rect 17 11533 56 11567
rect -25 11525 56 11533
rect 494 11525 500 11575
rect 19200 11567 19306 11575
rect 19200 11533 19233 11567
rect 19267 11533 19306 11567
rect 19200 11525 19306 11533
rect 19744 11567 19825 11575
rect 19744 11533 19783 11567
rect 19817 11533 19825 11567
rect 19744 11525 19825 11533
rect -25 11025 25 11525
rect 19225 11494 19275 11525
rect 19225 11025 19275 11056
rect 19775 11025 19825 11525
rect -25 11017 56 11025
rect -25 10983 -17 11017
rect 17 10983 56 11017
rect -25 10975 56 10983
rect 494 10975 500 11025
rect 19200 11017 19306 11025
rect 19200 10983 19233 11017
rect 19267 10983 19306 11017
rect 19200 10975 19306 10983
rect 19744 11017 19825 11025
rect 19744 10983 19783 11017
rect 19817 10983 19825 11017
rect 19744 10975 19825 10983
rect -25 10475 25 10975
rect 19225 10944 19275 10975
rect 19225 10475 19275 10506
rect 19775 10475 19825 10975
rect -25 10467 56 10475
rect -25 10433 -17 10467
rect 17 10433 56 10467
rect -25 10425 56 10433
rect 494 10425 500 10475
rect 19200 10467 19306 10475
rect 19200 10433 19233 10467
rect 19267 10433 19306 10467
rect 19200 10425 19306 10433
rect 19744 10467 19825 10475
rect 19744 10433 19783 10467
rect 19817 10433 19825 10467
rect 19744 10425 19825 10433
rect -25 9925 25 10425
rect 19225 10394 19275 10425
rect 19225 9925 19275 9956
rect 19775 9925 19825 10425
rect -25 9917 56 9925
rect -25 9883 -17 9917
rect 17 9883 56 9917
rect -25 9875 56 9883
rect 494 9875 500 9925
rect 19200 9917 19306 9925
rect 19200 9883 19233 9917
rect 19267 9883 19306 9917
rect 19200 9875 19306 9883
rect 19744 9917 19825 9925
rect 19744 9883 19783 9917
rect 19817 9883 19825 9917
rect 19744 9875 19825 9883
rect -25 9375 25 9875
rect 19225 9844 19275 9875
rect 19225 9375 19275 9406
rect 19775 9375 19825 9875
rect -25 9367 56 9375
rect -25 9333 -17 9367
rect 17 9333 56 9367
rect -25 9325 56 9333
rect 494 9325 500 9375
rect 19200 9367 19306 9375
rect 19200 9333 19233 9367
rect 19267 9333 19306 9367
rect 19200 9325 19306 9333
rect 19744 9367 19825 9375
rect 19744 9333 19783 9367
rect 19817 9333 19825 9367
rect 19744 9325 19825 9333
rect -25 8825 25 9325
rect 19225 9294 19275 9325
rect 19225 8825 19275 8856
rect 19775 8825 19825 9325
rect -25 8817 56 8825
rect -25 8783 -17 8817
rect 17 8783 56 8817
rect -25 8775 56 8783
rect 494 8775 500 8825
rect 19200 8817 19306 8825
rect 19200 8783 19233 8817
rect 19267 8783 19306 8817
rect 19200 8775 19306 8783
rect 19744 8817 19825 8825
rect 19744 8783 19783 8817
rect 19817 8783 19825 8817
rect 19744 8775 19825 8783
rect -25 8275 25 8775
rect 19225 8744 19275 8775
rect 19225 8275 19275 8306
rect 19775 8275 19825 8775
rect -25 8267 56 8275
rect -25 8233 -17 8267
rect 17 8233 56 8267
rect -25 8225 56 8233
rect 494 8225 500 8275
rect 19200 8267 19306 8275
rect 19200 8233 19233 8267
rect 19267 8233 19306 8267
rect 19200 8225 19306 8233
rect 19744 8267 19825 8275
rect 19744 8233 19783 8267
rect 19817 8233 19825 8267
rect 19744 8225 19825 8233
rect -25 7725 25 8225
rect 19225 8194 19275 8225
rect 19225 7725 19275 7756
rect 19775 7725 19825 8225
rect -25 7717 56 7725
rect -25 7683 -17 7717
rect 17 7683 56 7717
rect -25 7675 56 7683
rect 494 7675 500 7725
rect 19200 7717 19306 7725
rect 19200 7683 19233 7717
rect 19267 7683 19306 7717
rect 19200 7675 19306 7683
rect 19744 7717 19825 7725
rect 19744 7683 19783 7717
rect 19817 7683 19825 7717
rect 19744 7675 19825 7683
rect -25 7175 25 7675
rect 19225 7644 19275 7675
rect 19225 7175 19275 7206
rect 19775 7175 19825 7675
rect -25 7167 56 7175
rect -25 7133 -17 7167
rect 17 7133 56 7167
rect -25 7125 56 7133
rect 494 7125 500 7175
rect 19200 7167 19306 7175
rect 19200 7133 19233 7167
rect 19267 7133 19306 7167
rect 19200 7125 19306 7133
rect 19744 7167 19825 7175
rect 19744 7133 19783 7167
rect 19817 7133 19825 7167
rect 19744 7125 19825 7133
rect -25 6625 25 7125
rect 19225 7094 19275 7125
rect 19225 6625 19275 6656
rect 19775 6625 19825 7125
rect -25 6617 56 6625
rect -25 6583 -17 6617
rect 17 6583 56 6617
rect -25 6575 56 6583
rect 494 6575 500 6625
rect 19200 6617 19306 6625
rect 19200 6583 19233 6617
rect 19267 6583 19306 6617
rect 19200 6575 19306 6583
rect 19744 6617 19825 6625
rect 19744 6583 19783 6617
rect 19817 6583 19825 6617
rect 19744 6575 19825 6583
rect -25 6075 25 6575
rect 19225 6544 19275 6575
rect 19225 6075 19275 6106
rect 19775 6075 19825 6575
rect -25 6067 56 6075
rect -25 6033 -17 6067
rect 17 6033 56 6067
rect -25 6025 56 6033
rect 494 6025 500 6075
rect 19200 6067 19306 6075
rect 19200 6033 19233 6067
rect 19267 6033 19306 6067
rect 19200 6025 19306 6033
rect 19744 6067 19825 6075
rect 19744 6033 19783 6067
rect 19817 6033 19825 6067
rect 19744 6025 19825 6033
rect -25 5525 25 6025
rect 19225 5994 19275 6025
rect 19225 5525 19275 5556
rect 19775 5525 19825 6025
rect -25 5517 56 5525
rect -25 5483 -17 5517
rect 17 5483 56 5517
rect -25 5475 56 5483
rect 494 5475 500 5525
rect 19200 5517 19306 5525
rect 19200 5483 19233 5517
rect 19267 5483 19306 5517
rect 19200 5475 19306 5483
rect 19744 5517 19825 5525
rect 19744 5483 19783 5517
rect 19817 5483 19825 5517
rect 19744 5475 19825 5483
rect -25 4975 25 5475
rect 19225 5444 19275 5475
rect 19225 4975 19275 5006
rect 19775 4975 19825 5475
rect -25 4967 56 4975
rect -25 4933 -17 4967
rect 17 4933 56 4967
rect -25 4925 56 4933
rect 494 4925 500 4975
rect 19200 4967 19306 4975
rect 19200 4933 19233 4967
rect 19267 4933 19306 4967
rect 19200 4925 19306 4933
rect 19744 4967 19825 4975
rect 19744 4933 19783 4967
rect 19817 4933 19825 4967
rect 19744 4925 19825 4933
rect -25 4425 25 4925
rect 19225 4894 19275 4925
rect 19225 4425 19275 4456
rect 19775 4425 19825 4925
rect -25 4417 56 4425
rect -25 4383 -17 4417
rect 17 4383 56 4417
rect -25 4375 56 4383
rect 494 4375 500 4425
rect 19200 4417 19306 4425
rect 19200 4383 19233 4417
rect 19267 4383 19306 4417
rect 19200 4375 19306 4383
rect 19744 4417 19825 4425
rect 19744 4383 19783 4417
rect 19817 4383 19825 4417
rect 19744 4375 19825 4383
rect -25 3875 25 4375
rect 19225 4344 19275 4375
rect 19225 3875 19275 3906
rect 19775 3875 19825 4375
rect -25 3867 56 3875
rect -25 3833 -17 3867
rect 17 3833 56 3867
rect -25 3825 56 3833
rect 494 3825 500 3875
rect 19200 3867 19306 3875
rect 19200 3833 19233 3867
rect 19267 3833 19306 3867
rect 19200 3825 19306 3833
rect 19744 3867 19825 3875
rect 19744 3833 19783 3867
rect 19817 3833 19825 3867
rect 19744 3825 19825 3833
rect -25 3325 25 3825
rect 19225 3794 19275 3825
rect 19225 3325 19275 3356
rect 19775 3325 19825 3825
rect -25 3317 56 3325
rect -25 3283 -17 3317
rect 17 3283 56 3317
rect -25 3275 56 3283
rect 494 3275 500 3325
rect 19200 3317 19306 3325
rect 19200 3283 19233 3317
rect 19267 3283 19306 3317
rect 19200 3275 19306 3283
rect 19744 3317 19825 3325
rect 19744 3283 19783 3317
rect 19817 3283 19825 3317
rect 19744 3275 19825 3283
rect -25 2775 25 3275
rect 19225 3244 19275 3275
rect 19225 2775 19275 2806
rect 19775 2775 19825 3275
rect -25 2767 56 2775
rect -25 2733 -17 2767
rect 17 2733 56 2767
rect -25 2725 56 2733
rect 494 2725 500 2775
rect 19200 2767 19306 2775
rect 19200 2733 19233 2767
rect 19267 2733 19306 2767
rect 19200 2725 19306 2733
rect 19744 2767 19825 2775
rect 19744 2733 19783 2767
rect 19817 2733 19825 2767
rect 19744 2725 19825 2733
rect -25 2225 25 2725
rect 19225 2694 19275 2725
rect 19225 2225 19275 2256
rect 19775 2225 19825 2725
rect -25 2217 56 2225
rect -25 2183 -17 2217
rect 17 2183 56 2217
rect -25 2175 56 2183
rect 494 2175 500 2225
rect 19200 2217 19306 2225
rect 19200 2183 19233 2217
rect 19267 2183 19306 2217
rect 19200 2175 19306 2183
rect 19744 2217 19825 2225
rect 19744 2183 19783 2217
rect 19817 2183 19825 2217
rect 19744 2175 19825 2183
rect -25 1675 25 2175
rect 19225 2144 19275 2175
rect 19225 1675 19275 1706
rect 19775 1675 19825 2175
rect -25 1667 56 1675
rect -25 1633 -17 1667
rect 17 1633 56 1667
rect -25 1625 56 1633
rect 494 1625 500 1675
rect 19200 1667 19306 1675
rect 19200 1633 19233 1667
rect 19267 1633 19306 1667
rect 19200 1625 19306 1633
rect 19744 1667 19825 1675
rect 19744 1633 19783 1667
rect 19817 1633 19825 1667
rect 19744 1625 19825 1633
rect -25 1125 25 1625
rect 19225 1594 19275 1625
rect 19225 1125 19275 1156
rect 19775 1125 19825 1625
rect -25 1117 56 1125
rect -25 1083 -17 1117
rect 17 1083 56 1117
rect -25 1075 56 1083
rect 494 1075 500 1125
rect 19200 1117 19306 1125
rect 19200 1083 19233 1117
rect 19267 1083 19306 1117
rect 19200 1075 19306 1083
rect 19744 1117 19825 1125
rect 19744 1083 19783 1117
rect 19817 1083 19825 1117
rect 19744 1075 19825 1083
rect -25 575 25 1075
rect 19225 1044 19275 1075
rect 19225 575 19275 606
rect 19775 575 19825 1075
rect -25 567 56 575
rect -25 533 -17 567
rect 17 533 56 567
rect -25 525 56 533
rect 494 525 500 575
rect 19200 567 19306 575
rect 19200 533 19233 567
rect 19267 533 19306 567
rect 19200 525 19306 533
rect 19744 567 19825 575
rect 19744 533 19783 567
rect 19817 533 19825 567
rect 19744 525 19825 533
rect -25 25 25 525
rect 525 494 575 500
rect 1075 494 1125 500
rect 1625 494 1675 500
rect 2175 494 2225 500
rect 2725 494 2775 500
rect 3275 494 3325 500
rect 3825 494 3875 500
rect 4375 494 4425 500
rect 4925 494 4975 500
rect 5475 494 5525 500
rect 6025 494 6075 500
rect 6575 494 6625 500
rect 7125 494 7175 500
rect 7675 494 7725 500
rect 8225 494 8275 500
rect 8775 494 8825 500
rect 9325 494 9375 500
rect 9875 494 9925 500
rect 10425 494 10475 500
rect 10975 494 11025 500
rect 11525 494 11575 500
rect 12075 494 12125 500
rect 12625 494 12675 500
rect 13175 494 13225 500
rect 13725 494 13775 500
rect 14275 494 14325 500
rect 14825 494 14875 500
rect 15375 494 15425 500
rect 15925 494 15975 500
rect 16475 494 16525 500
rect 17025 494 17075 500
rect 17575 494 17625 500
rect 18125 494 18175 500
rect 18675 494 18725 500
rect 19225 494 19275 525
rect 525 25 575 56
rect 1075 25 1125 56
rect 1625 25 1675 56
rect 2175 25 2225 56
rect 2725 25 2775 56
rect 3275 25 3325 56
rect 3825 25 3875 56
rect 4375 25 4425 56
rect 4925 25 4975 56
rect 5475 25 5525 56
rect 6025 25 6075 56
rect 6575 25 6625 56
rect 7125 25 7175 56
rect 7675 25 7725 56
rect 8225 25 8275 56
rect 8775 25 8825 56
rect 9325 25 9375 56
rect 9875 25 9925 56
rect 10425 25 10475 56
rect 10975 25 11025 56
rect 11525 25 11575 56
rect 12075 25 12125 56
rect 12625 25 12675 56
rect 13175 25 13225 56
rect 13725 25 13775 56
rect 14275 25 14325 56
rect 14825 25 14875 56
rect 15375 25 15425 56
rect 15925 25 15975 56
rect 16475 25 16525 56
rect 17025 25 17075 56
rect 17575 25 17625 56
rect 18125 25 18175 56
rect 18675 25 18725 56
rect 19225 25 19275 56
rect 19775 25 19825 525
rect -25 17 19825 25
rect -25 -17 -17 17
rect 17 -17 533 17
rect 567 -17 1083 17
rect 1117 -17 1633 17
rect 1667 -17 2183 17
rect 2217 -17 2733 17
rect 2767 -17 3283 17
rect 3317 -17 3833 17
rect 3867 -17 4383 17
rect 4417 -17 4933 17
rect 4967 -17 5483 17
rect 5517 -17 6033 17
rect 6067 -17 6583 17
rect 6617 -17 7133 17
rect 7167 -17 7683 17
rect 7717 -17 8233 17
rect 8267 -17 8783 17
rect 8817 -17 9333 17
rect 9367 -17 9883 17
rect 9917 -17 10433 17
rect 10467 -17 10983 17
rect 11017 -17 11533 17
rect 11567 -17 12083 17
rect 12117 -17 12633 17
rect 12667 -17 13183 17
rect 13217 -17 13733 17
rect 13767 -17 14283 17
rect 14317 -17 14833 17
rect 14867 -17 15383 17
rect 15417 -17 15933 17
rect 15967 -17 16483 17
rect 16517 -17 17033 17
rect 17067 -17 17583 17
rect 17617 -17 18133 17
rect 18167 -17 18683 17
rect 18717 -17 19233 17
rect 19267 -17 19783 17
rect 19817 -17 19825 17
rect -25 -25 19825 -17
<< polycont >>
rect -17 19783 17 19817
rect 533 19783 567 19817
rect 1083 19783 1117 19817
rect 1633 19783 1667 19817
rect 2183 19783 2217 19817
rect 2733 19783 2767 19817
rect 3283 19783 3317 19817
rect 3833 19783 3867 19817
rect 4383 19783 4417 19817
rect 4933 19783 4967 19817
rect 5483 19783 5517 19817
rect 6033 19783 6067 19817
rect 6583 19783 6617 19817
rect 7133 19783 7167 19817
rect 7683 19783 7717 19817
rect 8233 19783 8267 19817
rect 8783 19783 8817 19817
rect 9333 19783 9367 19817
rect 9883 19783 9917 19817
rect 10433 19783 10467 19817
rect 10983 19783 11017 19817
rect 11533 19783 11567 19817
rect 12083 19783 12117 19817
rect 12633 19783 12667 19817
rect 13183 19783 13217 19817
rect 13733 19783 13767 19817
rect 14283 19783 14317 19817
rect 14833 19783 14867 19817
rect 15383 19783 15417 19817
rect 15933 19783 15967 19817
rect 16483 19783 16517 19817
rect 17033 19783 17067 19817
rect 17583 19783 17617 19817
rect 18133 19783 18167 19817
rect 18683 19783 18717 19817
rect 19233 19783 19267 19817
rect 19783 19783 19817 19817
rect -17 19233 17 19267
rect 533 19233 567 19267
rect 1083 19233 1117 19267
rect 1633 19233 1667 19267
rect 2183 19233 2217 19267
rect 2733 19233 2767 19267
rect 3283 19233 3317 19267
rect 3833 19233 3867 19267
rect 4383 19233 4417 19267
rect 4933 19233 4967 19267
rect 5483 19233 5517 19267
rect 6033 19233 6067 19267
rect 6583 19233 6617 19267
rect 7133 19233 7167 19267
rect 7683 19233 7717 19267
rect 8233 19233 8267 19267
rect 8783 19233 8817 19267
rect 9333 19233 9367 19267
rect 9883 19233 9917 19267
rect 10433 19233 10467 19267
rect 10983 19233 11017 19267
rect 11533 19233 11567 19267
rect 12083 19233 12117 19267
rect 12633 19233 12667 19267
rect 13183 19233 13217 19267
rect 13733 19233 13767 19267
rect 14283 19233 14317 19267
rect 14833 19233 14867 19267
rect 15383 19233 15417 19267
rect 15933 19233 15967 19267
rect 16483 19233 16517 19267
rect 17033 19233 17067 19267
rect 17583 19233 17617 19267
rect 18133 19233 18167 19267
rect 18683 19233 18717 19267
rect 19233 19233 19267 19267
rect 19783 19233 19817 19267
rect -17 18683 17 18717
rect 19233 18683 19267 18717
rect 19783 18683 19817 18717
rect -17 18133 17 18167
rect 19233 18133 19267 18167
rect 19783 18133 19817 18167
rect -17 17583 17 17617
rect 19233 17583 19267 17617
rect 19783 17583 19817 17617
rect -17 17033 17 17067
rect 19233 17033 19267 17067
rect 19783 17033 19817 17067
rect -17 16483 17 16517
rect 19233 16483 19267 16517
rect 19783 16483 19817 16517
rect -17 15933 17 15967
rect 19233 15933 19267 15967
rect 19783 15933 19817 15967
rect -17 15383 17 15417
rect 19233 15383 19267 15417
rect 19783 15383 19817 15417
rect -17 14833 17 14867
rect 19233 14833 19267 14867
rect 19783 14833 19817 14867
rect -17 14283 17 14317
rect 19233 14283 19267 14317
rect 19783 14283 19817 14317
rect -17 13733 17 13767
rect 19233 13733 19267 13767
rect 19783 13733 19817 13767
rect -17 13183 17 13217
rect 19233 13183 19267 13217
rect 19783 13183 19817 13217
rect -17 12633 17 12667
rect 19233 12633 19267 12667
rect 19783 12633 19817 12667
rect -17 12083 17 12117
rect 19233 12083 19267 12117
rect 19783 12083 19817 12117
rect -17 11533 17 11567
rect 19233 11533 19267 11567
rect 19783 11533 19817 11567
rect -17 10983 17 11017
rect 19233 10983 19267 11017
rect 19783 10983 19817 11017
rect -17 10433 17 10467
rect 19233 10433 19267 10467
rect 19783 10433 19817 10467
rect -17 9883 17 9917
rect 19233 9883 19267 9917
rect 19783 9883 19817 9917
rect -17 9333 17 9367
rect 19233 9333 19267 9367
rect 19783 9333 19817 9367
rect -17 8783 17 8817
rect 19233 8783 19267 8817
rect 19783 8783 19817 8817
rect -17 8233 17 8267
rect 19233 8233 19267 8267
rect 19783 8233 19817 8267
rect -17 7683 17 7717
rect 19233 7683 19267 7717
rect 19783 7683 19817 7717
rect -17 7133 17 7167
rect 19233 7133 19267 7167
rect 19783 7133 19817 7167
rect -17 6583 17 6617
rect 19233 6583 19267 6617
rect 19783 6583 19817 6617
rect -17 6033 17 6067
rect 19233 6033 19267 6067
rect 19783 6033 19817 6067
rect -17 5483 17 5517
rect 19233 5483 19267 5517
rect 19783 5483 19817 5517
rect -17 4933 17 4967
rect 19233 4933 19267 4967
rect 19783 4933 19817 4967
rect -17 4383 17 4417
rect 19233 4383 19267 4417
rect 19783 4383 19817 4417
rect -17 3833 17 3867
rect 19233 3833 19267 3867
rect 19783 3833 19817 3867
rect -17 3283 17 3317
rect 19233 3283 19267 3317
rect 19783 3283 19817 3317
rect -17 2733 17 2767
rect 19233 2733 19267 2767
rect 19783 2733 19817 2767
rect -17 2183 17 2217
rect 19233 2183 19267 2217
rect 19783 2183 19817 2217
rect -17 1633 17 1667
rect 19233 1633 19267 1667
rect 19783 1633 19817 1667
rect -17 1083 17 1117
rect 19233 1083 19267 1117
rect 19783 1083 19817 1117
rect -17 533 17 567
rect 19233 533 19267 567
rect 19783 533 19817 567
rect -17 -17 17 17
rect 533 -17 567 17
rect 1083 -17 1117 17
rect 1633 -17 1667 17
rect 2183 -17 2217 17
rect 2733 -17 2767 17
rect 3283 -17 3317 17
rect 3833 -17 3867 17
rect 4383 -17 4417 17
rect 4933 -17 4967 17
rect 5483 -17 5517 17
rect 6033 -17 6067 17
rect 6583 -17 6617 17
rect 7133 -17 7167 17
rect 7683 -17 7717 17
rect 8233 -17 8267 17
rect 8783 -17 8817 17
rect 9333 -17 9367 17
rect 9883 -17 9917 17
rect 10433 -17 10467 17
rect 10983 -17 11017 17
rect 11533 -17 11567 17
rect 12083 -17 12117 17
rect 12633 -17 12667 17
rect 13183 -17 13217 17
rect 13733 -17 13767 17
rect 14283 -17 14317 17
rect 14833 -17 14867 17
rect 15383 -17 15417 17
rect 15933 -17 15967 17
rect 16483 -17 16517 17
rect 17033 -17 17067 17
rect 17583 -17 17617 17
rect 18133 -17 18167 17
rect 18683 -17 18717 17
rect 19233 -17 19267 17
rect 19783 -17 19817 17
<< locali >>
rect -5000 24788 24800 24800
rect -5000 -4988 -4988 24788
rect -1012 20800 20812 20812
rect -1012 -1000 -1000 20800
rect -500 20288 20300 20300
rect -500 -488 -488 20288
rect -212 20000 20012 20012
rect -212 -200 -200 20000
rect -25 19817 25 19825
rect -25 19783 -17 19817
rect 17 19783 25 19817
rect -25 19775 25 19783
rect 525 19817 575 19825
rect 525 19783 533 19817
rect 567 19783 575 19817
rect 525 19775 575 19783
rect 1075 19817 1125 19825
rect 1075 19783 1083 19817
rect 1117 19783 1125 19817
rect 1075 19775 1125 19783
rect 1625 19817 1675 19825
rect 1625 19783 1633 19817
rect 1667 19783 1675 19817
rect 1625 19775 1675 19783
rect 2175 19817 2225 19825
rect 2175 19783 2183 19817
rect 2217 19783 2225 19817
rect 2175 19775 2225 19783
rect 2725 19817 2775 19825
rect 2725 19783 2733 19817
rect 2767 19783 2775 19817
rect 2725 19775 2775 19783
rect 3275 19817 3325 19825
rect 3275 19783 3283 19817
rect 3317 19783 3325 19817
rect 3275 19775 3325 19783
rect 3825 19817 3875 19825
rect 3825 19783 3833 19817
rect 3867 19783 3875 19817
rect 3825 19775 3875 19783
rect 4375 19817 4425 19825
rect 4375 19783 4383 19817
rect 4417 19783 4425 19817
rect 4375 19775 4425 19783
rect 4925 19817 4975 19825
rect 4925 19783 4933 19817
rect 4967 19783 4975 19817
rect 4925 19775 4975 19783
rect 5475 19817 5525 19825
rect 5475 19783 5483 19817
rect 5517 19783 5525 19817
rect 5475 19775 5525 19783
rect 6025 19817 6075 19825
rect 6025 19783 6033 19817
rect 6067 19783 6075 19817
rect 6025 19775 6075 19783
rect 6575 19817 6625 19825
rect 6575 19783 6583 19817
rect 6617 19783 6625 19817
rect 6575 19775 6625 19783
rect 7125 19817 7175 19825
rect 7125 19783 7133 19817
rect 7167 19783 7175 19817
rect 7125 19775 7175 19783
rect 7675 19817 7725 19825
rect 7675 19783 7683 19817
rect 7717 19783 7725 19817
rect 7675 19775 7725 19783
rect 8225 19817 8275 19825
rect 8225 19783 8233 19817
rect 8267 19783 8275 19817
rect 8225 19775 8275 19783
rect 8775 19817 8825 19825
rect 8775 19783 8783 19817
rect 8817 19783 8825 19817
rect 8775 19775 8825 19783
rect 9325 19817 9375 19825
rect 9325 19783 9333 19817
rect 9367 19783 9375 19817
rect 9325 19775 9375 19783
rect 9875 19817 9925 19825
rect 9875 19783 9883 19817
rect 9917 19783 9925 19817
rect 9875 19775 9925 19783
rect 10425 19817 10475 19825
rect 10425 19783 10433 19817
rect 10467 19783 10475 19817
rect 10425 19775 10475 19783
rect 10975 19817 11025 19825
rect 10975 19783 10983 19817
rect 11017 19783 11025 19817
rect 10975 19775 11025 19783
rect 11525 19817 11575 19825
rect 11525 19783 11533 19817
rect 11567 19783 11575 19817
rect 11525 19775 11575 19783
rect 12075 19817 12125 19825
rect 12075 19783 12083 19817
rect 12117 19783 12125 19817
rect 12075 19775 12125 19783
rect 12625 19817 12675 19825
rect 12625 19783 12633 19817
rect 12667 19783 12675 19817
rect 12625 19775 12675 19783
rect 13175 19817 13225 19825
rect 13175 19783 13183 19817
rect 13217 19783 13225 19817
rect 13175 19775 13225 19783
rect 13725 19817 13775 19825
rect 13725 19783 13733 19817
rect 13767 19783 13775 19817
rect 13725 19775 13775 19783
rect 14275 19817 14325 19825
rect 14275 19783 14283 19817
rect 14317 19783 14325 19817
rect 14275 19775 14325 19783
rect 14825 19817 14875 19825
rect 14825 19783 14833 19817
rect 14867 19783 14875 19817
rect 14825 19775 14875 19783
rect 15375 19817 15425 19825
rect 15375 19783 15383 19817
rect 15417 19783 15425 19817
rect 15375 19775 15425 19783
rect 15925 19817 15975 19825
rect 15925 19783 15933 19817
rect 15967 19783 15975 19817
rect 15925 19775 15975 19783
rect 16475 19817 16525 19825
rect 16475 19783 16483 19817
rect 16517 19783 16525 19817
rect 16475 19775 16525 19783
rect 17025 19817 17075 19825
rect 17025 19783 17033 19817
rect 17067 19783 17075 19817
rect 17025 19775 17075 19783
rect 17575 19817 17625 19825
rect 17575 19783 17583 19817
rect 17617 19783 17625 19817
rect 17575 19775 17625 19783
rect 18125 19817 18175 19825
rect 18125 19783 18133 19817
rect 18167 19783 18175 19817
rect 18125 19775 18175 19783
rect 18675 19817 18725 19825
rect 18675 19783 18683 19817
rect 18717 19783 18725 19817
rect 18675 19775 18725 19783
rect 19225 19817 19275 19825
rect 19225 19783 19233 19817
rect 19267 19783 19275 19817
rect 19225 19775 19275 19783
rect 19775 19817 19825 19825
rect 19775 19783 19783 19817
rect 19817 19783 19825 19817
rect 19775 19775 19825 19783
rect 598 19746 1052 19752
rect 1698 19746 2152 19752
rect 2798 19746 3252 19752
rect 3898 19746 4352 19752
rect 4998 19746 5452 19752
rect 6098 19746 6552 19752
rect 7198 19746 7652 19752
rect 8298 19746 8752 19752
rect 9398 19746 9852 19752
rect 10498 19746 10952 19752
rect 11598 19746 12052 19752
rect 12698 19746 13152 19752
rect 13798 19746 14252 19752
rect 14898 19746 15352 19752
rect 15998 19746 16452 19752
rect 17098 19746 17552 19752
rect 18198 19746 18652 19752
rect 19298 19746 19752 19752
rect 502 19738 519 19746
rect 461 19312 502 19339
rect 461 19304 519 19312
rect 581 19738 1069 19746
rect 598 19690 1052 19738
rect 598 19360 660 19690
rect 990 19360 1052 19690
rect 598 19312 1052 19360
rect 581 19304 1069 19312
rect 1131 19738 1148 19746
rect 1602 19738 1619 19746
rect 1148 19312 1189 19339
rect 1131 19304 1189 19312
rect 461 19298 496 19304
rect 598 19298 1052 19304
rect 1154 19298 1189 19304
rect 1561 19312 1602 19339
rect 1561 19304 1619 19312
rect 1681 19738 2169 19746
rect 1698 19690 2152 19738
rect 1698 19360 1760 19690
rect 2090 19360 2152 19690
rect 1698 19312 2152 19360
rect 1681 19304 2169 19312
rect 2231 19738 2248 19746
rect 2702 19738 2719 19746
rect 2248 19312 2289 19339
rect 2231 19304 2289 19312
rect 1561 19298 1596 19304
rect 1698 19298 2152 19304
rect 2254 19298 2289 19304
rect 2661 19312 2702 19339
rect 2661 19304 2719 19312
rect 2781 19738 3269 19746
rect 2798 19690 3252 19738
rect 2798 19360 2860 19690
rect 3190 19360 3252 19690
rect 2798 19312 3252 19360
rect 2781 19304 3269 19312
rect 3331 19738 3348 19746
rect 3802 19738 3819 19746
rect 3348 19312 3389 19339
rect 3331 19304 3389 19312
rect 2661 19298 2696 19304
rect 2798 19298 3252 19304
rect 3354 19298 3389 19304
rect 3761 19312 3802 19339
rect 3761 19304 3819 19312
rect 3881 19738 4369 19746
rect 3898 19690 4352 19738
rect 3898 19360 3960 19690
rect 4290 19360 4352 19690
rect 3898 19312 4352 19360
rect 3881 19304 4369 19312
rect 4431 19738 4448 19746
rect 4902 19738 4919 19746
rect 4448 19312 4489 19339
rect 4431 19304 4489 19312
rect 3761 19298 3796 19304
rect 3898 19298 4352 19304
rect 4454 19298 4489 19304
rect 4861 19312 4902 19339
rect 4861 19304 4919 19312
rect 4981 19738 5469 19746
rect 4998 19690 5452 19738
rect 4998 19360 5060 19690
rect 5390 19360 5452 19690
rect 4998 19312 5452 19360
rect 4981 19304 5469 19312
rect 5531 19738 5548 19746
rect 6002 19738 6019 19746
rect 5548 19312 5589 19339
rect 5531 19304 5589 19312
rect 4861 19298 4896 19304
rect 4998 19298 5452 19304
rect 5554 19298 5589 19304
rect 5961 19312 6002 19339
rect 5961 19304 6019 19312
rect 6081 19738 6569 19746
rect 6098 19690 6552 19738
rect 6098 19360 6160 19690
rect 6490 19360 6552 19690
rect 6098 19312 6552 19360
rect 6081 19304 6569 19312
rect 6631 19738 6648 19746
rect 7102 19738 7119 19746
rect 6648 19312 6689 19339
rect 6631 19304 6689 19312
rect 5961 19298 5996 19304
rect 6098 19298 6552 19304
rect 6654 19298 6689 19304
rect 7061 19312 7102 19339
rect 7061 19304 7119 19312
rect 7181 19738 7669 19746
rect 7198 19690 7652 19738
rect 7198 19360 7260 19690
rect 7590 19360 7652 19690
rect 7198 19312 7652 19360
rect 7181 19304 7669 19312
rect 7731 19738 7748 19746
rect 8202 19738 8219 19746
rect 7748 19312 7789 19339
rect 7731 19304 7789 19312
rect 7061 19298 7096 19304
rect 7198 19298 7652 19304
rect 7754 19298 7789 19304
rect 8161 19312 8202 19339
rect 8161 19304 8219 19312
rect 8281 19738 8769 19746
rect 8298 19690 8752 19738
rect 8298 19360 8360 19690
rect 8690 19360 8752 19690
rect 8298 19312 8752 19360
rect 8281 19304 8769 19312
rect 8831 19738 8848 19746
rect 9302 19738 9319 19746
rect 8848 19312 8889 19339
rect 8831 19304 8889 19312
rect 8161 19298 8196 19304
rect 8298 19298 8752 19304
rect 8854 19298 8889 19304
rect 9261 19312 9302 19339
rect 9261 19304 9319 19312
rect 9381 19738 9869 19746
rect 9398 19690 9852 19738
rect 9398 19360 9460 19690
rect 9790 19360 9852 19690
rect 9398 19312 9852 19360
rect 9381 19304 9869 19312
rect 9931 19738 9948 19746
rect 10402 19738 10419 19746
rect 9948 19312 9989 19339
rect 9931 19304 9989 19312
rect 9261 19298 9296 19304
rect 9398 19298 9852 19304
rect 9954 19298 9989 19304
rect 10361 19312 10402 19339
rect 10361 19304 10419 19312
rect 10481 19738 10969 19746
rect 10498 19690 10952 19738
rect 10498 19360 10560 19690
rect 10890 19360 10952 19690
rect 10498 19312 10952 19360
rect 10481 19304 10969 19312
rect 11031 19738 11048 19746
rect 11502 19738 11519 19746
rect 11048 19312 11089 19339
rect 11031 19304 11089 19312
rect 10361 19298 10396 19304
rect 10498 19298 10952 19304
rect 11054 19298 11089 19304
rect 11461 19312 11502 19339
rect 11461 19304 11519 19312
rect 11581 19738 12069 19746
rect 11598 19690 12052 19738
rect 11598 19360 11660 19690
rect 11990 19360 12052 19690
rect 11598 19312 12052 19360
rect 11581 19304 12069 19312
rect 12131 19738 12148 19746
rect 12602 19738 12619 19746
rect 12148 19312 12189 19339
rect 12131 19304 12189 19312
rect 11461 19298 11496 19304
rect 11598 19298 12052 19304
rect 12154 19298 12189 19304
rect 12561 19312 12602 19339
rect 12561 19304 12619 19312
rect 12681 19738 13169 19746
rect 12698 19690 13152 19738
rect 12698 19360 12760 19690
rect 13090 19360 13152 19690
rect 12698 19312 13152 19360
rect 12681 19304 13169 19312
rect 13231 19738 13248 19746
rect 13702 19738 13719 19746
rect 13248 19312 13289 19339
rect 13231 19304 13289 19312
rect 12561 19298 12596 19304
rect 12698 19298 13152 19304
rect 13254 19298 13289 19304
rect 13661 19312 13702 19339
rect 13661 19304 13719 19312
rect 13781 19738 14269 19746
rect 13798 19690 14252 19738
rect 13798 19360 13860 19690
rect 14190 19360 14252 19690
rect 13798 19312 14252 19360
rect 13781 19304 14269 19312
rect 14331 19738 14348 19746
rect 14802 19738 14819 19746
rect 14348 19312 14389 19339
rect 14331 19304 14389 19312
rect 13661 19298 13696 19304
rect 13798 19298 14252 19304
rect 14354 19298 14389 19304
rect 14761 19312 14802 19339
rect 14761 19304 14819 19312
rect 14881 19738 15369 19746
rect 14898 19690 15352 19738
rect 14898 19360 14960 19690
rect 15290 19360 15352 19690
rect 14898 19312 15352 19360
rect 14881 19304 15369 19312
rect 15431 19738 15448 19746
rect 15902 19738 15919 19746
rect 15448 19312 15489 19339
rect 15431 19304 15489 19312
rect 14761 19298 14796 19304
rect 14898 19298 15352 19304
rect 15454 19298 15489 19304
rect 15861 19312 15902 19339
rect 15861 19304 15919 19312
rect 15981 19738 16469 19746
rect 15998 19690 16452 19738
rect 15998 19360 16060 19690
rect 16390 19360 16452 19690
rect 15998 19312 16452 19360
rect 15981 19304 16469 19312
rect 16531 19738 16548 19746
rect 17002 19738 17019 19746
rect 16548 19312 16589 19339
rect 16531 19304 16589 19312
rect 15861 19298 15896 19304
rect 15998 19298 16452 19304
rect 16554 19298 16589 19304
rect 16961 19312 17002 19339
rect 16961 19304 17019 19312
rect 17081 19738 17569 19746
rect 17098 19690 17552 19738
rect 17098 19360 17160 19690
rect 17490 19360 17552 19690
rect 17098 19312 17552 19360
rect 17081 19304 17569 19312
rect 17631 19738 17648 19746
rect 18102 19738 18119 19746
rect 17648 19312 17689 19339
rect 17631 19304 17689 19312
rect 16961 19298 16996 19304
rect 17098 19298 17552 19304
rect 17654 19298 17689 19304
rect 18061 19312 18102 19339
rect 18061 19304 18119 19312
rect 18181 19738 18669 19746
rect 18198 19690 18652 19738
rect 18198 19360 18260 19690
rect 18590 19360 18652 19690
rect 18198 19312 18652 19360
rect 18181 19304 18669 19312
rect 18731 19738 18748 19746
rect 19202 19738 19219 19746
rect 18748 19312 18789 19339
rect 18731 19304 18789 19312
rect 18061 19298 18096 19304
rect 18198 19298 18652 19304
rect 18754 19298 18789 19304
rect 19161 19312 19202 19339
rect 19161 19304 19219 19312
rect 19281 19738 19752 19746
rect 19298 19690 19752 19738
rect 19298 19360 19360 19690
rect 19690 19360 19752 19690
rect 19298 19312 19752 19360
rect 19281 19304 19752 19312
rect 19161 19298 19196 19304
rect 19298 19298 19752 19304
rect 54 19281 62 19298
rect 488 19281 496 19298
rect 604 19281 612 19298
rect 1038 19281 1046 19298
rect 1154 19281 1162 19298
rect 1588 19281 1596 19298
rect 1704 19281 1712 19298
rect 2138 19281 2146 19298
rect 2254 19281 2262 19298
rect 2688 19281 2696 19298
rect 2804 19281 2812 19298
rect 3238 19281 3246 19298
rect 3354 19281 3362 19298
rect 3788 19281 3796 19298
rect 3904 19281 3912 19298
rect 4338 19281 4346 19298
rect 4454 19281 4462 19298
rect 4888 19281 4896 19298
rect 5004 19281 5012 19298
rect 5438 19281 5446 19298
rect 5554 19281 5562 19298
rect 5988 19281 5996 19298
rect 6104 19281 6112 19298
rect 6538 19281 6546 19298
rect 6654 19281 6662 19298
rect 7088 19281 7096 19298
rect 7204 19281 7212 19298
rect 7638 19281 7646 19298
rect 7754 19281 7762 19298
rect 8188 19281 8196 19298
rect 8304 19281 8312 19298
rect 8738 19281 8746 19298
rect 8854 19281 8862 19298
rect 9288 19281 9296 19298
rect 9404 19281 9412 19298
rect 9838 19281 9846 19298
rect 9954 19281 9962 19298
rect 10388 19281 10396 19298
rect 10504 19281 10512 19298
rect 10938 19281 10946 19298
rect 11054 19281 11062 19298
rect 11488 19281 11496 19298
rect 11604 19281 11612 19298
rect 12038 19281 12046 19298
rect 12154 19281 12162 19298
rect 12588 19281 12596 19298
rect 12704 19281 12712 19298
rect 13138 19281 13146 19298
rect 13254 19281 13262 19298
rect 13688 19281 13696 19298
rect 13804 19281 13812 19298
rect 14238 19281 14246 19298
rect 14354 19281 14362 19298
rect 14788 19281 14796 19298
rect 14904 19281 14912 19298
rect 15338 19281 15346 19298
rect 15454 19281 15462 19298
rect 15888 19281 15896 19298
rect 16004 19281 16012 19298
rect 16438 19281 16446 19298
rect 16554 19281 16562 19298
rect 16988 19281 16996 19298
rect 17104 19281 17112 19298
rect 17538 19281 17546 19298
rect 17654 19281 17662 19298
rect 18088 19281 18096 19298
rect 18204 19281 18212 19298
rect 18638 19281 18646 19298
rect 18754 19281 18762 19298
rect 19188 19281 19196 19298
rect 19304 19281 19312 19298
rect 19738 19281 19746 19298
rect -25 19267 25 19275
rect -25 19233 -17 19267
rect 17 19233 25 19267
rect -25 19225 25 19233
rect 525 19267 575 19275
rect 525 19233 533 19267
rect 567 19233 575 19267
rect 525 19225 575 19233
rect 1075 19267 1125 19275
rect 1075 19233 1083 19267
rect 1117 19233 1125 19267
rect 1075 19225 1125 19233
rect 1625 19267 1675 19275
rect 1625 19233 1633 19267
rect 1667 19233 1675 19267
rect 1625 19225 1675 19233
rect 2175 19267 2225 19275
rect 2175 19233 2183 19267
rect 2217 19233 2225 19267
rect 2175 19225 2225 19233
rect 2725 19267 2775 19275
rect 2725 19233 2733 19267
rect 2767 19233 2775 19267
rect 2725 19225 2775 19233
rect 3275 19267 3325 19275
rect 3275 19233 3283 19267
rect 3317 19233 3325 19267
rect 3275 19225 3325 19233
rect 3825 19267 3875 19275
rect 3825 19233 3833 19267
rect 3867 19233 3875 19267
rect 3825 19225 3875 19233
rect 4375 19267 4425 19275
rect 4375 19233 4383 19267
rect 4417 19233 4425 19267
rect 4375 19225 4425 19233
rect 4925 19267 4975 19275
rect 4925 19233 4933 19267
rect 4967 19233 4975 19267
rect 4925 19225 4975 19233
rect 5475 19267 5525 19275
rect 5475 19233 5483 19267
rect 5517 19233 5525 19267
rect 5475 19225 5525 19233
rect 6025 19267 6075 19275
rect 6025 19233 6033 19267
rect 6067 19233 6075 19267
rect 6025 19225 6075 19233
rect 6575 19267 6625 19275
rect 6575 19233 6583 19267
rect 6617 19233 6625 19267
rect 6575 19225 6625 19233
rect 7125 19267 7175 19275
rect 7125 19233 7133 19267
rect 7167 19233 7175 19267
rect 7125 19225 7175 19233
rect 7675 19267 7725 19275
rect 7675 19233 7683 19267
rect 7717 19233 7725 19267
rect 7675 19225 7725 19233
rect 8225 19267 8275 19275
rect 8225 19233 8233 19267
rect 8267 19233 8275 19267
rect 8225 19225 8275 19233
rect 8775 19267 8825 19275
rect 8775 19233 8783 19267
rect 8817 19233 8825 19267
rect 8775 19225 8825 19233
rect 9325 19267 9375 19275
rect 9325 19233 9333 19267
rect 9367 19233 9375 19267
rect 9325 19225 9375 19233
rect 9875 19267 9925 19275
rect 9875 19233 9883 19267
rect 9917 19233 9925 19267
rect 9875 19225 9925 19233
rect 10425 19267 10475 19275
rect 10425 19233 10433 19267
rect 10467 19233 10475 19267
rect 10425 19225 10475 19233
rect 10975 19267 11025 19275
rect 10975 19233 10983 19267
rect 11017 19233 11025 19267
rect 10975 19225 11025 19233
rect 11525 19267 11575 19275
rect 11525 19233 11533 19267
rect 11567 19233 11575 19267
rect 11525 19225 11575 19233
rect 12075 19267 12125 19275
rect 12075 19233 12083 19267
rect 12117 19233 12125 19267
rect 12075 19225 12125 19233
rect 12625 19267 12675 19275
rect 12625 19233 12633 19267
rect 12667 19233 12675 19267
rect 12625 19225 12675 19233
rect 13175 19267 13225 19275
rect 13175 19233 13183 19267
rect 13217 19233 13225 19267
rect 13175 19225 13225 19233
rect 13725 19267 13775 19275
rect 13725 19233 13733 19267
rect 13767 19233 13775 19267
rect 13725 19225 13775 19233
rect 14275 19267 14325 19275
rect 14275 19233 14283 19267
rect 14317 19233 14325 19267
rect 14275 19225 14325 19233
rect 14825 19267 14875 19275
rect 14825 19233 14833 19267
rect 14867 19233 14875 19267
rect 14825 19225 14875 19233
rect 15375 19267 15425 19275
rect 15375 19233 15383 19267
rect 15417 19233 15425 19267
rect 15375 19225 15425 19233
rect 15925 19267 15975 19275
rect 15925 19233 15933 19267
rect 15967 19233 15975 19267
rect 15925 19225 15975 19233
rect 16475 19267 16525 19275
rect 16475 19233 16483 19267
rect 16517 19233 16525 19267
rect 16475 19225 16525 19233
rect 17025 19267 17075 19275
rect 17025 19233 17033 19267
rect 17067 19233 17075 19267
rect 17025 19225 17075 19233
rect 17575 19267 17625 19275
rect 17575 19233 17583 19267
rect 17617 19233 17625 19267
rect 17575 19225 17625 19233
rect 18125 19267 18175 19275
rect 18125 19233 18133 19267
rect 18167 19233 18175 19267
rect 18125 19225 18175 19233
rect 18675 19267 18725 19275
rect 18675 19233 18683 19267
rect 18717 19233 18725 19267
rect 18675 19225 18725 19233
rect 19225 19267 19275 19275
rect 19225 19233 19233 19267
rect 19267 19233 19275 19267
rect 19225 19225 19275 19233
rect 19775 19267 19825 19275
rect 19775 19233 19783 19267
rect 19817 19233 19825 19267
rect 19775 19225 19825 19233
rect 54 19202 62 19219
rect 488 19202 496 19219
rect 604 19202 612 19219
rect 1038 19202 1046 19219
rect 1154 19202 1162 19219
rect 1588 19202 1596 19219
rect 1704 19202 1712 19219
rect 2138 19202 2146 19219
rect 2254 19202 2262 19219
rect 2688 19202 2696 19219
rect 2804 19202 2812 19219
rect 3238 19202 3246 19219
rect 3354 19202 3362 19219
rect 3788 19202 3796 19219
rect 3904 19202 3912 19219
rect 4338 19202 4346 19219
rect 4454 19202 4462 19219
rect 4888 19202 4896 19219
rect 5004 19202 5012 19219
rect 5438 19202 5446 19219
rect 5554 19202 5562 19219
rect 5988 19202 5996 19219
rect 6104 19202 6112 19219
rect 6538 19202 6546 19219
rect 6654 19202 6662 19219
rect 7088 19202 7096 19219
rect 7204 19202 7212 19219
rect 7638 19202 7646 19219
rect 7754 19202 7762 19219
rect 8188 19202 8196 19219
rect 8304 19202 8312 19219
rect 8738 19202 8746 19219
rect 8854 19202 8862 19219
rect 9288 19202 9296 19219
rect 9404 19202 9412 19219
rect 9838 19202 9846 19219
rect 9954 19202 9962 19219
rect 10388 19202 10396 19219
rect 10504 19202 10512 19219
rect 10938 19202 10946 19219
rect 11054 19202 11062 19219
rect 11488 19202 11496 19219
rect 11604 19202 11612 19219
rect 12038 19202 12046 19219
rect 12154 19202 12162 19219
rect 12588 19202 12596 19219
rect 12704 19202 12712 19219
rect 13138 19202 13146 19219
rect 13254 19202 13262 19219
rect 13688 19202 13696 19219
rect 13804 19202 13812 19219
rect 14238 19202 14246 19219
rect 14354 19202 14362 19219
rect 14788 19202 14796 19219
rect 14904 19202 14912 19219
rect 15338 19202 15346 19219
rect 15454 19202 15462 19219
rect 15888 19202 15896 19219
rect 16004 19202 16012 19219
rect 16438 19202 16446 19219
rect 16554 19202 16562 19219
rect 16988 19202 16996 19219
rect 17104 19202 17112 19219
rect 17538 19202 17546 19219
rect 17654 19202 17662 19219
rect 18088 19202 18096 19219
rect 18204 19202 18212 19219
rect 18638 19202 18646 19219
rect 18754 19202 18762 19219
rect 19188 19202 19196 19219
rect 19304 19202 19312 19219
rect 19738 19202 19746 19219
rect 48 19200 502 19202
rect 604 19200 639 19202
rect 1011 19200 1046 19202
rect 1148 19200 1602 19202
rect 1704 19200 1739 19202
rect 2111 19200 2146 19202
rect 2248 19200 2702 19202
rect 2804 19200 2839 19202
rect 3211 19200 3246 19202
rect 3348 19200 3802 19202
rect 3904 19200 3939 19202
rect 4311 19200 4346 19202
rect 4448 19200 4902 19202
rect 5004 19200 5039 19202
rect 5411 19200 5446 19202
rect 5548 19200 6002 19202
rect 6104 19200 6139 19202
rect 6511 19200 6546 19202
rect 6648 19200 7102 19202
rect 7204 19200 7239 19202
rect 7611 19200 7646 19202
rect 7748 19200 8202 19202
rect 8304 19200 8339 19202
rect 8711 19200 8746 19202
rect 8848 19200 9302 19202
rect 9404 19200 9439 19202
rect 9811 19200 9846 19202
rect 9948 19200 10402 19202
rect 10504 19200 10539 19202
rect 10911 19200 10946 19202
rect 11048 19200 11502 19202
rect 11604 19200 11639 19202
rect 12011 19200 12046 19202
rect 12148 19200 12602 19202
rect 12704 19200 12739 19202
rect 13111 19200 13146 19202
rect 13248 19200 13702 19202
rect 13804 19200 13839 19202
rect 14211 19200 14246 19202
rect 14348 19200 14802 19202
rect 14904 19200 14939 19202
rect 15311 19200 15346 19202
rect 15448 19200 15902 19202
rect 16004 19200 16039 19202
rect 16411 19200 16446 19202
rect 16548 19200 17002 19202
rect 17104 19200 17139 19202
rect 17511 19200 17546 19202
rect 17648 19200 18102 19202
rect 18204 19200 18239 19202
rect 18611 19200 18646 19202
rect 18748 19200 19202 19202
rect 48 19140 500 19200
rect 48 18810 110 19140
rect 440 18810 500 19140
rect 48 18748 500 18810
rect 19200 19196 19202 19200
rect 19304 19196 19339 19202
rect 19200 19188 19219 19196
rect 19200 18762 19202 19188
rect 19200 18754 19219 18762
rect 19281 19188 19339 19196
rect 19298 19161 19339 19188
rect 19298 18762 19339 18789
rect 19281 18754 19339 18762
rect 19200 18748 19202 18754
rect 19304 18748 19339 18754
rect 54 18731 62 18748
rect 488 18731 496 18748
rect 19304 18731 19312 18748
rect 19738 18731 19746 18748
rect -25 18717 25 18725
rect -25 18683 -17 18717
rect 17 18683 25 18717
rect -25 18675 25 18683
rect 19225 18717 19275 18725
rect 19225 18683 19233 18717
rect 19267 18683 19275 18717
rect 19225 18675 19275 18683
rect 19775 18717 19825 18725
rect 19775 18683 19783 18717
rect 19817 18683 19825 18717
rect 19775 18675 19825 18683
rect 54 18652 62 18669
rect 488 18652 496 18669
rect 19304 18652 19312 18669
rect 19738 18652 19746 18669
rect 461 18646 496 18652
rect 19298 18646 19752 18652
rect 461 18611 500 18646
rect 19200 18638 19219 18646
rect 19200 18611 19202 18638
rect 461 18204 500 18239
rect 19200 18212 19202 18239
rect 19200 18204 19219 18212
rect 19281 18638 19752 18646
rect 19298 18590 19752 18638
rect 19298 18260 19360 18590
rect 19690 18260 19752 18590
rect 19298 18212 19752 18260
rect 19281 18204 19752 18212
rect 461 18198 496 18204
rect 19298 18198 19752 18204
rect 54 18181 62 18198
rect 488 18181 496 18198
rect 19304 18181 19312 18198
rect 19738 18181 19746 18198
rect -25 18167 25 18175
rect -25 18133 -17 18167
rect 17 18133 25 18167
rect -25 18125 25 18133
rect 19225 18167 19275 18175
rect 19225 18133 19233 18167
rect 19267 18133 19275 18167
rect 19225 18125 19275 18133
rect 19775 18167 19825 18175
rect 19775 18133 19783 18167
rect 19817 18133 19825 18167
rect 19775 18125 19825 18133
rect 54 18102 62 18119
rect 488 18102 496 18119
rect 19304 18102 19312 18119
rect 19738 18102 19746 18119
rect 48 18040 500 18102
rect 48 17710 110 18040
rect 440 17710 500 18040
rect 48 17648 500 17710
rect 19200 18096 19202 18102
rect 19304 18096 19339 18102
rect 19200 18088 19219 18096
rect 19200 17662 19202 18088
rect 19200 17654 19219 17662
rect 19281 18088 19339 18096
rect 19298 18061 19339 18088
rect 19298 17662 19339 17689
rect 19281 17654 19339 17662
rect 19200 17648 19202 17654
rect 19304 17648 19339 17654
rect 54 17631 62 17648
rect 488 17631 496 17648
rect 19304 17631 19312 17648
rect 19738 17631 19746 17648
rect -25 17617 25 17625
rect -25 17583 -17 17617
rect 17 17583 25 17617
rect -25 17575 25 17583
rect 19225 17617 19275 17625
rect 19225 17583 19233 17617
rect 19267 17583 19275 17617
rect 19225 17575 19275 17583
rect 19775 17617 19825 17625
rect 19775 17583 19783 17617
rect 19817 17583 19825 17617
rect 19775 17575 19825 17583
rect 54 17552 62 17569
rect 488 17552 496 17569
rect 19304 17552 19312 17569
rect 19738 17552 19746 17569
rect 461 17546 496 17552
rect 19298 17546 19752 17552
rect 461 17511 500 17546
rect 19200 17538 19219 17546
rect 19200 17511 19202 17538
rect 461 17104 500 17139
rect 19200 17112 19202 17139
rect 19200 17104 19219 17112
rect 19281 17538 19752 17546
rect 19298 17490 19752 17538
rect 19298 17160 19360 17490
rect 19690 17160 19752 17490
rect 19298 17112 19752 17160
rect 19281 17104 19752 17112
rect 461 17098 496 17104
rect 19298 17098 19752 17104
rect 54 17081 62 17098
rect 488 17081 496 17098
rect 19304 17081 19312 17098
rect 19738 17081 19746 17098
rect -25 17067 25 17075
rect -25 17033 -17 17067
rect 17 17033 25 17067
rect -25 17025 25 17033
rect 19225 17067 19275 17075
rect 19225 17033 19233 17067
rect 19267 17033 19275 17067
rect 19225 17025 19275 17033
rect 19775 17067 19825 17075
rect 19775 17033 19783 17067
rect 19817 17033 19825 17067
rect 19775 17025 19825 17033
rect 54 17002 62 17019
rect 488 17002 496 17019
rect 19304 17002 19312 17019
rect 19738 17002 19746 17019
rect 48 16940 500 17002
rect 48 16610 110 16940
rect 440 16610 500 16940
rect 48 16548 500 16610
rect 19200 16996 19202 17002
rect 19304 16996 19339 17002
rect 19200 16988 19219 16996
rect 19200 16562 19202 16988
rect 19200 16554 19219 16562
rect 19281 16988 19339 16996
rect 19298 16961 19339 16988
rect 19298 16562 19339 16589
rect 19281 16554 19339 16562
rect 19200 16548 19202 16554
rect 19304 16548 19339 16554
rect 54 16531 62 16548
rect 488 16531 496 16548
rect 19304 16531 19312 16548
rect 19738 16531 19746 16548
rect -25 16517 25 16525
rect -25 16483 -17 16517
rect 17 16483 25 16517
rect -25 16475 25 16483
rect 19225 16517 19275 16525
rect 19225 16483 19233 16517
rect 19267 16483 19275 16517
rect 19225 16475 19275 16483
rect 19775 16517 19825 16525
rect 19775 16483 19783 16517
rect 19817 16483 19825 16517
rect 19775 16475 19825 16483
rect 54 16452 62 16469
rect 488 16452 496 16469
rect 19304 16452 19312 16469
rect 19738 16452 19746 16469
rect 461 16446 496 16452
rect 19298 16446 19752 16452
rect 461 16411 500 16446
rect 19200 16438 19219 16446
rect 19200 16411 19202 16438
rect 461 16004 500 16039
rect 19200 16012 19202 16039
rect 19200 16004 19219 16012
rect 19281 16438 19752 16446
rect 19298 16390 19752 16438
rect 19298 16060 19360 16390
rect 19690 16060 19752 16390
rect 19298 16012 19752 16060
rect 19281 16004 19752 16012
rect 461 15998 496 16004
rect 19298 15998 19752 16004
rect 54 15981 62 15998
rect 488 15981 496 15998
rect 19304 15981 19312 15998
rect 19738 15981 19746 15998
rect -25 15967 25 15975
rect -25 15933 -17 15967
rect 17 15933 25 15967
rect -25 15925 25 15933
rect 19225 15967 19275 15975
rect 19225 15933 19233 15967
rect 19267 15933 19275 15967
rect 19225 15925 19275 15933
rect 19775 15967 19825 15975
rect 19775 15933 19783 15967
rect 19817 15933 19825 15967
rect 19775 15925 19825 15933
rect 54 15902 62 15919
rect 488 15902 496 15919
rect 19304 15902 19312 15919
rect 19738 15902 19746 15919
rect 48 15840 500 15902
rect 48 15510 110 15840
rect 440 15510 500 15840
rect 48 15448 500 15510
rect 19200 15896 19202 15902
rect 19304 15896 19339 15902
rect 19200 15888 19219 15896
rect 19200 15462 19202 15888
rect 19200 15454 19219 15462
rect 19281 15888 19339 15896
rect 19298 15861 19339 15888
rect 19298 15462 19339 15489
rect 19281 15454 19339 15462
rect 19200 15448 19202 15454
rect 19304 15448 19339 15454
rect 54 15431 62 15448
rect 488 15431 496 15448
rect 19304 15431 19312 15448
rect 19738 15431 19746 15448
rect -25 15417 25 15425
rect -25 15383 -17 15417
rect 17 15383 25 15417
rect -25 15375 25 15383
rect 19225 15417 19275 15425
rect 19225 15383 19233 15417
rect 19267 15383 19275 15417
rect 19225 15375 19275 15383
rect 19775 15417 19825 15425
rect 19775 15383 19783 15417
rect 19817 15383 19825 15417
rect 19775 15375 19825 15383
rect 54 15352 62 15369
rect 488 15352 496 15369
rect 19304 15352 19312 15369
rect 19738 15352 19746 15369
rect 461 15346 496 15352
rect 19298 15346 19752 15352
rect 461 15311 500 15346
rect 19200 15338 19219 15346
rect 19200 15311 19202 15338
rect 461 14904 500 14939
rect 19200 14912 19202 14939
rect 19200 14904 19219 14912
rect 19281 15338 19752 15346
rect 19298 15290 19752 15338
rect 19298 14960 19360 15290
rect 19690 14960 19752 15290
rect 19298 14912 19752 14960
rect 19281 14904 19752 14912
rect 461 14898 496 14904
rect 19298 14898 19752 14904
rect 54 14881 62 14898
rect 488 14881 496 14898
rect 19304 14881 19312 14898
rect 19738 14881 19746 14898
rect -25 14867 25 14875
rect -25 14833 -17 14867
rect 17 14833 25 14867
rect -25 14825 25 14833
rect 19225 14867 19275 14875
rect 19225 14833 19233 14867
rect 19267 14833 19275 14867
rect 19225 14825 19275 14833
rect 19775 14867 19825 14875
rect 19775 14833 19783 14867
rect 19817 14833 19825 14867
rect 19775 14825 19825 14833
rect 54 14802 62 14819
rect 488 14802 496 14819
rect 19304 14802 19312 14819
rect 19738 14802 19746 14819
rect 48 14740 500 14802
rect 48 14410 110 14740
rect 440 14410 500 14740
rect 48 14348 500 14410
rect 19200 14796 19202 14802
rect 19304 14796 19339 14802
rect 19200 14788 19219 14796
rect 19200 14362 19202 14788
rect 19200 14354 19219 14362
rect 19281 14788 19339 14796
rect 19298 14761 19339 14788
rect 19298 14362 19339 14389
rect 19281 14354 19339 14362
rect 19200 14348 19202 14354
rect 19304 14348 19339 14354
rect 54 14331 62 14348
rect 488 14331 496 14348
rect 19304 14331 19312 14348
rect 19738 14331 19746 14348
rect -25 14317 25 14325
rect -25 14283 -17 14317
rect 17 14283 25 14317
rect -25 14275 25 14283
rect 19225 14317 19275 14325
rect 19225 14283 19233 14317
rect 19267 14283 19275 14317
rect 19225 14275 19275 14283
rect 19775 14317 19825 14325
rect 19775 14283 19783 14317
rect 19817 14283 19825 14317
rect 19775 14275 19825 14283
rect 54 14252 62 14269
rect 488 14252 496 14269
rect 19304 14252 19312 14269
rect 19738 14252 19746 14269
rect 461 14246 496 14252
rect 19298 14246 19752 14252
rect 461 14211 500 14246
rect 19200 14238 19219 14246
rect 19200 14211 19202 14238
rect 461 13804 500 13839
rect 19200 13812 19202 13839
rect 19200 13804 19219 13812
rect 19281 14238 19752 14246
rect 19298 14190 19752 14238
rect 19298 13860 19360 14190
rect 19690 13860 19752 14190
rect 19298 13812 19752 13860
rect 19281 13804 19752 13812
rect 461 13798 496 13804
rect 19298 13798 19752 13804
rect 54 13781 62 13798
rect 488 13781 496 13798
rect 19304 13781 19312 13798
rect 19738 13781 19746 13798
rect -25 13767 25 13775
rect -25 13733 -17 13767
rect 17 13733 25 13767
rect -25 13725 25 13733
rect 19225 13767 19275 13775
rect 19225 13733 19233 13767
rect 19267 13733 19275 13767
rect 19225 13725 19275 13733
rect 19775 13767 19825 13775
rect 19775 13733 19783 13767
rect 19817 13733 19825 13767
rect 19775 13725 19825 13733
rect 54 13702 62 13719
rect 488 13702 496 13719
rect 19304 13702 19312 13719
rect 19738 13702 19746 13719
rect 48 13640 500 13702
rect 48 13310 110 13640
rect 440 13310 500 13640
rect 48 13248 500 13310
rect 19200 13696 19202 13702
rect 19304 13696 19339 13702
rect 19200 13688 19219 13696
rect 19200 13262 19202 13688
rect 19200 13254 19219 13262
rect 19281 13688 19339 13696
rect 19298 13661 19339 13688
rect 19298 13262 19339 13289
rect 19281 13254 19339 13262
rect 19200 13248 19202 13254
rect 19304 13248 19339 13254
rect 54 13231 62 13248
rect 488 13231 496 13248
rect 19304 13231 19312 13248
rect 19738 13231 19746 13248
rect -25 13217 25 13225
rect -25 13183 -17 13217
rect 17 13183 25 13217
rect -25 13175 25 13183
rect 19225 13217 19275 13225
rect 19225 13183 19233 13217
rect 19267 13183 19275 13217
rect 19225 13175 19275 13183
rect 19775 13217 19825 13225
rect 19775 13183 19783 13217
rect 19817 13183 19825 13217
rect 19775 13175 19825 13183
rect 54 13152 62 13169
rect 488 13152 496 13169
rect 19304 13152 19312 13169
rect 19738 13152 19746 13169
rect 461 13146 496 13152
rect 19298 13146 19752 13152
rect 461 13111 500 13146
rect 19200 13138 19219 13146
rect 19200 13111 19202 13138
rect 461 12704 500 12739
rect 19200 12712 19202 12739
rect 19200 12704 19219 12712
rect 19281 13138 19752 13146
rect 19298 13090 19752 13138
rect 19298 12760 19360 13090
rect 19690 12760 19752 13090
rect 19298 12712 19752 12760
rect 19281 12704 19752 12712
rect 461 12698 496 12704
rect 19298 12698 19752 12704
rect 54 12681 62 12698
rect 488 12681 496 12698
rect 19304 12681 19312 12698
rect 19738 12681 19746 12698
rect -25 12667 25 12675
rect -25 12633 -17 12667
rect 17 12633 25 12667
rect -25 12625 25 12633
rect 19225 12667 19275 12675
rect 19225 12633 19233 12667
rect 19267 12633 19275 12667
rect 19225 12625 19275 12633
rect 19775 12667 19825 12675
rect 19775 12633 19783 12667
rect 19817 12633 19825 12667
rect 19775 12625 19825 12633
rect 54 12602 62 12619
rect 488 12602 496 12619
rect 19304 12602 19312 12619
rect 19738 12602 19746 12619
rect 48 12540 500 12602
rect 48 12210 110 12540
rect 440 12210 500 12540
rect 48 12148 500 12210
rect 19200 12596 19202 12602
rect 19304 12596 19339 12602
rect 19200 12588 19219 12596
rect 19200 12162 19202 12588
rect 19200 12154 19219 12162
rect 19281 12588 19339 12596
rect 19298 12561 19339 12588
rect 19298 12162 19339 12189
rect 19281 12154 19339 12162
rect 19200 12148 19202 12154
rect 19304 12148 19339 12154
rect 54 12131 62 12148
rect 488 12131 496 12148
rect 19304 12131 19312 12148
rect 19738 12131 19746 12148
rect -25 12117 25 12125
rect -25 12083 -17 12117
rect 17 12083 25 12117
rect -25 12075 25 12083
rect 19225 12117 19275 12125
rect 19225 12083 19233 12117
rect 19267 12083 19275 12117
rect 19225 12075 19275 12083
rect 19775 12117 19825 12125
rect 19775 12083 19783 12117
rect 19817 12083 19825 12117
rect 19775 12075 19825 12083
rect 54 12052 62 12069
rect 488 12052 496 12069
rect 19304 12052 19312 12069
rect 19738 12052 19746 12069
rect 461 12046 496 12052
rect 19298 12046 19752 12052
rect 461 12011 500 12046
rect 19200 12038 19219 12046
rect 19200 12011 19202 12038
rect 461 11604 500 11639
rect 19200 11612 19202 11639
rect 19200 11604 19219 11612
rect 19281 12038 19752 12046
rect 19298 11990 19752 12038
rect 19298 11660 19360 11990
rect 19690 11660 19752 11990
rect 19298 11612 19752 11660
rect 19281 11604 19752 11612
rect 461 11598 496 11604
rect 19298 11598 19752 11604
rect 54 11581 62 11598
rect 488 11581 496 11598
rect 19304 11581 19312 11598
rect 19738 11581 19746 11598
rect -25 11567 25 11575
rect -25 11533 -17 11567
rect 17 11533 25 11567
rect -25 11525 25 11533
rect 19225 11567 19275 11575
rect 19225 11533 19233 11567
rect 19267 11533 19275 11567
rect 19225 11525 19275 11533
rect 19775 11567 19825 11575
rect 19775 11533 19783 11567
rect 19817 11533 19825 11567
rect 19775 11525 19825 11533
rect 54 11502 62 11519
rect 488 11502 496 11519
rect 19304 11502 19312 11519
rect 19738 11502 19746 11519
rect 48 11440 500 11502
rect 48 11110 110 11440
rect 440 11110 500 11440
rect 48 11048 500 11110
rect 19200 11496 19202 11502
rect 19304 11496 19339 11502
rect 19200 11488 19219 11496
rect 19200 11062 19202 11488
rect 19200 11054 19219 11062
rect 19281 11488 19339 11496
rect 19298 11461 19339 11488
rect 19298 11062 19339 11089
rect 19281 11054 19339 11062
rect 19200 11048 19202 11054
rect 19304 11048 19339 11054
rect 54 11031 62 11048
rect 488 11031 496 11048
rect 19304 11031 19312 11048
rect 19738 11031 19746 11048
rect -25 11017 25 11025
rect -25 10983 -17 11017
rect 17 10983 25 11017
rect -25 10975 25 10983
rect 19225 11017 19275 11025
rect 19225 10983 19233 11017
rect 19267 10983 19275 11017
rect 19225 10975 19275 10983
rect 19775 11017 19825 11025
rect 19775 10983 19783 11017
rect 19817 10983 19825 11017
rect 19775 10975 19825 10983
rect 54 10952 62 10969
rect 488 10952 496 10969
rect 19304 10952 19312 10969
rect 19738 10952 19746 10969
rect 461 10946 496 10952
rect 19298 10946 19752 10952
rect 461 10911 500 10946
rect 19200 10938 19219 10946
rect 19200 10911 19202 10938
rect 461 10504 500 10539
rect 19200 10512 19202 10539
rect 19200 10504 19219 10512
rect 19281 10938 19752 10946
rect 19298 10890 19752 10938
rect 19298 10560 19360 10890
rect 19690 10560 19752 10890
rect 19298 10512 19752 10560
rect 19281 10504 19752 10512
rect 461 10498 496 10504
rect 19298 10498 19752 10504
rect 54 10481 62 10498
rect 488 10481 496 10498
rect 19304 10481 19312 10498
rect 19738 10481 19746 10498
rect -25 10467 25 10475
rect -25 10433 -17 10467
rect 17 10433 25 10467
rect -25 10425 25 10433
rect 19225 10467 19275 10475
rect 19225 10433 19233 10467
rect 19267 10433 19275 10467
rect 19225 10425 19275 10433
rect 19775 10467 19825 10475
rect 19775 10433 19783 10467
rect 19817 10433 19825 10467
rect 19775 10425 19825 10433
rect 54 10402 62 10419
rect 488 10402 496 10419
rect 19304 10402 19312 10419
rect 19738 10402 19746 10419
rect 48 10340 500 10402
rect 48 10010 110 10340
rect 440 10010 500 10340
rect 48 9948 500 10010
rect 19200 10396 19202 10402
rect 19304 10396 19339 10402
rect 19200 10388 19219 10396
rect 19200 9962 19202 10388
rect 19200 9954 19219 9962
rect 19281 10388 19339 10396
rect 19298 10361 19339 10388
rect 19298 9962 19339 9989
rect 19281 9954 19339 9962
rect 19200 9948 19202 9954
rect 19304 9948 19339 9954
rect 54 9931 62 9948
rect 488 9931 496 9948
rect 19304 9931 19312 9948
rect 19738 9931 19746 9948
rect -25 9917 25 9925
rect -25 9883 -17 9917
rect 17 9883 25 9917
rect -25 9875 25 9883
rect 19225 9917 19275 9925
rect 19225 9883 19233 9917
rect 19267 9883 19275 9917
rect 19225 9875 19275 9883
rect 19775 9917 19825 9925
rect 19775 9883 19783 9917
rect 19817 9883 19825 9917
rect 19775 9875 19825 9883
rect 54 9852 62 9869
rect 488 9852 496 9869
rect 19304 9852 19312 9869
rect 19738 9852 19746 9869
rect 461 9846 496 9852
rect 19298 9846 19752 9852
rect 461 9811 500 9846
rect 19200 9838 19219 9846
rect 19200 9811 19202 9838
rect 461 9404 500 9439
rect 19200 9412 19202 9439
rect 19200 9404 19219 9412
rect 19281 9838 19752 9846
rect 19298 9790 19752 9838
rect 19298 9460 19360 9790
rect 19690 9460 19752 9790
rect 19298 9412 19752 9460
rect 19281 9404 19752 9412
rect 461 9398 496 9404
rect 19298 9398 19752 9404
rect 54 9381 62 9398
rect 488 9381 496 9398
rect 19304 9381 19312 9398
rect 19738 9381 19746 9398
rect -25 9367 25 9375
rect -25 9333 -17 9367
rect 17 9333 25 9367
rect -25 9325 25 9333
rect 19225 9367 19275 9375
rect 19225 9333 19233 9367
rect 19267 9333 19275 9367
rect 19225 9325 19275 9333
rect 19775 9367 19825 9375
rect 19775 9333 19783 9367
rect 19817 9333 19825 9367
rect 19775 9325 19825 9333
rect 54 9302 62 9319
rect 488 9302 496 9319
rect 19304 9302 19312 9319
rect 19738 9302 19746 9319
rect 48 9240 500 9302
rect 48 8910 110 9240
rect 440 8910 500 9240
rect 48 8848 500 8910
rect 19200 9296 19202 9302
rect 19304 9296 19339 9302
rect 19200 9288 19219 9296
rect 19200 8862 19202 9288
rect 19200 8854 19219 8862
rect 19281 9288 19339 9296
rect 19298 9261 19339 9288
rect 19298 8862 19339 8889
rect 19281 8854 19339 8862
rect 19200 8848 19202 8854
rect 19304 8848 19339 8854
rect 54 8831 62 8848
rect 488 8831 496 8848
rect 19304 8831 19312 8848
rect 19738 8831 19746 8848
rect -25 8817 25 8825
rect -25 8783 -17 8817
rect 17 8783 25 8817
rect -25 8775 25 8783
rect 19225 8817 19275 8825
rect 19225 8783 19233 8817
rect 19267 8783 19275 8817
rect 19225 8775 19275 8783
rect 19775 8817 19825 8825
rect 19775 8783 19783 8817
rect 19817 8783 19825 8817
rect 19775 8775 19825 8783
rect 54 8752 62 8769
rect 488 8752 496 8769
rect 19304 8752 19312 8769
rect 19738 8752 19746 8769
rect 461 8746 496 8752
rect 19298 8746 19752 8752
rect 461 8711 500 8746
rect 19200 8738 19219 8746
rect 19200 8711 19202 8738
rect 461 8304 500 8339
rect 19200 8312 19202 8339
rect 19200 8304 19219 8312
rect 19281 8738 19752 8746
rect 19298 8690 19752 8738
rect 19298 8360 19360 8690
rect 19690 8360 19752 8690
rect 19298 8312 19752 8360
rect 19281 8304 19752 8312
rect 461 8298 496 8304
rect 19298 8298 19752 8304
rect 54 8281 62 8298
rect 488 8281 496 8298
rect 19304 8281 19312 8298
rect 19738 8281 19746 8298
rect -25 8267 25 8275
rect -25 8233 -17 8267
rect 17 8233 25 8267
rect -25 8225 25 8233
rect 19225 8267 19275 8275
rect 19225 8233 19233 8267
rect 19267 8233 19275 8267
rect 19225 8225 19275 8233
rect 19775 8267 19825 8275
rect 19775 8233 19783 8267
rect 19817 8233 19825 8267
rect 19775 8225 19825 8233
rect 54 8202 62 8219
rect 488 8202 496 8219
rect 19304 8202 19312 8219
rect 19738 8202 19746 8219
rect 48 8140 500 8202
rect 48 7810 110 8140
rect 440 7810 500 8140
rect 48 7748 500 7810
rect 19200 8196 19202 8202
rect 19304 8196 19339 8202
rect 19200 8188 19219 8196
rect 19200 7762 19202 8188
rect 19200 7754 19219 7762
rect 19281 8188 19339 8196
rect 19298 8161 19339 8188
rect 19298 7762 19339 7789
rect 19281 7754 19339 7762
rect 19200 7748 19202 7754
rect 19304 7748 19339 7754
rect 54 7731 62 7748
rect 488 7731 496 7748
rect 19304 7731 19312 7748
rect 19738 7731 19746 7748
rect -25 7717 25 7725
rect -25 7683 -17 7717
rect 17 7683 25 7717
rect -25 7675 25 7683
rect 19225 7717 19275 7725
rect 19225 7683 19233 7717
rect 19267 7683 19275 7717
rect 19225 7675 19275 7683
rect 19775 7717 19825 7725
rect 19775 7683 19783 7717
rect 19817 7683 19825 7717
rect 19775 7675 19825 7683
rect 54 7652 62 7669
rect 488 7652 496 7669
rect 19304 7652 19312 7669
rect 19738 7652 19746 7669
rect 461 7646 496 7652
rect 19298 7646 19752 7652
rect 461 7611 500 7646
rect 19200 7638 19219 7646
rect 19200 7611 19202 7638
rect 461 7204 500 7239
rect 19200 7212 19202 7239
rect 19200 7204 19219 7212
rect 19281 7638 19752 7646
rect 19298 7590 19752 7638
rect 19298 7260 19360 7590
rect 19690 7260 19752 7590
rect 19298 7212 19752 7260
rect 19281 7204 19752 7212
rect 461 7198 496 7204
rect 19298 7198 19752 7204
rect 54 7181 62 7198
rect 488 7181 496 7198
rect 19304 7181 19312 7198
rect 19738 7181 19746 7198
rect -25 7167 25 7175
rect -25 7133 -17 7167
rect 17 7133 25 7167
rect -25 7125 25 7133
rect 19225 7167 19275 7175
rect 19225 7133 19233 7167
rect 19267 7133 19275 7167
rect 19225 7125 19275 7133
rect 19775 7167 19825 7175
rect 19775 7133 19783 7167
rect 19817 7133 19825 7167
rect 19775 7125 19825 7133
rect 54 7102 62 7119
rect 488 7102 496 7119
rect 19304 7102 19312 7119
rect 19738 7102 19746 7119
rect 48 7040 500 7102
rect 48 6710 110 7040
rect 440 6710 500 7040
rect 48 6648 500 6710
rect 19200 7096 19202 7102
rect 19304 7096 19339 7102
rect 19200 7088 19219 7096
rect 19200 6662 19202 7088
rect 19200 6654 19219 6662
rect 19281 7088 19339 7096
rect 19298 7061 19339 7088
rect 19298 6662 19339 6689
rect 19281 6654 19339 6662
rect 19200 6648 19202 6654
rect 19304 6648 19339 6654
rect 54 6631 62 6648
rect 488 6631 496 6648
rect 19304 6631 19312 6648
rect 19738 6631 19746 6648
rect -25 6617 25 6625
rect -25 6583 -17 6617
rect 17 6583 25 6617
rect -25 6575 25 6583
rect 19225 6617 19275 6625
rect 19225 6583 19233 6617
rect 19267 6583 19275 6617
rect 19225 6575 19275 6583
rect 19775 6617 19825 6625
rect 19775 6583 19783 6617
rect 19817 6583 19825 6617
rect 19775 6575 19825 6583
rect 54 6552 62 6569
rect 488 6552 496 6569
rect 19304 6552 19312 6569
rect 19738 6552 19746 6569
rect 461 6546 496 6552
rect 19298 6546 19752 6552
rect 461 6511 500 6546
rect 19200 6538 19219 6546
rect 19200 6511 19202 6538
rect 461 6104 500 6139
rect 19200 6112 19202 6139
rect 19200 6104 19219 6112
rect 19281 6538 19752 6546
rect 19298 6490 19752 6538
rect 19298 6160 19360 6490
rect 19690 6160 19752 6490
rect 19298 6112 19752 6160
rect 19281 6104 19752 6112
rect 461 6098 496 6104
rect 19298 6098 19752 6104
rect 54 6081 62 6098
rect 488 6081 496 6098
rect 19304 6081 19312 6098
rect 19738 6081 19746 6098
rect -25 6067 25 6075
rect -25 6033 -17 6067
rect 17 6033 25 6067
rect -25 6025 25 6033
rect 19225 6067 19275 6075
rect 19225 6033 19233 6067
rect 19267 6033 19275 6067
rect 19225 6025 19275 6033
rect 19775 6067 19825 6075
rect 19775 6033 19783 6067
rect 19817 6033 19825 6067
rect 19775 6025 19825 6033
rect 54 6002 62 6019
rect 488 6002 496 6019
rect 19304 6002 19312 6019
rect 19738 6002 19746 6019
rect 48 5940 500 6002
rect 48 5610 110 5940
rect 440 5610 500 5940
rect 48 5548 500 5610
rect 19200 5996 19202 6002
rect 19304 5996 19339 6002
rect 19200 5988 19219 5996
rect 19200 5562 19202 5988
rect 19200 5554 19219 5562
rect 19281 5988 19339 5996
rect 19298 5961 19339 5988
rect 19298 5562 19339 5589
rect 19281 5554 19339 5562
rect 19200 5548 19202 5554
rect 19304 5548 19339 5554
rect 54 5531 62 5548
rect 488 5531 496 5548
rect 19304 5531 19312 5548
rect 19738 5531 19746 5548
rect -25 5517 25 5525
rect -25 5483 -17 5517
rect 17 5483 25 5517
rect -25 5475 25 5483
rect 19225 5517 19275 5525
rect 19225 5483 19233 5517
rect 19267 5483 19275 5517
rect 19225 5475 19275 5483
rect 19775 5517 19825 5525
rect 19775 5483 19783 5517
rect 19817 5483 19825 5517
rect 19775 5475 19825 5483
rect 54 5452 62 5469
rect 488 5452 496 5469
rect 19304 5452 19312 5469
rect 19738 5452 19746 5469
rect 461 5446 496 5452
rect 19298 5446 19752 5452
rect 461 5411 500 5446
rect 19200 5438 19219 5446
rect 19200 5411 19202 5438
rect 461 5004 500 5039
rect 19200 5012 19202 5039
rect 19200 5004 19219 5012
rect 19281 5438 19752 5446
rect 19298 5390 19752 5438
rect 19298 5060 19360 5390
rect 19690 5060 19752 5390
rect 19298 5012 19752 5060
rect 19281 5004 19752 5012
rect 461 4998 496 5004
rect 19298 4998 19752 5004
rect 54 4981 62 4998
rect 488 4981 496 4998
rect 19304 4981 19312 4998
rect 19738 4981 19746 4998
rect -25 4967 25 4975
rect -25 4933 -17 4967
rect 17 4933 25 4967
rect -25 4925 25 4933
rect 19225 4967 19275 4975
rect 19225 4933 19233 4967
rect 19267 4933 19275 4967
rect 19225 4925 19275 4933
rect 19775 4967 19825 4975
rect 19775 4933 19783 4967
rect 19817 4933 19825 4967
rect 19775 4925 19825 4933
rect 54 4902 62 4919
rect 488 4902 496 4919
rect 19304 4902 19312 4919
rect 19738 4902 19746 4919
rect 48 4840 500 4902
rect 48 4510 110 4840
rect 440 4510 500 4840
rect 48 4448 500 4510
rect 19200 4896 19202 4902
rect 19304 4896 19339 4902
rect 19200 4888 19219 4896
rect 19200 4462 19202 4888
rect 19200 4454 19219 4462
rect 19281 4888 19339 4896
rect 19298 4861 19339 4888
rect 19298 4462 19339 4489
rect 19281 4454 19339 4462
rect 19200 4448 19202 4454
rect 19304 4448 19339 4454
rect 54 4431 62 4448
rect 488 4431 496 4448
rect 19304 4431 19312 4448
rect 19738 4431 19746 4448
rect -25 4417 25 4425
rect -25 4383 -17 4417
rect 17 4383 25 4417
rect -25 4375 25 4383
rect 19225 4417 19275 4425
rect 19225 4383 19233 4417
rect 19267 4383 19275 4417
rect 19225 4375 19275 4383
rect 19775 4417 19825 4425
rect 19775 4383 19783 4417
rect 19817 4383 19825 4417
rect 19775 4375 19825 4383
rect 54 4352 62 4369
rect 488 4352 496 4369
rect 19304 4352 19312 4369
rect 19738 4352 19746 4369
rect 461 4346 496 4352
rect 19298 4346 19752 4352
rect 461 4311 500 4346
rect 19200 4338 19219 4346
rect 19200 4311 19202 4338
rect 461 3904 500 3939
rect 19200 3912 19202 3939
rect 19200 3904 19219 3912
rect 19281 4338 19752 4346
rect 19298 4290 19752 4338
rect 19298 3960 19360 4290
rect 19690 3960 19752 4290
rect 19298 3912 19752 3960
rect 19281 3904 19752 3912
rect 461 3898 496 3904
rect 19298 3898 19752 3904
rect 54 3881 62 3898
rect 488 3881 496 3898
rect 19304 3881 19312 3898
rect 19738 3881 19746 3898
rect -25 3867 25 3875
rect -25 3833 -17 3867
rect 17 3833 25 3867
rect -25 3825 25 3833
rect 19225 3867 19275 3875
rect 19225 3833 19233 3867
rect 19267 3833 19275 3867
rect 19225 3825 19275 3833
rect 19775 3867 19825 3875
rect 19775 3833 19783 3867
rect 19817 3833 19825 3867
rect 19775 3825 19825 3833
rect 54 3802 62 3819
rect 488 3802 496 3819
rect 19304 3802 19312 3819
rect 19738 3802 19746 3819
rect 48 3740 500 3802
rect 48 3410 110 3740
rect 440 3410 500 3740
rect 48 3348 500 3410
rect 19200 3796 19202 3802
rect 19304 3796 19339 3802
rect 19200 3788 19219 3796
rect 19200 3362 19202 3788
rect 19200 3354 19219 3362
rect 19281 3788 19339 3796
rect 19298 3761 19339 3788
rect 19298 3362 19339 3389
rect 19281 3354 19339 3362
rect 19200 3348 19202 3354
rect 19304 3348 19339 3354
rect 54 3331 62 3348
rect 488 3331 496 3348
rect 19304 3331 19312 3348
rect 19738 3331 19746 3348
rect -25 3317 25 3325
rect -25 3283 -17 3317
rect 17 3283 25 3317
rect -25 3275 25 3283
rect 19225 3317 19275 3325
rect 19225 3283 19233 3317
rect 19267 3283 19275 3317
rect 19225 3275 19275 3283
rect 19775 3317 19825 3325
rect 19775 3283 19783 3317
rect 19817 3283 19825 3317
rect 19775 3275 19825 3283
rect 54 3252 62 3269
rect 488 3252 496 3269
rect 19304 3252 19312 3269
rect 19738 3252 19746 3269
rect 461 3246 496 3252
rect 19298 3246 19752 3252
rect 461 3211 500 3246
rect 19200 3238 19219 3246
rect 19200 3211 19202 3238
rect 461 2804 500 2839
rect 19200 2812 19202 2839
rect 19200 2804 19219 2812
rect 19281 3238 19752 3246
rect 19298 3190 19752 3238
rect 19298 2860 19360 3190
rect 19690 2860 19752 3190
rect 19298 2812 19752 2860
rect 19281 2804 19752 2812
rect 461 2798 496 2804
rect 19298 2798 19752 2804
rect 54 2781 62 2798
rect 488 2781 496 2798
rect 19304 2781 19312 2798
rect 19738 2781 19746 2798
rect -25 2767 25 2775
rect -25 2733 -17 2767
rect 17 2733 25 2767
rect -25 2725 25 2733
rect 19225 2767 19275 2775
rect 19225 2733 19233 2767
rect 19267 2733 19275 2767
rect 19225 2725 19275 2733
rect 19775 2767 19825 2775
rect 19775 2733 19783 2767
rect 19817 2733 19825 2767
rect 19775 2725 19825 2733
rect 54 2702 62 2719
rect 488 2702 496 2719
rect 19304 2702 19312 2719
rect 19738 2702 19746 2719
rect 48 2640 500 2702
rect 48 2310 110 2640
rect 440 2310 500 2640
rect 48 2248 500 2310
rect 19200 2696 19202 2702
rect 19304 2696 19339 2702
rect 19200 2688 19219 2696
rect 19200 2262 19202 2688
rect 19200 2254 19219 2262
rect 19281 2688 19339 2696
rect 19298 2661 19339 2688
rect 19298 2262 19339 2289
rect 19281 2254 19339 2262
rect 19200 2248 19202 2254
rect 19304 2248 19339 2254
rect 54 2231 62 2248
rect 488 2231 496 2248
rect 19304 2231 19312 2248
rect 19738 2231 19746 2248
rect -25 2217 25 2225
rect -25 2183 -17 2217
rect 17 2183 25 2217
rect -25 2175 25 2183
rect 19225 2217 19275 2225
rect 19225 2183 19233 2217
rect 19267 2183 19275 2217
rect 19225 2175 19275 2183
rect 19775 2217 19825 2225
rect 19775 2183 19783 2217
rect 19817 2183 19825 2217
rect 19775 2175 19825 2183
rect 54 2152 62 2169
rect 488 2152 496 2169
rect 19304 2152 19312 2169
rect 19738 2152 19746 2169
rect 461 2146 496 2152
rect 19298 2146 19752 2152
rect 461 2111 500 2146
rect 19200 2138 19219 2146
rect 19200 2111 19202 2138
rect 461 1704 500 1739
rect 19200 1712 19202 1739
rect 19200 1704 19219 1712
rect 19281 2138 19752 2146
rect 19298 2090 19752 2138
rect 19298 1760 19360 2090
rect 19690 1760 19752 2090
rect 19298 1712 19752 1760
rect 19281 1704 19752 1712
rect 461 1698 496 1704
rect 19298 1698 19752 1704
rect 54 1681 62 1698
rect 488 1681 496 1698
rect 19304 1681 19312 1698
rect 19738 1681 19746 1698
rect -25 1667 25 1675
rect -25 1633 -17 1667
rect 17 1633 25 1667
rect -25 1625 25 1633
rect 19225 1667 19275 1675
rect 19225 1633 19233 1667
rect 19267 1633 19275 1667
rect 19225 1625 19275 1633
rect 19775 1667 19825 1675
rect 19775 1633 19783 1667
rect 19817 1633 19825 1667
rect 19775 1625 19825 1633
rect 54 1602 62 1619
rect 488 1602 496 1619
rect 19304 1602 19312 1619
rect 19738 1602 19746 1619
rect 48 1540 500 1602
rect 48 1210 110 1540
rect 440 1210 500 1540
rect 48 1148 500 1210
rect 19200 1596 19202 1602
rect 19304 1596 19339 1602
rect 19200 1588 19219 1596
rect 19200 1162 19202 1588
rect 19200 1154 19219 1162
rect 19281 1588 19339 1596
rect 19298 1561 19339 1588
rect 19298 1162 19339 1189
rect 19281 1154 19339 1162
rect 19200 1148 19202 1154
rect 19304 1148 19339 1154
rect 54 1131 62 1148
rect 488 1131 496 1148
rect 19304 1131 19312 1148
rect 19738 1131 19746 1148
rect -25 1117 25 1125
rect -25 1083 -17 1117
rect 17 1083 25 1117
rect -25 1075 25 1083
rect 19225 1117 19275 1125
rect 19225 1083 19233 1117
rect 19267 1083 19275 1117
rect 19225 1075 19275 1083
rect 19775 1117 19825 1125
rect 19775 1083 19783 1117
rect 19817 1083 19825 1117
rect 19775 1075 19825 1083
rect 54 1052 62 1069
rect 488 1052 496 1069
rect 19304 1052 19312 1069
rect 19738 1052 19746 1069
rect 461 1046 496 1052
rect 19298 1046 19752 1052
rect 461 1011 500 1046
rect 19200 1038 19219 1046
rect 19200 1011 19202 1038
rect 461 604 500 639
rect 19200 612 19202 639
rect 19200 604 19219 612
rect 19281 1038 19752 1046
rect 19298 990 19752 1038
rect 19298 660 19360 990
rect 19690 660 19752 990
rect 19298 612 19752 660
rect 19281 604 19752 612
rect 461 598 496 604
rect 19298 598 19752 604
rect 54 581 62 598
rect 488 581 496 598
rect 19304 581 19312 598
rect 19738 581 19746 598
rect -25 567 25 575
rect -25 533 -17 567
rect 17 533 25 567
rect -25 525 25 533
rect 19225 567 19275 575
rect 19225 533 19233 567
rect 19267 533 19275 567
rect 19225 525 19275 533
rect 19775 567 19825 575
rect 19775 533 19783 567
rect 19817 533 19825 567
rect 19775 525 19825 533
rect 54 502 62 519
rect 488 502 496 519
rect 19304 502 19312 519
rect 19738 502 19746 519
rect 48 500 500 502
rect 19200 500 19202 502
rect 48 496 502 500
rect 604 496 639 500
rect 48 488 519 496
rect 48 440 502 488
rect 48 110 110 440
rect 440 110 502 440
rect 48 62 502 110
rect 48 54 519 62
rect 581 488 639 496
rect 598 461 639 488
rect 1011 496 1046 500
rect 1148 496 1602 500
rect 1704 496 1739 500
rect 1011 488 1069 496
rect 1011 461 1052 488
rect 581 54 598 62
rect 1052 54 1069 62
rect 1131 488 1619 496
rect 1148 440 1602 488
rect 1148 110 1210 440
rect 1540 110 1602 440
rect 1148 62 1602 110
rect 1131 54 1619 62
rect 1681 488 1739 496
rect 1698 461 1739 488
rect 2111 496 2146 500
rect 2248 496 2702 500
rect 2804 496 2839 500
rect 2111 488 2169 496
rect 2111 461 2152 488
rect 1681 54 1698 62
rect 2152 54 2169 62
rect 2231 488 2719 496
rect 2248 440 2702 488
rect 2248 110 2310 440
rect 2640 110 2702 440
rect 2248 62 2702 110
rect 2231 54 2719 62
rect 2781 488 2839 496
rect 2798 461 2839 488
rect 3211 496 3246 500
rect 3348 496 3802 500
rect 3904 496 3939 500
rect 3211 488 3269 496
rect 3211 461 3252 488
rect 2781 54 2798 62
rect 3252 54 3269 62
rect 3331 488 3819 496
rect 3348 440 3802 488
rect 3348 110 3410 440
rect 3740 110 3802 440
rect 3348 62 3802 110
rect 3331 54 3819 62
rect 3881 488 3939 496
rect 3898 461 3939 488
rect 4311 496 4346 500
rect 4448 496 4902 500
rect 5004 496 5039 500
rect 4311 488 4369 496
rect 4311 461 4352 488
rect 3881 54 3898 62
rect 4352 54 4369 62
rect 4431 488 4919 496
rect 4448 440 4902 488
rect 4448 110 4510 440
rect 4840 110 4902 440
rect 4448 62 4902 110
rect 4431 54 4919 62
rect 4981 488 5039 496
rect 4998 461 5039 488
rect 5411 496 5446 500
rect 5548 496 6002 500
rect 6104 496 6139 500
rect 5411 488 5469 496
rect 5411 461 5452 488
rect 4981 54 4998 62
rect 5452 54 5469 62
rect 5531 488 6019 496
rect 5548 440 6002 488
rect 5548 110 5610 440
rect 5940 110 6002 440
rect 5548 62 6002 110
rect 5531 54 6019 62
rect 6081 488 6139 496
rect 6098 461 6139 488
rect 6511 496 6546 500
rect 6648 496 7102 500
rect 7204 496 7239 500
rect 6511 488 6569 496
rect 6511 461 6552 488
rect 6081 54 6098 62
rect 6552 54 6569 62
rect 6631 488 7119 496
rect 6648 440 7102 488
rect 6648 110 6710 440
rect 7040 110 7102 440
rect 6648 62 7102 110
rect 6631 54 7119 62
rect 7181 488 7239 496
rect 7198 461 7239 488
rect 7611 496 7646 500
rect 7748 496 8202 500
rect 8304 496 8339 500
rect 7611 488 7669 496
rect 7611 461 7652 488
rect 7181 54 7198 62
rect 7652 54 7669 62
rect 7731 488 8219 496
rect 7748 440 8202 488
rect 7748 110 7810 440
rect 8140 110 8202 440
rect 7748 62 8202 110
rect 7731 54 8219 62
rect 8281 488 8339 496
rect 8298 461 8339 488
rect 8711 496 8746 500
rect 8848 496 9302 500
rect 9404 496 9439 500
rect 8711 488 8769 496
rect 8711 461 8752 488
rect 8281 54 8298 62
rect 8752 54 8769 62
rect 8831 488 9319 496
rect 8848 440 9302 488
rect 8848 110 8910 440
rect 9240 110 9302 440
rect 8848 62 9302 110
rect 8831 54 9319 62
rect 9381 488 9439 496
rect 9398 461 9439 488
rect 9811 496 9846 500
rect 9948 496 10402 500
rect 10504 496 10539 500
rect 9811 488 9869 496
rect 9811 461 9852 488
rect 9381 54 9398 62
rect 9852 54 9869 62
rect 9931 488 10419 496
rect 9948 440 10402 488
rect 9948 110 10010 440
rect 10340 110 10402 440
rect 9948 62 10402 110
rect 9931 54 10419 62
rect 10481 488 10539 496
rect 10498 461 10539 488
rect 10911 496 10946 500
rect 11048 496 11502 500
rect 11604 496 11639 500
rect 10911 488 10969 496
rect 10911 461 10952 488
rect 10481 54 10498 62
rect 10952 54 10969 62
rect 11031 488 11519 496
rect 11048 440 11502 488
rect 11048 110 11110 440
rect 11440 110 11502 440
rect 11048 62 11502 110
rect 11031 54 11519 62
rect 11581 488 11639 496
rect 11598 461 11639 488
rect 12011 496 12046 500
rect 12148 496 12602 500
rect 12704 496 12739 500
rect 12011 488 12069 496
rect 12011 461 12052 488
rect 11581 54 11598 62
rect 12052 54 12069 62
rect 12131 488 12619 496
rect 12148 440 12602 488
rect 12148 110 12210 440
rect 12540 110 12602 440
rect 12148 62 12602 110
rect 12131 54 12619 62
rect 12681 488 12739 496
rect 12698 461 12739 488
rect 13111 496 13146 500
rect 13248 496 13702 500
rect 13804 496 13839 500
rect 13111 488 13169 496
rect 13111 461 13152 488
rect 12681 54 12698 62
rect 13152 54 13169 62
rect 13231 488 13719 496
rect 13248 440 13702 488
rect 13248 110 13310 440
rect 13640 110 13702 440
rect 13248 62 13702 110
rect 13231 54 13719 62
rect 13781 488 13839 496
rect 13798 461 13839 488
rect 14211 496 14246 500
rect 14348 496 14802 500
rect 14904 496 14939 500
rect 14211 488 14269 496
rect 14211 461 14252 488
rect 13781 54 13798 62
rect 14252 54 14269 62
rect 14331 488 14819 496
rect 14348 440 14802 488
rect 14348 110 14410 440
rect 14740 110 14802 440
rect 14348 62 14802 110
rect 14331 54 14819 62
rect 14881 488 14939 496
rect 14898 461 14939 488
rect 15311 496 15346 500
rect 15448 496 15902 500
rect 16004 496 16039 500
rect 15311 488 15369 496
rect 15311 461 15352 488
rect 14881 54 14898 62
rect 15352 54 15369 62
rect 15431 488 15919 496
rect 15448 440 15902 488
rect 15448 110 15510 440
rect 15840 110 15902 440
rect 15448 62 15902 110
rect 15431 54 15919 62
rect 15981 488 16039 496
rect 15998 461 16039 488
rect 16411 496 16446 500
rect 16548 496 17002 500
rect 17104 496 17139 500
rect 16411 488 16469 496
rect 16411 461 16452 488
rect 15981 54 15998 62
rect 16452 54 16469 62
rect 16531 488 17019 496
rect 16548 440 17002 488
rect 16548 110 16610 440
rect 16940 110 17002 440
rect 16548 62 17002 110
rect 16531 54 17019 62
rect 17081 488 17139 496
rect 17098 461 17139 488
rect 17511 496 17546 500
rect 17648 496 18102 500
rect 18204 496 18239 500
rect 17511 488 17569 496
rect 17511 461 17552 488
rect 17081 54 17098 62
rect 17552 54 17569 62
rect 17631 488 18119 496
rect 17648 440 18102 488
rect 17648 110 17710 440
rect 18040 110 18102 440
rect 17648 62 18102 110
rect 17631 54 18119 62
rect 18181 488 18239 496
rect 18198 461 18239 488
rect 18611 496 18646 500
rect 18748 496 19202 500
rect 19304 496 19339 502
rect 18611 488 18669 496
rect 18611 461 18652 488
rect 18181 54 18198 62
rect 18652 54 18669 62
rect 18731 488 19219 496
rect 18748 440 19202 488
rect 18748 110 18810 440
rect 19140 110 19202 440
rect 18748 62 19202 110
rect 18731 54 19219 62
rect 19281 488 19339 496
rect 19298 461 19339 488
rect 19281 54 19298 62
rect 48 48 502 54
rect 1148 48 1602 54
rect 2248 48 2702 54
rect 3348 48 3802 54
rect 4448 48 4902 54
rect 5548 48 6002 54
rect 6648 48 7102 54
rect 7748 48 8202 54
rect 8848 48 9302 54
rect 9948 48 10402 54
rect 11048 48 11502 54
rect 12148 48 12602 54
rect 13248 48 13702 54
rect 14348 48 14802 54
rect 15448 48 15902 54
rect 16548 48 17002 54
rect 17648 48 18102 54
rect 18748 48 19202 54
rect -25 17 25 25
rect -25 -17 -17 17
rect 17 -17 25 17
rect -25 -25 25 -17
rect 525 17 575 25
rect 525 -17 533 17
rect 567 -17 575 17
rect 525 -25 575 -17
rect 1075 17 1125 25
rect 1075 -17 1083 17
rect 1117 -17 1125 17
rect 1075 -25 1125 -17
rect 1625 17 1675 25
rect 1625 -17 1633 17
rect 1667 -17 1675 17
rect 1625 -25 1675 -17
rect 2175 17 2225 25
rect 2175 -17 2183 17
rect 2217 -17 2225 17
rect 2175 -25 2225 -17
rect 2725 17 2775 25
rect 2725 -17 2733 17
rect 2767 -17 2775 17
rect 2725 -25 2775 -17
rect 3275 17 3325 25
rect 3275 -17 3283 17
rect 3317 -17 3325 17
rect 3275 -25 3325 -17
rect 3825 17 3875 25
rect 3825 -17 3833 17
rect 3867 -17 3875 17
rect 3825 -25 3875 -17
rect 4375 17 4425 25
rect 4375 -17 4383 17
rect 4417 -17 4425 17
rect 4375 -25 4425 -17
rect 4925 17 4975 25
rect 4925 -17 4933 17
rect 4967 -17 4975 17
rect 4925 -25 4975 -17
rect 5475 17 5525 25
rect 5475 -17 5483 17
rect 5517 -17 5525 17
rect 5475 -25 5525 -17
rect 6025 17 6075 25
rect 6025 -17 6033 17
rect 6067 -17 6075 17
rect 6025 -25 6075 -17
rect 6575 17 6625 25
rect 6575 -17 6583 17
rect 6617 -17 6625 17
rect 6575 -25 6625 -17
rect 7125 17 7175 25
rect 7125 -17 7133 17
rect 7167 -17 7175 17
rect 7125 -25 7175 -17
rect 7675 17 7725 25
rect 7675 -17 7683 17
rect 7717 -17 7725 17
rect 7675 -25 7725 -17
rect 8225 17 8275 25
rect 8225 -17 8233 17
rect 8267 -17 8275 17
rect 8225 -25 8275 -17
rect 8775 17 8825 25
rect 8775 -17 8783 17
rect 8817 -17 8825 17
rect 8775 -25 8825 -17
rect 9325 17 9375 25
rect 9325 -17 9333 17
rect 9367 -17 9375 17
rect 9325 -25 9375 -17
rect 9875 17 9925 25
rect 9875 -17 9883 17
rect 9917 -17 9925 17
rect 9875 -25 9925 -17
rect 10425 17 10475 25
rect 10425 -17 10433 17
rect 10467 -17 10475 17
rect 10425 -25 10475 -17
rect 10975 17 11025 25
rect 10975 -17 10983 17
rect 11017 -17 11025 17
rect 10975 -25 11025 -17
rect 11525 17 11575 25
rect 11525 -17 11533 17
rect 11567 -17 11575 17
rect 11525 -25 11575 -17
rect 12075 17 12125 25
rect 12075 -17 12083 17
rect 12117 -17 12125 17
rect 12075 -25 12125 -17
rect 12625 17 12675 25
rect 12625 -17 12633 17
rect 12667 -17 12675 17
rect 12625 -25 12675 -17
rect 13175 17 13225 25
rect 13175 -17 13183 17
rect 13217 -17 13225 17
rect 13175 -25 13225 -17
rect 13725 17 13775 25
rect 13725 -17 13733 17
rect 13767 -17 13775 17
rect 13725 -25 13775 -17
rect 14275 17 14325 25
rect 14275 -17 14283 17
rect 14317 -17 14325 17
rect 14275 -25 14325 -17
rect 14825 17 14875 25
rect 14825 -17 14833 17
rect 14867 -17 14875 17
rect 14825 -25 14875 -17
rect 15375 17 15425 25
rect 15375 -17 15383 17
rect 15417 -17 15425 17
rect 15375 -25 15425 -17
rect 15925 17 15975 25
rect 15925 -17 15933 17
rect 15967 -17 15975 17
rect 15925 -25 15975 -17
rect 16475 17 16525 25
rect 16475 -17 16483 17
rect 16517 -17 16525 17
rect 16475 -25 16525 -17
rect 17025 17 17075 25
rect 17025 -17 17033 17
rect 17067 -17 17075 17
rect 17025 -25 17075 -17
rect 17575 17 17625 25
rect 17575 -17 17583 17
rect 17617 -17 17625 17
rect 17575 -25 17625 -17
rect 18125 17 18175 25
rect 18125 -17 18133 17
rect 18167 -17 18175 17
rect 18125 -25 18175 -17
rect 18675 17 18725 25
rect 18675 -17 18683 17
rect 18717 -17 18725 17
rect 18675 -25 18725 -17
rect 19225 17 19275 25
rect 19225 -17 19233 17
rect 19267 -17 19275 17
rect 19225 -25 19275 -17
rect 19775 17 19825 25
rect 19775 -17 19783 17
rect 19817 -17 19825 17
rect 19775 -25 19825 -17
rect 20000 -200 20012 20000
rect -212 -212 20012 -200
rect 20288 -488 20300 20288
rect -500 -500 20300 -488
rect 20800 -1000 20812 20800
rect -1012 -1012 20812 -1000
rect 24788 -4988 24800 24788
rect -5000 -5000 24800 -4988
<< viali >>
rect -4988 20812 24788 24788
rect -4988 -1012 -1012 20812
rect -488 20012 20288 20288
rect -488 -212 -212 20012
rect -17 19783 17 19817
rect 533 19783 567 19817
rect 1083 19783 1117 19817
rect 1633 19783 1667 19817
rect 2183 19783 2217 19817
rect 2733 19783 2767 19817
rect 3283 19783 3317 19817
rect 3833 19783 3867 19817
rect 4383 19783 4417 19817
rect 4933 19783 4967 19817
rect 5483 19783 5517 19817
rect 6033 19783 6067 19817
rect 6583 19783 6617 19817
rect 7133 19783 7167 19817
rect 7683 19783 7717 19817
rect 8233 19783 8267 19817
rect 8783 19783 8817 19817
rect 9333 19783 9367 19817
rect 9883 19783 9917 19817
rect 10433 19783 10467 19817
rect 10983 19783 11017 19817
rect 11533 19783 11567 19817
rect 12083 19783 12117 19817
rect 12633 19783 12667 19817
rect 13183 19783 13217 19817
rect 13733 19783 13767 19817
rect 14283 19783 14317 19817
rect 14833 19783 14867 19817
rect 15383 19783 15417 19817
rect 15933 19783 15967 19817
rect 16483 19783 16517 19817
rect 17033 19783 17067 19817
rect 17583 19783 17617 19817
rect 18133 19783 18167 19817
rect 18683 19783 18717 19817
rect 19233 19783 19267 19817
rect 19783 19783 19817 19817
rect 502 19312 519 19738
rect 581 19312 598 19738
rect 660 19678 990 19690
rect 660 19372 672 19678
rect 672 19372 978 19678
rect 978 19372 990 19678
rect 660 19360 990 19372
rect 1052 19312 1069 19738
rect 1131 19312 1148 19738
rect 1602 19312 1619 19738
rect 1681 19312 1698 19738
rect 1760 19678 2090 19690
rect 1760 19372 1772 19678
rect 1772 19372 2078 19678
rect 2078 19372 2090 19678
rect 1760 19360 2090 19372
rect 2152 19312 2169 19738
rect 2231 19312 2248 19738
rect 2702 19312 2719 19738
rect 2781 19312 2798 19738
rect 2860 19678 3190 19690
rect 2860 19372 2872 19678
rect 2872 19372 3178 19678
rect 3178 19372 3190 19678
rect 2860 19360 3190 19372
rect 3252 19312 3269 19738
rect 3331 19312 3348 19738
rect 3802 19312 3819 19738
rect 3881 19312 3898 19738
rect 3960 19678 4290 19690
rect 3960 19372 3972 19678
rect 3972 19372 4278 19678
rect 4278 19372 4290 19678
rect 3960 19360 4290 19372
rect 4352 19312 4369 19738
rect 4431 19312 4448 19738
rect 4902 19312 4919 19738
rect 4981 19312 4998 19738
rect 5060 19678 5390 19690
rect 5060 19372 5072 19678
rect 5072 19372 5378 19678
rect 5378 19372 5390 19678
rect 5060 19360 5390 19372
rect 5452 19312 5469 19738
rect 5531 19312 5548 19738
rect 6002 19312 6019 19738
rect 6081 19312 6098 19738
rect 6160 19678 6490 19690
rect 6160 19372 6172 19678
rect 6172 19372 6478 19678
rect 6478 19372 6490 19678
rect 6160 19360 6490 19372
rect 6552 19312 6569 19738
rect 6631 19312 6648 19738
rect 7102 19312 7119 19738
rect 7181 19312 7198 19738
rect 7260 19678 7590 19690
rect 7260 19372 7272 19678
rect 7272 19372 7578 19678
rect 7578 19372 7590 19678
rect 7260 19360 7590 19372
rect 7652 19312 7669 19738
rect 7731 19312 7748 19738
rect 8202 19312 8219 19738
rect 8281 19312 8298 19738
rect 8360 19678 8690 19690
rect 8360 19372 8372 19678
rect 8372 19372 8678 19678
rect 8678 19372 8690 19678
rect 8360 19360 8690 19372
rect 8752 19312 8769 19738
rect 8831 19312 8848 19738
rect 9302 19312 9319 19738
rect 9381 19312 9398 19738
rect 9460 19678 9790 19690
rect 9460 19372 9472 19678
rect 9472 19372 9778 19678
rect 9778 19372 9790 19678
rect 9460 19360 9790 19372
rect 9852 19312 9869 19738
rect 9931 19312 9948 19738
rect 10402 19312 10419 19738
rect 10481 19312 10498 19738
rect 10560 19678 10890 19690
rect 10560 19372 10572 19678
rect 10572 19372 10878 19678
rect 10878 19372 10890 19678
rect 10560 19360 10890 19372
rect 10952 19312 10969 19738
rect 11031 19312 11048 19738
rect 11502 19312 11519 19738
rect 11581 19312 11598 19738
rect 11660 19678 11990 19690
rect 11660 19372 11672 19678
rect 11672 19372 11978 19678
rect 11978 19372 11990 19678
rect 11660 19360 11990 19372
rect 12052 19312 12069 19738
rect 12131 19312 12148 19738
rect 12602 19312 12619 19738
rect 12681 19312 12698 19738
rect 12760 19678 13090 19690
rect 12760 19372 12772 19678
rect 12772 19372 13078 19678
rect 13078 19372 13090 19678
rect 12760 19360 13090 19372
rect 13152 19312 13169 19738
rect 13231 19312 13248 19738
rect 13702 19312 13719 19738
rect 13781 19312 13798 19738
rect 13860 19678 14190 19690
rect 13860 19372 13872 19678
rect 13872 19372 14178 19678
rect 14178 19372 14190 19678
rect 13860 19360 14190 19372
rect 14252 19312 14269 19738
rect 14331 19312 14348 19738
rect 14802 19312 14819 19738
rect 14881 19312 14898 19738
rect 14960 19678 15290 19690
rect 14960 19372 14972 19678
rect 14972 19372 15278 19678
rect 15278 19372 15290 19678
rect 14960 19360 15290 19372
rect 15352 19312 15369 19738
rect 15431 19312 15448 19738
rect 15902 19312 15919 19738
rect 15981 19312 15998 19738
rect 16060 19678 16390 19690
rect 16060 19372 16072 19678
rect 16072 19372 16378 19678
rect 16378 19372 16390 19678
rect 16060 19360 16390 19372
rect 16452 19312 16469 19738
rect 16531 19312 16548 19738
rect 17002 19312 17019 19738
rect 17081 19312 17098 19738
rect 17160 19678 17490 19690
rect 17160 19372 17172 19678
rect 17172 19372 17478 19678
rect 17478 19372 17490 19678
rect 17160 19360 17490 19372
rect 17552 19312 17569 19738
rect 17631 19312 17648 19738
rect 18102 19312 18119 19738
rect 18181 19312 18198 19738
rect 18260 19678 18590 19690
rect 18260 19372 18272 19678
rect 18272 19372 18578 19678
rect 18578 19372 18590 19678
rect 18260 19360 18590 19372
rect 18652 19312 18669 19738
rect 18731 19312 18748 19738
rect 19202 19312 19219 19738
rect 19281 19312 19298 19738
rect 19360 19678 19690 19690
rect 19360 19372 19372 19678
rect 19372 19372 19678 19678
rect 19678 19372 19690 19678
rect 19360 19360 19690 19372
rect 62 19281 488 19298
rect 612 19281 1038 19298
rect 1162 19281 1588 19298
rect 1712 19281 2138 19298
rect 2262 19281 2688 19298
rect 2812 19281 3238 19298
rect 3362 19281 3788 19298
rect 3912 19281 4338 19298
rect 4462 19281 4888 19298
rect 5012 19281 5438 19298
rect 5562 19281 5988 19298
rect 6112 19281 6538 19298
rect 6662 19281 7088 19298
rect 7212 19281 7638 19298
rect 7762 19281 8188 19298
rect 8312 19281 8738 19298
rect 8862 19281 9288 19298
rect 9412 19281 9838 19298
rect 9962 19281 10388 19298
rect 10512 19281 10938 19298
rect 11062 19281 11488 19298
rect 11612 19281 12038 19298
rect 12162 19281 12588 19298
rect 12712 19281 13138 19298
rect 13262 19281 13688 19298
rect 13812 19281 14238 19298
rect 14362 19281 14788 19298
rect 14912 19281 15338 19298
rect 15462 19281 15888 19298
rect 16012 19281 16438 19298
rect 16562 19281 16988 19298
rect 17112 19281 17538 19298
rect 17662 19281 18088 19298
rect 18212 19281 18638 19298
rect 18762 19281 19188 19298
rect 19312 19281 19738 19298
rect -17 19233 17 19267
rect 533 19233 567 19267
rect 1083 19233 1117 19267
rect 1633 19233 1667 19267
rect 2183 19233 2217 19267
rect 2733 19233 2767 19267
rect 3283 19233 3317 19267
rect 3833 19233 3867 19267
rect 4383 19233 4417 19267
rect 4933 19233 4967 19267
rect 5483 19233 5517 19267
rect 6033 19233 6067 19267
rect 6583 19233 6617 19267
rect 7133 19233 7167 19267
rect 7683 19233 7717 19267
rect 8233 19233 8267 19267
rect 8783 19233 8817 19267
rect 9333 19233 9367 19267
rect 9883 19233 9917 19267
rect 10433 19233 10467 19267
rect 10983 19233 11017 19267
rect 11533 19233 11567 19267
rect 12083 19233 12117 19267
rect 12633 19233 12667 19267
rect 13183 19233 13217 19267
rect 13733 19233 13767 19267
rect 14283 19233 14317 19267
rect 14833 19233 14867 19267
rect 15383 19233 15417 19267
rect 15933 19233 15967 19267
rect 16483 19233 16517 19267
rect 17033 19233 17067 19267
rect 17583 19233 17617 19267
rect 18133 19233 18167 19267
rect 18683 19233 18717 19267
rect 19233 19233 19267 19267
rect 19783 19233 19817 19267
rect 62 19202 488 19219
rect 612 19202 1038 19219
rect 1162 19202 1588 19219
rect 1712 19202 2138 19219
rect 2262 19202 2688 19219
rect 2812 19202 3238 19219
rect 3362 19202 3788 19219
rect 3912 19202 4338 19219
rect 4462 19202 4888 19219
rect 5012 19202 5438 19219
rect 5562 19202 5988 19219
rect 6112 19202 6538 19219
rect 6662 19202 7088 19219
rect 7212 19202 7638 19219
rect 7762 19202 8188 19219
rect 8312 19202 8738 19219
rect 8862 19202 9288 19219
rect 9412 19202 9838 19219
rect 9962 19202 10388 19219
rect 10512 19202 10938 19219
rect 11062 19202 11488 19219
rect 11612 19202 12038 19219
rect 12162 19202 12588 19219
rect 12712 19202 13138 19219
rect 13262 19202 13688 19219
rect 13812 19202 14238 19219
rect 14362 19202 14788 19219
rect 14912 19202 15338 19219
rect 15462 19202 15888 19219
rect 16012 19202 16438 19219
rect 16562 19202 16988 19219
rect 17112 19202 17538 19219
rect 17662 19202 18088 19219
rect 18212 19202 18638 19219
rect 18762 19202 19188 19219
rect 19312 19202 19738 19219
rect 110 19128 440 19140
rect 110 18822 122 19128
rect 122 18822 428 19128
rect 428 18822 440 19128
rect 110 18810 440 18822
rect 19202 18762 19219 19188
rect 19281 18762 19298 19188
rect 62 18731 488 18748
rect 19312 18731 19738 18748
rect -17 18683 17 18717
rect 19233 18683 19267 18717
rect 19783 18683 19817 18717
rect 62 18652 488 18669
rect 19312 18652 19738 18669
rect 19202 18212 19219 18638
rect 19281 18212 19298 18638
rect 19360 18578 19690 18590
rect 19360 18272 19372 18578
rect 19372 18272 19678 18578
rect 19678 18272 19690 18578
rect 19360 18260 19690 18272
rect 62 18181 488 18198
rect 19312 18181 19738 18198
rect -17 18133 17 18167
rect 19233 18133 19267 18167
rect 19783 18133 19817 18167
rect 62 18102 488 18119
rect 19312 18102 19738 18119
rect 110 18028 440 18040
rect 110 17722 122 18028
rect 122 17722 428 18028
rect 428 17722 440 18028
rect 110 17710 440 17722
rect 19202 17662 19219 18088
rect 19281 17662 19298 18088
rect 62 17631 488 17648
rect 19312 17631 19738 17648
rect -17 17583 17 17617
rect 19233 17583 19267 17617
rect 19783 17583 19817 17617
rect 62 17552 488 17569
rect 19312 17552 19738 17569
rect 19202 17112 19219 17538
rect 19281 17112 19298 17538
rect 19360 17478 19690 17490
rect 19360 17172 19372 17478
rect 19372 17172 19678 17478
rect 19678 17172 19690 17478
rect 19360 17160 19690 17172
rect 62 17081 488 17098
rect 19312 17081 19738 17098
rect -17 17033 17 17067
rect 19233 17033 19267 17067
rect 19783 17033 19817 17067
rect 62 17002 488 17019
rect 19312 17002 19738 17019
rect 110 16928 440 16940
rect 110 16622 122 16928
rect 122 16622 428 16928
rect 428 16622 440 16928
rect 110 16610 440 16622
rect 19202 16562 19219 16988
rect 19281 16562 19298 16988
rect 62 16531 488 16548
rect 19312 16531 19738 16548
rect -17 16483 17 16517
rect 19233 16483 19267 16517
rect 19783 16483 19817 16517
rect 62 16452 488 16469
rect 19312 16452 19738 16469
rect 19202 16012 19219 16438
rect 19281 16012 19298 16438
rect 19360 16378 19690 16390
rect 19360 16072 19372 16378
rect 19372 16072 19678 16378
rect 19678 16072 19690 16378
rect 19360 16060 19690 16072
rect 62 15981 488 15998
rect 19312 15981 19738 15998
rect -17 15933 17 15967
rect 19233 15933 19267 15967
rect 19783 15933 19817 15967
rect 62 15902 488 15919
rect 19312 15902 19738 15919
rect 110 15828 440 15840
rect 110 15522 122 15828
rect 122 15522 428 15828
rect 428 15522 440 15828
rect 110 15510 440 15522
rect 19202 15462 19219 15888
rect 19281 15462 19298 15888
rect 62 15431 488 15448
rect 19312 15431 19738 15448
rect -17 15383 17 15417
rect 19233 15383 19267 15417
rect 19783 15383 19817 15417
rect 62 15352 488 15369
rect 19312 15352 19738 15369
rect 19202 14912 19219 15338
rect 19281 14912 19298 15338
rect 19360 15278 19690 15290
rect 19360 14972 19372 15278
rect 19372 14972 19678 15278
rect 19678 14972 19690 15278
rect 19360 14960 19690 14972
rect 62 14881 488 14898
rect 19312 14881 19738 14898
rect -17 14833 17 14867
rect 19233 14833 19267 14867
rect 19783 14833 19817 14867
rect 62 14802 488 14819
rect 19312 14802 19738 14819
rect 110 14728 440 14740
rect 110 14422 122 14728
rect 122 14422 428 14728
rect 428 14422 440 14728
rect 110 14410 440 14422
rect 19202 14362 19219 14788
rect 19281 14362 19298 14788
rect 62 14331 488 14348
rect 19312 14331 19738 14348
rect -17 14283 17 14317
rect 19233 14283 19267 14317
rect 19783 14283 19817 14317
rect 62 14252 488 14269
rect 19312 14252 19738 14269
rect 19202 13812 19219 14238
rect 19281 13812 19298 14238
rect 19360 14178 19690 14190
rect 19360 13872 19372 14178
rect 19372 13872 19678 14178
rect 19678 13872 19690 14178
rect 19360 13860 19690 13872
rect 62 13781 488 13798
rect 19312 13781 19738 13798
rect -17 13733 17 13767
rect 19233 13733 19267 13767
rect 19783 13733 19817 13767
rect 62 13702 488 13719
rect 19312 13702 19738 13719
rect 110 13628 440 13640
rect 110 13322 122 13628
rect 122 13322 428 13628
rect 428 13322 440 13628
rect 110 13310 440 13322
rect 19202 13262 19219 13688
rect 19281 13262 19298 13688
rect 62 13231 488 13248
rect 19312 13231 19738 13248
rect -17 13183 17 13217
rect 19233 13183 19267 13217
rect 19783 13183 19817 13217
rect 62 13152 488 13169
rect 19312 13152 19738 13169
rect 19202 12712 19219 13138
rect 19281 12712 19298 13138
rect 19360 13078 19690 13090
rect 19360 12772 19372 13078
rect 19372 12772 19678 13078
rect 19678 12772 19690 13078
rect 19360 12760 19690 12772
rect 62 12681 488 12698
rect 19312 12681 19738 12698
rect -17 12633 17 12667
rect 19233 12633 19267 12667
rect 19783 12633 19817 12667
rect 62 12602 488 12619
rect 19312 12602 19738 12619
rect 110 12528 440 12540
rect 110 12222 122 12528
rect 122 12222 428 12528
rect 428 12222 440 12528
rect 110 12210 440 12222
rect 19202 12162 19219 12588
rect 19281 12162 19298 12588
rect 62 12131 488 12148
rect 19312 12131 19738 12148
rect -17 12083 17 12117
rect 19233 12083 19267 12117
rect 19783 12083 19817 12117
rect 62 12052 488 12069
rect 19312 12052 19738 12069
rect 19202 11612 19219 12038
rect 19281 11612 19298 12038
rect 19360 11978 19690 11990
rect 19360 11672 19372 11978
rect 19372 11672 19678 11978
rect 19678 11672 19690 11978
rect 19360 11660 19690 11672
rect 62 11581 488 11598
rect 19312 11581 19738 11598
rect -17 11533 17 11567
rect 19233 11533 19267 11567
rect 19783 11533 19817 11567
rect 62 11502 488 11519
rect 19312 11502 19738 11519
rect 110 11428 440 11440
rect 110 11122 122 11428
rect 122 11122 428 11428
rect 428 11122 440 11428
rect 110 11110 440 11122
rect 19202 11062 19219 11488
rect 19281 11062 19298 11488
rect 62 11031 488 11048
rect 19312 11031 19738 11048
rect -17 10983 17 11017
rect 19233 10983 19267 11017
rect 19783 10983 19817 11017
rect 62 10952 488 10969
rect 19312 10952 19738 10969
rect 19202 10512 19219 10938
rect 19281 10512 19298 10938
rect 19360 10878 19690 10890
rect 19360 10572 19372 10878
rect 19372 10572 19678 10878
rect 19678 10572 19690 10878
rect 19360 10560 19690 10572
rect 62 10481 488 10498
rect 19312 10481 19738 10498
rect -17 10433 17 10467
rect 19233 10433 19267 10467
rect 19783 10433 19817 10467
rect 62 10402 488 10419
rect 19312 10402 19738 10419
rect 110 10328 440 10340
rect 110 10022 122 10328
rect 122 10022 428 10328
rect 428 10022 440 10328
rect 110 10010 440 10022
rect 19202 9962 19219 10388
rect 19281 9962 19298 10388
rect 62 9931 488 9948
rect 19312 9931 19738 9948
rect -17 9883 17 9917
rect 19233 9883 19267 9917
rect 19783 9883 19817 9917
rect 62 9852 488 9869
rect 19312 9852 19738 9869
rect 19202 9412 19219 9838
rect 19281 9412 19298 9838
rect 19360 9778 19690 9790
rect 19360 9472 19372 9778
rect 19372 9472 19678 9778
rect 19678 9472 19690 9778
rect 19360 9460 19690 9472
rect 62 9381 488 9398
rect 19312 9381 19738 9398
rect -17 9333 17 9367
rect 19233 9333 19267 9367
rect 19783 9333 19817 9367
rect 62 9302 488 9319
rect 19312 9302 19738 9319
rect 110 9228 440 9240
rect 110 8922 122 9228
rect 122 8922 428 9228
rect 428 8922 440 9228
rect 110 8910 440 8922
rect 19202 8862 19219 9288
rect 19281 8862 19298 9288
rect 62 8831 488 8848
rect 19312 8831 19738 8848
rect -17 8783 17 8817
rect 19233 8783 19267 8817
rect 19783 8783 19817 8817
rect 62 8752 488 8769
rect 19312 8752 19738 8769
rect 19202 8312 19219 8738
rect 19281 8312 19298 8738
rect 19360 8678 19690 8690
rect 19360 8372 19372 8678
rect 19372 8372 19678 8678
rect 19678 8372 19690 8678
rect 19360 8360 19690 8372
rect 62 8281 488 8298
rect 19312 8281 19738 8298
rect -17 8233 17 8267
rect 19233 8233 19267 8267
rect 19783 8233 19817 8267
rect 62 8202 488 8219
rect 19312 8202 19738 8219
rect 110 8128 440 8140
rect 110 7822 122 8128
rect 122 7822 428 8128
rect 428 7822 440 8128
rect 110 7810 440 7822
rect 19202 7762 19219 8188
rect 19281 7762 19298 8188
rect 62 7731 488 7748
rect 19312 7731 19738 7748
rect -17 7683 17 7717
rect 19233 7683 19267 7717
rect 19783 7683 19817 7717
rect 62 7652 488 7669
rect 19312 7652 19738 7669
rect 19202 7212 19219 7638
rect 19281 7212 19298 7638
rect 19360 7578 19690 7590
rect 19360 7272 19372 7578
rect 19372 7272 19678 7578
rect 19678 7272 19690 7578
rect 19360 7260 19690 7272
rect 62 7181 488 7198
rect 19312 7181 19738 7198
rect -17 7133 17 7167
rect 19233 7133 19267 7167
rect 19783 7133 19817 7167
rect 62 7102 488 7119
rect 19312 7102 19738 7119
rect 110 7028 440 7040
rect 110 6722 122 7028
rect 122 6722 428 7028
rect 428 6722 440 7028
rect 110 6710 440 6722
rect 19202 6662 19219 7088
rect 19281 6662 19298 7088
rect 62 6631 488 6648
rect 19312 6631 19738 6648
rect -17 6583 17 6617
rect 19233 6583 19267 6617
rect 19783 6583 19817 6617
rect 62 6552 488 6569
rect 19312 6552 19738 6569
rect 19202 6112 19219 6538
rect 19281 6112 19298 6538
rect 19360 6478 19690 6490
rect 19360 6172 19372 6478
rect 19372 6172 19678 6478
rect 19678 6172 19690 6478
rect 19360 6160 19690 6172
rect 62 6081 488 6098
rect 19312 6081 19738 6098
rect -17 6033 17 6067
rect 19233 6033 19267 6067
rect 19783 6033 19817 6067
rect 62 6002 488 6019
rect 19312 6002 19738 6019
rect 110 5928 440 5940
rect 110 5622 122 5928
rect 122 5622 428 5928
rect 428 5622 440 5928
rect 110 5610 440 5622
rect 19202 5562 19219 5988
rect 19281 5562 19298 5988
rect 62 5531 488 5548
rect 19312 5531 19738 5548
rect -17 5483 17 5517
rect 19233 5483 19267 5517
rect 19783 5483 19817 5517
rect 62 5452 488 5469
rect 19312 5452 19738 5469
rect 19202 5012 19219 5438
rect 19281 5012 19298 5438
rect 19360 5378 19690 5390
rect 19360 5072 19372 5378
rect 19372 5072 19678 5378
rect 19678 5072 19690 5378
rect 19360 5060 19690 5072
rect 62 4981 488 4998
rect 19312 4981 19738 4998
rect -17 4933 17 4967
rect 19233 4933 19267 4967
rect 19783 4933 19817 4967
rect 62 4902 488 4919
rect 19312 4902 19738 4919
rect 110 4828 440 4840
rect 110 4522 122 4828
rect 122 4522 428 4828
rect 428 4522 440 4828
rect 110 4510 440 4522
rect 19202 4462 19219 4888
rect 19281 4462 19298 4888
rect 62 4431 488 4448
rect 19312 4431 19738 4448
rect -17 4383 17 4417
rect 19233 4383 19267 4417
rect 19783 4383 19817 4417
rect 62 4352 488 4369
rect 19312 4352 19738 4369
rect 19202 3912 19219 4338
rect 19281 3912 19298 4338
rect 19360 4278 19690 4290
rect 19360 3972 19372 4278
rect 19372 3972 19678 4278
rect 19678 3972 19690 4278
rect 19360 3960 19690 3972
rect 62 3881 488 3898
rect 19312 3881 19738 3898
rect -17 3833 17 3867
rect 19233 3833 19267 3867
rect 19783 3833 19817 3867
rect 62 3802 488 3819
rect 19312 3802 19738 3819
rect 110 3728 440 3740
rect 110 3422 122 3728
rect 122 3422 428 3728
rect 428 3422 440 3728
rect 110 3410 440 3422
rect 19202 3362 19219 3788
rect 19281 3362 19298 3788
rect 62 3331 488 3348
rect 19312 3331 19738 3348
rect -17 3283 17 3317
rect 19233 3283 19267 3317
rect 19783 3283 19817 3317
rect 62 3252 488 3269
rect 19312 3252 19738 3269
rect 19202 2812 19219 3238
rect 19281 2812 19298 3238
rect 19360 3178 19690 3190
rect 19360 2872 19372 3178
rect 19372 2872 19678 3178
rect 19678 2872 19690 3178
rect 19360 2860 19690 2872
rect 62 2781 488 2798
rect 19312 2781 19738 2798
rect -17 2733 17 2767
rect 19233 2733 19267 2767
rect 19783 2733 19817 2767
rect 62 2702 488 2719
rect 19312 2702 19738 2719
rect 110 2628 440 2640
rect 110 2322 122 2628
rect 122 2322 428 2628
rect 428 2322 440 2628
rect 110 2310 440 2322
rect 19202 2262 19219 2688
rect 19281 2262 19298 2688
rect 62 2231 488 2248
rect 19312 2231 19738 2248
rect -17 2183 17 2217
rect 19233 2183 19267 2217
rect 19783 2183 19817 2217
rect 62 2152 488 2169
rect 19312 2152 19738 2169
rect 19202 1712 19219 2138
rect 19281 1712 19298 2138
rect 19360 2078 19690 2090
rect 19360 1772 19372 2078
rect 19372 1772 19678 2078
rect 19678 1772 19690 2078
rect 19360 1760 19690 1772
rect 62 1681 488 1698
rect 19312 1681 19738 1698
rect -17 1633 17 1667
rect 19233 1633 19267 1667
rect 19783 1633 19817 1667
rect 62 1602 488 1619
rect 19312 1602 19738 1619
rect 110 1528 440 1540
rect 110 1222 122 1528
rect 122 1222 428 1528
rect 428 1222 440 1528
rect 110 1210 440 1222
rect 19202 1162 19219 1588
rect 19281 1162 19298 1588
rect 62 1131 488 1148
rect 19312 1131 19738 1148
rect -17 1083 17 1117
rect 19233 1083 19267 1117
rect 19783 1083 19817 1117
rect 62 1052 488 1069
rect 19312 1052 19738 1069
rect 19202 612 19219 1038
rect 19281 612 19298 1038
rect 19360 978 19690 990
rect 19360 672 19372 978
rect 19372 672 19678 978
rect 19678 672 19690 978
rect 19360 660 19690 672
rect 62 581 488 598
rect 19312 581 19738 598
rect -17 533 17 567
rect 19233 533 19267 567
rect 19783 533 19817 567
rect 62 502 488 519
rect 19312 502 19738 519
rect 110 428 440 440
rect 110 122 122 428
rect 122 122 428 428
rect 428 122 440 428
rect 110 110 440 122
rect 502 62 519 488
rect 581 62 598 488
rect 1052 62 1069 488
rect 1131 62 1148 488
rect 1210 428 1540 440
rect 1210 122 1222 428
rect 1222 122 1528 428
rect 1528 122 1540 428
rect 1210 110 1540 122
rect 1602 62 1619 488
rect 1681 62 1698 488
rect 2152 62 2169 488
rect 2231 62 2248 488
rect 2310 428 2640 440
rect 2310 122 2322 428
rect 2322 122 2628 428
rect 2628 122 2640 428
rect 2310 110 2640 122
rect 2702 62 2719 488
rect 2781 62 2798 488
rect 3252 62 3269 488
rect 3331 62 3348 488
rect 3410 428 3740 440
rect 3410 122 3422 428
rect 3422 122 3728 428
rect 3728 122 3740 428
rect 3410 110 3740 122
rect 3802 62 3819 488
rect 3881 62 3898 488
rect 4352 62 4369 488
rect 4431 62 4448 488
rect 4510 428 4840 440
rect 4510 122 4522 428
rect 4522 122 4828 428
rect 4828 122 4840 428
rect 4510 110 4840 122
rect 4902 62 4919 488
rect 4981 62 4998 488
rect 5452 62 5469 488
rect 5531 62 5548 488
rect 5610 428 5940 440
rect 5610 122 5622 428
rect 5622 122 5928 428
rect 5928 122 5940 428
rect 5610 110 5940 122
rect 6002 62 6019 488
rect 6081 62 6098 488
rect 6552 62 6569 488
rect 6631 62 6648 488
rect 6710 428 7040 440
rect 6710 122 6722 428
rect 6722 122 7028 428
rect 7028 122 7040 428
rect 6710 110 7040 122
rect 7102 62 7119 488
rect 7181 62 7198 488
rect 7652 62 7669 488
rect 7731 62 7748 488
rect 7810 428 8140 440
rect 7810 122 7822 428
rect 7822 122 8128 428
rect 8128 122 8140 428
rect 7810 110 8140 122
rect 8202 62 8219 488
rect 8281 62 8298 488
rect 8752 62 8769 488
rect 8831 62 8848 488
rect 8910 428 9240 440
rect 8910 122 8922 428
rect 8922 122 9228 428
rect 9228 122 9240 428
rect 8910 110 9240 122
rect 9302 62 9319 488
rect 9381 62 9398 488
rect 9852 62 9869 488
rect 9931 62 9948 488
rect 10010 428 10340 440
rect 10010 122 10022 428
rect 10022 122 10328 428
rect 10328 122 10340 428
rect 10010 110 10340 122
rect 10402 62 10419 488
rect 10481 62 10498 488
rect 10952 62 10969 488
rect 11031 62 11048 488
rect 11110 428 11440 440
rect 11110 122 11122 428
rect 11122 122 11428 428
rect 11428 122 11440 428
rect 11110 110 11440 122
rect 11502 62 11519 488
rect 11581 62 11598 488
rect 12052 62 12069 488
rect 12131 62 12148 488
rect 12210 428 12540 440
rect 12210 122 12222 428
rect 12222 122 12528 428
rect 12528 122 12540 428
rect 12210 110 12540 122
rect 12602 62 12619 488
rect 12681 62 12698 488
rect 13152 62 13169 488
rect 13231 62 13248 488
rect 13310 428 13640 440
rect 13310 122 13322 428
rect 13322 122 13628 428
rect 13628 122 13640 428
rect 13310 110 13640 122
rect 13702 62 13719 488
rect 13781 62 13798 488
rect 14252 62 14269 488
rect 14331 62 14348 488
rect 14410 428 14740 440
rect 14410 122 14422 428
rect 14422 122 14728 428
rect 14728 122 14740 428
rect 14410 110 14740 122
rect 14802 62 14819 488
rect 14881 62 14898 488
rect 15352 62 15369 488
rect 15431 62 15448 488
rect 15510 428 15840 440
rect 15510 122 15522 428
rect 15522 122 15828 428
rect 15828 122 15840 428
rect 15510 110 15840 122
rect 15902 62 15919 488
rect 15981 62 15998 488
rect 16452 62 16469 488
rect 16531 62 16548 488
rect 16610 428 16940 440
rect 16610 122 16622 428
rect 16622 122 16928 428
rect 16928 122 16940 428
rect 16610 110 16940 122
rect 17002 62 17019 488
rect 17081 62 17098 488
rect 17552 62 17569 488
rect 17631 62 17648 488
rect 17710 428 18040 440
rect 17710 122 17722 428
rect 17722 122 18028 428
rect 18028 122 18040 428
rect 17710 110 18040 122
rect 18102 62 18119 488
rect 18181 62 18198 488
rect 18652 62 18669 488
rect 18731 62 18748 488
rect 18810 428 19140 440
rect 18810 122 18822 428
rect 18822 122 19128 428
rect 19128 122 19140 428
rect 18810 110 19140 122
rect 19202 62 19219 488
rect 19281 62 19298 488
rect -17 -17 17 17
rect 533 -17 567 17
rect 1083 -17 1117 17
rect 1633 -17 1667 17
rect 2183 -17 2217 17
rect 2733 -17 2767 17
rect 3283 -17 3317 17
rect 3833 -17 3867 17
rect 4383 -17 4417 17
rect 4933 -17 4967 17
rect 5483 -17 5517 17
rect 6033 -17 6067 17
rect 6583 -17 6617 17
rect 7133 -17 7167 17
rect 7683 -17 7717 17
rect 8233 -17 8267 17
rect 8783 -17 8817 17
rect 9333 -17 9367 17
rect 9883 -17 9917 17
rect 10433 -17 10467 17
rect 10983 -17 11017 17
rect 11533 -17 11567 17
rect 12083 -17 12117 17
rect 12633 -17 12667 17
rect 13183 -17 13217 17
rect 13733 -17 13767 17
rect 14283 -17 14317 17
rect 14833 -17 14867 17
rect 15383 -17 15417 17
rect 15933 -17 15967 17
rect 16483 -17 16517 17
rect 17033 -17 17067 17
rect 17583 -17 17617 17
rect 18133 -17 18167 17
rect 18683 -17 18717 17
rect 19233 -17 19267 17
rect 19783 -17 19817 17
rect 20012 -212 20288 20012
rect -488 -488 20288 -212
rect 20812 -1012 24788 20812
rect -4988 -4988 24788 -1012
<< metal1 >>
rect -5000 24788 24800 24800
rect -5000 -4988 -4988 24788
rect -1012 20800 20812 20812
rect -1012 -1000 -1000 20800
rect -500 20288 20300 20300
rect -500 -488 -488 20288
rect -212 20000 20012 20012
rect -212 -200 -200 20000
rect -25 19817 25 19825
rect -25 19783 -17 19817
rect 17 19783 25 19817
rect -25 19775 25 19783
rect 525 19817 575 19825
rect 525 19783 533 19817
rect 567 19783 575 19817
rect 525 19775 575 19783
rect 1075 19817 1125 19825
rect 1075 19783 1083 19817
rect 1117 19783 1125 19817
rect 1075 19775 1125 19783
rect 1625 19817 1675 19825
rect 1625 19783 1633 19817
rect 1667 19783 1675 19817
rect 1625 19775 1675 19783
rect 2175 19817 2225 19825
rect 2175 19783 2183 19817
rect 2217 19783 2225 19817
rect 2175 19775 2225 19783
rect 2725 19817 2775 19825
rect 2725 19783 2733 19817
rect 2767 19783 2775 19817
rect 2725 19775 2775 19783
rect 3275 19817 3325 19825
rect 3275 19783 3283 19817
rect 3317 19783 3325 19817
rect 3275 19775 3325 19783
rect 3825 19817 3875 19825
rect 3825 19783 3833 19817
rect 3867 19783 3875 19817
rect 3825 19775 3875 19783
rect 4375 19817 4425 19825
rect 4375 19783 4383 19817
rect 4417 19783 4425 19817
rect 4375 19775 4425 19783
rect 4925 19817 4975 19825
rect 4925 19783 4933 19817
rect 4967 19783 4975 19817
rect 4925 19775 4975 19783
rect 5475 19817 5525 19825
rect 5475 19783 5483 19817
rect 5517 19783 5525 19817
rect 5475 19775 5525 19783
rect 6025 19817 6075 19825
rect 6025 19783 6033 19817
rect 6067 19783 6075 19817
rect 6025 19775 6075 19783
rect 6575 19817 6625 19825
rect 6575 19783 6583 19817
rect 6617 19783 6625 19817
rect 6575 19775 6625 19783
rect 7125 19817 7175 19825
rect 7125 19783 7133 19817
rect 7167 19783 7175 19817
rect 7125 19775 7175 19783
rect 7675 19817 7725 19825
rect 7675 19783 7683 19817
rect 7717 19783 7725 19817
rect 7675 19775 7725 19783
rect 8225 19817 8275 19825
rect 8225 19783 8233 19817
rect 8267 19783 8275 19817
rect 8225 19775 8275 19783
rect 8775 19817 8825 19825
rect 8775 19783 8783 19817
rect 8817 19783 8825 19817
rect 8775 19775 8825 19783
rect 9325 19817 9375 19825
rect 9325 19783 9333 19817
rect 9367 19783 9375 19817
rect 9325 19775 9375 19783
rect 9875 19817 9925 19825
rect 9875 19783 9883 19817
rect 9917 19783 9925 19817
rect 9875 19775 9925 19783
rect 10425 19817 10475 19825
rect 10425 19783 10433 19817
rect 10467 19783 10475 19817
rect 10425 19775 10475 19783
rect 10975 19817 11025 19825
rect 10975 19783 10983 19817
rect 11017 19783 11025 19817
rect 10975 19775 11025 19783
rect 11525 19817 11575 19825
rect 11525 19783 11533 19817
rect 11567 19783 11575 19817
rect 11525 19775 11575 19783
rect 12075 19817 12125 19825
rect 12075 19783 12083 19817
rect 12117 19783 12125 19817
rect 12075 19775 12125 19783
rect 12625 19817 12675 19825
rect 12625 19783 12633 19817
rect 12667 19783 12675 19817
rect 12625 19775 12675 19783
rect 13175 19817 13225 19825
rect 13175 19783 13183 19817
rect 13217 19783 13225 19817
rect 13175 19775 13225 19783
rect 13725 19817 13775 19825
rect 13725 19783 13733 19817
rect 13767 19783 13775 19817
rect 13725 19775 13775 19783
rect 14275 19817 14325 19825
rect 14275 19783 14283 19817
rect 14317 19783 14325 19817
rect 14275 19775 14325 19783
rect 14825 19817 14875 19825
rect 14825 19783 14833 19817
rect 14867 19783 14875 19817
rect 14825 19775 14875 19783
rect 15375 19817 15425 19825
rect 15375 19783 15383 19817
rect 15417 19783 15425 19817
rect 15375 19775 15425 19783
rect 15925 19817 15975 19825
rect 15925 19783 15933 19817
rect 15967 19783 15975 19817
rect 15925 19775 15975 19783
rect 16475 19817 16525 19825
rect 16475 19783 16483 19817
rect 16517 19783 16525 19817
rect 16475 19775 16525 19783
rect 17025 19817 17075 19825
rect 17025 19783 17033 19817
rect 17067 19783 17075 19817
rect 17025 19775 17075 19783
rect 17575 19817 17625 19825
rect 17575 19783 17583 19817
rect 17617 19783 17625 19817
rect 17575 19775 17625 19783
rect 18125 19817 18175 19825
rect 18125 19783 18133 19817
rect 18167 19783 18175 19817
rect 18125 19775 18175 19783
rect 18675 19817 18725 19825
rect 18675 19783 18683 19817
rect 18717 19783 18725 19817
rect 18675 19775 18725 19783
rect 19225 19817 19275 19825
rect 19225 19783 19233 19817
rect 19267 19783 19275 19817
rect 19225 19775 19275 19783
rect 19775 19817 19825 19825
rect 19775 19783 19783 19817
rect 19817 19783 19825 19817
rect 19775 19775 19825 19783
rect 51 19744 499 19749
rect 601 19744 1049 19749
rect 1151 19744 1599 19749
rect 1701 19744 2149 19749
rect 2251 19744 2699 19749
rect 2801 19744 3249 19749
rect 3351 19744 3799 19749
rect 3901 19744 4349 19749
rect 4451 19744 4899 19749
rect 5001 19744 5449 19749
rect 5551 19744 5999 19749
rect 6101 19744 6549 19749
rect 6651 19744 7099 19749
rect 7201 19744 7649 19749
rect 7751 19744 8199 19749
rect 8301 19744 8749 19749
rect 8851 19744 9299 19749
rect 9401 19744 9849 19749
rect 9951 19744 10399 19749
rect 10501 19744 10949 19749
rect 11051 19744 11499 19749
rect 11601 19744 12049 19749
rect 12151 19744 12599 19749
rect 12701 19744 13149 19749
rect 13251 19744 13699 19749
rect 13801 19744 14249 19749
rect 14351 19744 14799 19749
rect 14901 19744 15349 19749
rect 15451 19744 15899 19749
rect 16001 19744 16449 19749
rect 16551 19744 16999 19749
rect 17101 19744 17549 19749
rect 17651 19744 18099 19749
rect 18201 19744 18649 19749
rect 18751 19744 19199 19749
rect 19301 19744 19749 19749
rect 51 19738 522 19744
rect 51 19690 502 19738
rect 51 19360 110 19690
rect 440 19360 502 19690
rect 51 19312 502 19360
rect 519 19312 522 19738
rect 51 19306 522 19312
rect 578 19738 1072 19744
rect 578 19312 581 19738
rect 598 19690 1052 19738
rect 598 19360 660 19690
rect 990 19360 1052 19690
rect 598 19312 1052 19360
rect 1069 19312 1072 19738
rect 578 19306 1072 19312
rect 1128 19738 1622 19744
rect 1128 19312 1131 19738
rect 1148 19690 1602 19738
rect 1148 19360 1210 19690
rect 1540 19360 1602 19690
rect 1148 19312 1602 19360
rect 1619 19312 1622 19738
rect 1128 19306 1622 19312
rect 1678 19738 2172 19744
rect 1678 19312 1681 19738
rect 1698 19690 2152 19738
rect 1698 19360 1760 19690
rect 2090 19360 2152 19690
rect 1698 19312 2152 19360
rect 2169 19312 2172 19738
rect 1678 19306 2172 19312
rect 2228 19738 2722 19744
rect 2228 19312 2231 19738
rect 2248 19690 2702 19738
rect 2248 19360 2310 19690
rect 2640 19360 2702 19690
rect 2248 19312 2702 19360
rect 2719 19312 2722 19738
rect 2228 19306 2722 19312
rect 2778 19738 3272 19744
rect 2778 19312 2781 19738
rect 2798 19690 3252 19738
rect 2798 19360 2860 19690
rect 3190 19360 3252 19690
rect 2798 19312 3252 19360
rect 3269 19312 3272 19738
rect 2778 19306 3272 19312
rect 3328 19738 3822 19744
rect 3328 19312 3331 19738
rect 3348 19690 3802 19738
rect 3348 19360 3410 19690
rect 3740 19360 3802 19690
rect 3348 19312 3802 19360
rect 3819 19312 3822 19738
rect 3328 19306 3822 19312
rect 3878 19738 4372 19744
rect 3878 19312 3881 19738
rect 3898 19690 4352 19738
rect 3898 19360 3960 19690
rect 4290 19360 4352 19690
rect 3898 19312 4352 19360
rect 4369 19312 4372 19738
rect 3878 19306 4372 19312
rect 4428 19738 4922 19744
rect 4428 19312 4431 19738
rect 4448 19690 4902 19738
rect 4448 19360 4510 19690
rect 4840 19360 4902 19690
rect 4448 19312 4902 19360
rect 4919 19312 4922 19738
rect 4428 19306 4922 19312
rect 4978 19738 5472 19744
rect 4978 19312 4981 19738
rect 4998 19690 5452 19738
rect 4998 19360 5060 19690
rect 5390 19360 5452 19690
rect 4998 19312 5452 19360
rect 5469 19312 5472 19738
rect 4978 19306 5472 19312
rect 5528 19738 6022 19744
rect 5528 19312 5531 19738
rect 5548 19690 6002 19738
rect 5548 19360 5610 19690
rect 5940 19360 6002 19690
rect 5548 19312 6002 19360
rect 6019 19312 6022 19738
rect 5528 19306 6022 19312
rect 6078 19738 6572 19744
rect 6078 19312 6081 19738
rect 6098 19690 6552 19738
rect 6098 19360 6160 19690
rect 6490 19360 6552 19690
rect 6098 19312 6552 19360
rect 6569 19312 6572 19738
rect 6078 19306 6572 19312
rect 6628 19738 7122 19744
rect 6628 19312 6631 19738
rect 6648 19690 7102 19738
rect 6648 19360 6710 19690
rect 7040 19360 7102 19690
rect 6648 19312 7102 19360
rect 7119 19312 7122 19738
rect 6628 19306 7122 19312
rect 7178 19738 7672 19744
rect 7178 19312 7181 19738
rect 7198 19690 7652 19738
rect 7198 19360 7260 19690
rect 7590 19360 7652 19690
rect 7198 19312 7652 19360
rect 7669 19312 7672 19738
rect 7178 19306 7672 19312
rect 7728 19738 8222 19744
rect 7728 19312 7731 19738
rect 7748 19690 8202 19738
rect 7748 19360 7810 19690
rect 8140 19360 8202 19690
rect 7748 19312 8202 19360
rect 8219 19312 8222 19738
rect 7728 19306 8222 19312
rect 8278 19738 8772 19744
rect 8278 19312 8281 19738
rect 8298 19690 8752 19738
rect 8298 19360 8360 19690
rect 8690 19360 8752 19690
rect 8298 19312 8752 19360
rect 8769 19312 8772 19738
rect 8278 19306 8772 19312
rect 8828 19738 9322 19744
rect 8828 19312 8831 19738
rect 8848 19690 9302 19738
rect 8848 19360 8910 19690
rect 9240 19360 9302 19690
rect 8848 19312 9302 19360
rect 9319 19312 9322 19738
rect 8828 19306 9322 19312
rect 9378 19738 9872 19744
rect 9378 19312 9381 19738
rect 9398 19690 9852 19738
rect 9398 19360 9460 19690
rect 9790 19360 9852 19690
rect 9398 19312 9852 19360
rect 9869 19312 9872 19738
rect 9378 19306 9872 19312
rect 9928 19738 10422 19744
rect 9928 19312 9931 19738
rect 9948 19690 10402 19738
rect 9948 19360 10010 19690
rect 10340 19360 10402 19690
rect 9948 19312 10402 19360
rect 10419 19312 10422 19738
rect 9928 19306 10422 19312
rect 10478 19738 10972 19744
rect 10478 19312 10481 19738
rect 10498 19690 10952 19738
rect 10498 19360 10560 19690
rect 10890 19360 10952 19690
rect 10498 19312 10952 19360
rect 10969 19312 10972 19738
rect 10478 19306 10972 19312
rect 11028 19738 11522 19744
rect 11028 19312 11031 19738
rect 11048 19690 11502 19738
rect 11048 19360 11110 19690
rect 11440 19360 11502 19690
rect 11048 19312 11502 19360
rect 11519 19312 11522 19738
rect 11028 19306 11522 19312
rect 11578 19738 12072 19744
rect 11578 19312 11581 19738
rect 11598 19690 12052 19738
rect 11598 19360 11660 19690
rect 11990 19360 12052 19690
rect 11598 19312 12052 19360
rect 12069 19312 12072 19738
rect 11578 19306 12072 19312
rect 12128 19738 12622 19744
rect 12128 19312 12131 19738
rect 12148 19690 12602 19738
rect 12148 19360 12210 19690
rect 12540 19360 12602 19690
rect 12148 19312 12602 19360
rect 12619 19312 12622 19738
rect 12128 19306 12622 19312
rect 12678 19738 13172 19744
rect 12678 19312 12681 19738
rect 12698 19690 13152 19738
rect 12698 19360 12760 19690
rect 13090 19360 13152 19690
rect 12698 19312 13152 19360
rect 13169 19312 13172 19738
rect 12678 19306 13172 19312
rect 13228 19738 13722 19744
rect 13228 19312 13231 19738
rect 13248 19690 13702 19738
rect 13248 19360 13310 19690
rect 13640 19360 13702 19690
rect 13248 19312 13702 19360
rect 13719 19312 13722 19738
rect 13228 19306 13722 19312
rect 13778 19738 14272 19744
rect 13778 19312 13781 19738
rect 13798 19690 14252 19738
rect 13798 19360 13860 19690
rect 14190 19360 14252 19690
rect 13798 19312 14252 19360
rect 14269 19312 14272 19738
rect 13778 19306 14272 19312
rect 14328 19738 14822 19744
rect 14328 19312 14331 19738
rect 14348 19690 14802 19738
rect 14348 19360 14410 19690
rect 14740 19360 14802 19690
rect 14348 19312 14802 19360
rect 14819 19312 14822 19738
rect 14328 19306 14822 19312
rect 14878 19738 15372 19744
rect 14878 19312 14881 19738
rect 14898 19690 15352 19738
rect 14898 19360 14960 19690
rect 15290 19360 15352 19690
rect 14898 19312 15352 19360
rect 15369 19312 15372 19738
rect 14878 19306 15372 19312
rect 15428 19738 15922 19744
rect 15428 19312 15431 19738
rect 15448 19690 15902 19738
rect 15448 19360 15510 19690
rect 15840 19360 15902 19690
rect 15448 19312 15902 19360
rect 15919 19312 15922 19738
rect 15428 19306 15922 19312
rect 15978 19738 16472 19744
rect 15978 19312 15981 19738
rect 15998 19690 16452 19738
rect 15998 19360 16060 19690
rect 16390 19360 16452 19690
rect 15998 19312 16452 19360
rect 16469 19312 16472 19738
rect 15978 19306 16472 19312
rect 16528 19738 17022 19744
rect 16528 19312 16531 19738
rect 16548 19690 17002 19738
rect 16548 19360 16610 19690
rect 16940 19360 17002 19690
rect 16548 19312 17002 19360
rect 17019 19312 17022 19738
rect 16528 19306 17022 19312
rect 17078 19738 17572 19744
rect 17078 19312 17081 19738
rect 17098 19690 17552 19738
rect 17098 19360 17160 19690
rect 17490 19360 17552 19690
rect 17098 19312 17552 19360
rect 17569 19312 17572 19738
rect 17078 19306 17572 19312
rect 17628 19738 18122 19744
rect 17628 19312 17631 19738
rect 17648 19690 18102 19738
rect 17648 19360 17710 19690
rect 18040 19360 18102 19690
rect 17648 19312 18102 19360
rect 18119 19312 18122 19738
rect 17628 19306 18122 19312
rect 18178 19738 18672 19744
rect 18178 19312 18181 19738
rect 18198 19690 18652 19738
rect 18198 19360 18260 19690
rect 18590 19360 18652 19690
rect 18198 19312 18652 19360
rect 18669 19312 18672 19738
rect 18178 19306 18672 19312
rect 18728 19738 19222 19744
rect 18728 19312 18731 19738
rect 18748 19690 19202 19738
rect 18748 19360 18810 19690
rect 19140 19360 19202 19690
rect 18748 19312 19202 19360
rect 19219 19312 19222 19738
rect 18728 19306 19222 19312
rect 19278 19738 19749 19744
rect 19278 19312 19281 19738
rect 19298 19690 19749 19738
rect 19298 19360 19360 19690
rect 19690 19360 19749 19690
rect 19298 19312 19749 19360
rect 19278 19306 19749 19312
rect 51 19301 499 19306
rect 601 19301 1049 19306
rect 1151 19301 1599 19306
rect 1701 19301 2149 19306
rect 2251 19301 2699 19306
rect 2801 19301 3249 19306
rect 3351 19301 3799 19306
rect 3901 19301 4349 19306
rect 4451 19301 4899 19306
rect 5001 19301 5449 19306
rect 5551 19301 5999 19306
rect 6101 19301 6549 19306
rect 6651 19301 7099 19306
rect 7201 19301 7649 19306
rect 7751 19301 8199 19306
rect 8301 19301 8749 19306
rect 8851 19301 9299 19306
rect 9401 19301 9849 19306
rect 9951 19301 10399 19306
rect 10501 19301 10949 19306
rect 11051 19301 11499 19306
rect 11601 19301 12049 19306
rect 12151 19301 12599 19306
rect 12701 19301 13149 19306
rect 13251 19301 13699 19306
rect 13801 19301 14249 19306
rect 14351 19301 14799 19306
rect 14901 19301 15349 19306
rect 15451 19301 15899 19306
rect 16001 19301 16449 19306
rect 16551 19301 16999 19306
rect 17101 19301 17549 19306
rect 17651 19301 18099 19306
rect 18201 19301 18649 19306
rect 18751 19301 19199 19306
rect 19301 19301 19749 19306
rect 56 19298 494 19301
rect 56 19281 62 19298
rect 488 19281 494 19298
rect 56 19278 494 19281
rect 606 19298 1044 19301
rect 606 19281 612 19298
rect 1038 19281 1044 19298
rect 606 19278 1044 19281
rect 1156 19298 1594 19301
rect 1156 19281 1162 19298
rect 1588 19281 1594 19298
rect 1156 19278 1594 19281
rect 1706 19298 2144 19301
rect 1706 19281 1712 19298
rect 2138 19281 2144 19298
rect 1706 19278 2144 19281
rect 2256 19298 2694 19301
rect 2256 19281 2262 19298
rect 2688 19281 2694 19298
rect 2256 19278 2694 19281
rect 2806 19298 3244 19301
rect 2806 19281 2812 19298
rect 3238 19281 3244 19298
rect 2806 19278 3244 19281
rect 3356 19298 3794 19301
rect 3356 19281 3362 19298
rect 3788 19281 3794 19298
rect 3356 19278 3794 19281
rect 3906 19298 4344 19301
rect 3906 19281 3912 19298
rect 4338 19281 4344 19298
rect 3906 19278 4344 19281
rect 4456 19298 4894 19301
rect 4456 19281 4462 19298
rect 4888 19281 4894 19298
rect 4456 19278 4894 19281
rect 5006 19298 5444 19301
rect 5006 19281 5012 19298
rect 5438 19281 5444 19298
rect 5006 19278 5444 19281
rect 5556 19298 5994 19301
rect 5556 19281 5562 19298
rect 5988 19281 5994 19298
rect 5556 19278 5994 19281
rect 6106 19298 6544 19301
rect 6106 19281 6112 19298
rect 6538 19281 6544 19298
rect 6106 19278 6544 19281
rect 6656 19298 7094 19301
rect 6656 19281 6662 19298
rect 7088 19281 7094 19298
rect 6656 19278 7094 19281
rect 7206 19298 7644 19301
rect 7206 19281 7212 19298
rect 7638 19281 7644 19298
rect 7206 19278 7644 19281
rect 7756 19298 8194 19301
rect 7756 19281 7762 19298
rect 8188 19281 8194 19298
rect 7756 19278 8194 19281
rect 8306 19298 8744 19301
rect 8306 19281 8312 19298
rect 8738 19281 8744 19298
rect 8306 19278 8744 19281
rect 8856 19298 9294 19301
rect 8856 19281 8862 19298
rect 9288 19281 9294 19298
rect 8856 19278 9294 19281
rect 9406 19298 9844 19301
rect 9406 19281 9412 19298
rect 9838 19281 9844 19298
rect 9406 19278 9844 19281
rect 9956 19298 10394 19301
rect 9956 19281 9962 19298
rect 10388 19281 10394 19298
rect 9956 19278 10394 19281
rect 10506 19298 10944 19301
rect 10506 19281 10512 19298
rect 10938 19281 10944 19298
rect 10506 19278 10944 19281
rect 11056 19298 11494 19301
rect 11056 19281 11062 19298
rect 11488 19281 11494 19298
rect 11056 19278 11494 19281
rect 11606 19298 12044 19301
rect 11606 19281 11612 19298
rect 12038 19281 12044 19298
rect 11606 19278 12044 19281
rect 12156 19298 12594 19301
rect 12156 19281 12162 19298
rect 12588 19281 12594 19298
rect 12156 19278 12594 19281
rect 12706 19298 13144 19301
rect 12706 19281 12712 19298
rect 13138 19281 13144 19298
rect 12706 19278 13144 19281
rect 13256 19298 13694 19301
rect 13256 19281 13262 19298
rect 13688 19281 13694 19298
rect 13256 19278 13694 19281
rect 13806 19298 14244 19301
rect 13806 19281 13812 19298
rect 14238 19281 14244 19298
rect 13806 19278 14244 19281
rect 14356 19298 14794 19301
rect 14356 19281 14362 19298
rect 14788 19281 14794 19298
rect 14356 19278 14794 19281
rect 14906 19298 15344 19301
rect 14906 19281 14912 19298
rect 15338 19281 15344 19298
rect 14906 19278 15344 19281
rect 15456 19298 15894 19301
rect 15456 19281 15462 19298
rect 15888 19281 15894 19298
rect 15456 19278 15894 19281
rect 16006 19298 16444 19301
rect 16006 19281 16012 19298
rect 16438 19281 16444 19298
rect 16006 19278 16444 19281
rect 16556 19298 16994 19301
rect 16556 19281 16562 19298
rect 16988 19281 16994 19298
rect 16556 19278 16994 19281
rect 17106 19298 17544 19301
rect 17106 19281 17112 19298
rect 17538 19281 17544 19298
rect 17106 19278 17544 19281
rect 17656 19298 18094 19301
rect 17656 19281 17662 19298
rect 18088 19281 18094 19298
rect 17656 19278 18094 19281
rect 18206 19298 18644 19301
rect 18206 19281 18212 19298
rect 18638 19281 18644 19298
rect 18206 19278 18644 19281
rect 18756 19298 19194 19301
rect 18756 19281 18762 19298
rect 19188 19281 19194 19298
rect 18756 19278 19194 19281
rect 19306 19298 19744 19301
rect 19306 19281 19312 19298
rect 19738 19281 19744 19298
rect 19306 19278 19744 19281
rect -25 19267 25 19275
rect -25 19233 -17 19267
rect 17 19233 25 19267
rect -25 19225 25 19233
rect 525 19267 575 19275
rect 525 19233 533 19267
rect 567 19233 575 19267
rect 525 19225 575 19233
rect 1075 19267 1125 19275
rect 1075 19233 1083 19267
rect 1117 19233 1125 19267
rect 1075 19225 1125 19233
rect 1625 19267 1675 19275
rect 1625 19233 1633 19267
rect 1667 19233 1675 19267
rect 1625 19225 1675 19233
rect 2175 19267 2225 19275
rect 2175 19233 2183 19267
rect 2217 19233 2225 19267
rect 2175 19225 2225 19233
rect 2725 19267 2775 19275
rect 2725 19233 2733 19267
rect 2767 19233 2775 19267
rect 2725 19225 2775 19233
rect 3275 19267 3325 19275
rect 3275 19233 3283 19267
rect 3317 19233 3325 19267
rect 3275 19225 3325 19233
rect 3825 19267 3875 19275
rect 3825 19233 3833 19267
rect 3867 19233 3875 19267
rect 3825 19225 3875 19233
rect 4375 19267 4425 19275
rect 4375 19233 4383 19267
rect 4417 19233 4425 19267
rect 4375 19225 4425 19233
rect 4925 19267 4975 19275
rect 4925 19233 4933 19267
rect 4967 19233 4975 19267
rect 4925 19225 4975 19233
rect 5475 19267 5525 19275
rect 5475 19233 5483 19267
rect 5517 19233 5525 19267
rect 5475 19225 5525 19233
rect 6025 19267 6075 19275
rect 6025 19233 6033 19267
rect 6067 19233 6075 19267
rect 6025 19225 6075 19233
rect 6575 19267 6625 19275
rect 6575 19233 6583 19267
rect 6617 19233 6625 19267
rect 6575 19225 6625 19233
rect 7125 19267 7175 19275
rect 7125 19233 7133 19267
rect 7167 19233 7175 19267
rect 7125 19225 7175 19233
rect 7675 19267 7725 19275
rect 7675 19233 7683 19267
rect 7717 19233 7725 19267
rect 7675 19225 7725 19233
rect 8225 19267 8275 19275
rect 8225 19233 8233 19267
rect 8267 19233 8275 19267
rect 8225 19225 8275 19233
rect 8775 19267 8825 19275
rect 8775 19233 8783 19267
rect 8817 19233 8825 19267
rect 8775 19225 8825 19233
rect 9325 19267 9375 19275
rect 9325 19233 9333 19267
rect 9367 19233 9375 19267
rect 9325 19225 9375 19233
rect 9875 19267 9925 19275
rect 9875 19233 9883 19267
rect 9917 19233 9925 19267
rect 9875 19225 9925 19233
rect 10425 19267 10475 19275
rect 10425 19233 10433 19267
rect 10467 19233 10475 19267
rect 10425 19225 10475 19233
rect 10975 19267 11025 19275
rect 10975 19233 10983 19267
rect 11017 19233 11025 19267
rect 10975 19225 11025 19233
rect 11525 19267 11575 19275
rect 11525 19233 11533 19267
rect 11567 19233 11575 19267
rect 11525 19225 11575 19233
rect 12075 19267 12125 19275
rect 12075 19233 12083 19267
rect 12117 19233 12125 19267
rect 12075 19225 12125 19233
rect 12625 19267 12675 19275
rect 12625 19233 12633 19267
rect 12667 19233 12675 19267
rect 12625 19225 12675 19233
rect 13175 19267 13225 19275
rect 13175 19233 13183 19267
rect 13217 19233 13225 19267
rect 13175 19225 13225 19233
rect 13725 19267 13775 19275
rect 13725 19233 13733 19267
rect 13767 19233 13775 19267
rect 13725 19225 13775 19233
rect 14275 19267 14325 19275
rect 14275 19233 14283 19267
rect 14317 19233 14325 19267
rect 14275 19225 14325 19233
rect 14825 19267 14875 19275
rect 14825 19233 14833 19267
rect 14867 19233 14875 19267
rect 14825 19225 14875 19233
rect 15375 19267 15425 19275
rect 15375 19233 15383 19267
rect 15417 19233 15425 19267
rect 15375 19225 15425 19233
rect 15925 19267 15975 19275
rect 15925 19233 15933 19267
rect 15967 19233 15975 19267
rect 15925 19225 15975 19233
rect 16475 19267 16525 19275
rect 16475 19233 16483 19267
rect 16517 19233 16525 19267
rect 16475 19225 16525 19233
rect 17025 19267 17075 19275
rect 17025 19233 17033 19267
rect 17067 19233 17075 19267
rect 17025 19225 17075 19233
rect 17575 19267 17625 19275
rect 17575 19233 17583 19267
rect 17617 19233 17625 19267
rect 17575 19225 17625 19233
rect 18125 19267 18175 19275
rect 18125 19233 18133 19267
rect 18167 19233 18175 19267
rect 18125 19225 18175 19233
rect 18675 19267 18725 19275
rect 18675 19233 18683 19267
rect 18717 19233 18725 19267
rect 18675 19225 18725 19233
rect 19225 19267 19275 19275
rect 19225 19233 19233 19267
rect 19267 19233 19275 19267
rect 19225 19225 19275 19233
rect 19775 19267 19825 19275
rect 19775 19233 19783 19267
rect 19817 19233 19825 19267
rect 19775 19225 19825 19233
rect 56 19219 494 19222
rect 56 19202 62 19219
rect 488 19202 494 19219
rect 56 19199 494 19202
rect 606 19219 1044 19222
rect 606 19202 612 19219
rect 1038 19202 1044 19219
rect 606 19200 1044 19202
rect 1156 19219 1594 19222
rect 1156 19202 1162 19219
rect 1588 19202 1594 19219
rect 1156 19200 1594 19202
rect 1706 19219 2144 19222
rect 1706 19202 1712 19219
rect 2138 19202 2144 19219
rect 1706 19200 2144 19202
rect 2256 19219 2694 19222
rect 2256 19202 2262 19219
rect 2688 19202 2694 19219
rect 2256 19200 2694 19202
rect 2806 19219 3244 19222
rect 2806 19202 2812 19219
rect 3238 19202 3244 19219
rect 2806 19200 3244 19202
rect 3356 19219 3794 19222
rect 3356 19202 3362 19219
rect 3788 19202 3794 19219
rect 3356 19200 3794 19202
rect 3906 19219 4344 19222
rect 3906 19202 3912 19219
rect 4338 19202 4344 19219
rect 3906 19200 4344 19202
rect 4456 19219 4894 19222
rect 4456 19202 4462 19219
rect 4888 19202 4894 19219
rect 4456 19200 4894 19202
rect 5006 19219 5444 19222
rect 5006 19202 5012 19219
rect 5438 19202 5444 19219
rect 5006 19200 5444 19202
rect 5556 19219 5994 19222
rect 5556 19202 5562 19219
rect 5988 19202 5994 19219
rect 5556 19200 5994 19202
rect 6106 19219 6544 19222
rect 6106 19202 6112 19219
rect 6538 19202 6544 19219
rect 6106 19200 6544 19202
rect 6656 19219 7094 19222
rect 6656 19202 6662 19219
rect 7088 19202 7094 19219
rect 6656 19200 7094 19202
rect 7206 19219 7644 19222
rect 7206 19202 7212 19219
rect 7638 19202 7644 19219
rect 7206 19200 7644 19202
rect 7756 19219 8194 19222
rect 7756 19202 7762 19219
rect 8188 19202 8194 19219
rect 7756 19200 8194 19202
rect 8306 19219 8744 19222
rect 8306 19202 8312 19219
rect 8738 19202 8744 19219
rect 8306 19200 8744 19202
rect 8856 19219 9294 19222
rect 8856 19202 8862 19219
rect 9288 19202 9294 19219
rect 8856 19200 9294 19202
rect 9406 19219 9844 19222
rect 9406 19202 9412 19219
rect 9838 19202 9844 19219
rect 9406 19200 9844 19202
rect 9956 19219 10394 19222
rect 9956 19202 9962 19219
rect 10388 19202 10394 19219
rect 9956 19200 10394 19202
rect 10506 19219 10944 19222
rect 10506 19202 10512 19219
rect 10938 19202 10944 19219
rect 10506 19200 10944 19202
rect 11056 19219 11494 19222
rect 11056 19202 11062 19219
rect 11488 19202 11494 19219
rect 11056 19200 11494 19202
rect 11606 19219 12044 19222
rect 11606 19202 11612 19219
rect 12038 19202 12044 19219
rect 11606 19200 12044 19202
rect 12156 19219 12594 19222
rect 12156 19202 12162 19219
rect 12588 19202 12594 19219
rect 12156 19200 12594 19202
rect 12706 19219 13144 19222
rect 12706 19202 12712 19219
rect 13138 19202 13144 19219
rect 12706 19200 13144 19202
rect 13256 19219 13694 19222
rect 13256 19202 13262 19219
rect 13688 19202 13694 19219
rect 13256 19200 13694 19202
rect 13806 19219 14244 19222
rect 13806 19202 13812 19219
rect 14238 19202 14244 19219
rect 13806 19200 14244 19202
rect 14356 19219 14794 19222
rect 14356 19202 14362 19219
rect 14788 19202 14794 19219
rect 14356 19200 14794 19202
rect 14906 19219 15344 19222
rect 14906 19202 14912 19219
rect 15338 19202 15344 19219
rect 14906 19200 15344 19202
rect 15456 19219 15894 19222
rect 15456 19202 15462 19219
rect 15888 19202 15894 19219
rect 15456 19200 15894 19202
rect 16006 19219 16444 19222
rect 16006 19202 16012 19219
rect 16438 19202 16444 19219
rect 16006 19200 16444 19202
rect 16556 19219 16994 19222
rect 16556 19202 16562 19219
rect 16988 19202 16994 19219
rect 16556 19200 16994 19202
rect 17106 19219 17544 19222
rect 17106 19202 17112 19219
rect 17538 19202 17544 19219
rect 17106 19200 17544 19202
rect 17656 19219 18094 19222
rect 17656 19202 17662 19219
rect 18088 19202 18094 19219
rect 17656 19200 18094 19202
rect 18206 19219 18644 19222
rect 18206 19202 18212 19219
rect 18638 19202 18644 19219
rect 18206 19200 18644 19202
rect 18756 19219 19194 19222
rect 18756 19202 18762 19219
rect 19188 19202 19194 19219
rect 18756 19200 19194 19202
rect 19306 19219 19744 19222
rect 19306 19202 19312 19219
rect 19738 19202 19744 19219
rect 19306 19199 19744 19202
rect 51 19194 499 19199
rect 19301 19194 19749 19199
rect 51 19140 500 19194
rect 51 18810 110 19140
rect 440 18810 500 19140
rect 51 18756 500 18810
rect 19200 19188 19222 19194
rect 19200 18762 19202 19188
rect 19219 18762 19222 19188
rect 19200 18756 19222 18762
rect 19278 19188 19749 19194
rect 19278 18762 19281 19188
rect 19298 19140 19749 19188
rect 19298 18810 19360 19140
rect 19690 18810 19749 19140
rect 19298 18762 19749 18810
rect 19278 18756 19749 18762
rect 51 18751 499 18756
rect 19301 18751 19749 18756
rect 56 18748 494 18751
rect 56 18731 62 18748
rect 488 18731 494 18748
rect 56 18728 494 18731
rect 19306 18748 19744 18751
rect 19306 18731 19312 18748
rect 19738 18731 19744 18748
rect 19306 18728 19744 18731
rect -25 18717 25 18725
rect -25 18683 -17 18717
rect 17 18683 25 18717
rect -25 18675 25 18683
rect 19225 18717 19275 18725
rect 19225 18683 19233 18717
rect 19267 18683 19275 18717
rect 19225 18675 19275 18683
rect 19775 18717 19825 18725
rect 19775 18683 19783 18717
rect 19817 18683 19825 18717
rect 19775 18675 19825 18683
rect 56 18669 494 18672
rect 56 18652 62 18669
rect 488 18652 494 18669
rect 56 18649 494 18652
rect 19306 18669 19744 18672
rect 19306 18652 19312 18669
rect 19738 18652 19744 18669
rect 19306 18649 19744 18652
rect 51 18644 499 18649
rect 19301 18644 19749 18649
rect 51 18590 500 18644
rect 51 18260 110 18590
rect 440 18260 500 18590
rect 51 18206 500 18260
rect 19200 18638 19222 18644
rect 19200 18212 19202 18638
rect 19219 18212 19222 18638
rect 19200 18206 19222 18212
rect 19278 18638 19749 18644
rect 19278 18212 19281 18638
rect 19298 18590 19749 18638
rect 19298 18260 19360 18590
rect 19690 18260 19749 18590
rect 19298 18212 19749 18260
rect 19278 18206 19749 18212
rect 51 18201 499 18206
rect 19301 18201 19749 18206
rect 56 18198 494 18201
rect 56 18181 62 18198
rect 488 18181 494 18198
rect 56 18178 494 18181
rect 19306 18198 19744 18201
rect 19306 18181 19312 18198
rect 19738 18181 19744 18198
rect 19306 18178 19744 18181
rect -25 18167 25 18175
rect -25 18133 -17 18167
rect 17 18133 25 18167
rect -25 18125 25 18133
rect 19225 18167 19275 18175
rect 19225 18133 19233 18167
rect 19267 18133 19275 18167
rect 19225 18125 19275 18133
rect 19775 18167 19825 18175
rect 19775 18133 19783 18167
rect 19817 18133 19825 18167
rect 19775 18125 19825 18133
rect 56 18119 494 18122
rect 56 18102 62 18119
rect 488 18102 494 18119
rect 56 18099 494 18102
rect 19306 18119 19744 18122
rect 19306 18102 19312 18119
rect 19738 18102 19744 18119
rect 19306 18099 19744 18102
rect 51 18094 499 18099
rect 19301 18094 19749 18099
rect 51 18040 500 18094
rect 51 17710 110 18040
rect 440 17710 500 18040
rect 51 17656 500 17710
rect 19200 18088 19222 18094
rect 19200 17662 19202 18088
rect 19219 17662 19222 18088
rect 19200 17656 19222 17662
rect 19278 18088 19749 18094
rect 19278 17662 19281 18088
rect 19298 18040 19749 18088
rect 19298 17710 19360 18040
rect 19690 17710 19749 18040
rect 19298 17662 19749 17710
rect 19278 17656 19749 17662
rect 51 17651 499 17656
rect 19301 17651 19749 17656
rect 56 17648 494 17651
rect 56 17631 62 17648
rect 488 17631 494 17648
rect 56 17628 494 17631
rect 19306 17648 19744 17651
rect 19306 17631 19312 17648
rect 19738 17631 19744 17648
rect 19306 17628 19744 17631
rect -25 17617 25 17625
rect -25 17583 -17 17617
rect 17 17583 25 17617
rect -25 17575 25 17583
rect 19225 17617 19275 17625
rect 19225 17583 19233 17617
rect 19267 17583 19275 17617
rect 19225 17575 19275 17583
rect 19775 17617 19825 17625
rect 19775 17583 19783 17617
rect 19817 17583 19825 17617
rect 19775 17575 19825 17583
rect 56 17569 494 17572
rect 56 17552 62 17569
rect 488 17552 494 17569
rect 56 17549 494 17552
rect 19306 17569 19744 17572
rect 19306 17552 19312 17569
rect 19738 17552 19744 17569
rect 19306 17549 19744 17552
rect 51 17544 499 17549
rect 19301 17544 19749 17549
rect 51 17490 500 17544
rect 51 17160 110 17490
rect 440 17160 500 17490
rect 51 17106 500 17160
rect 19200 17538 19222 17544
rect 19200 17112 19202 17538
rect 19219 17112 19222 17538
rect 19200 17106 19222 17112
rect 19278 17538 19749 17544
rect 19278 17112 19281 17538
rect 19298 17490 19749 17538
rect 19298 17160 19360 17490
rect 19690 17160 19749 17490
rect 19298 17112 19749 17160
rect 19278 17106 19749 17112
rect 51 17101 499 17106
rect 19301 17101 19749 17106
rect 56 17098 494 17101
rect 56 17081 62 17098
rect 488 17081 494 17098
rect 56 17078 494 17081
rect 19306 17098 19744 17101
rect 19306 17081 19312 17098
rect 19738 17081 19744 17098
rect 19306 17078 19744 17081
rect -25 17067 25 17075
rect -25 17033 -17 17067
rect 17 17033 25 17067
rect -25 17025 25 17033
rect 19225 17067 19275 17075
rect 19225 17033 19233 17067
rect 19267 17033 19275 17067
rect 19225 17025 19275 17033
rect 19775 17067 19825 17075
rect 19775 17033 19783 17067
rect 19817 17033 19825 17067
rect 19775 17025 19825 17033
rect 56 17019 494 17022
rect 56 17002 62 17019
rect 488 17002 494 17019
rect 56 16999 494 17002
rect 19306 17019 19744 17022
rect 19306 17002 19312 17019
rect 19738 17002 19744 17019
rect 19306 16999 19744 17002
rect 51 16994 499 16999
rect 19301 16994 19749 16999
rect 51 16940 500 16994
rect 51 16610 110 16940
rect 440 16610 500 16940
rect 51 16556 500 16610
rect 19200 16988 19222 16994
rect 19200 16562 19202 16988
rect 19219 16562 19222 16988
rect 19200 16556 19222 16562
rect 19278 16988 19749 16994
rect 19278 16562 19281 16988
rect 19298 16940 19749 16988
rect 19298 16610 19360 16940
rect 19690 16610 19749 16940
rect 19298 16562 19749 16610
rect 19278 16556 19749 16562
rect 51 16551 499 16556
rect 19301 16551 19749 16556
rect 56 16548 494 16551
rect 56 16531 62 16548
rect 488 16531 494 16548
rect 56 16528 494 16531
rect 19306 16548 19744 16551
rect 19306 16531 19312 16548
rect 19738 16531 19744 16548
rect 19306 16528 19744 16531
rect -25 16517 25 16525
rect -25 16483 -17 16517
rect 17 16483 25 16517
rect -25 16475 25 16483
rect 19225 16517 19275 16525
rect 19225 16483 19233 16517
rect 19267 16483 19275 16517
rect 19225 16475 19275 16483
rect 19775 16517 19825 16525
rect 19775 16483 19783 16517
rect 19817 16483 19825 16517
rect 19775 16475 19825 16483
rect 56 16469 494 16472
rect 56 16452 62 16469
rect 488 16452 494 16469
rect 56 16449 494 16452
rect 19306 16469 19744 16472
rect 19306 16452 19312 16469
rect 19738 16452 19744 16469
rect 19306 16449 19744 16452
rect 51 16444 499 16449
rect 19301 16444 19749 16449
rect 51 16390 500 16444
rect 51 16060 110 16390
rect 440 16060 500 16390
rect 51 16006 500 16060
rect 19200 16438 19222 16444
rect 19200 16012 19202 16438
rect 19219 16012 19222 16438
rect 19200 16006 19222 16012
rect 19278 16438 19749 16444
rect 19278 16012 19281 16438
rect 19298 16390 19749 16438
rect 19298 16060 19360 16390
rect 19690 16060 19749 16390
rect 19298 16012 19749 16060
rect 19278 16006 19749 16012
rect 51 16001 499 16006
rect 19301 16001 19749 16006
rect 56 15998 494 16001
rect 56 15981 62 15998
rect 488 15981 494 15998
rect 56 15978 494 15981
rect 19306 15998 19744 16001
rect 19306 15981 19312 15998
rect 19738 15981 19744 15998
rect 19306 15978 19744 15981
rect -25 15967 25 15975
rect -25 15933 -17 15967
rect 17 15933 25 15967
rect -25 15925 25 15933
rect 19225 15967 19275 15975
rect 19225 15933 19233 15967
rect 19267 15933 19275 15967
rect 19225 15925 19275 15933
rect 19775 15967 19825 15975
rect 19775 15933 19783 15967
rect 19817 15933 19825 15967
rect 19775 15925 19825 15933
rect 56 15919 494 15922
rect 56 15902 62 15919
rect 488 15902 494 15919
rect 56 15899 494 15902
rect 19306 15919 19744 15922
rect 19306 15902 19312 15919
rect 19738 15902 19744 15919
rect 19306 15899 19744 15902
rect 51 15894 499 15899
rect 19301 15894 19749 15899
rect 51 15840 500 15894
rect 51 15510 110 15840
rect 440 15510 500 15840
rect 51 15456 500 15510
rect 19200 15888 19222 15894
rect 19200 15462 19202 15888
rect 19219 15462 19222 15888
rect 19200 15456 19222 15462
rect 19278 15888 19749 15894
rect 19278 15462 19281 15888
rect 19298 15840 19749 15888
rect 19298 15510 19360 15840
rect 19690 15510 19749 15840
rect 19298 15462 19749 15510
rect 19278 15456 19749 15462
rect 51 15451 499 15456
rect 19301 15451 19749 15456
rect 56 15448 494 15451
rect 56 15431 62 15448
rect 488 15431 494 15448
rect 56 15428 494 15431
rect 19306 15448 19744 15451
rect 19306 15431 19312 15448
rect 19738 15431 19744 15448
rect 19306 15428 19744 15431
rect -25 15417 25 15425
rect -25 15383 -17 15417
rect 17 15383 25 15417
rect -25 15375 25 15383
rect 19225 15417 19275 15425
rect 19225 15383 19233 15417
rect 19267 15383 19275 15417
rect 19225 15375 19275 15383
rect 19775 15417 19825 15425
rect 19775 15383 19783 15417
rect 19817 15383 19825 15417
rect 19775 15375 19825 15383
rect 56 15369 494 15372
rect 56 15352 62 15369
rect 488 15352 494 15369
rect 56 15349 494 15352
rect 19306 15369 19744 15372
rect 19306 15352 19312 15369
rect 19738 15352 19744 15369
rect 19306 15349 19744 15352
rect 51 15344 499 15349
rect 19301 15344 19749 15349
rect 51 15290 500 15344
rect 51 14960 110 15290
rect 440 14960 500 15290
rect 51 14906 500 14960
rect 19200 15338 19222 15344
rect 19200 14912 19202 15338
rect 19219 14912 19222 15338
rect 19200 14906 19222 14912
rect 19278 15338 19749 15344
rect 19278 14912 19281 15338
rect 19298 15290 19749 15338
rect 19298 14960 19360 15290
rect 19690 14960 19749 15290
rect 19298 14912 19749 14960
rect 19278 14906 19749 14912
rect 51 14901 499 14906
rect 19301 14901 19749 14906
rect 56 14898 494 14901
rect 56 14881 62 14898
rect 488 14881 494 14898
rect 56 14878 494 14881
rect 19306 14898 19744 14901
rect 19306 14881 19312 14898
rect 19738 14881 19744 14898
rect 19306 14878 19744 14881
rect -25 14867 25 14875
rect -25 14833 -17 14867
rect 17 14833 25 14867
rect -25 14825 25 14833
rect 19225 14867 19275 14875
rect 19225 14833 19233 14867
rect 19267 14833 19275 14867
rect 19225 14825 19275 14833
rect 19775 14867 19825 14875
rect 19775 14833 19783 14867
rect 19817 14833 19825 14867
rect 19775 14825 19825 14833
rect 56 14819 494 14822
rect 56 14802 62 14819
rect 488 14802 494 14819
rect 56 14799 494 14802
rect 19306 14819 19744 14822
rect 19306 14802 19312 14819
rect 19738 14802 19744 14819
rect 19306 14799 19744 14802
rect 51 14794 499 14799
rect 19301 14794 19749 14799
rect 51 14740 500 14794
rect 51 14410 110 14740
rect 440 14410 500 14740
rect 51 14356 500 14410
rect 19200 14788 19222 14794
rect 19200 14362 19202 14788
rect 19219 14362 19222 14788
rect 19200 14356 19222 14362
rect 19278 14788 19749 14794
rect 19278 14362 19281 14788
rect 19298 14740 19749 14788
rect 19298 14410 19360 14740
rect 19690 14410 19749 14740
rect 19298 14362 19749 14410
rect 19278 14356 19749 14362
rect 51 14351 499 14356
rect 19301 14351 19749 14356
rect 56 14348 494 14351
rect 56 14331 62 14348
rect 488 14331 494 14348
rect 56 14328 494 14331
rect 19306 14348 19744 14351
rect 19306 14331 19312 14348
rect 19738 14331 19744 14348
rect 19306 14328 19744 14331
rect -25 14317 25 14325
rect -25 14283 -17 14317
rect 17 14283 25 14317
rect -25 14275 25 14283
rect 19225 14317 19275 14325
rect 19225 14283 19233 14317
rect 19267 14283 19275 14317
rect 19225 14275 19275 14283
rect 19775 14317 19825 14325
rect 19775 14283 19783 14317
rect 19817 14283 19825 14317
rect 19775 14275 19825 14283
rect 56 14269 494 14272
rect 56 14252 62 14269
rect 488 14252 494 14269
rect 56 14249 494 14252
rect 19306 14269 19744 14272
rect 19306 14252 19312 14269
rect 19738 14252 19744 14269
rect 19306 14249 19744 14252
rect 51 14244 499 14249
rect 19301 14244 19749 14249
rect 51 14190 500 14244
rect 51 13860 110 14190
rect 440 13860 500 14190
rect 51 13806 500 13860
rect 19200 14238 19222 14244
rect 19200 13812 19202 14238
rect 19219 13812 19222 14238
rect 19200 13806 19222 13812
rect 19278 14238 19749 14244
rect 19278 13812 19281 14238
rect 19298 14190 19749 14238
rect 19298 13860 19360 14190
rect 19690 13860 19749 14190
rect 19298 13812 19749 13860
rect 19278 13806 19749 13812
rect 51 13801 499 13806
rect 19301 13801 19749 13806
rect 56 13798 494 13801
rect 56 13781 62 13798
rect 488 13781 494 13798
rect 56 13778 494 13781
rect 19306 13798 19744 13801
rect 19306 13781 19312 13798
rect 19738 13781 19744 13798
rect 19306 13778 19744 13781
rect -25 13767 25 13775
rect -25 13733 -17 13767
rect 17 13733 25 13767
rect -25 13725 25 13733
rect 19225 13767 19275 13775
rect 19225 13733 19233 13767
rect 19267 13733 19275 13767
rect 19225 13725 19275 13733
rect 19775 13767 19825 13775
rect 19775 13733 19783 13767
rect 19817 13733 19825 13767
rect 19775 13725 19825 13733
rect 56 13719 494 13722
rect 56 13702 62 13719
rect 488 13702 494 13719
rect 56 13699 494 13702
rect 19306 13719 19744 13722
rect 19306 13702 19312 13719
rect 19738 13702 19744 13719
rect 19306 13699 19744 13702
rect 51 13694 499 13699
rect 19301 13694 19749 13699
rect 51 13640 500 13694
rect 51 13310 110 13640
rect 440 13310 500 13640
rect 51 13256 500 13310
rect 19200 13688 19222 13694
rect 19200 13262 19202 13688
rect 19219 13262 19222 13688
rect 19200 13256 19222 13262
rect 19278 13688 19749 13694
rect 19278 13262 19281 13688
rect 19298 13640 19749 13688
rect 19298 13310 19360 13640
rect 19690 13310 19749 13640
rect 19298 13262 19749 13310
rect 19278 13256 19749 13262
rect 51 13251 499 13256
rect 19301 13251 19749 13256
rect 56 13248 494 13251
rect 56 13231 62 13248
rect 488 13231 494 13248
rect 56 13228 494 13231
rect 19306 13248 19744 13251
rect 19306 13231 19312 13248
rect 19738 13231 19744 13248
rect 19306 13228 19744 13231
rect -25 13217 25 13225
rect -25 13183 -17 13217
rect 17 13183 25 13217
rect -25 13175 25 13183
rect 19225 13217 19275 13225
rect 19225 13183 19233 13217
rect 19267 13183 19275 13217
rect 19225 13175 19275 13183
rect 19775 13217 19825 13225
rect 19775 13183 19783 13217
rect 19817 13183 19825 13217
rect 19775 13175 19825 13183
rect 56 13169 494 13172
rect 56 13152 62 13169
rect 488 13152 494 13169
rect 56 13149 494 13152
rect 19306 13169 19744 13172
rect 19306 13152 19312 13169
rect 19738 13152 19744 13169
rect 19306 13149 19744 13152
rect 51 13144 499 13149
rect 19301 13144 19749 13149
rect 51 13090 500 13144
rect 51 12760 110 13090
rect 440 12760 500 13090
rect 51 12706 500 12760
rect 19200 13138 19222 13144
rect 19200 12712 19202 13138
rect 19219 12712 19222 13138
rect 19200 12706 19222 12712
rect 19278 13138 19749 13144
rect 19278 12712 19281 13138
rect 19298 13090 19749 13138
rect 19298 12760 19360 13090
rect 19690 12760 19749 13090
rect 19298 12712 19749 12760
rect 19278 12706 19749 12712
rect 51 12701 499 12706
rect 19301 12701 19749 12706
rect 56 12698 494 12701
rect 56 12681 62 12698
rect 488 12681 494 12698
rect 56 12678 494 12681
rect 19306 12698 19744 12701
rect 19306 12681 19312 12698
rect 19738 12681 19744 12698
rect 19306 12678 19744 12681
rect -25 12667 25 12675
rect -25 12633 -17 12667
rect 17 12633 25 12667
rect -25 12625 25 12633
rect 19225 12667 19275 12675
rect 19225 12633 19233 12667
rect 19267 12633 19275 12667
rect 19225 12625 19275 12633
rect 19775 12667 19825 12675
rect 19775 12633 19783 12667
rect 19817 12633 19825 12667
rect 19775 12625 19825 12633
rect 56 12619 494 12622
rect 56 12602 62 12619
rect 488 12602 494 12619
rect 56 12599 494 12602
rect 19306 12619 19744 12622
rect 19306 12602 19312 12619
rect 19738 12602 19744 12619
rect 19306 12599 19744 12602
rect 51 12594 499 12599
rect 19301 12594 19749 12599
rect 51 12540 500 12594
rect 51 12210 110 12540
rect 440 12210 500 12540
rect 51 12156 500 12210
rect 19200 12588 19222 12594
rect 19200 12162 19202 12588
rect 19219 12162 19222 12588
rect 19200 12156 19222 12162
rect 19278 12588 19749 12594
rect 19278 12162 19281 12588
rect 19298 12540 19749 12588
rect 19298 12210 19360 12540
rect 19690 12210 19749 12540
rect 19298 12162 19749 12210
rect 19278 12156 19749 12162
rect 51 12151 499 12156
rect 19301 12151 19749 12156
rect 56 12148 494 12151
rect 56 12131 62 12148
rect 488 12131 494 12148
rect 56 12128 494 12131
rect 19306 12148 19744 12151
rect 19306 12131 19312 12148
rect 19738 12131 19744 12148
rect 19306 12128 19744 12131
rect -25 12117 25 12125
rect -25 12083 -17 12117
rect 17 12083 25 12117
rect -25 12075 25 12083
rect 19225 12117 19275 12125
rect 19225 12083 19233 12117
rect 19267 12083 19275 12117
rect 19225 12075 19275 12083
rect 19775 12117 19825 12125
rect 19775 12083 19783 12117
rect 19817 12083 19825 12117
rect 19775 12075 19825 12083
rect 56 12069 494 12072
rect 56 12052 62 12069
rect 488 12052 494 12069
rect 56 12049 494 12052
rect 19306 12069 19744 12072
rect 19306 12052 19312 12069
rect 19738 12052 19744 12069
rect 19306 12049 19744 12052
rect 51 12044 499 12049
rect 19301 12044 19749 12049
rect 51 11990 500 12044
rect 51 11660 110 11990
rect 440 11660 500 11990
rect 51 11606 500 11660
rect 19200 12038 19222 12044
rect 19200 11612 19202 12038
rect 19219 11612 19222 12038
rect 19200 11606 19222 11612
rect 19278 12038 19749 12044
rect 19278 11612 19281 12038
rect 19298 11990 19749 12038
rect 19298 11660 19360 11990
rect 19690 11660 19749 11990
rect 19298 11612 19749 11660
rect 19278 11606 19749 11612
rect 51 11601 499 11606
rect 19301 11601 19749 11606
rect 56 11598 494 11601
rect 56 11581 62 11598
rect 488 11581 494 11598
rect 56 11578 494 11581
rect 19306 11598 19744 11601
rect 19306 11581 19312 11598
rect 19738 11581 19744 11598
rect 19306 11578 19744 11581
rect -25 11567 25 11575
rect -25 11533 -17 11567
rect 17 11533 25 11567
rect -25 11525 25 11533
rect 19225 11567 19275 11575
rect 19225 11533 19233 11567
rect 19267 11533 19275 11567
rect 19225 11525 19275 11533
rect 19775 11567 19825 11575
rect 19775 11533 19783 11567
rect 19817 11533 19825 11567
rect 19775 11525 19825 11533
rect 56 11519 494 11522
rect 56 11502 62 11519
rect 488 11502 494 11519
rect 56 11499 494 11502
rect 19306 11519 19744 11522
rect 19306 11502 19312 11519
rect 19738 11502 19744 11519
rect 19306 11499 19744 11502
rect 51 11494 499 11499
rect 19301 11494 19749 11499
rect 51 11440 500 11494
rect 51 11110 110 11440
rect 440 11110 500 11440
rect 51 11056 500 11110
rect 19200 11488 19222 11494
rect 19200 11062 19202 11488
rect 19219 11062 19222 11488
rect 19200 11056 19222 11062
rect 19278 11488 19749 11494
rect 19278 11062 19281 11488
rect 19298 11440 19749 11488
rect 19298 11110 19360 11440
rect 19690 11110 19749 11440
rect 19298 11062 19749 11110
rect 19278 11056 19749 11062
rect 51 11051 499 11056
rect 19301 11051 19749 11056
rect 56 11048 494 11051
rect 56 11031 62 11048
rect 488 11031 494 11048
rect 56 11028 494 11031
rect 19306 11048 19744 11051
rect 19306 11031 19312 11048
rect 19738 11031 19744 11048
rect 19306 11028 19744 11031
rect -25 11017 25 11025
rect -25 10983 -17 11017
rect 17 10983 25 11017
rect -25 10975 25 10983
rect 19225 11017 19275 11025
rect 19225 10983 19233 11017
rect 19267 10983 19275 11017
rect 19225 10975 19275 10983
rect 19775 11017 19825 11025
rect 19775 10983 19783 11017
rect 19817 10983 19825 11017
rect 19775 10975 19825 10983
rect 56 10969 494 10972
rect 56 10952 62 10969
rect 488 10952 494 10969
rect 56 10949 494 10952
rect 19306 10969 19744 10972
rect 19306 10952 19312 10969
rect 19738 10952 19744 10969
rect 19306 10949 19744 10952
rect 51 10944 499 10949
rect 19301 10944 19749 10949
rect 51 10890 500 10944
rect 51 10560 110 10890
rect 440 10560 500 10890
rect 51 10506 500 10560
rect 19200 10938 19222 10944
rect 19200 10512 19202 10938
rect 19219 10512 19222 10938
rect 19200 10506 19222 10512
rect 19278 10938 19749 10944
rect 19278 10512 19281 10938
rect 19298 10890 19749 10938
rect 19298 10560 19360 10890
rect 19690 10560 19749 10890
rect 19298 10512 19749 10560
rect 19278 10506 19749 10512
rect 51 10501 499 10506
rect 19301 10501 19749 10506
rect 56 10498 494 10501
rect 56 10481 62 10498
rect 488 10481 494 10498
rect 56 10478 494 10481
rect 19306 10498 19744 10501
rect 19306 10481 19312 10498
rect 19738 10481 19744 10498
rect 19306 10478 19744 10481
rect -25 10467 25 10475
rect -25 10433 -17 10467
rect 17 10433 25 10467
rect -25 10425 25 10433
rect 19225 10467 19275 10475
rect 19225 10433 19233 10467
rect 19267 10433 19275 10467
rect 19225 10425 19275 10433
rect 19775 10467 19825 10475
rect 19775 10433 19783 10467
rect 19817 10433 19825 10467
rect 19775 10425 19825 10433
rect 56 10419 494 10422
rect 56 10402 62 10419
rect 488 10402 494 10419
rect 56 10399 494 10402
rect 19306 10419 19744 10422
rect 19306 10402 19312 10419
rect 19738 10402 19744 10419
rect 19306 10399 19744 10402
rect 51 10394 499 10399
rect 19301 10394 19749 10399
rect 51 10340 500 10394
rect 51 10010 110 10340
rect 440 10010 500 10340
rect 51 9956 500 10010
rect 19200 10388 19222 10394
rect 19200 9962 19202 10388
rect 19219 9962 19222 10388
rect 19200 9956 19222 9962
rect 19278 10388 19749 10394
rect 19278 9962 19281 10388
rect 19298 10340 19749 10388
rect 19298 10010 19360 10340
rect 19690 10010 19749 10340
rect 19298 9962 19749 10010
rect 19278 9956 19749 9962
rect 51 9951 499 9956
rect 19301 9951 19749 9956
rect 56 9948 494 9951
rect 56 9931 62 9948
rect 488 9931 494 9948
rect 56 9928 494 9931
rect 19306 9948 19744 9951
rect 19306 9931 19312 9948
rect 19738 9931 19744 9948
rect 19306 9928 19744 9931
rect -25 9917 25 9925
rect -25 9883 -17 9917
rect 17 9883 25 9917
rect -25 9875 25 9883
rect 19225 9917 19275 9925
rect 19225 9883 19233 9917
rect 19267 9883 19275 9917
rect 19225 9875 19275 9883
rect 19775 9917 19825 9925
rect 19775 9883 19783 9917
rect 19817 9883 19825 9917
rect 19775 9875 19825 9883
rect 56 9869 494 9872
rect 56 9852 62 9869
rect 488 9852 494 9869
rect 56 9849 494 9852
rect 19306 9869 19744 9872
rect 19306 9852 19312 9869
rect 19738 9852 19744 9869
rect 19306 9849 19744 9852
rect 51 9844 499 9849
rect 19301 9844 19749 9849
rect 51 9790 500 9844
rect 51 9460 110 9790
rect 440 9460 500 9790
rect 51 9406 500 9460
rect 19200 9838 19222 9844
rect 19200 9412 19202 9838
rect 19219 9412 19222 9838
rect 19200 9406 19222 9412
rect 19278 9838 19749 9844
rect 19278 9412 19281 9838
rect 19298 9790 19749 9838
rect 19298 9460 19360 9790
rect 19690 9460 19749 9790
rect 19298 9412 19749 9460
rect 19278 9406 19749 9412
rect 51 9401 499 9406
rect 19301 9401 19749 9406
rect 56 9398 494 9401
rect 56 9381 62 9398
rect 488 9381 494 9398
rect 56 9378 494 9381
rect 19306 9398 19744 9401
rect 19306 9381 19312 9398
rect 19738 9381 19744 9398
rect 19306 9378 19744 9381
rect -25 9367 25 9375
rect -25 9333 -17 9367
rect 17 9333 25 9367
rect -25 9325 25 9333
rect 19225 9367 19275 9375
rect 19225 9333 19233 9367
rect 19267 9333 19275 9367
rect 19225 9325 19275 9333
rect 19775 9367 19825 9375
rect 19775 9333 19783 9367
rect 19817 9333 19825 9367
rect 19775 9325 19825 9333
rect 56 9319 494 9322
rect 56 9302 62 9319
rect 488 9302 494 9319
rect 56 9299 494 9302
rect 19306 9319 19744 9322
rect 19306 9302 19312 9319
rect 19738 9302 19744 9319
rect 19306 9299 19744 9302
rect 51 9294 499 9299
rect 19301 9294 19749 9299
rect 51 9240 500 9294
rect 51 8910 110 9240
rect 440 8910 500 9240
rect 51 8856 500 8910
rect 19200 9288 19222 9294
rect 19200 8862 19202 9288
rect 19219 8862 19222 9288
rect 19200 8856 19222 8862
rect 19278 9288 19749 9294
rect 19278 8862 19281 9288
rect 19298 9240 19749 9288
rect 19298 8910 19360 9240
rect 19690 8910 19749 9240
rect 19298 8862 19749 8910
rect 19278 8856 19749 8862
rect 51 8851 499 8856
rect 19301 8851 19749 8856
rect 56 8848 494 8851
rect 56 8831 62 8848
rect 488 8831 494 8848
rect 56 8828 494 8831
rect 19306 8848 19744 8851
rect 19306 8831 19312 8848
rect 19738 8831 19744 8848
rect 19306 8828 19744 8831
rect -25 8817 25 8825
rect -25 8783 -17 8817
rect 17 8783 25 8817
rect -25 8775 25 8783
rect 19225 8817 19275 8825
rect 19225 8783 19233 8817
rect 19267 8783 19275 8817
rect 19225 8775 19275 8783
rect 19775 8817 19825 8825
rect 19775 8783 19783 8817
rect 19817 8783 19825 8817
rect 19775 8775 19825 8783
rect 56 8769 494 8772
rect 56 8752 62 8769
rect 488 8752 494 8769
rect 56 8749 494 8752
rect 19306 8769 19744 8772
rect 19306 8752 19312 8769
rect 19738 8752 19744 8769
rect 19306 8749 19744 8752
rect 51 8744 499 8749
rect 19301 8744 19749 8749
rect 51 8690 500 8744
rect 51 8360 110 8690
rect 440 8360 500 8690
rect 51 8306 500 8360
rect 19200 8738 19222 8744
rect 19200 8312 19202 8738
rect 19219 8312 19222 8738
rect 19200 8306 19222 8312
rect 19278 8738 19749 8744
rect 19278 8312 19281 8738
rect 19298 8690 19749 8738
rect 19298 8360 19360 8690
rect 19690 8360 19749 8690
rect 19298 8312 19749 8360
rect 19278 8306 19749 8312
rect 51 8301 499 8306
rect 19301 8301 19749 8306
rect 56 8298 494 8301
rect 56 8281 62 8298
rect 488 8281 494 8298
rect 56 8278 494 8281
rect 19306 8298 19744 8301
rect 19306 8281 19312 8298
rect 19738 8281 19744 8298
rect 19306 8278 19744 8281
rect -25 8267 25 8275
rect -25 8233 -17 8267
rect 17 8233 25 8267
rect -25 8225 25 8233
rect 19225 8267 19275 8275
rect 19225 8233 19233 8267
rect 19267 8233 19275 8267
rect 19225 8225 19275 8233
rect 19775 8267 19825 8275
rect 19775 8233 19783 8267
rect 19817 8233 19825 8267
rect 19775 8225 19825 8233
rect 56 8219 494 8222
rect 56 8202 62 8219
rect 488 8202 494 8219
rect 56 8199 494 8202
rect 19306 8219 19744 8222
rect 19306 8202 19312 8219
rect 19738 8202 19744 8219
rect 19306 8199 19744 8202
rect 51 8194 499 8199
rect 19301 8194 19749 8199
rect 51 8140 500 8194
rect 51 7810 110 8140
rect 440 7810 500 8140
rect 51 7756 500 7810
rect 19200 8188 19222 8194
rect 19200 7762 19202 8188
rect 19219 7762 19222 8188
rect 19200 7756 19222 7762
rect 19278 8188 19749 8194
rect 19278 7762 19281 8188
rect 19298 8140 19749 8188
rect 19298 7810 19360 8140
rect 19690 7810 19749 8140
rect 19298 7762 19749 7810
rect 19278 7756 19749 7762
rect 51 7751 499 7756
rect 19301 7751 19749 7756
rect 56 7748 494 7751
rect 56 7731 62 7748
rect 488 7731 494 7748
rect 56 7728 494 7731
rect 19306 7748 19744 7751
rect 19306 7731 19312 7748
rect 19738 7731 19744 7748
rect 19306 7728 19744 7731
rect -25 7717 25 7725
rect -25 7683 -17 7717
rect 17 7683 25 7717
rect -25 7675 25 7683
rect 19225 7717 19275 7725
rect 19225 7683 19233 7717
rect 19267 7683 19275 7717
rect 19225 7675 19275 7683
rect 19775 7717 19825 7725
rect 19775 7683 19783 7717
rect 19817 7683 19825 7717
rect 19775 7675 19825 7683
rect 56 7669 494 7672
rect 56 7652 62 7669
rect 488 7652 494 7669
rect 56 7649 494 7652
rect 19306 7669 19744 7672
rect 19306 7652 19312 7669
rect 19738 7652 19744 7669
rect 19306 7649 19744 7652
rect 51 7644 499 7649
rect 19301 7644 19749 7649
rect 51 7590 500 7644
rect 51 7260 110 7590
rect 440 7260 500 7590
rect 51 7206 500 7260
rect 19200 7638 19222 7644
rect 19200 7212 19202 7638
rect 19219 7212 19222 7638
rect 19200 7206 19222 7212
rect 19278 7638 19749 7644
rect 19278 7212 19281 7638
rect 19298 7590 19749 7638
rect 19298 7260 19360 7590
rect 19690 7260 19749 7590
rect 19298 7212 19749 7260
rect 19278 7206 19749 7212
rect 51 7201 499 7206
rect 19301 7201 19749 7206
rect 56 7198 494 7201
rect 56 7181 62 7198
rect 488 7181 494 7198
rect 56 7178 494 7181
rect 19306 7198 19744 7201
rect 19306 7181 19312 7198
rect 19738 7181 19744 7198
rect 19306 7178 19744 7181
rect -25 7167 25 7175
rect -25 7133 -17 7167
rect 17 7133 25 7167
rect -25 7125 25 7133
rect 19225 7167 19275 7175
rect 19225 7133 19233 7167
rect 19267 7133 19275 7167
rect 19225 7125 19275 7133
rect 19775 7167 19825 7175
rect 19775 7133 19783 7167
rect 19817 7133 19825 7167
rect 19775 7125 19825 7133
rect 56 7119 494 7122
rect 56 7102 62 7119
rect 488 7102 494 7119
rect 56 7099 494 7102
rect 19306 7119 19744 7122
rect 19306 7102 19312 7119
rect 19738 7102 19744 7119
rect 19306 7099 19744 7102
rect 51 7094 499 7099
rect 19301 7094 19749 7099
rect 51 7040 500 7094
rect 51 6710 110 7040
rect 440 6710 500 7040
rect 51 6656 500 6710
rect 19200 7088 19222 7094
rect 19200 6662 19202 7088
rect 19219 6662 19222 7088
rect 19200 6656 19222 6662
rect 19278 7088 19749 7094
rect 19278 6662 19281 7088
rect 19298 7040 19749 7088
rect 19298 6710 19360 7040
rect 19690 6710 19749 7040
rect 19298 6662 19749 6710
rect 19278 6656 19749 6662
rect 51 6651 499 6656
rect 19301 6651 19749 6656
rect 56 6648 494 6651
rect 56 6631 62 6648
rect 488 6631 494 6648
rect 56 6628 494 6631
rect 19306 6648 19744 6651
rect 19306 6631 19312 6648
rect 19738 6631 19744 6648
rect 19306 6628 19744 6631
rect -25 6617 25 6625
rect -25 6583 -17 6617
rect 17 6583 25 6617
rect -25 6575 25 6583
rect 19225 6617 19275 6625
rect 19225 6583 19233 6617
rect 19267 6583 19275 6617
rect 19225 6575 19275 6583
rect 19775 6617 19825 6625
rect 19775 6583 19783 6617
rect 19817 6583 19825 6617
rect 19775 6575 19825 6583
rect 56 6569 494 6572
rect 56 6552 62 6569
rect 488 6552 494 6569
rect 56 6549 494 6552
rect 19306 6569 19744 6572
rect 19306 6552 19312 6569
rect 19738 6552 19744 6569
rect 19306 6549 19744 6552
rect 51 6544 499 6549
rect 19301 6544 19749 6549
rect 51 6490 500 6544
rect 51 6160 110 6490
rect 440 6160 500 6490
rect 51 6106 500 6160
rect 19200 6538 19222 6544
rect 19200 6112 19202 6538
rect 19219 6112 19222 6538
rect 19200 6106 19222 6112
rect 19278 6538 19749 6544
rect 19278 6112 19281 6538
rect 19298 6490 19749 6538
rect 19298 6160 19360 6490
rect 19690 6160 19749 6490
rect 19298 6112 19749 6160
rect 19278 6106 19749 6112
rect 51 6101 499 6106
rect 19301 6101 19749 6106
rect 56 6098 494 6101
rect 56 6081 62 6098
rect 488 6081 494 6098
rect 56 6078 494 6081
rect 19306 6098 19744 6101
rect 19306 6081 19312 6098
rect 19738 6081 19744 6098
rect 19306 6078 19744 6081
rect -25 6067 25 6075
rect -25 6033 -17 6067
rect 17 6033 25 6067
rect -25 6025 25 6033
rect 19225 6067 19275 6075
rect 19225 6033 19233 6067
rect 19267 6033 19275 6067
rect 19225 6025 19275 6033
rect 19775 6067 19825 6075
rect 19775 6033 19783 6067
rect 19817 6033 19825 6067
rect 19775 6025 19825 6033
rect 56 6019 494 6022
rect 56 6002 62 6019
rect 488 6002 494 6019
rect 56 5999 494 6002
rect 19306 6019 19744 6022
rect 19306 6002 19312 6019
rect 19738 6002 19744 6019
rect 19306 5999 19744 6002
rect 51 5994 499 5999
rect 19301 5994 19749 5999
rect 51 5940 500 5994
rect 51 5610 110 5940
rect 440 5610 500 5940
rect 51 5556 500 5610
rect 19200 5988 19222 5994
rect 19200 5562 19202 5988
rect 19219 5562 19222 5988
rect 19200 5556 19222 5562
rect 19278 5988 19749 5994
rect 19278 5562 19281 5988
rect 19298 5940 19749 5988
rect 19298 5610 19360 5940
rect 19690 5610 19749 5940
rect 19298 5562 19749 5610
rect 19278 5556 19749 5562
rect 51 5551 499 5556
rect 19301 5551 19749 5556
rect 56 5548 494 5551
rect 56 5531 62 5548
rect 488 5531 494 5548
rect 56 5528 494 5531
rect 19306 5548 19744 5551
rect 19306 5531 19312 5548
rect 19738 5531 19744 5548
rect 19306 5528 19744 5531
rect -25 5517 25 5525
rect -25 5483 -17 5517
rect 17 5483 25 5517
rect -25 5475 25 5483
rect 19225 5517 19275 5525
rect 19225 5483 19233 5517
rect 19267 5483 19275 5517
rect 19225 5475 19275 5483
rect 19775 5517 19825 5525
rect 19775 5483 19783 5517
rect 19817 5483 19825 5517
rect 19775 5475 19825 5483
rect 56 5469 494 5472
rect 56 5452 62 5469
rect 488 5452 494 5469
rect 56 5449 494 5452
rect 19306 5469 19744 5472
rect 19306 5452 19312 5469
rect 19738 5452 19744 5469
rect 19306 5449 19744 5452
rect 51 5444 499 5449
rect 19301 5444 19749 5449
rect 51 5390 500 5444
rect 51 5060 110 5390
rect 440 5060 500 5390
rect 51 5006 500 5060
rect 19200 5438 19222 5444
rect 19200 5012 19202 5438
rect 19219 5012 19222 5438
rect 19200 5006 19222 5012
rect 19278 5438 19749 5444
rect 19278 5012 19281 5438
rect 19298 5390 19749 5438
rect 19298 5060 19360 5390
rect 19690 5060 19749 5390
rect 19298 5012 19749 5060
rect 19278 5006 19749 5012
rect 51 5001 499 5006
rect 19301 5001 19749 5006
rect 56 4998 494 5001
rect 56 4981 62 4998
rect 488 4981 494 4998
rect 56 4978 494 4981
rect 19306 4998 19744 5001
rect 19306 4981 19312 4998
rect 19738 4981 19744 4998
rect 19306 4978 19744 4981
rect -25 4967 25 4975
rect -25 4933 -17 4967
rect 17 4933 25 4967
rect -25 4925 25 4933
rect 19225 4967 19275 4975
rect 19225 4933 19233 4967
rect 19267 4933 19275 4967
rect 19225 4925 19275 4933
rect 19775 4967 19825 4975
rect 19775 4933 19783 4967
rect 19817 4933 19825 4967
rect 19775 4925 19825 4933
rect 56 4919 494 4922
rect 56 4902 62 4919
rect 488 4902 494 4919
rect 56 4899 494 4902
rect 19306 4919 19744 4922
rect 19306 4902 19312 4919
rect 19738 4902 19744 4919
rect 19306 4899 19744 4902
rect 51 4894 499 4899
rect 19301 4894 19749 4899
rect 51 4840 500 4894
rect 51 4510 110 4840
rect 440 4510 500 4840
rect 51 4456 500 4510
rect 19200 4888 19222 4894
rect 19200 4462 19202 4888
rect 19219 4462 19222 4888
rect 19200 4456 19222 4462
rect 19278 4888 19749 4894
rect 19278 4462 19281 4888
rect 19298 4840 19749 4888
rect 19298 4510 19360 4840
rect 19690 4510 19749 4840
rect 19298 4462 19749 4510
rect 19278 4456 19749 4462
rect 51 4451 499 4456
rect 19301 4451 19749 4456
rect 56 4448 494 4451
rect 56 4431 62 4448
rect 488 4431 494 4448
rect 56 4428 494 4431
rect 19306 4448 19744 4451
rect 19306 4431 19312 4448
rect 19738 4431 19744 4448
rect 19306 4428 19744 4431
rect -25 4417 25 4425
rect -25 4383 -17 4417
rect 17 4383 25 4417
rect -25 4375 25 4383
rect 19225 4417 19275 4425
rect 19225 4383 19233 4417
rect 19267 4383 19275 4417
rect 19225 4375 19275 4383
rect 19775 4417 19825 4425
rect 19775 4383 19783 4417
rect 19817 4383 19825 4417
rect 19775 4375 19825 4383
rect 56 4369 494 4372
rect 56 4352 62 4369
rect 488 4352 494 4369
rect 56 4349 494 4352
rect 19306 4369 19744 4372
rect 19306 4352 19312 4369
rect 19738 4352 19744 4369
rect 19306 4349 19744 4352
rect 51 4344 499 4349
rect 19301 4344 19749 4349
rect 51 4290 500 4344
rect 51 3960 110 4290
rect 440 3960 500 4290
rect 51 3906 500 3960
rect 19200 4338 19222 4344
rect 19200 3912 19202 4338
rect 19219 3912 19222 4338
rect 19200 3906 19222 3912
rect 19278 4338 19749 4344
rect 19278 3912 19281 4338
rect 19298 4290 19749 4338
rect 19298 3960 19360 4290
rect 19690 3960 19749 4290
rect 19298 3912 19749 3960
rect 19278 3906 19749 3912
rect 51 3901 499 3906
rect 19301 3901 19749 3906
rect 56 3898 494 3901
rect 56 3881 62 3898
rect 488 3881 494 3898
rect 56 3878 494 3881
rect 19306 3898 19744 3901
rect 19306 3881 19312 3898
rect 19738 3881 19744 3898
rect 19306 3878 19744 3881
rect -25 3867 25 3875
rect -25 3833 -17 3867
rect 17 3833 25 3867
rect -25 3825 25 3833
rect 19225 3867 19275 3875
rect 19225 3833 19233 3867
rect 19267 3833 19275 3867
rect 19225 3825 19275 3833
rect 19775 3867 19825 3875
rect 19775 3833 19783 3867
rect 19817 3833 19825 3867
rect 19775 3825 19825 3833
rect 56 3819 494 3822
rect 56 3802 62 3819
rect 488 3802 494 3819
rect 56 3799 494 3802
rect 19306 3819 19744 3822
rect 19306 3802 19312 3819
rect 19738 3802 19744 3819
rect 19306 3799 19744 3802
rect 51 3794 499 3799
rect 19301 3794 19749 3799
rect 51 3740 500 3794
rect 51 3410 110 3740
rect 440 3410 500 3740
rect 51 3356 500 3410
rect 19200 3788 19222 3794
rect 19200 3362 19202 3788
rect 19219 3362 19222 3788
rect 19200 3356 19222 3362
rect 19278 3788 19749 3794
rect 19278 3362 19281 3788
rect 19298 3740 19749 3788
rect 19298 3410 19360 3740
rect 19690 3410 19749 3740
rect 19298 3362 19749 3410
rect 19278 3356 19749 3362
rect 51 3351 499 3356
rect 19301 3351 19749 3356
rect 56 3348 494 3351
rect 56 3331 62 3348
rect 488 3331 494 3348
rect 56 3328 494 3331
rect 19306 3348 19744 3351
rect 19306 3331 19312 3348
rect 19738 3331 19744 3348
rect 19306 3328 19744 3331
rect -25 3317 25 3325
rect -25 3283 -17 3317
rect 17 3283 25 3317
rect -25 3275 25 3283
rect 19225 3317 19275 3325
rect 19225 3283 19233 3317
rect 19267 3283 19275 3317
rect 19225 3275 19275 3283
rect 19775 3317 19825 3325
rect 19775 3283 19783 3317
rect 19817 3283 19825 3317
rect 19775 3275 19825 3283
rect 56 3269 494 3272
rect 56 3252 62 3269
rect 488 3252 494 3269
rect 56 3249 494 3252
rect 19306 3269 19744 3272
rect 19306 3252 19312 3269
rect 19738 3252 19744 3269
rect 19306 3249 19744 3252
rect 51 3244 499 3249
rect 19301 3244 19749 3249
rect 51 3190 500 3244
rect 51 2860 110 3190
rect 440 2860 500 3190
rect 51 2806 500 2860
rect 19200 3238 19222 3244
rect 19200 2812 19202 3238
rect 19219 2812 19222 3238
rect 19200 2806 19222 2812
rect 19278 3238 19749 3244
rect 19278 2812 19281 3238
rect 19298 3190 19749 3238
rect 19298 2860 19360 3190
rect 19690 2860 19749 3190
rect 19298 2812 19749 2860
rect 19278 2806 19749 2812
rect 51 2801 499 2806
rect 19301 2801 19749 2806
rect 56 2798 494 2801
rect 56 2781 62 2798
rect 488 2781 494 2798
rect 56 2778 494 2781
rect 19306 2798 19744 2801
rect 19306 2781 19312 2798
rect 19738 2781 19744 2798
rect 19306 2778 19744 2781
rect -25 2767 25 2775
rect -25 2733 -17 2767
rect 17 2733 25 2767
rect -25 2725 25 2733
rect 19225 2767 19275 2775
rect 19225 2733 19233 2767
rect 19267 2733 19275 2767
rect 19225 2725 19275 2733
rect 19775 2767 19825 2775
rect 19775 2733 19783 2767
rect 19817 2733 19825 2767
rect 19775 2725 19825 2733
rect 56 2719 494 2722
rect 56 2702 62 2719
rect 488 2702 494 2719
rect 56 2699 494 2702
rect 19306 2719 19744 2722
rect 19306 2702 19312 2719
rect 19738 2702 19744 2719
rect 19306 2699 19744 2702
rect 51 2694 499 2699
rect 19301 2694 19749 2699
rect 51 2640 500 2694
rect 51 2310 110 2640
rect 440 2310 500 2640
rect 51 2256 500 2310
rect 19200 2688 19222 2694
rect 19200 2262 19202 2688
rect 19219 2262 19222 2688
rect 19200 2256 19222 2262
rect 19278 2688 19749 2694
rect 19278 2262 19281 2688
rect 19298 2640 19749 2688
rect 19298 2310 19360 2640
rect 19690 2310 19749 2640
rect 19298 2262 19749 2310
rect 19278 2256 19749 2262
rect 51 2251 499 2256
rect 19301 2251 19749 2256
rect 56 2248 494 2251
rect 56 2231 62 2248
rect 488 2231 494 2248
rect 56 2228 494 2231
rect 19306 2248 19744 2251
rect 19306 2231 19312 2248
rect 19738 2231 19744 2248
rect 19306 2228 19744 2231
rect -25 2217 25 2225
rect -25 2183 -17 2217
rect 17 2183 25 2217
rect -25 2175 25 2183
rect 19225 2217 19275 2225
rect 19225 2183 19233 2217
rect 19267 2183 19275 2217
rect 19225 2175 19275 2183
rect 19775 2217 19825 2225
rect 19775 2183 19783 2217
rect 19817 2183 19825 2217
rect 19775 2175 19825 2183
rect 56 2169 494 2172
rect 56 2152 62 2169
rect 488 2152 494 2169
rect 56 2149 494 2152
rect 19306 2169 19744 2172
rect 19306 2152 19312 2169
rect 19738 2152 19744 2169
rect 19306 2149 19744 2152
rect 51 2144 499 2149
rect 19301 2144 19749 2149
rect 51 2090 500 2144
rect 51 1760 110 2090
rect 440 1760 500 2090
rect 51 1706 500 1760
rect 19200 2138 19222 2144
rect 19200 1712 19202 2138
rect 19219 1712 19222 2138
rect 19200 1706 19222 1712
rect 19278 2138 19749 2144
rect 19278 1712 19281 2138
rect 19298 2090 19749 2138
rect 19298 1760 19360 2090
rect 19690 1760 19749 2090
rect 19298 1712 19749 1760
rect 19278 1706 19749 1712
rect 51 1701 499 1706
rect 19301 1701 19749 1706
rect 56 1698 494 1701
rect 56 1681 62 1698
rect 488 1681 494 1698
rect 56 1678 494 1681
rect 19306 1698 19744 1701
rect 19306 1681 19312 1698
rect 19738 1681 19744 1698
rect 19306 1678 19744 1681
rect -25 1667 25 1675
rect -25 1633 -17 1667
rect 17 1633 25 1667
rect -25 1625 25 1633
rect 19225 1667 19275 1675
rect 19225 1633 19233 1667
rect 19267 1633 19275 1667
rect 19225 1625 19275 1633
rect 19775 1667 19825 1675
rect 19775 1633 19783 1667
rect 19817 1633 19825 1667
rect 19775 1625 19825 1633
rect 56 1619 494 1622
rect 56 1602 62 1619
rect 488 1602 494 1619
rect 56 1599 494 1602
rect 19306 1619 19744 1622
rect 19306 1602 19312 1619
rect 19738 1602 19744 1619
rect 19306 1599 19744 1602
rect 51 1594 499 1599
rect 19301 1594 19749 1599
rect 51 1540 500 1594
rect 51 1210 110 1540
rect 440 1210 500 1540
rect 51 1156 500 1210
rect 19200 1588 19222 1594
rect 19200 1162 19202 1588
rect 19219 1162 19222 1588
rect 19200 1156 19222 1162
rect 19278 1588 19749 1594
rect 19278 1162 19281 1588
rect 19298 1540 19749 1588
rect 19298 1210 19360 1540
rect 19690 1210 19749 1540
rect 19298 1162 19749 1210
rect 19278 1156 19749 1162
rect 51 1151 499 1156
rect 19301 1151 19749 1156
rect 56 1148 494 1151
rect 56 1131 62 1148
rect 488 1131 494 1148
rect 56 1128 494 1131
rect 19306 1148 19744 1151
rect 19306 1131 19312 1148
rect 19738 1131 19744 1148
rect 19306 1128 19744 1131
rect -25 1117 25 1125
rect -25 1083 -17 1117
rect 17 1083 25 1117
rect -25 1075 25 1083
rect 19225 1117 19275 1125
rect 19225 1083 19233 1117
rect 19267 1083 19275 1117
rect 19225 1075 19275 1083
rect 19775 1117 19825 1125
rect 19775 1083 19783 1117
rect 19817 1083 19825 1117
rect 19775 1075 19825 1083
rect 56 1069 494 1072
rect 56 1052 62 1069
rect 488 1052 494 1069
rect 56 1049 494 1052
rect 19306 1069 19744 1072
rect 19306 1052 19312 1069
rect 19738 1052 19744 1069
rect 19306 1049 19744 1052
rect 51 1044 499 1049
rect 19301 1044 19749 1049
rect 51 990 500 1044
rect 51 660 110 990
rect 440 660 500 990
rect 51 606 500 660
rect 19200 1038 19222 1044
rect 19200 612 19202 1038
rect 19219 612 19222 1038
rect 19200 606 19222 612
rect 19278 1038 19749 1044
rect 19278 612 19281 1038
rect 19298 990 19749 1038
rect 19298 660 19360 990
rect 19690 660 19749 990
rect 19298 612 19749 660
rect 19278 606 19749 612
rect 51 601 499 606
rect 19301 601 19749 606
rect 56 598 494 601
rect 56 581 62 598
rect 488 581 494 598
rect 56 578 494 581
rect 19306 598 19744 601
rect 19306 581 19312 598
rect 19738 581 19744 598
rect 19306 578 19744 581
rect -25 567 25 575
rect -25 533 -17 567
rect 17 533 25 567
rect -25 525 25 533
rect 19225 567 19275 575
rect 19225 533 19233 567
rect 19267 533 19275 567
rect 19225 525 19275 533
rect 19775 567 19825 575
rect 19775 533 19783 567
rect 19817 533 19825 567
rect 19775 525 19825 533
rect 56 519 494 522
rect 56 502 62 519
rect 488 502 494 519
rect 56 499 494 502
rect 19306 519 19744 522
rect 19306 502 19312 519
rect 19738 502 19744 519
rect 606 499 1044 500
rect 1156 499 1594 500
rect 1706 499 2144 500
rect 2256 499 2694 500
rect 2806 499 3244 500
rect 3356 499 3794 500
rect 3906 499 4344 500
rect 4456 499 4894 500
rect 5006 499 5444 500
rect 5556 499 5994 500
rect 6106 499 6544 500
rect 6656 499 7094 500
rect 7206 499 7644 500
rect 7756 499 8194 500
rect 8306 499 8744 500
rect 8856 499 9294 500
rect 9406 499 9844 500
rect 9956 499 10394 500
rect 10506 499 10944 500
rect 11056 499 11494 500
rect 11606 499 12044 500
rect 12156 499 12594 500
rect 12706 499 13144 500
rect 13256 499 13694 500
rect 13806 499 14244 500
rect 14356 499 14794 500
rect 14906 499 15344 500
rect 15456 499 15894 500
rect 16006 499 16444 500
rect 16556 499 16994 500
rect 17106 499 17544 500
rect 17656 499 18094 500
rect 18206 499 18644 500
rect 18756 499 19194 500
rect 19306 499 19744 502
rect 51 494 499 499
rect 601 494 1049 499
rect 1151 494 1599 499
rect 1701 494 2149 499
rect 2251 494 2699 499
rect 2801 494 3249 499
rect 3351 494 3799 499
rect 3901 494 4349 499
rect 4451 494 4899 499
rect 5001 494 5449 499
rect 5551 494 5999 499
rect 6101 494 6549 499
rect 6651 494 7099 499
rect 7201 494 7649 499
rect 7751 494 8199 499
rect 8301 494 8749 499
rect 8851 494 9299 499
rect 9401 494 9849 499
rect 9951 494 10399 499
rect 10501 494 10949 499
rect 11051 494 11499 499
rect 11601 494 12049 499
rect 12151 494 12599 499
rect 12701 494 13149 499
rect 13251 494 13699 499
rect 13801 494 14249 499
rect 14351 494 14799 499
rect 14901 494 15349 499
rect 15451 494 15899 499
rect 16001 494 16449 499
rect 16551 494 16999 499
rect 17101 494 17549 499
rect 17651 494 18099 499
rect 18201 494 18649 499
rect 18751 494 19199 499
rect 19301 494 19749 499
rect 51 488 522 494
rect 51 440 502 488
rect 51 110 110 440
rect 440 110 502 440
rect 51 62 502 110
rect 519 62 522 488
rect 51 56 522 62
rect 578 488 1072 494
rect 578 62 581 488
rect 598 440 1052 488
rect 598 110 660 440
rect 990 110 1052 440
rect 598 62 1052 110
rect 1069 62 1072 488
rect 578 56 1072 62
rect 1128 488 1622 494
rect 1128 62 1131 488
rect 1148 440 1602 488
rect 1148 110 1210 440
rect 1540 110 1602 440
rect 1148 62 1602 110
rect 1619 62 1622 488
rect 1128 56 1622 62
rect 1678 488 2172 494
rect 1678 62 1681 488
rect 1698 440 2152 488
rect 1698 110 1760 440
rect 2090 110 2152 440
rect 1698 62 2152 110
rect 2169 62 2172 488
rect 1678 56 2172 62
rect 2228 488 2722 494
rect 2228 62 2231 488
rect 2248 440 2702 488
rect 2248 110 2310 440
rect 2640 110 2702 440
rect 2248 62 2702 110
rect 2719 62 2722 488
rect 2228 56 2722 62
rect 2778 488 3272 494
rect 2778 62 2781 488
rect 2798 440 3252 488
rect 2798 110 2860 440
rect 3190 110 3252 440
rect 2798 62 3252 110
rect 3269 62 3272 488
rect 2778 56 3272 62
rect 3328 488 3822 494
rect 3328 62 3331 488
rect 3348 440 3802 488
rect 3348 110 3410 440
rect 3740 110 3802 440
rect 3348 62 3802 110
rect 3819 62 3822 488
rect 3328 56 3822 62
rect 3878 488 4372 494
rect 3878 62 3881 488
rect 3898 440 4352 488
rect 3898 110 3960 440
rect 4290 110 4352 440
rect 3898 62 4352 110
rect 4369 62 4372 488
rect 3878 56 4372 62
rect 4428 488 4922 494
rect 4428 62 4431 488
rect 4448 440 4902 488
rect 4448 110 4510 440
rect 4840 110 4902 440
rect 4448 62 4902 110
rect 4919 62 4922 488
rect 4428 56 4922 62
rect 4978 488 5472 494
rect 4978 62 4981 488
rect 4998 440 5452 488
rect 4998 110 5060 440
rect 5390 110 5452 440
rect 4998 62 5452 110
rect 5469 62 5472 488
rect 4978 56 5472 62
rect 5528 488 6022 494
rect 5528 62 5531 488
rect 5548 440 6002 488
rect 5548 110 5610 440
rect 5940 110 6002 440
rect 5548 62 6002 110
rect 6019 62 6022 488
rect 5528 56 6022 62
rect 6078 488 6572 494
rect 6078 62 6081 488
rect 6098 440 6552 488
rect 6098 110 6160 440
rect 6490 110 6552 440
rect 6098 62 6552 110
rect 6569 62 6572 488
rect 6078 56 6572 62
rect 6628 488 7122 494
rect 6628 62 6631 488
rect 6648 440 7102 488
rect 6648 110 6710 440
rect 7040 110 7102 440
rect 6648 62 7102 110
rect 7119 62 7122 488
rect 6628 56 7122 62
rect 7178 488 7672 494
rect 7178 62 7181 488
rect 7198 440 7652 488
rect 7198 110 7260 440
rect 7590 110 7652 440
rect 7198 62 7652 110
rect 7669 62 7672 488
rect 7178 56 7672 62
rect 7728 488 8222 494
rect 7728 62 7731 488
rect 7748 440 8202 488
rect 7748 110 7810 440
rect 8140 110 8202 440
rect 7748 62 8202 110
rect 8219 62 8222 488
rect 7728 56 8222 62
rect 8278 488 8772 494
rect 8278 62 8281 488
rect 8298 440 8752 488
rect 8298 110 8360 440
rect 8690 110 8752 440
rect 8298 62 8752 110
rect 8769 62 8772 488
rect 8278 56 8772 62
rect 8828 488 9322 494
rect 8828 62 8831 488
rect 8848 440 9302 488
rect 8848 110 8910 440
rect 9240 110 9302 440
rect 8848 62 9302 110
rect 9319 62 9322 488
rect 8828 56 9322 62
rect 9378 488 9872 494
rect 9378 62 9381 488
rect 9398 440 9852 488
rect 9398 110 9460 440
rect 9790 110 9852 440
rect 9398 62 9852 110
rect 9869 62 9872 488
rect 9378 56 9872 62
rect 9928 488 10422 494
rect 9928 62 9931 488
rect 9948 440 10402 488
rect 9948 110 10010 440
rect 10340 110 10402 440
rect 9948 62 10402 110
rect 10419 62 10422 488
rect 9928 56 10422 62
rect 10478 488 10972 494
rect 10478 62 10481 488
rect 10498 440 10952 488
rect 10498 110 10560 440
rect 10890 110 10952 440
rect 10498 62 10952 110
rect 10969 62 10972 488
rect 10478 56 10972 62
rect 11028 488 11522 494
rect 11028 62 11031 488
rect 11048 440 11502 488
rect 11048 110 11110 440
rect 11440 110 11502 440
rect 11048 62 11502 110
rect 11519 62 11522 488
rect 11028 56 11522 62
rect 11578 488 12072 494
rect 11578 62 11581 488
rect 11598 440 12052 488
rect 11598 110 11660 440
rect 11990 110 12052 440
rect 11598 62 12052 110
rect 12069 62 12072 488
rect 11578 56 12072 62
rect 12128 488 12622 494
rect 12128 62 12131 488
rect 12148 440 12602 488
rect 12148 110 12210 440
rect 12540 110 12602 440
rect 12148 62 12602 110
rect 12619 62 12622 488
rect 12128 56 12622 62
rect 12678 488 13172 494
rect 12678 62 12681 488
rect 12698 440 13152 488
rect 12698 110 12760 440
rect 13090 110 13152 440
rect 12698 62 13152 110
rect 13169 62 13172 488
rect 12678 56 13172 62
rect 13228 488 13722 494
rect 13228 62 13231 488
rect 13248 440 13702 488
rect 13248 110 13310 440
rect 13640 110 13702 440
rect 13248 62 13702 110
rect 13719 62 13722 488
rect 13228 56 13722 62
rect 13778 488 14272 494
rect 13778 62 13781 488
rect 13798 440 14252 488
rect 13798 110 13860 440
rect 14190 110 14252 440
rect 13798 62 14252 110
rect 14269 62 14272 488
rect 13778 56 14272 62
rect 14328 488 14822 494
rect 14328 62 14331 488
rect 14348 440 14802 488
rect 14348 110 14410 440
rect 14740 110 14802 440
rect 14348 62 14802 110
rect 14819 62 14822 488
rect 14328 56 14822 62
rect 14878 488 15372 494
rect 14878 62 14881 488
rect 14898 440 15352 488
rect 14898 110 14960 440
rect 15290 110 15352 440
rect 14898 62 15352 110
rect 15369 62 15372 488
rect 14878 56 15372 62
rect 15428 488 15922 494
rect 15428 62 15431 488
rect 15448 440 15902 488
rect 15448 110 15510 440
rect 15840 110 15902 440
rect 15448 62 15902 110
rect 15919 62 15922 488
rect 15428 56 15922 62
rect 15978 488 16472 494
rect 15978 62 15981 488
rect 15998 440 16452 488
rect 15998 110 16060 440
rect 16390 110 16452 440
rect 15998 62 16452 110
rect 16469 62 16472 488
rect 15978 56 16472 62
rect 16528 488 17022 494
rect 16528 62 16531 488
rect 16548 440 17002 488
rect 16548 110 16610 440
rect 16940 110 17002 440
rect 16548 62 17002 110
rect 17019 62 17022 488
rect 16528 56 17022 62
rect 17078 488 17572 494
rect 17078 62 17081 488
rect 17098 440 17552 488
rect 17098 110 17160 440
rect 17490 110 17552 440
rect 17098 62 17552 110
rect 17569 62 17572 488
rect 17078 56 17572 62
rect 17628 488 18122 494
rect 17628 62 17631 488
rect 17648 440 18102 488
rect 17648 110 17710 440
rect 18040 110 18102 440
rect 17648 62 18102 110
rect 18119 62 18122 488
rect 17628 56 18122 62
rect 18178 488 18672 494
rect 18178 62 18181 488
rect 18198 440 18652 488
rect 18198 110 18260 440
rect 18590 110 18652 440
rect 18198 62 18652 110
rect 18669 62 18672 488
rect 18178 56 18672 62
rect 18728 488 19222 494
rect 18728 62 18731 488
rect 18748 440 19202 488
rect 18748 110 18810 440
rect 19140 110 19202 440
rect 18748 62 19202 110
rect 19219 62 19222 488
rect 18728 56 19222 62
rect 19278 488 19749 494
rect 19278 62 19281 488
rect 19298 440 19749 488
rect 19298 110 19360 440
rect 19690 110 19749 440
rect 19298 62 19749 110
rect 19278 56 19749 62
rect 51 51 499 56
rect 601 51 1049 56
rect 1151 51 1599 56
rect 1701 51 2149 56
rect 2251 51 2699 56
rect 2801 51 3249 56
rect 3351 51 3799 56
rect 3901 51 4349 56
rect 4451 51 4899 56
rect 5001 51 5449 56
rect 5551 51 5999 56
rect 6101 51 6549 56
rect 6651 51 7099 56
rect 7201 51 7649 56
rect 7751 51 8199 56
rect 8301 51 8749 56
rect 8851 51 9299 56
rect 9401 51 9849 56
rect 9951 51 10399 56
rect 10501 51 10949 56
rect 11051 51 11499 56
rect 11601 51 12049 56
rect 12151 51 12599 56
rect 12701 51 13149 56
rect 13251 51 13699 56
rect 13801 51 14249 56
rect 14351 51 14799 56
rect 14901 51 15349 56
rect 15451 51 15899 56
rect 16001 51 16449 56
rect 16551 51 16999 56
rect 17101 51 17549 56
rect 17651 51 18099 56
rect 18201 51 18649 56
rect 18751 51 19199 56
rect 19301 51 19749 56
rect -25 17 25 25
rect -25 -17 -17 17
rect 17 -17 25 17
rect -25 -25 25 -17
rect 525 17 575 25
rect 525 -17 533 17
rect 567 -17 575 17
rect 525 -25 575 -17
rect 1075 17 1125 25
rect 1075 -17 1083 17
rect 1117 -17 1125 17
rect 1075 -25 1125 -17
rect 1625 17 1675 25
rect 1625 -17 1633 17
rect 1667 -17 1675 17
rect 1625 -25 1675 -17
rect 2175 17 2225 25
rect 2175 -17 2183 17
rect 2217 -17 2225 17
rect 2175 -25 2225 -17
rect 2725 17 2775 25
rect 2725 -17 2733 17
rect 2767 -17 2775 17
rect 2725 -25 2775 -17
rect 3275 17 3325 25
rect 3275 -17 3283 17
rect 3317 -17 3325 17
rect 3275 -25 3325 -17
rect 3825 17 3875 25
rect 3825 -17 3833 17
rect 3867 -17 3875 17
rect 3825 -25 3875 -17
rect 4375 17 4425 25
rect 4375 -17 4383 17
rect 4417 -17 4425 17
rect 4375 -25 4425 -17
rect 4925 17 4975 25
rect 4925 -17 4933 17
rect 4967 -17 4975 17
rect 4925 -25 4975 -17
rect 5475 17 5525 25
rect 5475 -17 5483 17
rect 5517 -17 5525 17
rect 5475 -25 5525 -17
rect 6025 17 6075 25
rect 6025 -17 6033 17
rect 6067 -17 6075 17
rect 6025 -25 6075 -17
rect 6575 17 6625 25
rect 6575 -17 6583 17
rect 6617 -17 6625 17
rect 6575 -25 6625 -17
rect 7125 17 7175 25
rect 7125 -17 7133 17
rect 7167 -17 7175 17
rect 7125 -25 7175 -17
rect 7675 17 7725 25
rect 7675 -17 7683 17
rect 7717 -17 7725 17
rect 7675 -25 7725 -17
rect 8225 17 8275 25
rect 8225 -17 8233 17
rect 8267 -17 8275 17
rect 8225 -25 8275 -17
rect 8775 17 8825 25
rect 8775 -17 8783 17
rect 8817 -17 8825 17
rect 8775 -25 8825 -17
rect 9325 17 9375 25
rect 9325 -17 9333 17
rect 9367 -17 9375 17
rect 9325 -25 9375 -17
rect 9875 17 9925 25
rect 9875 -17 9883 17
rect 9917 -17 9925 17
rect 9875 -25 9925 -17
rect 10425 17 10475 25
rect 10425 -17 10433 17
rect 10467 -17 10475 17
rect 10425 -25 10475 -17
rect 10975 17 11025 25
rect 10975 -17 10983 17
rect 11017 -17 11025 17
rect 10975 -25 11025 -17
rect 11525 17 11575 25
rect 11525 -17 11533 17
rect 11567 -17 11575 17
rect 11525 -25 11575 -17
rect 12075 17 12125 25
rect 12075 -17 12083 17
rect 12117 -17 12125 17
rect 12075 -25 12125 -17
rect 12625 17 12675 25
rect 12625 -17 12633 17
rect 12667 -17 12675 17
rect 12625 -25 12675 -17
rect 13175 17 13225 25
rect 13175 -17 13183 17
rect 13217 -17 13225 17
rect 13175 -25 13225 -17
rect 13725 17 13775 25
rect 13725 -17 13733 17
rect 13767 -17 13775 17
rect 13725 -25 13775 -17
rect 14275 17 14325 25
rect 14275 -17 14283 17
rect 14317 -17 14325 17
rect 14275 -25 14325 -17
rect 14825 17 14875 25
rect 14825 -17 14833 17
rect 14867 -17 14875 17
rect 14825 -25 14875 -17
rect 15375 17 15425 25
rect 15375 -17 15383 17
rect 15417 -17 15425 17
rect 15375 -25 15425 -17
rect 15925 17 15975 25
rect 15925 -17 15933 17
rect 15967 -17 15975 17
rect 15925 -25 15975 -17
rect 16475 17 16525 25
rect 16475 -17 16483 17
rect 16517 -17 16525 17
rect 16475 -25 16525 -17
rect 17025 17 17075 25
rect 17025 -17 17033 17
rect 17067 -17 17075 17
rect 17025 -25 17075 -17
rect 17575 17 17625 25
rect 17575 -17 17583 17
rect 17617 -17 17625 17
rect 17575 -25 17625 -17
rect 18125 17 18175 25
rect 18125 -17 18133 17
rect 18167 -17 18175 17
rect 18125 -25 18175 -17
rect 18675 17 18725 25
rect 18675 -17 18683 17
rect 18717 -17 18725 17
rect 18675 -25 18725 -17
rect 19225 17 19275 25
rect 19225 -17 19233 17
rect 19267 -17 19275 17
rect 19225 -25 19275 -17
rect 19775 17 19825 25
rect 19775 -17 19783 17
rect 19817 -17 19825 17
rect 19775 -25 19825 -17
rect 20000 -200 20012 20000
rect -212 -212 20012 -200
rect 20288 -488 20300 20288
rect -500 -500 20300 -488
rect 20800 -1000 20812 20800
rect -1012 -1012 20812 -1000
rect 24788 -4988 24800 24788
rect -5000 -5000 24800 -4988
<< via1 >>
rect -4988 20812 24788 24788
rect -4988 1680 -1012 20812
rect 613 20100 713 20200
rect 1713 20100 1813 20200
rect 2813 20100 2913 20200
rect 3913 20100 4013 20200
rect 5013 20100 5113 20200
rect 6113 20100 6213 20200
rect 7213 20100 7313 20200
rect 8313 20100 8413 20200
rect 9413 20100 9513 20200
rect 10513 20100 10613 20200
rect 11613 20100 11713 20200
rect 12713 20100 12813 20200
rect 13813 20100 13913 20200
rect 14913 20100 15013 20200
rect 16013 20100 16113 20200
rect 17113 20100 17213 20200
rect 18213 20100 18313 20200
rect 19313 20100 19413 20200
rect -400 19087 -300 19187
rect -400 17987 -300 18087
rect -400 16887 -300 16987
rect -400 15787 -300 15887
rect -400 14687 -300 14787
rect -400 13587 -300 13687
rect -400 12487 -300 12587
rect -400 11387 -300 11487
rect -400 10287 -300 10387
rect -400 9187 -300 9287
rect -400 8087 -300 8187
rect -400 6987 -300 7087
rect -400 5887 -300 5987
rect -400 4787 -300 4887
rect -400 3687 -300 3787
rect -400 2587 -300 2687
rect -400 1487 -300 1587
rect -400 387 -300 487
rect -17 19783 17 19817
rect 533 19783 567 19817
rect 1083 19783 1117 19817
rect 1633 19783 1667 19817
rect 2183 19783 2217 19817
rect 2733 19783 2767 19817
rect 3283 19783 3317 19817
rect 3833 19783 3867 19817
rect 4383 19783 4417 19817
rect 4933 19783 4967 19817
rect 5483 19783 5517 19817
rect 6033 19783 6067 19817
rect 6583 19783 6617 19817
rect 7133 19783 7167 19817
rect 7683 19783 7717 19817
rect 8233 19783 8267 19817
rect 8783 19783 8817 19817
rect 9333 19783 9367 19817
rect 9883 19783 9917 19817
rect 10433 19783 10467 19817
rect 10983 19783 11017 19817
rect 11533 19783 11567 19817
rect 12083 19783 12117 19817
rect 12633 19783 12667 19817
rect 13183 19783 13217 19817
rect 13733 19783 13767 19817
rect 14283 19783 14317 19817
rect 14833 19783 14867 19817
rect 15383 19783 15417 19817
rect 15933 19783 15967 19817
rect 16483 19783 16517 19817
rect 17033 19783 17067 19817
rect 17583 19783 17617 19817
rect 18133 19783 18167 19817
rect 18683 19783 18717 19817
rect 19233 19783 19267 19817
rect 19783 19783 19817 19817
rect 110 19360 440 19690
rect 660 19360 990 19690
rect 1210 19360 1540 19690
rect 1760 19360 2090 19690
rect 2310 19360 2640 19690
rect 2860 19360 3190 19690
rect 3410 19360 3740 19690
rect 3960 19360 4290 19690
rect 4510 19360 4840 19690
rect 5060 19360 5390 19690
rect 5610 19360 5940 19690
rect 6160 19360 6490 19690
rect 6710 19360 7040 19690
rect 7260 19360 7590 19690
rect 7810 19360 8140 19690
rect 8360 19360 8690 19690
rect 8910 19360 9240 19690
rect 9460 19360 9790 19690
rect 10010 19360 10340 19690
rect 10560 19360 10890 19690
rect 11110 19360 11440 19690
rect 11660 19360 11990 19690
rect 12210 19360 12540 19690
rect 12760 19360 13090 19690
rect 13310 19360 13640 19690
rect 13860 19360 14190 19690
rect 14410 19360 14740 19690
rect 14960 19360 15290 19690
rect 15510 19360 15840 19690
rect 16060 19360 16390 19690
rect 16610 19360 16940 19690
rect 17160 19360 17490 19690
rect 17710 19360 18040 19690
rect 18260 19360 18590 19690
rect 18810 19360 19140 19690
rect 19360 19360 19690 19690
rect -17 19233 17 19267
rect 533 19233 567 19267
rect 1083 19233 1117 19267
rect 1633 19233 1667 19267
rect 2183 19233 2217 19267
rect 2733 19233 2767 19267
rect 3283 19233 3317 19267
rect 3833 19233 3867 19267
rect 4383 19233 4417 19267
rect 4933 19233 4967 19267
rect 5483 19233 5517 19267
rect 6033 19233 6067 19267
rect 6583 19233 6617 19267
rect 7133 19233 7167 19267
rect 7683 19233 7717 19267
rect 8233 19233 8267 19267
rect 8783 19233 8817 19267
rect 9333 19233 9367 19267
rect 9883 19233 9917 19267
rect 10433 19233 10467 19267
rect 10983 19233 11017 19267
rect 11533 19233 11567 19267
rect 12083 19233 12117 19267
rect 12633 19233 12667 19267
rect 13183 19233 13217 19267
rect 13733 19233 13767 19267
rect 14283 19233 14317 19267
rect 14833 19233 14867 19267
rect 15383 19233 15417 19267
rect 15933 19233 15967 19267
rect 16483 19233 16517 19267
rect 17033 19233 17067 19267
rect 17583 19233 17617 19267
rect 18133 19233 18167 19267
rect 18683 19233 18717 19267
rect 19233 19233 19267 19267
rect 19783 19233 19817 19267
rect 110 18810 440 19140
rect 19360 18810 19690 19140
rect -17 18683 17 18717
rect 19233 18683 19267 18717
rect 19783 18683 19817 18717
rect 110 18260 440 18590
rect 19360 18260 19690 18590
rect -17 18133 17 18167
rect 19233 18133 19267 18167
rect 19783 18133 19817 18167
rect 110 17710 440 18040
rect 19360 17710 19690 18040
rect -17 17583 17 17617
rect 19233 17583 19267 17617
rect 19783 17583 19817 17617
rect 110 17160 440 17490
rect 19360 17160 19690 17490
rect -17 17033 17 17067
rect 19233 17033 19267 17067
rect 19783 17033 19817 17067
rect 110 16610 440 16940
rect 19360 16610 19690 16940
rect -17 16483 17 16517
rect 19233 16483 19267 16517
rect 19783 16483 19817 16517
rect 110 16060 440 16390
rect 19360 16060 19690 16390
rect -17 15933 17 15967
rect 19233 15933 19267 15967
rect 19783 15933 19817 15967
rect 110 15510 440 15840
rect 19360 15510 19690 15840
rect -17 15383 17 15417
rect 19233 15383 19267 15417
rect 19783 15383 19817 15417
rect 110 14960 440 15290
rect 19360 14960 19690 15290
rect -17 14833 17 14867
rect 19233 14833 19267 14867
rect 19783 14833 19817 14867
rect 110 14410 440 14740
rect 19360 14410 19690 14740
rect -17 14283 17 14317
rect 19233 14283 19267 14317
rect 19783 14283 19817 14317
rect 110 13860 440 14190
rect 19360 13860 19690 14190
rect -17 13733 17 13767
rect 19233 13733 19267 13767
rect 19783 13733 19817 13767
rect 110 13310 440 13640
rect 19360 13310 19690 13640
rect -17 13183 17 13217
rect 19233 13183 19267 13217
rect 19783 13183 19817 13217
rect 110 12760 440 13090
rect 19360 12760 19690 13090
rect -17 12633 17 12667
rect 19233 12633 19267 12667
rect 19783 12633 19817 12667
rect 110 12210 440 12540
rect 19360 12210 19690 12540
rect -17 12083 17 12117
rect 19233 12083 19267 12117
rect 19783 12083 19817 12117
rect 110 11660 440 11990
rect 19360 11660 19690 11990
rect -17 11533 17 11567
rect 19233 11533 19267 11567
rect 19783 11533 19817 11567
rect 110 11110 440 11440
rect 19360 11110 19690 11440
rect -17 10983 17 11017
rect 19233 10983 19267 11017
rect 19783 10983 19817 11017
rect 110 10560 440 10890
rect 19360 10560 19690 10890
rect -17 10433 17 10467
rect 19233 10433 19267 10467
rect 19783 10433 19817 10467
rect 110 10010 440 10340
rect 19360 10010 19690 10340
rect -17 9883 17 9917
rect 19233 9883 19267 9917
rect 19783 9883 19817 9917
rect 110 9460 440 9790
rect 19360 9460 19690 9790
rect -17 9333 17 9367
rect 19233 9333 19267 9367
rect 19783 9333 19817 9367
rect 110 8910 440 9240
rect 19360 8910 19690 9240
rect -17 8783 17 8817
rect 19233 8783 19267 8817
rect 19783 8783 19817 8817
rect 110 8360 440 8690
rect 19360 8360 19690 8690
rect -17 8233 17 8267
rect 19233 8233 19267 8267
rect 19783 8233 19817 8267
rect 110 7810 440 8140
rect 19360 7810 19690 8140
rect -17 7683 17 7717
rect 19233 7683 19267 7717
rect 19783 7683 19817 7717
rect 110 7260 440 7590
rect 19360 7260 19690 7590
rect -17 7133 17 7167
rect 19233 7133 19267 7167
rect 19783 7133 19817 7167
rect 110 6710 440 7040
rect 19360 6710 19690 7040
rect -17 6583 17 6617
rect 19233 6583 19267 6617
rect 19783 6583 19817 6617
rect 110 6160 440 6490
rect 19360 6160 19690 6490
rect -17 6033 17 6067
rect 19233 6033 19267 6067
rect 19783 6033 19817 6067
rect 110 5610 440 5940
rect 19360 5610 19690 5940
rect -17 5483 17 5517
rect 19233 5483 19267 5517
rect 19783 5483 19817 5517
rect 110 5060 440 5390
rect 19360 5060 19690 5390
rect -17 4933 17 4967
rect 19233 4933 19267 4967
rect 19783 4933 19817 4967
rect 110 4510 440 4840
rect 19360 4510 19690 4840
rect -17 4383 17 4417
rect 19233 4383 19267 4417
rect 19783 4383 19817 4417
rect 110 3960 440 4290
rect 19360 3960 19690 4290
rect -17 3833 17 3867
rect 19233 3833 19267 3867
rect 19783 3833 19817 3867
rect 110 3410 440 3740
rect 19360 3410 19690 3740
rect -17 3283 17 3317
rect 19233 3283 19267 3317
rect 19783 3283 19817 3317
rect 110 2860 440 3190
rect 19360 2860 19690 3190
rect -17 2733 17 2767
rect 19233 2733 19267 2767
rect 19783 2733 19817 2767
rect 110 2310 440 2640
rect 19360 2310 19690 2640
rect -17 2183 17 2217
rect 19233 2183 19267 2217
rect 19783 2183 19817 2217
rect 110 1760 440 2090
rect 19360 1760 19690 2090
rect -17 1633 17 1667
rect 19233 1633 19267 1667
rect 19783 1633 19817 1667
rect 110 1210 440 1540
rect 19360 1210 19690 1540
rect -17 1083 17 1117
rect 19233 1083 19267 1117
rect 19783 1083 19817 1117
rect 110 660 440 990
rect 19360 660 19690 990
rect -17 533 17 567
rect 19233 533 19267 567
rect 19783 533 19817 567
rect 110 110 440 440
rect 660 110 990 440
rect 1210 110 1540 440
rect 1760 110 2090 440
rect 2310 110 2640 440
rect 2860 110 3190 440
rect 3410 110 3740 440
rect 3960 110 4290 440
rect 4510 110 4840 440
rect 5060 110 5390 440
rect 5610 110 5940 440
rect 6160 110 6490 440
rect 6710 110 7040 440
rect 7260 110 7590 440
rect 7810 110 8140 440
rect 8360 110 8690 440
rect 8910 110 9240 440
rect 9460 110 9790 440
rect 10010 110 10340 440
rect 10560 110 10890 440
rect 11110 110 11440 440
rect 11660 110 11990 440
rect 12210 110 12540 440
rect 12760 110 13090 440
rect 13310 110 13640 440
rect 13860 110 14190 440
rect 14410 110 14740 440
rect 14960 110 15290 440
rect 15510 110 15840 440
rect 16060 110 16390 440
rect 16610 110 16940 440
rect 17160 110 17490 440
rect 17710 110 18040 440
rect 18260 110 18590 440
rect 18810 110 19140 440
rect 19360 110 19690 440
rect -17 -17 17 17
rect 533 -17 567 17
rect 1083 -17 1117 17
rect 1633 -17 1667 17
rect 2183 -17 2217 17
rect 2733 -17 2767 17
rect 3283 -17 3317 17
rect 3833 -17 3867 17
rect 4383 -17 4417 17
rect 4933 -17 4967 17
rect 5483 -17 5517 17
rect 6033 -17 6067 17
rect 6583 -17 6617 17
rect 7133 -17 7167 17
rect 7683 -17 7717 17
rect 8233 -17 8267 17
rect 8783 -17 8817 17
rect 9333 -17 9367 17
rect 9883 -17 9917 17
rect 10433 -17 10467 17
rect 10983 -17 11017 17
rect 11533 -17 11567 17
rect 12083 -17 12117 17
rect 12633 -17 12667 17
rect 13183 -17 13217 17
rect 13733 -17 13767 17
rect 14283 -17 14317 17
rect 14833 -17 14867 17
rect 15383 -17 15417 17
rect 15933 -17 15967 17
rect 16483 -17 16517 17
rect 17033 -17 17067 17
rect 17583 -17 17617 17
rect 18133 -17 18167 17
rect 18683 -17 18717 17
rect 19233 -17 19267 17
rect 19783 -17 19817 17
rect 20100 19313 20200 19413
rect 20100 18213 20200 18313
rect 20100 17113 20200 17213
rect 20100 16013 20200 16113
rect 20100 14913 20200 15013
rect 20100 13813 20200 13913
rect 20100 12713 20200 12813
rect 20100 11613 20200 11713
rect 20100 10513 20200 10613
rect 20100 9413 20200 9513
rect 20100 8313 20200 8413
rect 20100 7213 20200 7313
rect 20100 6113 20200 6213
rect 20100 5013 20200 5113
rect 20100 3913 20200 4013
rect 20100 2813 20200 2913
rect 20100 1713 20200 1813
rect 20100 613 20200 713
rect 387 -400 487 -300
rect 1487 -400 1587 -300
rect 2587 -400 2687 -300
rect 3687 -400 3787 -300
rect 4787 -400 4887 -300
rect 5887 -400 5987 -300
rect 6987 -400 7087 -300
rect 8087 -400 8187 -300
rect 9187 -400 9287 -300
rect 10287 -400 10387 -300
rect 11387 -400 11487 -300
rect 12487 -400 12587 -300
rect 13587 -400 13687 -300
rect 14687 -400 14787 -300
rect 15787 -400 15887 -300
rect 16887 -400 16987 -300
rect 17987 -400 18087 -300
rect 19087 -400 19187 -300
rect 20812 -1012 24788 20812
rect 30 -4988 24788 -1012
<< metal2 >>
rect -5000 24788 24800 24800
rect -5000 1680 -4988 24788
rect -1012 20800 20812 20812
rect -1012 1680 -1000 20800
rect 603 20200 723 20210
rect 603 20100 613 20200
rect 713 20100 723 20200
rect 603 20090 723 20100
rect 1703 20200 1823 20210
rect 1703 20100 1713 20200
rect 1813 20100 1823 20200
rect 1703 20090 1823 20100
rect 2803 20200 2923 20210
rect 2803 20100 2813 20200
rect 2913 20100 2923 20200
rect 2803 20090 2923 20100
rect 3903 20200 4023 20210
rect 3903 20100 3913 20200
rect 4013 20100 4023 20200
rect 3903 20090 4023 20100
rect 5003 20200 5123 20210
rect 5003 20100 5013 20200
rect 5113 20100 5123 20200
rect 5003 20090 5123 20100
rect 6103 20200 6223 20210
rect 6103 20100 6113 20200
rect 6213 20100 6223 20200
rect 6103 20090 6223 20100
rect 7203 20200 7323 20210
rect 7203 20100 7213 20200
rect 7313 20100 7323 20200
rect 7203 20090 7323 20100
rect 8303 20200 8423 20210
rect 8303 20100 8313 20200
rect 8413 20100 8423 20200
rect 8303 20090 8423 20100
rect 9403 20200 9523 20210
rect 9403 20100 9413 20200
rect 9513 20100 9523 20200
rect 9403 20090 9523 20100
rect 10503 20200 10623 20210
rect 10503 20100 10513 20200
rect 10613 20100 10623 20200
rect 10503 20090 10623 20100
rect 11603 20200 11723 20210
rect 11603 20100 11613 20200
rect 11713 20100 11723 20200
rect 11603 20090 11723 20100
rect 12703 20200 12823 20210
rect 12703 20100 12713 20200
rect 12813 20100 12823 20200
rect 12703 20090 12823 20100
rect 13803 20200 13923 20210
rect 13803 20100 13813 20200
rect 13913 20100 13923 20200
rect 13803 20090 13923 20100
rect 14903 20200 15023 20210
rect 14903 20100 14913 20200
rect 15013 20100 15023 20200
rect 14903 20090 15023 20100
rect 16003 20200 16123 20210
rect 16003 20100 16013 20200
rect 16113 20100 16123 20200
rect 16003 20090 16123 20100
rect 17103 20200 17223 20210
rect 17103 20100 17113 20200
rect 17213 20100 17223 20200
rect 17103 20090 17223 20100
rect 18203 20200 18323 20210
rect 18203 20100 18213 20200
rect 18313 20100 18323 20200
rect 18203 20090 18323 20100
rect 19303 20200 19423 20210
rect 19303 20100 19313 20200
rect 19413 20100 19423 20200
rect 19303 20090 19423 20100
rect -200 19817 20000 20000
rect -200 19783 -17 19817
rect 17 19783 533 19817
rect 567 19783 1083 19817
rect 1117 19783 1633 19817
rect 1667 19783 2183 19817
rect 2217 19783 2733 19817
rect 2767 19783 3283 19817
rect 3317 19783 3833 19817
rect 3867 19783 4383 19817
rect 4417 19783 4933 19817
rect 4967 19783 5483 19817
rect 5517 19783 6033 19817
rect 6067 19783 6583 19817
rect 6617 19783 7133 19817
rect 7167 19783 7683 19817
rect 7717 19783 8233 19817
rect 8267 19783 8783 19817
rect 8817 19783 9333 19817
rect 9367 19783 9883 19817
rect 9917 19783 10433 19817
rect 10467 19783 10983 19817
rect 11017 19783 11533 19817
rect 11567 19783 12083 19817
rect 12117 19783 12633 19817
rect 12667 19783 13183 19817
rect 13217 19783 13733 19817
rect 13767 19783 14283 19817
rect 14317 19783 14833 19817
rect 14867 19783 15383 19817
rect 15417 19783 15933 19817
rect 15967 19783 16483 19817
rect 16517 19783 17033 19817
rect 17067 19783 17583 19817
rect 17617 19783 18133 19817
rect 18167 19783 18683 19817
rect 18717 19783 19233 19817
rect 19267 19783 19783 19817
rect 19817 19783 20000 19817
rect -200 19775 20000 19783
rect -200 19275 25 19775
rect 100 19690 450 19700
rect 100 19360 110 19690
rect 440 19360 450 19690
rect 100 19350 450 19360
rect 525 19275 575 19775
rect 650 19690 1000 19700
rect 650 19360 660 19690
rect 990 19360 1000 19690
rect 650 19350 1000 19360
rect 1075 19275 1125 19775
rect 1200 19690 1550 19700
rect 1200 19360 1210 19690
rect 1540 19360 1550 19690
rect 1200 19350 1550 19360
rect 1625 19275 1675 19775
rect 1750 19690 2100 19700
rect 1750 19360 1760 19690
rect 2090 19360 2100 19690
rect 1750 19350 2100 19360
rect 2175 19275 2225 19775
rect 2300 19690 2650 19700
rect 2300 19360 2310 19690
rect 2640 19360 2650 19690
rect 2300 19350 2650 19360
rect 2725 19275 2775 19775
rect 2850 19690 3200 19700
rect 2850 19360 2860 19690
rect 3190 19360 3200 19690
rect 2850 19350 3200 19360
rect 3275 19275 3325 19775
rect 3400 19690 3750 19700
rect 3400 19360 3410 19690
rect 3740 19360 3750 19690
rect 3400 19350 3750 19360
rect 3825 19275 3875 19775
rect 3950 19690 4300 19700
rect 3950 19360 3960 19690
rect 4290 19360 4300 19690
rect 3950 19350 4300 19360
rect 4375 19275 4425 19775
rect 4500 19690 4850 19700
rect 4500 19360 4510 19690
rect 4840 19360 4850 19690
rect 4500 19350 4850 19360
rect 4925 19275 4975 19775
rect 5050 19690 5400 19700
rect 5050 19360 5060 19690
rect 5390 19360 5400 19690
rect 5050 19350 5400 19360
rect 5475 19275 5525 19775
rect 5600 19690 5950 19700
rect 5600 19360 5610 19690
rect 5940 19360 5950 19690
rect 5600 19350 5950 19360
rect 6025 19275 6075 19775
rect 6150 19690 6500 19700
rect 6150 19360 6160 19690
rect 6490 19360 6500 19690
rect 6150 19350 6500 19360
rect 6575 19275 6625 19775
rect 6700 19690 7050 19700
rect 6700 19360 6710 19690
rect 7040 19360 7050 19690
rect 6700 19350 7050 19360
rect 7125 19275 7175 19775
rect 7250 19690 7600 19700
rect 7250 19360 7260 19690
rect 7590 19360 7600 19690
rect 7250 19350 7600 19360
rect 7675 19275 7725 19775
rect 7800 19690 8150 19700
rect 7800 19360 7810 19690
rect 8140 19360 8150 19690
rect 7800 19350 8150 19360
rect 8225 19275 8275 19775
rect 8350 19690 8700 19700
rect 8350 19360 8360 19690
rect 8690 19360 8700 19690
rect 8350 19350 8700 19360
rect 8775 19275 8825 19775
rect 8900 19690 9250 19700
rect 8900 19360 8910 19690
rect 9240 19360 9250 19690
rect 8900 19350 9250 19360
rect 9325 19275 9375 19775
rect 9450 19690 9800 19700
rect 9450 19360 9460 19690
rect 9790 19360 9800 19690
rect 9450 19350 9800 19360
rect 9875 19275 9925 19775
rect 10000 19690 10350 19700
rect 10000 19360 10010 19690
rect 10340 19360 10350 19690
rect 10000 19350 10350 19360
rect 10425 19275 10475 19775
rect 10550 19690 10900 19700
rect 10550 19360 10560 19690
rect 10890 19360 10900 19690
rect 10550 19350 10900 19360
rect 10975 19275 11025 19775
rect 11100 19690 11450 19700
rect 11100 19360 11110 19690
rect 11440 19360 11450 19690
rect 11100 19350 11450 19360
rect 11525 19275 11575 19775
rect 11650 19690 12000 19700
rect 11650 19360 11660 19690
rect 11990 19360 12000 19690
rect 11650 19350 12000 19360
rect 12075 19275 12125 19775
rect 12200 19690 12550 19700
rect 12200 19360 12210 19690
rect 12540 19360 12550 19690
rect 12200 19350 12550 19360
rect 12625 19275 12675 19775
rect 12750 19690 13100 19700
rect 12750 19360 12760 19690
rect 13090 19360 13100 19690
rect 12750 19350 13100 19360
rect 13175 19275 13225 19775
rect 13300 19690 13650 19700
rect 13300 19360 13310 19690
rect 13640 19360 13650 19690
rect 13300 19350 13650 19360
rect 13725 19275 13775 19775
rect 13850 19690 14200 19700
rect 13850 19360 13860 19690
rect 14190 19360 14200 19690
rect 13850 19350 14200 19360
rect 14275 19275 14325 19775
rect 14400 19690 14750 19700
rect 14400 19360 14410 19690
rect 14740 19360 14750 19690
rect 14400 19350 14750 19360
rect 14825 19275 14875 19775
rect 14950 19690 15300 19700
rect 14950 19360 14960 19690
rect 15290 19360 15300 19690
rect 14950 19350 15300 19360
rect 15375 19275 15425 19775
rect 15500 19690 15850 19700
rect 15500 19360 15510 19690
rect 15840 19360 15850 19690
rect 15500 19350 15850 19360
rect 15925 19275 15975 19775
rect 16050 19690 16400 19700
rect 16050 19360 16060 19690
rect 16390 19360 16400 19690
rect 16050 19350 16400 19360
rect 16475 19275 16525 19775
rect 16600 19690 16950 19700
rect 16600 19360 16610 19690
rect 16940 19360 16950 19690
rect 16600 19350 16950 19360
rect 17025 19275 17075 19775
rect 17150 19690 17500 19700
rect 17150 19360 17160 19690
rect 17490 19360 17500 19690
rect 17150 19350 17500 19360
rect 17575 19275 17625 19775
rect 17700 19690 18050 19700
rect 17700 19360 17710 19690
rect 18040 19360 18050 19690
rect 17700 19350 18050 19360
rect 18125 19275 18175 19775
rect 18250 19690 18600 19700
rect 18250 19360 18260 19690
rect 18590 19360 18600 19690
rect 18250 19350 18600 19360
rect 18675 19275 18725 19775
rect 18800 19690 19150 19700
rect 18800 19360 18810 19690
rect 19140 19360 19150 19690
rect 18800 19350 19150 19360
rect 19225 19275 19275 19775
rect 19350 19690 19700 19700
rect 19350 19360 19360 19690
rect 19690 19360 19700 19690
rect 19350 19350 19700 19360
rect 19775 19275 20000 19775
rect 20090 19413 20210 19423
rect 20090 19313 20100 19413
rect 20200 19313 20210 19413
rect 20090 19303 20210 19313
rect -200 19267 20000 19275
rect -200 19233 -17 19267
rect 17 19233 533 19267
rect 567 19233 1083 19267
rect 1117 19233 1633 19267
rect 1667 19233 2183 19267
rect 2217 19233 2733 19267
rect 2767 19233 3283 19267
rect 3317 19233 3833 19267
rect 3867 19233 4383 19267
rect 4417 19233 4933 19267
rect 4967 19233 5483 19267
rect 5517 19233 6033 19267
rect 6067 19233 6583 19267
rect 6617 19233 7133 19267
rect 7167 19233 7683 19267
rect 7717 19233 8233 19267
rect 8267 19233 8783 19267
rect 8817 19233 9333 19267
rect 9367 19233 9883 19267
rect 9917 19233 10433 19267
rect 10467 19233 10983 19267
rect 11017 19233 11533 19267
rect 11567 19233 12083 19267
rect 12117 19233 12633 19267
rect 12667 19233 13183 19267
rect 13217 19233 13733 19267
rect 13767 19233 14283 19267
rect 14317 19233 14833 19267
rect 14867 19233 15383 19267
rect 15417 19233 15933 19267
rect 15967 19233 16483 19267
rect 16517 19233 17033 19267
rect 17067 19233 17583 19267
rect 17617 19233 18133 19267
rect 18167 19233 18683 19267
rect 18717 19233 19233 19267
rect 19267 19233 19783 19267
rect 19817 19233 20000 19267
rect -200 19225 20000 19233
rect -410 19187 -290 19197
rect -410 19087 -400 19187
rect -300 19087 -290 19187
rect -410 19077 -290 19087
rect -200 18725 25 19225
rect 525 19200 575 19225
rect 1075 19200 1125 19225
rect 1625 19200 1675 19225
rect 2175 19200 2225 19225
rect 2725 19200 2775 19225
rect 3275 19200 3325 19225
rect 3825 19200 3875 19225
rect 4375 19200 4425 19225
rect 4925 19200 4975 19225
rect 5475 19200 5525 19225
rect 6025 19200 6075 19225
rect 6575 19200 6625 19225
rect 7125 19200 7175 19225
rect 7675 19200 7725 19225
rect 8225 19200 8275 19225
rect 8775 19200 8825 19225
rect 9325 19200 9375 19225
rect 9875 19200 9925 19225
rect 10425 19200 10475 19225
rect 10975 19200 11025 19225
rect 11525 19200 11575 19225
rect 12075 19200 12125 19225
rect 12625 19200 12675 19225
rect 13175 19200 13225 19225
rect 13725 19200 13775 19225
rect 14275 19200 14325 19225
rect 14825 19200 14875 19225
rect 15375 19200 15425 19225
rect 15925 19200 15975 19225
rect 16475 19200 16525 19225
rect 17025 19200 17075 19225
rect 17575 19200 17625 19225
rect 18125 19200 18175 19225
rect 18675 19200 18725 19225
rect 100 19140 450 19150
rect 100 18810 110 19140
rect 440 18810 450 19140
rect 100 18800 450 18810
rect 19225 18725 19275 19225
rect 19350 19140 19700 19150
rect 19350 18810 19360 19140
rect 19690 18810 19700 19140
rect 19350 18800 19700 18810
rect 19775 18725 20000 19225
rect -200 18717 500 18725
rect -200 18683 -17 18717
rect 17 18683 500 18717
rect -200 18675 500 18683
rect 19200 18717 20000 18725
rect 19200 18683 19233 18717
rect 19267 18683 19783 18717
rect 19817 18683 20000 18717
rect 19200 18675 20000 18683
rect -200 18175 25 18675
rect 100 18590 450 18600
rect 100 18260 110 18590
rect 440 18260 450 18590
rect 100 18250 450 18260
rect 19225 18175 19275 18675
rect 19350 18590 19700 18600
rect 19350 18260 19360 18590
rect 19690 18260 19700 18590
rect 19350 18250 19700 18260
rect 19775 18175 20000 18675
rect 20090 18313 20210 18323
rect 20090 18213 20100 18313
rect 20200 18213 20210 18313
rect 20090 18203 20210 18213
rect -200 18167 500 18175
rect -200 18133 -17 18167
rect 17 18133 500 18167
rect -200 18125 500 18133
rect 19200 18167 20000 18175
rect 19200 18133 19233 18167
rect 19267 18133 19783 18167
rect 19817 18133 20000 18167
rect 19200 18125 20000 18133
rect -410 18087 -290 18097
rect -410 17987 -400 18087
rect -300 17987 -290 18087
rect -410 17977 -290 17987
rect -200 17625 25 18125
rect 100 18040 450 18050
rect 100 17710 110 18040
rect 440 17710 450 18040
rect 100 17700 450 17710
rect 19225 17625 19275 18125
rect 19350 18040 19700 18050
rect 19350 17710 19360 18040
rect 19690 17710 19700 18040
rect 19350 17700 19700 17710
rect 19775 17625 20000 18125
rect -200 17617 500 17625
rect -200 17583 -17 17617
rect 17 17583 500 17617
rect -200 17575 500 17583
rect 19200 17617 20000 17625
rect 19200 17583 19233 17617
rect 19267 17583 19783 17617
rect 19817 17583 20000 17617
rect 19200 17575 20000 17583
rect -200 17075 25 17575
rect 100 17490 450 17500
rect 100 17160 110 17490
rect 440 17160 450 17490
rect 100 17150 450 17160
rect 19225 17075 19275 17575
rect 19350 17490 19700 17500
rect 19350 17160 19360 17490
rect 19690 17160 19700 17490
rect 19350 17150 19700 17160
rect 19775 17075 20000 17575
rect 20090 17213 20210 17223
rect 20090 17113 20100 17213
rect 20200 17113 20210 17213
rect 20090 17103 20210 17113
rect -200 17067 500 17075
rect -200 17033 -17 17067
rect 17 17033 500 17067
rect -200 17025 500 17033
rect 19200 17067 20000 17075
rect 19200 17033 19233 17067
rect 19267 17033 19783 17067
rect 19817 17033 20000 17067
rect 19200 17025 20000 17033
rect -410 16987 -290 16997
rect -410 16887 -400 16987
rect -300 16887 -290 16987
rect -410 16877 -290 16887
rect -200 16525 25 17025
rect 100 16940 450 16950
rect 100 16610 110 16940
rect 440 16610 450 16940
rect 100 16600 450 16610
rect 19225 16525 19275 17025
rect 19350 16940 19700 16950
rect 19350 16610 19360 16940
rect 19690 16610 19700 16940
rect 19350 16600 19700 16610
rect 19775 16525 20000 17025
rect -200 16517 500 16525
rect -200 16483 -17 16517
rect 17 16483 500 16517
rect -200 16475 500 16483
rect 19200 16517 20000 16525
rect 19200 16483 19233 16517
rect 19267 16483 19783 16517
rect 19817 16483 20000 16517
rect 19200 16475 20000 16483
rect -200 15975 25 16475
rect 100 16390 450 16400
rect 100 16060 110 16390
rect 440 16060 450 16390
rect 100 16050 450 16060
rect 19225 15975 19275 16475
rect 19350 16390 19700 16400
rect 19350 16060 19360 16390
rect 19690 16060 19700 16390
rect 19350 16050 19700 16060
rect 19775 15975 20000 16475
rect 20090 16113 20210 16123
rect 20090 16013 20100 16113
rect 20200 16013 20210 16113
rect 20090 16003 20210 16013
rect -200 15967 500 15975
rect -200 15933 -17 15967
rect 17 15933 500 15967
rect -200 15925 500 15933
rect 19200 15967 20000 15975
rect 19200 15933 19233 15967
rect 19267 15933 19783 15967
rect 19817 15933 20000 15967
rect 19200 15925 20000 15933
rect -410 15887 -290 15897
rect -410 15787 -400 15887
rect -300 15787 -290 15887
rect -410 15777 -290 15787
rect -200 15425 25 15925
rect 100 15840 450 15850
rect 100 15510 110 15840
rect 440 15510 450 15840
rect 100 15500 450 15510
rect 19225 15425 19275 15925
rect 19350 15840 19700 15850
rect 19350 15510 19360 15840
rect 19690 15510 19700 15840
rect 19350 15500 19700 15510
rect 19775 15425 20000 15925
rect -200 15417 500 15425
rect -200 15383 -17 15417
rect 17 15383 500 15417
rect -200 15375 500 15383
rect 19200 15417 20000 15425
rect 19200 15383 19233 15417
rect 19267 15383 19783 15417
rect 19817 15383 20000 15417
rect 19200 15375 20000 15383
rect -200 14875 25 15375
rect 100 15290 450 15300
rect 100 14960 110 15290
rect 440 14960 450 15290
rect 100 14950 450 14960
rect 19225 14875 19275 15375
rect 19350 15290 19700 15300
rect 19350 14960 19360 15290
rect 19690 14960 19700 15290
rect 19350 14950 19700 14960
rect 19775 14875 20000 15375
rect 20090 15013 20210 15023
rect 20090 14913 20100 15013
rect 20200 14913 20210 15013
rect 20090 14903 20210 14913
rect -200 14867 500 14875
rect -200 14833 -17 14867
rect 17 14833 500 14867
rect -200 14825 500 14833
rect 19200 14867 20000 14875
rect 19200 14833 19233 14867
rect 19267 14833 19783 14867
rect 19817 14833 20000 14867
rect 19200 14825 20000 14833
rect -410 14787 -290 14797
rect -410 14687 -400 14787
rect -300 14687 -290 14787
rect -410 14677 -290 14687
rect -200 14325 25 14825
rect 100 14740 450 14750
rect 100 14410 110 14740
rect 440 14410 450 14740
rect 100 14400 450 14410
rect 19225 14325 19275 14825
rect 19350 14740 19700 14750
rect 19350 14410 19360 14740
rect 19690 14410 19700 14740
rect 19350 14400 19700 14410
rect 19775 14325 20000 14825
rect -200 14317 500 14325
rect -200 14283 -17 14317
rect 17 14283 500 14317
rect -200 14275 500 14283
rect 19200 14317 20000 14325
rect 19200 14283 19233 14317
rect 19267 14283 19783 14317
rect 19817 14283 20000 14317
rect 19200 14275 20000 14283
rect -200 13775 25 14275
rect 100 14190 450 14200
rect 100 13860 110 14190
rect 440 13860 450 14190
rect 100 13850 450 13860
rect 19225 13775 19275 14275
rect 19350 14190 19700 14200
rect 19350 13860 19360 14190
rect 19690 13860 19700 14190
rect 19350 13850 19700 13860
rect 19775 13775 20000 14275
rect 20090 13913 20210 13923
rect 20090 13813 20100 13913
rect 20200 13813 20210 13913
rect 20090 13803 20210 13813
rect -200 13767 500 13775
rect -200 13733 -17 13767
rect 17 13733 500 13767
rect -200 13725 500 13733
rect 19200 13767 20000 13775
rect 19200 13733 19233 13767
rect 19267 13733 19783 13767
rect 19817 13733 20000 13767
rect 19200 13725 20000 13733
rect -410 13687 -290 13697
rect -410 13587 -400 13687
rect -300 13587 -290 13687
rect -410 13577 -290 13587
rect -200 13225 25 13725
rect 100 13640 450 13650
rect 100 13310 110 13640
rect 440 13310 450 13640
rect 100 13300 450 13310
rect 19225 13225 19275 13725
rect 19350 13640 19700 13650
rect 19350 13310 19360 13640
rect 19690 13310 19700 13640
rect 19350 13300 19700 13310
rect 19775 13225 20000 13725
rect -200 13217 500 13225
rect -200 13183 -17 13217
rect 17 13183 500 13217
rect -200 13175 500 13183
rect 19200 13217 20000 13225
rect 19200 13183 19233 13217
rect 19267 13183 19783 13217
rect 19817 13183 20000 13217
rect 19200 13175 20000 13183
rect -200 12675 25 13175
rect 100 13090 450 13100
rect 100 12760 110 13090
rect 440 12760 450 13090
rect 100 12750 450 12760
rect 19225 12675 19275 13175
rect 19350 13090 19700 13100
rect 19350 12760 19360 13090
rect 19690 12760 19700 13090
rect 19350 12750 19700 12760
rect 19775 12675 20000 13175
rect 20090 12813 20210 12823
rect 20090 12713 20100 12813
rect 20200 12713 20210 12813
rect 20090 12703 20210 12713
rect -200 12667 500 12675
rect -200 12633 -17 12667
rect 17 12633 500 12667
rect -200 12625 500 12633
rect 19200 12667 20000 12675
rect 19200 12633 19233 12667
rect 19267 12633 19783 12667
rect 19817 12633 20000 12667
rect 19200 12625 20000 12633
rect -410 12587 -290 12597
rect -410 12487 -400 12587
rect -300 12487 -290 12587
rect -410 12477 -290 12487
rect -200 12125 25 12625
rect 100 12540 450 12550
rect 100 12210 110 12540
rect 440 12210 450 12540
rect 100 12200 450 12210
rect 19225 12125 19275 12625
rect 19350 12540 19700 12550
rect 19350 12210 19360 12540
rect 19690 12210 19700 12540
rect 19350 12200 19700 12210
rect 19775 12125 20000 12625
rect -200 12117 500 12125
rect -200 12083 -17 12117
rect 17 12083 500 12117
rect -200 12075 500 12083
rect 19200 12117 20000 12125
rect 19200 12083 19233 12117
rect 19267 12083 19783 12117
rect 19817 12083 20000 12117
rect 19200 12075 20000 12083
rect -200 11575 25 12075
rect 100 11990 450 12000
rect 100 11660 110 11990
rect 440 11660 450 11990
rect 100 11650 450 11660
rect 19225 11575 19275 12075
rect 19350 11990 19700 12000
rect 19350 11660 19360 11990
rect 19690 11660 19700 11990
rect 19350 11650 19700 11660
rect 19775 11575 20000 12075
rect 20090 11713 20210 11723
rect 20090 11613 20100 11713
rect 20200 11613 20210 11713
rect 20090 11603 20210 11613
rect -200 11567 500 11575
rect -200 11533 -17 11567
rect 17 11533 500 11567
rect -200 11525 500 11533
rect 19200 11567 20000 11575
rect 19200 11533 19233 11567
rect 19267 11533 19783 11567
rect 19817 11533 20000 11567
rect 19200 11525 20000 11533
rect -410 11487 -290 11497
rect -410 11387 -400 11487
rect -300 11387 -290 11487
rect -410 11377 -290 11387
rect -200 11025 25 11525
rect 100 11440 450 11450
rect 100 11110 110 11440
rect 440 11110 450 11440
rect 100 11100 450 11110
rect 19225 11025 19275 11525
rect 19350 11440 19700 11450
rect 19350 11110 19360 11440
rect 19690 11110 19700 11440
rect 19350 11100 19700 11110
rect 19775 11025 20000 11525
rect -200 11017 500 11025
rect -200 10983 -17 11017
rect 17 10983 500 11017
rect -200 10975 500 10983
rect 19200 11017 20000 11025
rect 19200 10983 19233 11017
rect 19267 10983 19783 11017
rect 19817 10983 20000 11017
rect 19200 10975 20000 10983
rect -200 10475 25 10975
rect 100 10890 450 10900
rect 100 10560 110 10890
rect 440 10560 450 10890
rect 100 10550 450 10560
rect 19225 10475 19275 10975
rect 19350 10890 19700 10900
rect 19350 10560 19360 10890
rect 19690 10560 19700 10890
rect 19350 10550 19700 10560
rect 19775 10475 20000 10975
rect 20090 10613 20210 10623
rect 20090 10513 20100 10613
rect 20200 10513 20210 10613
rect 20090 10503 20210 10513
rect -200 10467 500 10475
rect -200 10433 -17 10467
rect 17 10433 500 10467
rect -200 10425 500 10433
rect 19200 10467 20000 10475
rect 19200 10433 19233 10467
rect 19267 10433 19783 10467
rect 19817 10433 20000 10467
rect 19200 10425 20000 10433
rect -410 10387 -290 10397
rect -410 10287 -400 10387
rect -300 10287 -290 10387
rect -410 10277 -290 10287
rect -200 9925 25 10425
rect 100 10340 450 10350
rect 100 10010 110 10340
rect 440 10010 450 10340
rect 100 10000 450 10010
rect 19225 9925 19275 10425
rect 19350 10340 19700 10350
rect 19350 10010 19360 10340
rect 19690 10010 19700 10340
rect 19350 10000 19700 10010
rect 19775 9925 20000 10425
rect -200 9917 500 9925
rect -200 9883 -17 9917
rect 17 9883 500 9917
rect -200 9875 500 9883
rect 19200 9917 20000 9925
rect 19200 9883 19233 9917
rect 19267 9883 19783 9917
rect 19817 9883 20000 9917
rect 19200 9875 20000 9883
rect -200 9375 25 9875
rect 100 9790 450 9800
rect 100 9460 110 9790
rect 440 9460 450 9790
rect 100 9450 450 9460
rect 19225 9375 19275 9875
rect 19350 9790 19700 9800
rect 19350 9460 19360 9790
rect 19690 9460 19700 9790
rect 19350 9450 19700 9460
rect 19775 9375 20000 9875
rect 20090 9513 20210 9523
rect 20090 9413 20100 9513
rect 20200 9413 20210 9513
rect 20090 9403 20210 9413
rect -200 9367 500 9375
rect -200 9333 -17 9367
rect 17 9333 500 9367
rect -200 9325 500 9333
rect 19200 9367 20000 9375
rect 19200 9333 19233 9367
rect 19267 9333 19783 9367
rect 19817 9333 20000 9367
rect 19200 9325 20000 9333
rect -410 9287 -290 9297
rect -410 9187 -400 9287
rect -300 9187 -290 9287
rect -410 9177 -290 9187
rect -200 8825 25 9325
rect 100 9240 450 9250
rect 100 8910 110 9240
rect 440 8910 450 9240
rect 100 8900 450 8910
rect 19225 8825 19275 9325
rect 19350 9240 19700 9250
rect 19350 8910 19360 9240
rect 19690 8910 19700 9240
rect 19350 8900 19700 8910
rect 19775 8825 20000 9325
rect -200 8817 500 8825
rect -200 8783 -17 8817
rect 17 8783 500 8817
rect -200 8775 500 8783
rect 19200 8817 20000 8825
rect 19200 8783 19233 8817
rect 19267 8783 19783 8817
rect 19817 8783 20000 8817
rect 19200 8775 20000 8783
rect -200 8275 25 8775
rect 100 8690 450 8700
rect 100 8360 110 8690
rect 440 8360 450 8690
rect 100 8350 450 8360
rect 19225 8275 19275 8775
rect 19350 8690 19700 8700
rect 19350 8360 19360 8690
rect 19690 8360 19700 8690
rect 19350 8350 19700 8360
rect 19775 8275 20000 8775
rect 20090 8413 20210 8423
rect 20090 8313 20100 8413
rect 20200 8313 20210 8413
rect 20090 8303 20210 8313
rect -200 8267 500 8275
rect -200 8233 -17 8267
rect 17 8233 500 8267
rect -200 8225 500 8233
rect 19200 8267 20000 8275
rect 19200 8233 19233 8267
rect 19267 8233 19783 8267
rect 19817 8233 20000 8267
rect 19200 8225 20000 8233
rect -410 8187 -290 8197
rect -410 8087 -400 8187
rect -300 8087 -290 8187
rect -410 8077 -290 8087
rect -200 7725 25 8225
rect 100 8140 450 8150
rect 100 7810 110 8140
rect 440 7810 450 8140
rect 100 7800 450 7810
rect 19225 7725 19275 8225
rect 19350 8140 19700 8150
rect 19350 7810 19360 8140
rect 19690 7810 19700 8140
rect 19350 7800 19700 7810
rect 19775 7725 20000 8225
rect -200 7717 500 7725
rect -200 7683 -17 7717
rect 17 7683 500 7717
rect -200 7675 500 7683
rect 19200 7717 20000 7725
rect 19200 7683 19233 7717
rect 19267 7683 19783 7717
rect 19817 7683 20000 7717
rect 19200 7675 20000 7683
rect -200 7175 25 7675
rect 100 7590 450 7600
rect 100 7260 110 7590
rect 440 7260 450 7590
rect 100 7250 450 7260
rect 19225 7175 19275 7675
rect 19350 7590 19700 7600
rect 19350 7260 19360 7590
rect 19690 7260 19700 7590
rect 19350 7250 19700 7260
rect 19775 7175 20000 7675
rect 20090 7313 20210 7323
rect 20090 7213 20100 7313
rect 20200 7213 20210 7313
rect 20090 7203 20210 7213
rect -200 7167 500 7175
rect -200 7133 -17 7167
rect 17 7133 500 7167
rect -200 7125 500 7133
rect 19200 7167 20000 7175
rect 19200 7133 19233 7167
rect 19267 7133 19783 7167
rect 19817 7133 20000 7167
rect 19200 7125 20000 7133
rect -410 7087 -290 7097
rect -410 6987 -400 7087
rect -300 6987 -290 7087
rect -410 6977 -290 6987
rect -200 6625 25 7125
rect 100 7040 450 7050
rect 100 6710 110 7040
rect 440 6710 450 7040
rect 100 6700 450 6710
rect 19225 6625 19275 7125
rect 19350 7040 19700 7050
rect 19350 6710 19360 7040
rect 19690 6710 19700 7040
rect 19350 6700 19700 6710
rect 19775 6625 20000 7125
rect -200 6617 500 6625
rect -200 6583 -17 6617
rect 17 6583 500 6617
rect -200 6575 500 6583
rect 19200 6617 20000 6625
rect 19200 6583 19233 6617
rect 19267 6583 19783 6617
rect 19817 6583 20000 6617
rect 19200 6575 20000 6583
rect -200 6075 25 6575
rect 100 6490 450 6500
rect 100 6160 110 6490
rect 440 6160 450 6490
rect 100 6150 450 6160
rect 19225 6075 19275 6575
rect 19350 6490 19700 6500
rect 19350 6160 19360 6490
rect 19690 6160 19700 6490
rect 19350 6150 19700 6160
rect 19775 6075 20000 6575
rect 20090 6213 20210 6223
rect 20090 6113 20100 6213
rect 20200 6113 20210 6213
rect 20090 6103 20210 6113
rect -200 6067 500 6075
rect -200 6033 -17 6067
rect 17 6033 500 6067
rect -200 6025 500 6033
rect 19200 6067 20000 6075
rect 19200 6033 19233 6067
rect 19267 6033 19783 6067
rect 19817 6033 20000 6067
rect 19200 6025 20000 6033
rect -410 5987 -290 5997
rect -410 5887 -400 5987
rect -300 5887 -290 5987
rect -410 5877 -290 5887
rect -200 5525 25 6025
rect 100 5940 450 5950
rect 100 5610 110 5940
rect 440 5610 450 5940
rect 100 5600 450 5610
rect 19225 5525 19275 6025
rect 19350 5940 19700 5950
rect 19350 5610 19360 5940
rect 19690 5610 19700 5940
rect 19350 5600 19700 5610
rect 19775 5525 20000 6025
rect -200 5517 500 5525
rect -200 5483 -17 5517
rect 17 5483 500 5517
rect -200 5475 500 5483
rect 19200 5517 20000 5525
rect 19200 5483 19233 5517
rect 19267 5483 19783 5517
rect 19817 5483 20000 5517
rect 19200 5475 20000 5483
rect -200 4975 25 5475
rect 100 5390 450 5400
rect 100 5060 110 5390
rect 440 5060 450 5390
rect 100 5050 450 5060
rect 19225 4975 19275 5475
rect 19350 5390 19700 5400
rect 19350 5060 19360 5390
rect 19690 5060 19700 5390
rect 19350 5050 19700 5060
rect 19775 4975 20000 5475
rect 20090 5113 20210 5123
rect 20090 5013 20100 5113
rect 20200 5013 20210 5113
rect 20090 5003 20210 5013
rect -200 4967 500 4975
rect -200 4933 -17 4967
rect 17 4933 500 4967
rect -200 4925 500 4933
rect 19200 4967 20000 4975
rect 19200 4933 19233 4967
rect 19267 4933 19783 4967
rect 19817 4933 20000 4967
rect 19200 4925 20000 4933
rect -410 4887 -290 4897
rect -410 4787 -400 4887
rect -300 4787 -290 4887
rect -410 4777 -290 4787
rect -200 4425 25 4925
rect 100 4840 450 4850
rect 100 4510 110 4840
rect 440 4510 450 4840
rect 100 4500 450 4510
rect 19225 4425 19275 4925
rect 19350 4840 19700 4850
rect 19350 4510 19360 4840
rect 19690 4510 19700 4840
rect 19350 4500 19700 4510
rect 19775 4425 20000 4925
rect -200 4417 500 4425
rect -200 4383 -17 4417
rect 17 4383 500 4417
rect -200 4375 500 4383
rect 19200 4417 20000 4425
rect 19200 4383 19233 4417
rect 19267 4383 19783 4417
rect 19817 4383 20000 4417
rect 19200 4375 20000 4383
rect -200 3875 25 4375
rect 100 4290 450 4300
rect 100 3960 110 4290
rect 440 3960 450 4290
rect 100 3950 450 3960
rect 19225 3875 19275 4375
rect 19350 4290 19700 4300
rect 19350 3960 19360 4290
rect 19690 3960 19700 4290
rect 19350 3950 19700 3960
rect 19775 3875 20000 4375
rect 20090 4013 20210 4023
rect 20090 3913 20100 4013
rect 20200 3913 20210 4013
rect 20090 3903 20210 3913
rect -200 3867 500 3875
rect -200 3833 -17 3867
rect 17 3833 500 3867
rect -200 3825 500 3833
rect 19200 3867 20000 3875
rect 19200 3833 19233 3867
rect 19267 3833 19783 3867
rect 19817 3833 20000 3867
rect 19200 3825 20000 3833
rect -410 3787 -290 3797
rect -410 3687 -400 3787
rect -300 3687 -290 3787
rect -410 3677 -290 3687
rect -200 3325 25 3825
rect 100 3740 450 3750
rect 100 3410 110 3740
rect 440 3410 450 3740
rect 100 3400 450 3410
rect 19225 3325 19275 3825
rect 19350 3740 19700 3750
rect 19350 3410 19360 3740
rect 19690 3410 19700 3740
rect 19350 3400 19700 3410
rect 19775 3325 20000 3825
rect -200 3317 500 3325
rect -200 3283 -17 3317
rect 17 3283 500 3317
rect -200 3275 500 3283
rect 19200 3317 20000 3325
rect 19200 3283 19233 3317
rect 19267 3283 19783 3317
rect 19817 3283 20000 3317
rect 19200 3275 20000 3283
rect -200 2775 25 3275
rect 100 3190 450 3200
rect 100 2860 110 3190
rect 440 2860 450 3190
rect 100 2850 450 2860
rect 19225 2775 19275 3275
rect 19350 3190 19700 3200
rect 19350 2860 19360 3190
rect 19690 2860 19700 3190
rect 19350 2850 19700 2860
rect 19775 2775 20000 3275
rect 20090 2913 20210 2923
rect 20090 2813 20100 2913
rect 20200 2813 20210 2913
rect 20090 2803 20210 2813
rect -200 2767 500 2775
rect -200 2733 -17 2767
rect 17 2733 500 2767
rect -200 2725 500 2733
rect 19200 2767 20000 2775
rect 19200 2733 19233 2767
rect 19267 2733 19783 2767
rect 19817 2733 20000 2767
rect 19200 2725 20000 2733
rect -410 2687 -290 2697
rect -410 2587 -400 2687
rect -300 2587 -290 2687
rect -410 2577 -290 2587
rect -200 2225 25 2725
rect 100 2640 450 2650
rect 100 2310 110 2640
rect 440 2310 450 2640
rect 100 2300 450 2310
rect 19225 2225 19275 2725
rect 19350 2640 19700 2650
rect 19350 2310 19360 2640
rect 19690 2310 19700 2640
rect 19350 2300 19700 2310
rect 19775 2225 20000 2725
rect -200 2217 500 2225
rect -200 2183 -17 2217
rect 17 2183 500 2217
rect -200 2175 500 2183
rect 19200 2217 20000 2225
rect 19200 2183 19233 2217
rect 19267 2183 19783 2217
rect 19817 2183 20000 2217
rect 19200 2175 20000 2183
rect -200 1675 25 2175
rect 100 2090 450 2100
rect 100 1760 110 2090
rect 440 1760 450 2090
rect 100 1750 450 1760
rect 19225 1675 19275 2175
rect 19350 2090 19700 2100
rect 19350 1760 19360 2090
rect 19690 1760 19700 2090
rect 19350 1750 19700 1760
rect 19775 1675 20000 2175
rect 20090 1813 20210 1823
rect 20090 1713 20100 1813
rect 20200 1713 20210 1813
rect 20090 1703 20210 1713
rect -200 1667 500 1675
rect -200 1633 -17 1667
rect 17 1633 500 1667
rect -200 1625 500 1633
rect 19200 1667 20000 1675
rect 19200 1633 19233 1667
rect 19267 1633 19783 1667
rect 19817 1633 20000 1667
rect 19200 1625 20000 1633
rect -410 1587 -290 1597
rect -410 1487 -400 1587
rect -300 1487 -290 1587
rect -410 1477 -290 1487
rect -200 1125 25 1625
rect 100 1540 450 1550
rect 100 1210 110 1540
rect 440 1210 450 1540
rect 100 1200 450 1210
rect 19225 1125 19275 1625
rect 19350 1540 19700 1550
rect 19350 1210 19360 1540
rect 19690 1210 19700 1540
rect 19350 1200 19700 1210
rect 19775 1125 20000 1625
rect -200 1117 500 1125
rect -200 1083 -17 1117
rect 17 1083 500 1117
rect -200 1075 500 1083
rect 19200 1117 20000 1125
rect 19200 1083 19233 1117
rect 19267 1083 19783 1117
rect 19817 1083 20000 1117
rect 19200 1075 20000 1083
rect -200 575 25 1075
rect 100 990 450 1000
rect 100 660 110 990
rect 440 660 450 990
rect 100 650 450 660
rect 19225 575 19275 1075
rect 19350 990 19700 1000
rect 19350 660 19360 990
rect 19690 660 19700 990
rect 19350 650 19700 660
rect 19775 575 20000 1075
rect 20090 713 20210 723
rect 20090 613 20100 713
rect 20200 613 20210 713
rect 20090 603 20210 613
rect -200 567 500 575
rect -200 533 -17 567
rect 17 533 500 567
rect -200 525 500 533
rect 19200 567 20000 575
rect 19200 533 19233 567
rect 19267 533 19783 567
rect 19817 533 20000 567
rect 19200 525 20000 533
rect -410 487 -290 497
rect -410 387 -400 487
rect -300 387 -290 487
rect -410 377 -290 387
rect -200 25 25 525
rect 100 440 450 450
rect 100 110 110 440
rect 440 110 450 440
rect 100 100 450 110
rect 525 25 575 500
rect 650 440 1000 450
rect 650 110 660 440
rect 990 110 1000 440
rect 650 100 1000 110
rect 1075 25 1125 500
rect 1200 440 1550 450
rect 1200 110 1210 440
rect 1540 110 1550 440
rect 1200 100 1550 110
rect 1625 25 1675 500
rect 1750 440 2100 450
rect 1750 110 1760 440
rect 2090 110 2100 440
rect 1750 100 2100 110
rect 2175 25 2225 500
rect 2300 440 2650 450
rect 2300 110 2310 440
rect 2640 110 2650 440
rect 2300 100 2650 110
rect 2725 25 2775 500
rect 2850 440 3200 450
rect 2850 110 2860 440
rect 3190 110 3200 440
rect 2850 100 3200 110
rect 3275 25 3325 500
rect 3400 440 3750 450
rect 3400 110 3410 440
rect 3740 110 3750 440
rect 3400 100 3750 110
rect 3825 25 3875 500
rect 3950 440 4300 450
rect 3950 110 3960 440
rect 4290 110 4300 440
rect 3950 100 4300 110
rect 4375 25 4425 500
rect 4500 440 4850 450
rect 4500 110 4510 440
rect 4840 110 4850 440
rect 4500 100 4850 110
rect 4925 25 4975 500
rect 5050 440 5400 450
rect 5050 110 5060 440
rect 5390 110 5400 440
rect 5050 100 5400 110
rect 5475 25 5525 500
rect 5600 440 5950 450
rect 5600 110 5610 440
rect 5940 110 5950 440
rect 5600 100 5950 110
rect 6025 25 6075 500
rect 6150 440 6500 450
rect 6150 110 6160 440
rect 6490 110 6500 440
rect 6150 100 6500 110
rect 6575 25 6625 500
rect 6700 440 7050 450
rect 6700 110 6710 440
rect 7040 110 7050 440
rect 6700 100 7050 110
rect 7125 25 7175 500
rect 7250 440 7600 450
rect 7250 110 7260 440
rect 7590 110 7600 440
rect 7250 100 7600 110
rect 7675 25 7725 500
rect 7800 440 8150 450
rect 7800 110 7810 440
rect 8140 110 8150 440
rect 7800 100 8150 110
rect 8225 25 8275 500
rect 8350 440 8700 450
rect 8350 110 8360 440
rect 8690 110 8700 440
rect 8350 100 8700 110
rect 8775 25 8825 500
rect 8900 440 9250 450
rect 8900 110 8910 440
rect 9240 110 9250 440
rect 8900 100 9250 110
rect 9325 25 9375 500
rect 9450 440 9800 450
rect 9450 110 9460 440
rect 9790 110 9800 440
rect 9450 100 9800 110
rect 9875 25 9925 500
rect 10000 440 10350 450
rect 10000 110 10010 440
rect 10340 110 10350 440
rect 10000 100 10350 110
rect 10425 25 10475 500
rect 10550 440 10900 450
rect 10550 110 10560 440
rect 10890 110 10900 440
rect 10550 100 10900 110
rect 10975 25 11025 500
rect 11100 440 11450 450
rect 11100 110 11110 440
rect 11440 110 11450 440
rect 11100 100 11450 110
rect 11525 25 11575 500
rect 11650 440 12000 450
rect 11650 110 11660 440
rect 11990 110 12000 440
rect 11650 100 12000 110
rect 12075 25 12125 500
rect 12200 440 12550 450
rect 12200 110 12210 440
rect 12540 110 12550 440
rect 12200 100 12550 110
rect 12625 25 12675 500
rect 12750 440 13100 450
rect 12750 110 12760 440
rect 13090 110 13100 440
rect 12750 100 13100 110
rect 13175 25 13225 500
rect 13300 440 13650 450
rect 13300 110 13310 440
rect 13640 110 13650 440
rect 13300 100 13650 110
rect 13725 25 13775 500
rect 13850 440 14200 450
rect 13850 110 13860 440
rect 14190 110 14200 440
rect 13850 100 14200 110
rect 14275 25 14325 500
rect 14400 440 14750 450
rect 14400 110 14410 440
rect 14740 110 14750 440
rect 14400 100 14750 110
rect 14825 25 14875 500
rect 14950 440 15300 450
rect 14950 110 14960 440
rect 15290 110 15300 440
rect 14950 100 15300 110
rect 15375 25 15425 500
rect 15500 440 15850 450
rect 15500 110 15510 440
rect 15840 110 15850 440
rect 15500 100 15850 110
rect 15925 25 15975 500
rect 16050 440 16400 450
rect 16050 110 16060 440
rect 16390 110 16400 440
rect 16050 100 16400 110
rect 16475 25 16525 500
rect 16600 440 16950 450
rect 16600 110 16610 440
rect 16940 110 16950 440
rect 16600 100 16950 110
rect 17025 25 17075 500
rect 17150 440 17500 450
rect 17150 110 17160 440
rect 17490 110 17500 440
rect 17150 100 17500 110
rect 17575 25 17625 500
rect 17700 440 18050 450
rect 17700 110 17710 440
rect 18040 110 18050 440
rect 17700 100 18050 110
rect 18125 25 18175 500
rect 18250 440 18600 450
rect 18250 110 18260 440
rect 18590 110 18600 440
rect 18250 100 18600 110
rect 18675 25 18725 500
rect 18800 440 19150 450
rect 18800 110 18810 440
rect 19140 110 19150 440
rect 18800 100 19150 110
rect 19225 25 19275 525
rect 19350 440 19700 450
rect 19350 110 19360 440
rect 19690 110 19700 440
rect 19350 100 19700 110
rect 19775 25 20000 525
rect -200 17 20000 25
rect -200 -17 -17 17
rect 17 -17 533 17
rect 567 -17 1083 17
rect 1117 -17 1633 17
rect 1667 -17 2183 17
rect 2217 -17 2733 17
rect 2767 -17 3283 17
rect 3317 -17 3833 17
rect 3867 -17 4383 17
rect 4417 -17 4933 17
rect 4967 -17 5483 17
rect 5517 -17 6033 17
rect 6067 -17 6583 17
rect 6617 -17 7133 17
rect 7167 -17 7683 17
rect 7717 -17 8233 17
rect 8267 -17 8783 17
rect 8817 -17 9333 17
rect 9367 -17 9883 17
rect 9917 -17 10433 17
rect 10467 -17 10983 17
rect 11017 -17 11533 17
rect 11567 -17 12083 17
rect 12117 -17 12633 17
rect 12667 -17 13183 17
rect 13217 -17 13733 17
rect 13767 -17 14283 17
rect 14317 -17 14833 17
rect 14867 -17 15383 17
rect 15417 -17 15933 17
rect 15967 -17 16483 17
rect 16517 -17 17033 17
rect 17067 -17 17583 17
rect 17617 -17 18133 17
rect 18167 -17 18683 17
rect 18717 -17 19233 17
rect 19267 -17 19783 17
rect 19817 -17 20000 17
rect -200 -200 20000 -17
rect 377 -300 497 -290
rect 377 -400 387 -300
rect 487 -400 497 -300
rect 377 -410 497 -400
rect 1477 -300 1597 -290
rect 1477 -400 1487 -300
rect 1587 -400 1597 -300
rect 1477 -410 1597 -400
rect 2577 -300 2697 -290
rect 2577 -400 2587 -300
rect 2687 -400 2697 -300
rect 2577 -410 2697 -400
rect 3677 -300 3797 -290
rect 3677 -400 3687 -300
rect 3787 -400 3797 -300
rect 3677 -410 3797 -400
rect 4777 -300 4897 -290
rect 4777 -400 4787 -300
rect 4887 -400 4897 -300
rect 4777 -410 4897 -400
rect 5877 -300 5997 -290
rect 5877 -400 5887 -300
rect 5987 -400 5997 -300
rect 5877 -410 5997 -400
rect 6977 -300 7097 -290
rect 6977 -400 6987 -300
rect 7087 -400 7097 -300
rect 6977 -410 7097 -400
rect 8077 -300 8197 -290
rect 8077 -400 8087 -300
rect 8187 -400 8197 -300
rect 8077 -410 8197 -400
rect 9177 -300 9297 -290
rect 9177 -400 9187 -300
rect 9287 -400 9297 -300
rect 9177 -410 9297 -400
rect 10277 -300 10397 -290
rect 10277 -400 10287 -300
rect 10387 -400 10397 -300
rect 10277 -410 10397 -400
rect 11377 -300 11497 -290
rect 11377 -400 11387 -300
rect 11487 -400 11497 -300
rect 11377 -410 11497 -400
rect 12477 -300 12597 -290
rect 12477 -400 12487 -300
rect 12587 -400 12597 -300
rect 12477 -410 12597 -400
rect 13577 -300 13697 -290
rect 13577 -400 13587 -300
rect 13687 -400 13697 -300
rect 13577 -410 13697 -400
rect 14677 -300 14797 -290
rect 14677 -400 14687 -300
rect 14787 -400 14797 -300
rect 14677 -410 14797 -400
rect 15777 -300 15897 -290
rect 15777 -400 15787 -300
rect 15887 -400 15897 -300
rect 15777 -410 15897 -400
rect 16877 -300 16997 -290
rect 16877 -400 16887 -300
rect 16987 -400 16997 -300
rect 16877 -410 16997 -400
rect 17977 -300 18097 -290
rect 17977 -400 17987 -300
rect 18087 -400 18097 -300
rect 17977 -410 18097 -400
rect 19077 -300 19197 -290
rect 19077 -400 19087 -300
rect 19187 -400 19197 -300
rect 19077 -410 19197 -400
rect 20800 -1000 20812 20800
rect 30 -1012 20812 -1000
rect 24788 -4988 24800 24788
rect 30 -5000 24800 -4988
<< via2 >>
rect 613 20100 713 20200
rect 1713 20100 1813 20200
rect 2813 20100 2913 20200
rect 3913 20100 4013 20200
rect 5013 20100 5113 20200
rect 6113 20100 6213 20200
rect 7213 20100 7313 20200
rect 8313 20100 8413 20200
rect 9413 20100 9513 20200
rect 10513 20100 10613 20200
rect 11613 20100 11713 20200
rect 12713 20100 12813 20200
rect 13813 20100 13913 20200
rect 14913 20100 15013 20200
rect 16013 20100 16113 20200
rect 17113 20100 17213 20200
rect 18213 20100 18313 20200
rect 19313 20100 19413 20200
rect 215 19465 335 19585
rect 765 19465 885 19585
rect 1315 19465 1435 19585
rect 1865 19465 1985 19585
rect 2415 19465 2535 19585
rect 2965 19465 3085 19585
rect 3515 19465 3635 19585
rect 4065 19465 4185 19585
rect 4615 19465 4735 19585
rect 5165 19465 5285 19585
rect 5715 19465 5835 19585
rect 6265 19465 6385 19585
rect 6815 19465 6935 19585
rect 7365 19465 7485 19585
rect 7915 19465 8035 19585
rect 8465 19465 8585 19585
rect 9015 19465 9135 19585
rect 9565 19465 9685 19585
rect 10115 19465 10235 19585
rect 10665 19465 10785 19585
rect 11215 19465 11335 19585
rect 11765 19465 11885 19585
rect 12315 19465 12435 19585
rect 12865 19465 12985 19585
rect 13415 19465 13535 19585
rect 13965 19465 14085 19585
rect 14515 19465 14635 19585
rect 15065 19465 15185 19585
rect 15615 19465 15735 19585
rect 16165 19465 16285 19585
rect 16715 19465 16835 19585
rect 17265 19465 17385 19585
rect 17815 19465 17935 19585
rect 18365 19465 18485 19585
rect 18915 19465 19035 19585
rect 19465 19465 19585 19585
rect 20100 19313 20200 19413
rect -400 19087 -300 19187
rect 215 18915 335 19035
rect 19465 18915 19585 19035
rect 215 18365 335 18485
rect 19465 18365 19585 18485
rect 20100 18213 20200 18313
rect -400 17987 -300 18087
rect 215 17815 335 17935
rect 19465 17815 19585 17935
rect 215 17265 335 17385
rect 19465 17265 19585 17385
rect 20100 17113 20200 17213
rect -400 16887 -300 16987
rect 215 16715 335 16835
rect 19465 16715 19585 16835
rect 215 16165 335 16285
rect 19465 16165 19585 16285
rect 20100 16013 20200 16113
rect -400 15787 -300 15887
rect 215 15615 335 15735
rect 19465 15615 19585 15735
rect 215 15065 335 15185
rect 19465 15065 19585 15185
rect 20100 14913 20200 15013
rect -400 14687 -300 14787
rect 215 14515 335 14635
rect 19465 14515 19585 14635
rect 215 13965 335 14085
rect 19465 13965 19585 14085
rect 20100 13813 20200 13913
rect -400 13587 -300 13687
rect 215 13415 335 13535
rect 19465 13415 19585 13535
rect 215 12865 335 12985
rect 19465 12865 19585 12985
rect 20100 12713 20200 12813
rect -400 12487 -300 12587
rect 215 12315 335 12435
rect 19465 12315 19585 12435
rect 215 11765 335 11885
rect 19465 11765 19585 11885
rect 20100 11613 20200 11713
rect -400 11387 -300 11487
rect 215 11215 335 11335
rect 19465 11215 19585 11335
rect 215 10665 335 10785
rect 19465 10665 19585 10785
rect 20100 10513 20200 10613
rect -400 10287 -300 10387
rect 215 10115 335 10235
rect 19465 10115 19585 10235
rect 215 9565 335 9685
rect 19465 9565 19585 9685
rect 20100 9413 20200 9513
rect -400 9187 -300 9287
rect 215 9015 335 9135
rect 19465 9015 19585 9135
rect 215 8465 335 8585
rect 19465 8465 19585 8585
rect 20100 8313 20200 8413
rect -400 8087 -300 8187
rect 215 7915 335 8035
rect 19465 7915 19585 8035
rect 215 7365 335 7485
rect 19465 7365 19585 7485
rect 20100 7213 20200 7313
rect -400 6987 -300 7087
rect 215 6815 335 6935
rect 19465 6815 19585 6935
rect 215 6265 335 6385
rect 19465 6265 19585 6385
rect 20100 6113 20200 6213
rect -400 5887 -300 5987
rect 215 5715 335 5835
rect 19465 5715 19585 5835
rect 215 5165 335 5285
rect 19465 5165 19585 5285
rect 20100 5013 20200 5113
rect -400 4787 -300 4887
rect 215 4615 335 4735
rect 19465 4615 19585 4735
rect 215 4065 335 4185
rect 19465 4065 19585 4185
rect 20100 3913 20200 4013
rect -400 3687 -300 3787
rect 215 3515 335 3635
rect 19465 3515 19585 3635
rect 215 2965 335 3085
rect 19465 2965 19585 3085
rect 20100 2813 20200 2913
rect -400 2587 -300 2687
rect 215 2415 335 2535
rect 19465 2415 19585 2535
rect 215 1865 335 1985
rect 19465 1865 19585 1985
rect 20100 1713 20200 1813
rect -400 1487 -300 1587
rect 215 1315 335 1435
rect 19465 1315 19585 1435
rect 215 765 335 885
rect 19465 765 19585 885
rect 20100 613 20200 713
rect -400 387 -300 487
rect 215 215 335 335
rect 765 215 885 335
rect 1315 215 1435 335
rect 1865 215 1985 335
rect 2415 215 2535 335
rect 2965 215 3085 335
rect 3515 215 3635 335
rect 4065 215 4185 335
rect 4615 215 4735 335
rect 5165 215 5285 335
rect 5715 215 5835 335
rect 6265 215 6385 335
rect 6815 215 6935 335
rect 7365 215 7485 335
rect 7915 215 8035 335
rect 8465 215 8585 335
rect 9015 215 9135 335
rect 9565 215 9685 335
rect 10115 215 10235 335
rect 10665 215 10785 335
rect 11215 215 11335 335
rect 11765 215 11885 335
rect 12315 215 12435 335
rect 12865 215 12985 335
rect 13415 215 13535 335
rect 13965 215 14085 335
rect 14515 215 14635 335
rect 15065 215 15185 335
rect 15615 215 15735 335
rect 16165 215 16285 335
rect 16715 215 16835 335
rect 17265 215 17385 335
rect 17815 215 17935 335
rect 18365 215 18485 335
rect 18915 215 19035 335
rect 19465 215 19585 335
rect 387 -400 487 -300
rect 1487 -400 1587 -300
rect 2587 -400 2687 -300
rect 3687 -400 3787 -300
rect 4787 -400 4887 -300
rect 5887 -400 5987 -300
rect 6987 -400 7087 -300
rect 8087 -400 8187 -300
rect 9187 -400 9287 -300
rect 10287 -400 10387 -300
rect 11387 -400 11487 -300
rect 12487 -400 12587 -300
rect 13587 -400 13687 -300
rect 14687 -400 14787 -300
rect 15787 -400 15887 -300
rect 16887 -400 16987 -300
rect 17987 -400 18087 -300
rect 19087 -400 19187 -300
<< metal3 >>
rect -2000 20800 19800 21800
rect -2000 19913 -1000 20800
rect -113 19913 339 20800
rect -2000 19589 339 19913
rect 437 20200 889 20300
rect 437 20100 613 20200
rect 713 20100 889 20200
rect 437 19687 889 20100
rect 987 19687 1439 20800
rect 1537 20200 1989 20300
rect 1537 20100 1713 20200
rect 1813 20100 1989 20200
rect 1537 19687 1989 20100
rect 2087 19687 2539 20800
rect 2637 20200 3089 20300
rect 2637 20100 2813 20200
rect 2913 20100 3089 20200
rect 2637 19687 3089 20100
rect 3187 19687 3639 20800
rect 3737 20200 4189 20300
rect 3737 20100 3913 20200
rect 4013 20100 4189 20200
rect 3737 19687 4189 20100
rect 4287 19687 4739 20800
rect 4837 20200 5289 20300
rect 4837 20100 5013 20200
rect 5113 20100 5289 20200
rect 4837 19687 5289 20100
rect 5387 19687 5839 20800
rect 5937 20200 6389 20300
rect 5937 20100 6113 20200
rect 6213 20100 6389 20200
rect 5937 19687 6389 20100
rect 6487 19687 6939 20800
rect 7037 20200 7489 20300
rect 7037 20100 7213 20200
rect 7313 20100 7489 20200
rect 7037 19687 7489 20100
rect 7587 19687 8039 20800
rect 8137 20200 8589 20300
rect 8137 20100 8313 20200
rect 8413 20100 8589 20200
rect 8137 19687 8589 20100
rect 8687 19687 9139 20800
rect 9237 20200 9689 20300
rect 9237 20100 9413 20200
rect 9513 20100 9689 20200
rect 9237 19687 9689 20100
rect 9787 19687 10239 20800
rect 10337 20200 10789 20300
rect 10337 20100 10513 20200
rect 10613 20100 10789 20200
rect 10337 19687 10789 20100
rect 10887 19687 11339 20800
rect 11437 20200 11889 20300
rect 11437 20100 11613 20200
rect 11713 20100 11889 20200
rect 11437 19687 11889 20100
rect 11987 19687 12439 20800
rect 12537 20200 12989 20300
rect 12537 20100 12713 20200
rect 12813 20100 12989 20200
rect 12537 19687 12989 20100
rect 13087 19687 13539 20800
rect 13637 20200 14089 20300
rect 13637 20100 13813 20200
rect 13913 20100 14089 20200
rect 13637 19687 14089 20100
rect 14187 19687 14639 20800
rect 14737 20200 15189 20300
rect 14737 20100 14913 20200
rect 15013 20100 15189 20200
rect 14737 19687 15189 20100
rect 15287 19687 15739 20800
rect 15837 20200 16289 20300
rect 15837 20100 16013 20200
rect 16113 20100 16289 20200
rect 15837 19687 16289 20100
rect 16387 19687 16839 20800
rect 16937 20200 17389 20300
rect 16937 20100 17113 20200
rect 17213 20100 17389 20200
rect 16937 19687 17389 20100
rect 17487 19687 17939 20800
rect 18037 20200 18489 20300
rect 18037 20100 18213 20200
rect 18313 20100 18489 20200
rect 18037 19687 18489 20100
rect 18587 19687 19039 20800
rect 19137 20200 19589 20300
rect 19137 20100 19313 20200
rect 19413 20100 19589 20200
rect 19137 19687 19589 20100
tri 339 19589 437 19687 sw
tri 437 19589 535 19687 ne
rect 535 19589 889 19687
tri 889 19589 987 19687 sw
tri 987 19589 1085 19687 ne
rect 1085 19589 1439 19687
tri 1439 19589 1537 19687 sw
tri 1537 19589 1635 19687 ne
rect 1635 19589 1989 19687
tri 1989 19589 2087 19687 sw
tri 2087 19589 2185 19687 ne
rect 2185 19589 2539 19687
tri 2539 19589 2637 19687 sw
tri 2637 19589 2735 19687 ne
rect 2735 19589 3089 19687
tri 3089 19589 3187 19687 sw
tri 3187 19589 3285 19687 ne
rect 3285 19589 3639 19687
tri 3639 19589 3737 19687 sw
tri 3737 19589 3835 19687 ne
rect 3835 19589 4189 19687
tri 4189 19589 4287 19687 sw
tri 4287 19589 4385 19687 ne
rect 4385 19589 4739 19687
tri 4739 19589 4837 19687 sw
tri 4837 19589 4935 19687 ne
rect 4935 19589 5289 19687
tri 5289 19589 5387 19687 sw
tri 5387 19589 5485 19687 ne
rect 5485 19589 5839 19687
tri 5839 19589 5937 19687 sw
tri 5937 19589 6035 19687 ne
rect 6035 19589 6389 19687
tri 6389 19589 6487 19687 sw
tri 6487 19589 6585 19687 ne
rect 6585 19589 6939 19687
tri 6939 19589 7037 19687 sw
tri 7037 19589 7135 19687 ne
rect 7135 19589 7489 19687
tri 7489 19589 7587 19687 sw
tri 7587 19589 7685 19687 ne
rect 7685 19589 8039 19687
tri 8039 19589 8137 19687 sw
tri 8137 19589 8235 19687 ne
rect 8235 19589 8589 19687
tri 8589 19589 8687 19687 sw
tri 8687 19589 8785 19687 ne
rect 8785 19589 9139 19687
tri 9139 19589 9237 19687 sw
tri 9237 19589 9335 19687 ne
rect 9335 19589 9689 19687
tri 9689 19589 9787 19687 sw
tri 9787 19589 9885 19687 ne
rect 9885 19589 10239 19687
tri 10239 19589 10337 19687 sw
tri 10337 19589 10435 19687 ne
rect 10435 19589 10789 19687
tri 10789 19589 10887 19687 sw
tri 10887 19589 10985 19687 ne
rect 10985 19589 11339 19687
tri 11339 19589 11437 19687 sw
tri 11437 19589 11535 19687 ne
rect 11535 19589 11889 19687
tri 11889 19589 11987 19687 sw
tri 11987 19589 12085 19687 ne
rect 12085 19589 12439 19687
tri 12439 19589 12537 19687 sw
tri 12537 19589 12635 19687 ne
rect 12635 19589 12989 19687
tri 12989 19589 13087 19687 sw
tri 13087 19589 13185 19687 ne
rect 13185 19589 13539 19687
tri 13539 19589 13637 19687 sw
tri 13637 19589 13735 19687 ne
rect 13735 19589 14089 19687
tri 14089 19589 14187 19687 sw
tri 14187 19589 14285 19687 ne
rect 14285 19589 14639 19687
tri 14639 19589 14737 19687 sw
tri 14737 19589 14835 19687 ne
rect 14835 19589 15189 19687
tri 15189 19589 15287 19687 sw
tri 15287 19589 15385 19687 ne
rect 15385 19589 15739 19687
tri 15739 19589 15837 19687 sw
tri 15837 19589 15935 19687 ne
rect 15935 19589 16289 19687
tri 16289 19589 16387 19687 sw
tri 16387 19589 16485 19687 ne
rect 16485 19589 16839 19687
tri 16839 19589 16937 19687 sw
tri 16937 19589 17035 19687 ne
rect 17035 19589 17389 19687
tri 17389 19589 17487 19687 sw
tri 17487 19589 17585 19687 ne
rect 17585 19589 17939 19687
tri 17939 19589 18037 19687 sw
tri 18037 19589 18135 19687 ne
rect 18135 19589 18489 19687
tri 18489 19589 18587 19687 sw
tri 18587 19589 18685 19687 ne
rect 18685 19589 19039 19687
tri 19039 19589 19137 19687 sw
tri 19137 19589 19235 19687 ne
rect 19235 19589 19589 19687
tri 19589 19589 19687 19687 sw
rect 20800 19589 21800 19800
rect -2000 19585 437 19589
rect -2000 19465 215 19585
rect 335 19491 437 19585
tri 437 19491 535 19589 sw
tri 535 19491 633 19589 ne
rect 633 19585 987 19589
rect 633 19491 765 19585
rect 335 19465 535 19491
rect -2000 19461 535 19465
rect -2000 18813 -1000 19461
tri 113 19363 211 19461 ne
rect 211 19413 535 19461
tri 535 19413 613 19491 sw
tri 633 19413 711 19491 ne
rect 711 19465 765 19491
rect 885 19491 987 19585
tri 987 19491 1085 19589 sw
tri 1085 19491 1183 19589 ne
rect 1183 19585 1537 19589
rect 1183 19491 1315 19585
rect 885 19465 1085 19491
rect 711 19413 1085 19465
tri 1085 19413 1163 19491 sw
tri 1183 19413 1261 19491 ne
rect 1261 19465 1315 19491
rect 1435 19491 1537 19585
tri 1537 19491 1635 19589 sw
tri 1635 19491 1733 19589 ne
rect 1733 19585 2087 19589
rect 1733 19491 1865 19585
rect 1435 19465 1635 19491
rect 1261 19413 1635 19465
tri 1635 19413 1713 19491 sw
tri 1733 19413 1811 19491 ne
rect 1811 19465 1865 19491
rect 1985 19491 2087 19585
tri 2087 19491 2185 19589 sw
tri 2185 19491 2283 19589 ne
rect 2283 19585 2637 19589
rect 2283 19491 2415 19585
rect 1985 19465 2185 19491
rect 1811 19413 2185 19465
tri 2185 19413 2263 19491 sw
tri 2283 19413 2361 19491 ne
rect 2361 19465 2415 19491
rect 2535 19491 2637 19585
tri 2637 19491 2735 19589 sw
tri 2735 19491 2833 19589 ne
rect 2833 19585 3187 19589
rect 2833 19491 2965 19585
rect 2535 19465 2735 19491
rect 2361 19413 2735 19465
tri 2735 19413 2813 19491 sw
tri 2833 19413 2911 19491 ne
rect 2911 19465 2965 19491
rect 3085 19491 3187 19585
tri 3187 19491 3285 19589 sw
tri 3285 19491 3383 19589 ne
rect 3383 19585 3737 19589
rect 3383 19491 3515 19585
rect 3085 19465 3285 19491
rect 2911 19413 3285 19465
tri 3285 19413 3363 19491 sw
tri 3383 19413 3461 19491 ne
rect 3461 19465 3515 19491
rect 3635 19491 3737 19585
tri 3737 19491 3835 19589 sw
tri 3835 19491 3933 19589 ne
rect 3933 19585 4287 19589
rect 3933 19491 4065 19585
rect 3635 19465 3835 19491
rect 3461 19413 3835 19465
tri 3835 19413 3913 19491 sw
tri 3933 19413 4011 19491 ne
rect 4011 19465 4065 19491
rect 4185 19491 4287 19585
tri 4287 19491 4385 19589 sw
tri 4385 19491 4483 19589 ne
rect 4483 19585 4837 19589
rect 4483 19491 4615 19585
rect 4185 19465 4385 19491
rect 4011 19413 4385 19465
tri 4385 19413 4463 19491 sw
tri 4483 19413 4561 19491 ne
rect 4561 19465 4615 19491
rect 4735 19491 4837 19585
tri 4837 19491 4935 19589 sw
tri 4935 19491 5033 19589 ne
rect 5033 19585 5387 19589
rect 5033 19491 5165 19585
rect 4735 19465 4935 19491
rect 4561 19413 4935 19465
tri 4935 19413 5013 19491 sw
tri 5033 19413 5111 19491 ne
rect 5111 19465 5165 19491
rect 5285 19491 5387 19585
tri 5387 19491 5485 19589 sw
tri 5485 19491 5583 19589 ne
rect 5583 19585 5937 19589
rect 5583 19491 5715 19585
rect 5285 19465 5485 19491
rect 5111 19413 5485 19465
tri 5485 19413 5563 19491 sw
tri 5583 19413 5661 19491 ne
rect 5661 19465 5715 19491
rect 5835 19491 5937 19585
tri 5937 19491 6035 19589 sw
tri 6035 19491 6133 19589 ne
rect 6133 19585 6487 19589
rect 6133 19491 6265 19585
rect 5835 19465 6035 19491
rect 5661 19413 6035 19465
tri 6035 19413 6113 19491 sw
tri 6133 19413 6211 19491 ne
rect 6211 19465 6265 19491
rect 6385 19491 6487 19585
tri 6487 19491 6585 19589 sw
tri 6585 19491 6683 19589 ne
rect 6683 19585 7037 19589
rect 6683 19491 6815 19585
rect 6385 19465 6585 19491
rect 6211 19413 6585 19465
tri 6585 19413 6663 19491 sw
tri 6683 19413 6761 19491 ne
rect 6761 19465 6815 19491
rect 6935 19491 7037 19585
tri 7037 19491 7135 19589 sw
tri 7135 19491 7233 19589 ne
rect 7233 19585 7587 19589
rect 7233 19491 7365 19585
rect 6935 19465 7135 19491
rect 6761 19413 7135 19465
tri 7135 19413 7213 19491 sw
tri 7233 19413 7311 19491 ne
rect 7311 19465 7365 19491
rect 7485 19491 7587 19585
tri 7587 19491 7685 19589 sw
tri 7685 19491 7783 19589 ne
rect 7783 19585 8137 19589
rect 7783 19491 7915 19585
rect 7485 19465 7685 19491
rect 7311 19413 7685 19465
tri 7685 19413 7763 19491 sw
tri 7783 19413 7861 19491 ne
rect 7861 19465 7915 19491
rect 8035 19491 8137 19585
tri 8137 19491 8235 19589 sw
tri 8235 19491 8333 19589 ne
rect 8333 19585 8687 19589
rect 8333 19491 8465 19585
rect 8035 19465 8235 19491
rect 7861 19413 8235 19465
tri 8235 19413 8313 19491 sw
tri 8333 19413 8411 19491 ne
rect 8411 19465 8465 19491
rect 8585 19491 8687 19585
tri 8687 19491 8785 19589 sw
tri 8785 19491 8883 19589 ne
rect 8883 19585 9237 19589
rect 8883 19491 9015 19585
rect 8585 19465 8785 19491
rect 8411 19413 8785 19465
tri 8785 19413 8863 19491 sw
tri 8883 19413 8961 19491 ne
rect 8961 19465 9015 19491
rect 9135 19491 9237 19585
tri 9237 19491 9335 19589 sw
tri 9335 19491 9433 19589 ne
rect 9433 19585 9787 19589
rect 9433 19491 9565 19585
rect 9135 19465 9335 19491
rect 8961 19413 9335 19465
tri 9335 19413 9413 19491 sw
tri 9433 19413 9511 19491 ne
rect 9511 19465 9565 19491
rect 9685 19491 9787 19585
tri 9787 19491 9885 19589 sw
tri 9885 19491 9983 19589 ne
rect 9983 19585 10337 19589
rect 9983 19491 10115 19585
rect 9685 19465 9885 19491
rect 9511 19413 9885 19465
tri 9885 19413 9963 19491 sw
tri 9983 19413 10061 19491 ne
rect 10061 19465 10115 19491
rect 10235 19491 10337 19585
tri 10337 19491 10435 19589 sw
tri 10435 19491 10533 19589 ne
rect 10533 19585 10887 19589
rect 10533 19491 10665 19585
rect 10235 19465 10435 19491
rect 10061 19413 10435 19465
tri 10435 19413 10513 19491 sw
tri 10533 19413 10611 19491 ne
rect 10611 19465 10665 19491
rect 10785 19491 10887 19585
tri 10887 19491 10985 19589 sw
tri 10985 19491 11083 19589 ne
rect 11083 19585 11437 19589
rect 11083 19491 11215 19585
rect 10785 19465 10985 19491
rect 10611 19413 10985 19465
tri 10985 19413 11063 19491 sw
tri 11083 19413 11161 19491 ne
rect 11161 19465 11215 19491
rect 11335 19491 11437 19585
tri 11437 19491 11535 19589 sw
tri 11535 19491 11633 19589 ne
rect 11633 19585 11987 19589
rect 11633 19491 11765 19585
rect 11335 19465 11535 19491
rect 11161 19413 11535 19465
tri 11535 19413 11613 19491 sw
tri 11633 19413 11711 19491 ne
rect 11711 19465 11765 19491
rect 11885 19491 11987 19585
tri 11987 19491 12085 19589 sw
tri 12085 19491 12183 19589 ne
rect 12183 19585 12537 19589
rect 12183 19491 12315 19585
rect 11885 19465 12085 19491
rect 11711 19413 12085 19465
tri 12085 19413 12163 19491 sw
tri 12183 19413 12261 19491 ne
rect 12261 19465 12315 19491
rect 12435 19491 12537 19585
tri 12537 19491 12635 19589 sw
tri 12635 19491 12733 19589 ne
rect 12733 19585 13087 19589
rect 12733 19491 12865 19585
rect 12435 19465 12635 19491
rect 12261 19413 12635 19465
tri 12635 19413 12713 19491 sw
tri 12733 19413 12811 19491 ne
rect 12811 19465 12865 19491
rect 12985 19491 13087 19585
tri 13087 19491 13185 19589 sw
tri 13185 19491 13283 19589 ne
rect 13283 19585 13637 19589
rect 13283 19491 13415 19585
rect 12985 19465 13185 19491
rect 12811 19413 13185 19465
tri 13185 19413 13263 19491 sw
tri 13283 19413 13361 19491 ne
rect 13361 19465 13415 19491
rect 13535 19491 13637 19585
tri 13637 19491 13735 19589 sw
tri 13735 19491 13833 19589 ne
rect 13833 19585 14187 19589
rect 13833 19491 13965 19585
rect 13535 19465 13735 19491
rect 13361 19413 13735 19465
tri 13735 19413 13813 19491 sw
tri 13833 19413 13911 19491 ne
rect 13911 19465 13965 19491
rect 14085 19491 14187 19585
tri 14187 19491 14285 19589 sw
tri 14285 19491 14383 19589 ne
rect 14383 19585 14737 19589
rect 14383 19491 14515 19585
rect 14085 19465 14285 19491
rect 13911 19413 14285 19465
tri 14285 19413 14363 19491 sw
tri 14383 19413 14461 19491 ne
rect 14461 19465 14515 19491
rect 14635 19491 14737 19585
tri 14737 19491 14835 19589 sw
tri 14835 19491 14933 19589 ne
rect 14933 19585 15287 19589
rect 14933 19491 15065 19585
rect 14635 19465 14835 19491
rect 14461 19413 14835 19465
tri 14835 19413 14913 19491 sw
tri 14933 19413 15011 19491 ne
rect 15011 19465 15065 19491
rect 15185 19491 15287 19585
tri 15287 19491 15385 19589 sw
tri 15385 19491 15483 19589 ne
rect 15483 19585 15837 19589
rect 15483 19491 15615 19585
rect 15185 19465 15385 19491
rect 15011 19413 15385 19465
tri 15385 19413 15463 19491 sw
tri 15483 19413 15561 19491 ne
rect 15561 19465 15615 19491
rect 15735 19491 15837 19585
tri 15837 19491 15935 19589 sw
tri 15935 19491 16033 19589 ne
rect 16033 19585 16387 19589
rect 16033 19491 16165 19585
rect 15735 19465 15935 19491
rect 15561 19413 15935 19465
tri 15935 19413 16013 19491 sw
tri 16033 19413 16111 19491 ne
rect 16111 19465 16165 19491
rect 16285 19491 16387 19585
tri 16387 19491 16485 19589 sw
tri 16485 19491 16583 19589 ne
rect 16583 19585 16937 19589
rect 16583 19491 16715 19585
rect 16285 19465 16485 19491
rect 16111 19413 16485 19465
tri 16485 19413 16563 19491 sw
tri 16583 19413 16661 19491 ne
rect 16661 19465 16715 19491
rect 16835 19491 16937 19585
tri 16937 19491 17035 19589 sw
tri 17035 19491 17133 19589 ne
rect 17133 19585 17487 19589
rect 17133 19491 17265 19585
rect 16835 19465 17035 19491
rect 16661 19413 17035 19465
tri 17035 19413 17113 19491 sw
tri 17133 19413 17211 19491 ne
rect 17211 19465 17265 19491
rect 17385 19491 17487 19585
tri 17487 19491 17585 19589 sw
tri 17585 19491 17683 19589 ne
rect 17683 19585 18037 19589
rect 17683 19491 17815 19585
rect 17385 19465 17585 19491
rect 17211 19413 17585 19465
tri 17585 19413 17663 19491 sw
tri 17683 19413 17761 19491 ne
rect 17761 19465 17815 19491
rect 17935 19491 18037 19585
tri 18037 19491 18135 19589 sw
tri 18135 19491 18233 19589 ne
rect 18233 19585 18587 19589
rect 18233 19491 18365 19585
rect 17935 19465 18135 19491
rect 17761 19413 18135 19465
tri 18135 19413 18213 19491 sw
tri 18233 19413 18311 19491 ne
rect 18311 19465 18365 19491
rect 18485 19491 18587 19585
tri 18587 19491 18685 19589 sw
tri 18685 19491 18783 19589 ne
rect 18783 19585 19137 19589
rect 18783 19491 18915 19585
rect 18485 19465 18685 19491
rect 18311 19413 18685 19465
tri 18685 19413 18763 19491 sw
tri 18783 19413 18861 19491 ne
rect 18861 19465 18915 19491
rect 19035 19491 19137 19585
tri 19137 19491 19235 19589 sw
tri 19235 19491 19333 19589 ne
rect 19333 19585 21800 19589
rect 19333 19491 19465 19585
rect 19035 19465 19235 19491
rect 18861 19413 19235 19465
tri 19235 19413 19313 19491 sw
tri 19333 19413 19411 19491 ne
rect 19411 19465 19465 19491
rect 19585 19465 21800 19585
rect 19411 19413 21800 19465
rect 211 19363 613 19413
rect -500 19313 113 19363
tri 113 19313 163 19363 sw
tri 211 19313 261 19363 ne
rect 261 19333 613 19363
tri 613 19333 693 19413 sw
tri 711 19333 791 19413 ne
rect 791 19333 1163 19413
tri 1163 19333 1243 19413 sw
tri 1261 19333 1341 19413 ne
rect 1341 19333 1713 19413
tri 1713 19333 1793 19413 sw
tri 1811 19333 1891 19413 ne
rect 1891 19333 2263 19413
tri 2263 19333 2343 19413 sw
tri 2361 19333 2441 19413 ne
rect 2441 19333 2813 19413
tri 2813 19333 2893 19413 sw
tri 2911 19333 2991 19413 ne
rect 2991 19333 3363 19413
tri 3363 19333 3443 19413 sw
tri 3461 19333 3541 19413 ne
rect 3541 19333 3913 19413
tri 3913 19333 3993 19413 sw
tri 4011 19333 4091 19413 ne
rect 4091 19333 4463 19413
tri 4463 19333 4543 19413 sw
tri 4561 19333 4641 19413 ne
rect 4641 19333 5013 19413
tri 5013 19333 5093 19413 sw
tri 5111 19333 5191 19413 ne
rect 5191 19333 5563 19413
tri 5563 19333 5643 19413 sw
tri 5661 19333 5741 19413 ne
rect 5741 19333 6113 19413
tri 6113 19333 6193 19413 sw
tri 6211 19333 6291 19413 ne
rect 6291 19333 6663 19413
tri 6663 19333 6743 19413 sw
tri 6761 19333 6841 19413 ne
rect 6841 19333 7213 19413
tri 7213 19333 7293 19413 sw
tri 7311 19333 7391 19413 ne
rect 7391 19333 7763 19413
tri 7763 19333 7843 19413 sw
tri 7861 19333 7941 19413 ne
rect 7941 19333 8313 19413
tri 8313 19333 8393 19413 sw
tri 8411 19333 8491 19413 ne
rect 8491 19333 8863 19413
tri 8863 19333 8943 19413 sw
tri 8961 19333 9041 19413 ne
rect 9041 19333 9413 19413
tri 9413 19333 9493 19413 sw
tri 9511 19333 9591 19413 ne
rect 9591 19333 9963 19413
tri 9963 19333 10043 19413 sw
tri 10061 19333 10141 19413 ne
rect 10141 19333 10513 19413
tri 10513 19333 10593 19413 sw
tri 10611 19333 10691 19413 ne
rect 10691 19333 11063 19413
tri 11063 19333 11143 19413 sw
tri 11161 19333 11241 19413 ne
rect 11241 19333 11613 19413
tri 11613 19333 11693 19413 sw
tri 11711 19333 11791 19413 ne
rect 11791 19333 12163 19413
tri 12163 19333 12243 19413 sw
tri 12261 19333 12341 19413 ne
rect 12341 19333 12713 19413
tri 12713 19333 12793 19413 sw
tri 12811 19333 12891 19413 ne
rect 12891 19333 13263 19413
tri 13263 19333 13343 19413 sw
tri 13361 19333 13441 19413 ne
rect 13441 19333 13813 19413
tri 13813 19333 13893 19413 sw
tri 13911 19333 13991 19413 ne
rect 13991 19333 14363 19413
tri 14363 19333 14443 19413 sw
tri 14461 19333 14541 19413 ne
rect 14541 19333 14913 19413
tri 14913 19333 14993 19413 sw
tri 15011 19333 15091 19413 ne
rect 15091 19333 15463 19413
tri 15463 19333 15543 19413 sw
tri 15561 19333 15641 19413 ne
rect 15641 19333 16013 19413
tri 16013 19333 16093 19413 sw
tri 16111 19333 16191 19413 ne
rect 16191 19333 16563 19413
tri 16563 19333 16643 19413 sw
tri 16661 19333 16741 19413 ne
rect 16741 19333 17113 19413
tri 17113 19333 17193 19413 sw
tri 17211 19333 17291 19413 ne
rect 17291 19333 17663 19413
tri 17663 19333 17743 19413 sw
tri 17761 19333 17841 19413 ne
rect 17841 19333 18213 19413
tri 18213 19333 18293 19413 sw
tri 18311 19333 18391 19413 ne
rect 18391 19333 18763 19413
tri 18763 19333 18843 19413 sw
tri 18861 19333 18941 19413 ne
rect 18941 19333 19313 19413
tri 19313 19333 19393 19413 sw
tri 19411 19333 19491 19413 ne
rect 19491 19333 20100 19413
rect 261 19313 693 19333
rect -500 19235 163 19313
tri 163 19235 241 19313 sw
tri 261 19235 339 19313 ne
rect 339 19235 693 19313
tri 693 19235 791 19333 sw
tri 791 19235 889 19333 ne
rect 889 19235 1243 19333
tri 1243 19235 1341 19333 sw
tri 1341 19235 1439 19333 ne
rect 1439 19235 1793 19333
tri 1793 19235 1891 19333 sw
tri 1891 19235 1989 19333 ne
rect 1989 19235 2343 19333
tri 2343 19235 2441 19333 sw
tri 2441 19235 2539 19333 ne
rect 2539 19235 2893 19333
tri 2893 19235 2991 19333 sw
tri 2991 19235 3089 19333 ne
rect 3089 19235 3443 19333
tri 3443 19235 3541 19333 sw
tri 3541 19235 3639 19333 ne
rect 3639 19235 3993 19333
tri 3993 19235 4091 19333 sw
tri 4091 19235 4189 19333 ne
rect 4189 19235 4543 19333
tri 4543 19235 4641 19333 sw
tri 4641 19235 4739 19333 ne
rect 4739 19235 5093 19333
tri 5093 19235 5191 19333 sw
tri 5191 19235 5289 19333 ne
rect 5289 19235 5643 19333
tri 5643 19235 5741 19333 sw
tri 5741 19235 5839 19333 ne
rect 5839 19235 6193 19333
tri 6193 19235 6291 19333 sw
tri 6291 19235 6389 19333 ne
rect 6389 19235 6743 19333
tri 6743 19235 6841 19333 sw
tri 6841 19235 6939 19333 ne
rect 6939 19235 7293 19333
tri 7293 19235 7391 19333 sw
tri 7391 19235 7489 19333 ne
rect 7489 19235 7843 19333
tri 7843 19235 7941 19333 sw
tri 7941 19235 8039 19333 ne
rect 8039 19235 8393 19333
tri 8393 19235 8491 19333 sw
tri 8491 19235 8589 19333 ne
rect 8589 19235 8943 19333
tri 8943 19235 9041 19333 sw
tri 9041 19235 9139 19333 ne
rect 9139 19235 9493 19333
tri 9493 19235 9591 19333 sw
tri 9591 19235 9689 19333 ne
rect 9689 19235 10043 19333
tri 10043 19235 10141 19333 sw
tri 10141 19235 10239 19333 ne
rect 10239 19235 10593 19333
tri 10593 19235 10691 19333 sw
tri 10691 19235 10789 19333 ne
rect 10789 19235 11143 19333
tri 11143 19235 11241 19333 sw
tri 11241 19235 11339 19333 ne
rect 11339 19235 11693 19333
tri 11693 19235 11791 19333 sw
tri 11791 19235 11889 19333 ne
rect 11889 19235 12243 19333
tri 12243 19235 12341 19333 sw
tri 12341 19235 12439 19333 ne
rect 12439 19235 12793 19333
tri 12793 19235 12891 19333 sw
tri 12891 19235 12989 19333 ne
rect 12989 19235 13343 19333
tri 13343 19235 13441 19333 sw
tri 13441 19235 13539 19333 ne
rect 13539 19235 13893 19333
tri 13893 19235 13991 19333 sw
tri 13991 19235 14089 19333 ne
rect 14089 19235 14443 19333
tri 14443 19235 14541 19333 sw
tri 14541 19235 14639 19333 ne
rect 14639 19235 14993 19333
tri 14993 19235 15091 19333 sw
tri 15091 19235 15189 19333 ne
rect 15189 19235 15543 19333
tri 15543 19235 15641 19333 sw
tri 15641 19235 15739 19333 ne
rect 15739 19235 16093 19333
tri 16093 19235 16191 19333 sw
tri 16191 19235 16289 19333 ne
rect 16289 19235 16643 19333
tri 16643 19235 16741 19333 sw
tri 16741 19235 16839 19333 ne
rect 16839 19235 17193 19333
tri 17193 19235 17291 19333 sw
tri 17291 19235 17389 19333 ne
rect 17389 19235 17743 19333
tri 17743 19235 17841 19333 sw
tri 17841 19235 17939 19333 ne
rect 17939 19235 18293 19333
tri 18293 19235 18391 19333 sw
tri 18391 19235 18489 19333 ne
rect 18489 19235 18843 19333
tri 18843 19235 18941 19333 sw
tri 18941 19235 19039 19333 ne
rect 19039 19235 19393 19333
tri 19393 19235 19491 19333 sw
tri 19491 19235 19589 19333 ne
rect 19589 19313 20100 19333
rect 20200 19313 21800 19413
rect 19589 19235 21800 19313
rect -500 19187 241 19235
rect -500 19087 -400 19187
rect -300 19137 241 19187
tri 241 19137 339 19235 sw
tri 339 19137 437 19235 ne
rect 437 19137 791 19235
tri 791 19137 889 19235 sw
tri 889 19137 987 19235 ne
rect 987 19137 1341 19235
tri 1341 19137 1439 19235 sw
tri 1439 19137 1537 19235 ne
rect 1537 19137 1891 19235
tri 1891 19137 1989 19235 sw
tri 1989 19137 2087 19235 ne
rect 2087 19137 2441 19235
tri 2441 19137 2539 19235 sw
tri 2539 19137 2637 19235 ne
rect 2637 19137 2991 19235
tri 2991 19137 3089 19235 sw
tri 3089 19137 3187 19235 ne
rect 3187 19137 3541 19235
tri 3541 19137 3639 19235 sw
tri 3639 19137 3737 19235 ne
rect 3737 19137 4091 19235
tri 4091 19137 4189 19235 sw
tri 4189 19137 4287 19235 ne
rect 4287 19137 4641 19235
tri 4641 19137 4739 19235 sw
tri 4739 19137 4837 19235 ne
rect 4837 19137 5191 19235
tri 5191 19137 5289 19235 sw
tri 5289 19137 5387 19235 ne
rect 5387 19137 5741 19235
tri 5741 19137 5839 19235 sw
tri 5839 19137 5937 19235 ne
rect 5937 19137 6291 19235
tri 6291 19137 6389 19235 sw
tri 6389 19137 6487 19235 ne
rect 6487 19137 6841 19235
tri 6841 19137 6939 19235 sw
tri 6939 19137 7037 19235 ne
rect 7037 19137 7391 19235
tri 7391 19137 7489 19235 sw
tri 7489 19137 7587 19235 ne
rect 7587 19137 7941 19235
tri 7941 19137 8039 19235 sw
tri 8039 19137 8137 19235 ne
rect 8137 19137 8491 19235
tri 8491 19137 8589 19235 sw
tri 8589 19137 8687 19235 ne
rect 8687 19137 9041 19235
tri 9041 19137 9139 19235 sw
tri 9139 19137 9237 19235 ne
rect 9237 19137 9591 19235
tri 9591 19137 9689 19235 sw
tri 9689 19137 9787 19235 ne
rect 9787 19137 10141 19235
tri 10141 19137 10239 19235 sw
tri 10239 19137 10337 19235 ne
rect 10337 19137 10691 19235
tri 10691 19137 10789 19235 sw
tri 10789 19137 10887 19235 ne
rect 10887 19137 11241 19235
tri 11241 19137 11339 19235 sw
tri 11339 19137 11437 19235 ne
rect 11437 19137 11791 19235
tri 11791 19137 11889 19235 sw
tri 11889 19137 11987 19235 ne
rect 11987 19137 12341 19235
tri 12341 19137 12439 19235 sw
tri 12439 19137 12537 19235 ne
rect 12537 19137 12891 19235
tri 12891 19137 12989 19235 sw
tri 12989 19137 13087 19235 ne
rect 13087 19137 13441 19235
tri 13441 19137 13539 19235 sw
tri 13539 19137 13637 19235 ne
rect 13637 19137 13991 19235
tri 13991 19137 14089 19235 sw
tri 14089 19137 14187 19235 ne
rect 14187 19137 14541 19235
tri 14541 19137 14639 19235 sw
tri 14639 19137 14737 19235 ne
rect 14737 19137 15091 19235
tri 15091 19137 15189 19235 sw
tri 15189 19137 15287 19235 ne
rect 15287 19137 15641 19235
tri 15641 19137 15739 19235 sw
tri 15739 19137 15837 19235 ne
rect 15837 19137 16191 19235
tri 16191 19137 16289 19235 sw
tri 16289 19137 16387 19235 ne
rect 16387 19137 16741 19235
tri 16741 19137 16839 19235 sw
tri 16839 19137 16937 19235 ne
rect 16937 19137 17291 19235
tri 17291 19137 17389 19235 sw
tri 17389 19137 17487 19235 ne
rect 17487 19137 17841 19235
tri 17841 19137 17939 19235 sw
tri 17939 19137 18037 19235 ne
rect 18037 19137 18391 19235
tri 18391 19137 18489 19235 sw
tri 18489 19137 18587 19235 ne
rect 18587 19137 18941 19235
tri 18941 19137 19039 19235 sw
tri 19039 19137 19137 19235 ne
rect 19137 19137 19491 19235
tri 19491 19137 19589 19235 sw
tri 19589 19137 19687 19235 ne
rect 19687 19137 21800 19235
rect -300 19087 339 19137
rect -500 19039 339 19087
tri 339 19039 437 19137 sw
tri 437 19039 535 19137 ne
rect 535 19039 889 19137
tri 889 19039 987 19137 sw
tri 987 19039 1085 19137 ne
rect 1085 19039 1439 19137
tri 1439 19039 1537 19137 sw
tri 1537 19039 1635 19137 ne
rect 1635 19039 1989 19137
tri 1989 19039 2087 19137 sw
tri 2087 19039 2185 19137 ne
rect 2185 19039 2539 19137
tri 2539 19039 2637 19137 sw
tri 2637 19039 2735 19137 ne
rect 2735 19039 3089 19137
tri 3089 19039 3187 19137 sw
tri 3187 19039 3285 19137 ne
rect 3285 19039 3639 19137
tri 3639 19039 3737 19137 sw
tri 3737 19039 3835 19137 ne
rect 3835 19039 4189 19137
tri 4189 19039 4287 19137 sw
tri 4287 19039 4385 19137 ne
rect 4385 19039 4739 19137
tri 4739 19039 4837 19137 sw
tri 4837 19039 4935 19137 ne
rect 4935 19039 5289 19137
tri 5289 19039 5387 19137 sw
tri 5387 19039 5485 19137 ne
rect 5485 19039 5839 19137
tri 5839 19039 5937 19137 sw
tri 5937 19039 6035 19137 ne
rect 6035 19039 6389 19137
tri 6389 19039 6487 19137 sw
tri 6487 19039 6585 19137 ne
rect 6585 19039 6939 19137
tri 6939 19039 7037 19137 sw
tri 7037 19039 7135 19137 ne
rect 7135 19039 7489 19137
tri 7489 19039 7587 19137 sw
tri 7587 19039 7685 19137 ne
rect 7685 19039 8039 19137
tri 8039 19039 8137 19137 sw
tri 8137 19039 8235 19137 ne
rect 8235 19039 8589 19137
tri 8589 19039 8687 19137 sw
tri 8687 19039 8785 19137 ne
rect 8785 19039 9139 19137
tri 9139 19039 9237 19137 sw
tri 9237 19039 9335 19137 ne
rect 9335 19039 9689 19137
tri 9689 19039 9787 19137 sw
tri 9787 19039 9885 19137 ne
rect 9885 19039 10239 19137
tri 10239 19039 10337 19137 sw
tri 10337 19039 10435 19137 ne
rect 10435 19039 10789 19137
tri 10789 19039 10887 19137 sw
tri 10887 19039 10985 19137 ne
rect 10985 19039 11339 19137
tri 11339 19039 11437 19137 sw
tri 11437 19039 11535 19137 ne
rect 11535 19039 11889 19137
tri 11889 19039 11987 19137 sw
tri 11987 19039 12085 19137 ne
rect 12085 19039 12439 19137
tri 12439 19039 12537 19137 sw
tri 12537 19039 12635 19137 ne
rect 12635 19039 12989 19137
tri 12989 19039 13087 19137 sw
tri 13087 19039 13185 19137 ne
rect 13185 19039 13539 19137
tri 13539 19039 13637 19137 sw
tri 13637 19039 13735 19137 ne
rect 13735 19039 14089 19137
tri 14089 19039 14187 19137 sw
tri 14187 19039 14285 19137 ne
rect 14285 19039 14639 19137
tri 14639 19039 14737 19137 sw
tri 14737 19039 14835 19137 ne
rect 14835 19039 15189 19137
tri 15189 19039 15287 19137 sw
tri 15287 19039 15385 19137 ne
rect 15385 19039 15739 19137
tri 15739 19039 15837 19137 sw
tri 15837 19039 15935 19137 ne
rect 15935 19039 16289 19137
tri 16289 19039 16387 19137 sw
tri 16387 19039 16485 19137 ne
rect 16485 19039 16839 19137
tri 16839 19039 16937 19137 sw
tri 16937 19039 17035 19137 ne
rect 17035 19039 17389 19137
tri 17389 19039 17487 19137 sw
tri 17487 19039 17585 19137 ne
rect 17585 19039 17939 19137
tri 17939 19039 18037 19137 sw
tri 18037 19039 18135 19137 ne
rect 18135 19039 18489 19137
tri 18489 19039 18587 19137 sw
tri 18587 19039 18685 19137 ne
rect 18685 19039 19039 19137
tri 19039 19039 19137 19137 sw
tri 19137 19039 19235 19137 ne
rect 19235 19039 19589 19137
tri 19589 19039 19687 19137 sw
rect -500 19035 437 19039
rect -500 18915 215 19035
rect 335 18941 437 19035
tri 437 18941 535 19039 sw
tri 535 18941 633 19039 ne
rect 633 19035 987 19039
rect 633 18941 765 19035
rect 335 18915 535 18941
rect -500 18911 535 18915
tri 535 18911 565 18941 sw
tri 633 18911 663 18941 ne
rect 663 18915 765 18941
rect 885 18941 987 19035
tri 987 18941 1085 19039 sw
tri 1085 18941 1183 19039 ne
rect 1183 19035 1537 19039
rect 1183 18941 1315 19035
rect 885 18915 1085 18941
rect 663 18911 1085 18915
tri 1085 18911 1115 18941 sw
tri 1183 18911 1213 18941 ne
rect 1213 18915 1315 18941
rect 1435 18941 1537 19035
tri 1537 18941 1635 19039 sw
tri 1635 18941 1733 19039 ne
rect 1733 19035 2087 19039
rect 1733 18941 1865 19035
rect 1435 18915 1635 18941
rect 1213 18911 1635 18915
tri 1635 18911 1665 18941 sw
tri 1733 18911 1763 18941 ne
rect 1763 18915 1865 18941
rect 1985 18941 2087 19035
tri 2087 18941 2185 19039 sw
tri 2185 18941 2283 19039 ne
rect 2283 19035 2637 19039
rect 2283 18941 2415 19035
rect 1985 18915 2185 18941
rect 1763 18911 2185 18915
tri 2185 18911 2215 18941 sw
tri 2283 18911 2313 18941 ne
rect 2313 18915 2415 18941
rect 2535 18941 2637 19035
tri 2637 18941 2735 19039 sw
tri 2735 18941 2833 19039 ne
rect 2833 19035 3187 19039
rect 2833 18941 2965 19035
rect 2535 18915 2735 18941
rect 2313 18911 2735 18915
tri 2735 18911 2765 18941 sw
tri 2833 18911 2863 18941 ne
rect 2863 18915 2965 18941
rect 3085 18941 3187 19035
tri 3187 18941 3285 19039 sw
tri 3285 18941 3383 19039 ne
rect 3383 19035 3737 19039
rect 3383 18941 3515 19035
rect 3085 18915 3285 18941
rect 2863 18911 3285 18915
tri 3285 18911 3315 18941 sw
tri 3383 18911 3413 18941 ne
rect 3413 18915 3515 18941
rect 3635 18941 3737 19035
tri 3737 18941 3835 19039 sw
tri 3835 18941 3933 19039 ne
rect 3933 19035 4287 19039
rect 3933 18941 4065 19035
rect 3635 18915 3835 18941
rect 3413 18911 3835 18915
tri 3835 18911 3865 18941 sw
tri 3933 18911 3963 18941 ne
rect 3963 18915 4065 18941
rect 4185 18941 4287 19035
tri 4287 18941 4385 19039 sw
tri 4385 18941 4483 19039 ne
rect 4483 19035 4837 19039
rect 4483 18941 4615 19035
rect 4185 18915 4385 18941
rect 3963 18911 4385 18915
tri 4385 18911 4415 18941 sw
tri 4483 18911 4513 18941 ne
rect 4513 18915 4615 18941
rect 4735 18941 4837 19035
tri 4837 18941 4935 19039 sw
tri 4935 18941 5033 19039 ne
rect 5033 19035 5387 19039
rect 5033 18941 5165 19035
rect 4735 18915 4935 18941
rect 4513 18911 4935 18915
tri 4935 18911 4965 18941 sw
tri 5033 18911 5063 18941 ne
rect 5063 18915 5165 18941
rect 5285 18941 5387 19035
tri 5387 18941 5485 19039 sw
tri 5485 18941 5583 19039 ne
rect 5583 19035 5937 19039
rect 5583 18941 5715 19035
rect 5285 18915 5485 18941
rect 5063 18911 5485 18915
tri 5485 18911 5515 18941 sw
tri 5583 18911 5613 18941 ne
rect 5613 18915 5715 18941
rect 5835 18941 5937 19035
tri 5937 18941 6035 19039 sw
tri 6035 18941 6133 19039 ne
rect 6133 19035 6487 19039
rect 6133 18941 6265 19035
rect 5835 18915 6035 18941
rect 5613 18911 6035 18915
tri 6035 18911 6065 18941 sw
tri 6133 18911 6163 18941 ne
rect 6163 18915 6265 18941
rect 6385 18941 6487 19035
tri 6487 18941 6585 19039 sw
tri 6585 18941 6683 19039 ne
rect 6683 19035 7037 19039
rect 6683 18941 6815 19035
rect 6385 18915 6585 18941
rect 6163 18911 6585 18915
tri 6585 18911 6615 18941 sw
tri 6683 18911 6713 18941 ne
rect 6713 18915 6815 18941
rect 6935 18941 7037 19035
tri 7037 18941 7135 19039 sw
tri 7135 18941 7233 19039 ne
rect 7233 19035 7587 19039
rect 7233 18941 7365 19035
rect 6935 18915 7135 18941
rect 6713 18911 7135 18915
tri 7135 18911 7165 18941 sw
tri 7233 18911 7263 18941 ne
rect 7263 18915 7365 18941
rect 7485 18941 7587 19035
tri 7587 18941 7685 19039 sw
tri 7685 18941 7783 19039 ne
rect 7783 19035 8137 19039
rect 7783 18941 7915 19035
rect 7485 18915 7685 18941
rect 7263 18911 7685 18915
tri 7685 18911 7715 18941 sw
tri 7783 18911 7813 18941 ne
rect 7813 18915 7915 18941
rect 8035 18941 8137 19035
tri 8137 18941 8235 19039 sw
tri 8235 18941 8333 19039 ne
rect 8333 19035 8687 19039
rect 8333 18941 8465 19035
rect 8035 18915 8235 18941
rect 7813 18911 8235 18915
tri 8235 18911 8265 18941 sw
tri 8333 18911 8363 18941 ne
rect 8363 18915 8465 18941
rect 8585 18941 8687 19035
tri 8687 18941 8785 19039 sw
tri 8785 18941 8883 19039 ne
rect 8883 19035 9237 19039
rect 8883 18941 9015 19035
rect 8585 18915 8785 18941
rect 8363 18911 8785 18915
tri 8785 18911 8815 18941 sw
tri 8883 18911 8913 18941 ne
rect 8913 18915 9015 18941
rect 9135 18941 9237 19035
tri 9237 18941 9335 19039 sw
tri 9335 18941 9433 19039 ne
rect 9433 19035 9787 19039
rect 9433 18941 9565 19035
rect 9135 18915 9335 18941
rect 8913 18911 9335 18915
tri 9335 18911 9365 18941 sw
tri 9433 18911 9463 18941 ne
rect 9463 18915 9565 18941
rect 9685 18941 9787 19035
tri 9787 18941 9885 19039 sw
tri 9885 18941 9983 19039 ne
rect 9983 19035 10337 19039
rect 9983 18941 10115 19035
rect 9685 18915 9885 18941
rect 9463 18911 9885 18915
tri 9885 18911 9915 18941 sw
tri 9983 18911 10013 18941 ne
rect 10013 18915 10115 18941
rect 10235 18941 10337 19035
tri 10337 18941 10435 19039 sw
tri 10435 18941 10533 19039 ne
rect 10533 19035 10887 19039
rect 10533 18941 10665 19035
rect 10235 18915 10435 18941
rect 10013 18911 10435 18915
tri 10435 18911 10465 18941 sw
tri 10533 18911 10563 18941 ne
rect 10563 18915 10665 18941
rect 10785 18941 10887 19035
tri 10887 18941 10985 19039 sw
tri 10985 18941 11083 19039 ne
rect 11083 19035 11437 19039
rect 11083 18941 11215 19035
rect 10785 18915 10985 18941
rect 10563 18911 10985 18915
tri 10985 18911 11015 18941 sw
tri 11083 18911 11113 18941 ne
rect 11113 18915 11215 18941
rect 11335 18941 11437 19035
tri 11437 18941 11535 19039 sw
tri 11535 18941 11633 19039 ne
rect 11633 19035 11987 19039
rect 11633 18941 11765 19035
rect 11335 18915 11535 18941
rect 11113 18911 11535 18915
tri 11535 18911 11565 18941 sw
tri 11633 18911 11663 18941 ne
rect 11663 18915 11765 18941
rect 11885 18941 11987 19035
tri 11987 18941 12085 19039 sw
tri 12085 18941 12183 19039 ne
rect 12183 19035 12537 19039
rect 12183 18941 12315 19035
rect 11885 18915 12085 18941
rect 11663 18911 12085 18915
tri 12085 18911 12115 18941 sw
tri 12183 18911 12213 18941 ne
rect 12213 18915 12315 18941
rect 12435 18941 12537 19035
tri 12537 18941 12635 19039 sw
tri 12635 18941 12733 19039 ne
rect 12733 19035 13087 19039
rect 12733 18941 12865 19035
rect 12435 18915 12635 18941
rect 12213 18911 12635 18915
tri 12635 18911 12665 18941 sw
tri 12733 18911 12763 18941 ne
rect 12763 18915 12865 18941
rect 12985 18941 13087 19035
tri 13087 18941 13185 19039 sw
tri 13185 18941 13283 19039 ne
rect 13283 19035 13637 19039
rect 13283 18941 13415 19035
rect 12985 18915 13185 18941
rect 12763 18911 13185 18915
tri 13185 18911 13215 18941 sw
tri 13283 18911 13313 18941 ne
rect 13313 18915 13415 18941
rect 13535 18941 13637 19035
tri 13637 18941 13735 19039 sw
tri 13735 18941 13833 19039 ne
rect 13833 19035 14187 19039
rect 13833 18941 13965 19035
rect 13535 18915 13735 18941
rect 13313 18911 13735 18915
tri 13735 18911 13765 18941 sw
tri 13833 18911 13863 18941 ne
rect 13863 18915 13965 18941
rect 14085 18941 14187 19035
tri 14187 18941 14285 19039 sw
tri 14285 18941 14383 19039 ne
rect 14383 19035 14737 19039
rect 14383 18941 14515 19035
rect 14085 18915 14285 18941
rect 13863 18911 14285 18915
tri 14285 18911 14315 18941 sw
tri 14383 18911 14413 18941 ne
rect 14413 18915 14515 18941
rect 14635 18941 14737 19035
tri 14737 18941 14835 19039 sw
tri 14835 18941 14933 19039 ne
rect 14933 19035 15287 19039
rect 14933 18941 15065 19035
rect 14635 18915 14835 18941
rect 14413 18911 14835 18915
tri 14835 18911 14865 18941 sw
tri 14933 18911 14963 18941 ne
rect 14963 18915 15065 18941
rect 15185 18941 15287 19035
tri 15287 18941 15385 19039 sw
tri 15385 18941 15483 19039 ne
rect 15483 19035 15837 19039
rect 15483 18941 15615 19035
rect 15185 18915 15385 18941
rect 14963 18911 15385 18915
tri 15385 18911 15415 18941 sw
tri 15483 18911 15513 18941 ne
rect 15513 18915 15615 18941
rect 15735 18941 15837 19035
tri 15837 18941 15935 19039 sw
tri 15935 18941 16033 19039 ne
rect 16033 19035 16387 19039
rect 16033 18941 16165 19035
rect 15735 18915 15935 18941
rect 15513 18911 15935 18915
tri 15935 18911 15965 18941 sw
tri 16033 18911 16063 18941 ne
rect 16063 18915 16165 18941
rect 16285 18941 16387 19035
tri 16387 18941 16485 19039 sw
tri 16485 18941 16583 19039 ne
rect 16583 19035 16937 19039
rect 16583 18941 16715 19035
rect 16285 18915 16485 18941
rect 16063 18911 16485 18915
tri 16485 18911 16515 18941 sw
tri 16583 18911 16613 18941 ne
rect 16613 18915 16715 18941
rect 16835 18941 16937 19035
tri 16937 18941 17035 19039 sw
tri 17035 18941 17133 19039 ne
rect 17133 19035 17487 19039
rect 17133 18941 17265 19035
rect 16835 18915 17035 18941
rect 16613 18911 17035 18915
tri 17035 18911 17065 18941 sw
tri 17133 18911 17163 18941 ne
rect 17163 18915 17265 18941
rect 17385 18941 17487 19035
tri 17487 18941 17585 19039 sw
tri 17585 18941 17683 19039 ne
rect 17683 19035 18037 19039
rect 17683 18941 17815 19035
rect 17385 18915 17585 18941
rect 17163 18911 17585 18915
tri 17585 18911 17615 18941 sw
tri 17683 18911 17713 18941 ne
rect 17713 18915 17815 18941
rect 17935 18941 18037 19035
tri 18037 18941 18135 19039 sw
tri 18135 18941 18233 19039 ne
rect 18233 19035 18587 19039
rect 18233 18941 18365 19035
rect 17935 18915 18135 18941
rect 17713 18911 18135 18915
tri 18135 18911 18165 18941 sw
tri 18233 18911 18263 18941 ne
rect 18263 18915 18365 18941
rect 18485 18941 18587 19035
tri 18587 18941 18685 19039 sw
tri 18685 18941 18783 19039 ne
rect 18783 19035 19137 19039
rect 18783 18941 18915 19035
rect 18485 18915 18685 18941
rect 18263 18911 18685 18915
tri 18685 18911 18715 18941 sw
tri 18783 18911 18813 18941 ne
rect 18813 18915 18915 18941
rect 19035 18941 19137 19035
tri 19137 18941 19235 19039 sw
tri 19235 18941 19333 19039 ne
rect 19333 19035 20300 19039
rect 19333 18941 19465 19035
rect 19035 18915 19235 18941
rect 18813 18911 19235 18915
tri 19235 18911 19265 18941 sw
tri 19333 18911 19363 18941 ne
rect 19363 18915 19465 18941
rect 19585 18915 20300 19035
rect 19363 18911 20300 18915
tri 113 18813 211 18911 ne
rect 211 18813 565 18911
tri 565 18813 663 18911 sw
tri 663 18813 761 18911 ne
rect 761 18813 1115 18911
tri 1115 18813 1213 18911 sw
tri 1213 18813 1311 18911 ne
rect 1311 18813 1665 18911
tri 1665 18813 1763 18911 sw
tri 1763 18813 1861 18911 ne
rect 1861 18813 2215 18911
tri 2215 18813 2313 18911 sw
tri 2313 18813 2411 18911 ne
rect 2411 18813 2765 18911
tri 2765 18813 2863 18911 sw
tri 2863 18813 2961 18911 ne
rect 2961 18813 3315 18911
tri 3315 18813 3413 18911 sw
tri 3413 18813 3511 18911 ne
rect 3511 18813 3865 18911
tri 3865 18813 3963 18911 sw
tri 3963 18813 4061 18911 ne
rect 4061 18813 4415 18911
tri 4415 18813 4513 18911 sw
tri 4513 18813 4611 18911 ne
rect 4611 18813 4965 18911
tri 4965 18813 5063 18911 sw
tri 5063 18813 5161 18911 ne
rect 5161 18813 5515 18911
tri 5515 18813 5613 18911 sw
tri 5613 18813 5711 18911 ne
rect 5711 18813 6065 18911
tri 6065 18813 6163 18911 sw
tri 6163 18813 6261 18911 ne
rect 6261 18813 6615 18911
tri 6615 18813 6713 18911 sw
tri 6713 18813 6811 18911 ne
rect 6811 18813 7165 18911
tri 7165 18813 7263 18911 sw
tri 7263 18813 7361 18911 ne
rect 7361 18813 7715 18911
tri 7715 18813 7813 18911 sw
tri 7813 18813 7911 18911 ne
rect 7911 18813 8265 18911
tri 8265 18813 8363 18911 sw
tri 8363 18813 8461 18911 ne
rect 8461 18813 8815 18911
tri 8815 18813 8913 18911 sw
tri 8913 18813 9011 18911 ne
rect 9011 18813 9365 18911
tri 9365 18813 9463 18911 sw
tri 9463 18813 9561 18911 ne
rect 9561 18813 9915 18911
tri 9915 18813 10013 18911 sw
tri 10013 18813 10111 18911 ne
rect 10111 18813 10465 18911
tri 10465 18813 10563 18911 sw
tri 10563 18813 10661 18911 ne
rect 10661 18813 11015 18911
tri 11015 18813 11113 18911 sw
tri 11113 18813 11211 18911 ne
rect 11211 18813 11565 18911
tri 11565 18813 11663 18911 sw
tri 11663 18813 11761 18911 ne
rect 11761 18813 12115 18911
tri 12115 18813 12213 18911 sw
tri 12213 18813 12311 18911 ne
rect 12311 18813 12665 18911
tri 12665 18813 12763 18911 sw
tri 12763 18813 12861 18911 ne
rect 12861 18813 13215 18911
tri 13215 18813 13313 18911 sw
tri 13313 18813 13411 18911 ne
rect 13411 18813 13765 18911
tri 13765 18813 13863 18911 sw
tri 13863 18813 13961 18911 ne
rect 13961 18813 14315 18911
tri 14315 18813 14413 18911 sw
tri 14413 18813 14511 18911 ne
rect 14511 18813 14865 18911
tri 14865 18813 14963 18911 sw
tri 14963 18813 15061 18911 ne
rect 15061 18813 15415 18911
tri 15415 18813 15513 18911 sw
tri 15513 18813 15611 18911 ne
rect 15611 18813 15965 18911
tri 15965 18813 16063 18911 sw
tri 16063 18813 16161 18911 ne
rect 16161 18813 16515 18911
tri 16515 18813 16613 18911 sw
tri 16613 18813 16711 18911 ne
rect 16711 18813 17065 18911
tri 17065 18813 17163 18911 sw
tri 17163 18813 17261 18911 ne
rect 17261 18813 17615 18911
tri 17615 18813 17713 18911 sw
tri 17713 18813 17811 18911 ne
rect 17811 18813 18165 18911
tri 18165 18813 18263 18911 sw
tri 18263 18813 18361 18911 ne
rect 18361 18813 18715 18911
tri 18715 18813 18813 18911 sw
tri 18813 18813 18911 18911 ne
rect 18911 18813 19265 18911
tri 19265 18813 19363 18911 sw
tri 19363 18813 19461 18911 ne
rect 19461 18813 20300 18911
rect -2000 18783 113 18813
tri 113 18783 143 18813 sw
tri 211 18783 241 18813 ne
rect 241 18783 663 18813
tri 663 18783 693 18813 sw
tri 761 18783 791 18813 ne
rect 791 18783 1213 18813
tri 1213 18783 1243 18813 sw
tri 1311 18783 1341 18813 ne
rect 1341 18783 1763 18813
tri 1763 18783 1793 18813 sw
tri 1861 18783 1891 18813 ne
rect 1891 18783 2313 18813
tri 2313 18783 2343 18813 sw
tri 2411 18783 2441 18813 ne
rect 2441 18783 2863 18813
tri 2863 18783 2893 18813 sw
tri 2961 18783 2991 18813 ne
rect 2991 18783 3413 18813
tri 3413 18783 3443 18813 sw
tri 3511 18783 3541 18813 ne
rect 3541 18783 3963 18813
tri 3963 18783 3993 18813 sw
tri 4061 18783 4091 18813 ne
rect 4091 18783 4513 18813
tri 4513 18783 4543 18813 sw
tri 4611 18783 4641 18813 ne
rect 4641 18783 5063 18813
tri 5063 18783 5093 18813 sw
tri 5161 18783 5191 18813 ne
rect 5191 18783 5613 18813
tri 5613 18783 5643 18813 sw
tri 5711 18783 5741 18813 ne
rect 5741 18783 6163 18813
tri 6163 18783 6193 18813 sw
tri 6261 18783 6291 18813 ne
rect 6291 18783 6713 18813
tri 6713 18783 6743 18813 sw
tri 6811 18783 6841 18813 ne
rect 6841 18783 7263 18813
tri 7263 18783 7293 18813 sw
tri 7361 18783 7391 18813 ne
rect 7391 18783 7813 18813
tri 7813 18783 7843 18813 sw
tri 7911 18783 7941 18813 ne
rect 7941 18783 8363 18813
tri 8363 18783 8393 18813 sw
tri 8461 18783 8491 18813 ne
rect 8491 18783 8913 18813
tri 8913 18783 8943 18813 sw
tri 9011 18783 9041 18813 ne
rect 9041 18783 9463 18813
tri 9463 18783 9493 18813 sw
tri 9561 18783 9591 18813 ne
rect 9591 18783 10013 18813
tri 10013 18783 10043 18813 sw
tri 10111 18783 10141 18813 ne
rect 10141 18783 10563 18813
tri 10563 18783 10593 18813 sw
tri 10661 18783 10691 18813 ne
rect 10691 18783 11113 18813
tri 11113 18783 11143 18813 sw
tri 11211 18783 11241 18813 ne
rect 11241 18783 11663 18813
tri 11663 18783 11693 18813 sw
tri 11761 18783 11791 18813 ne
rect 11791 18783 12213 18813
tri 12213 18783 12243 18813 sw
tri 12311 18783 12341 18813 ne
rect 12341 18783 12763 18813
tri 12763 18783 12793 18813 sw
tri 12861 18783 12891 18813 ne
rect 12891 18783 13313 18813
tri 13313 18783 13343 18813 sw
tri 13411 18783 13441 18813 ne
rect 13441 18783 13863 18813
tri 13863 18783 13893 18813 sw
tri 13961 18783 13991 18813 ne
rect 13991 18783 14413 18813
tri 14413 18783 14443 18813 sw
tri 14511 18783 14541 18813 ne
rect 14541 18783 14963 18813
tri 14963 18783 14993 18813 sw
tri 15061 18783 15091 18813 ne
rect 15091 18783 15513 18813
tri 15513 18783 15543 18813 sw
tri 15611 18783 15641 18813 ne
rect 15641 18783 16063 18813
tri 16063 18783 16093 18813 sw
tri 16161 18783 16191 18813 ne
rect 16191 18783 16613 18813
tri 16613 18783 16643 18813 sw
tri 16711 18783 16741 18813 ne
rect 16741 18783 17163 18813
tri 17163 18783 17193 18813 sw
tri 17261 18783 17291 18813 ne
rect 17291 18783 17713 18813
tri 17713 18783 17743 18813 sw
tri 17811 18783 17841 18813 ne
rect 17841 18783 18263 18813
tri 18263 18783 18293 18813 sw
tri 18361 18783 18391 18813 ne
rect 18391 18783 18813 18813
tri 18813 18783 18843 18813 sw
tri 18911 18783 18941 18813 ne
rect 18941 18783 19363 18813
tri 19363 18783 19393 18813 sw
tri 19461 18783 19491 18813 ne
rect 19491 18783 20300 18813
rect -2000 18685 143 18783
tri 143 18685 241 18783 sw
tri 241 18685 339 18783 ne
rect 339 18685 693 18783
tri 693 18685 791 18783 sw
tri 791 18685 889 18783 ne
rect 889 18685 1243 18783
tri 1243 18685 1341 18783 sw
tri 1341 18685 1439 18783 ne
rect 1439 18685 1793 18783
tri 1793 18685 1891 18783 sw
tri 1891 18685 1989 18783 ne
rect 1989 18685 2343 18783
tri 2343 18685 2441 18783 sw
tri 2441 18685 2539 18783 ne
rect 2539 18685 2893 18783
tri 2893 18685 2991 18783 sw
tri 2991 18685 3089 18783 ne
rect 3089 18685 3443 18783
tri 3443 18685 3541 18783 sw
tri 3541 18685 3639 18783 ne
rect 3639 18685 3993 18783
tri 3993 18685 4091 18783 sw
tri 4091 18685 4189 18783 ne
rect 4189 18685 4543 18783
tri 4543 18685 4641 18783 sw
tri 4641 18685 4739 18783 ne
rect 4739 18685 5093 18783
tri 5093 18685 5191 18783 sw
tri 5191 18685 5289 18783 ne
rect 5289 18685 5643 18783
tri 5643 18685 5741 18783 sw
tri 5741 18685 5839 18783 ne
rect 5839 18685 6193 18783
tri 6193 18685 6291 18783 sw
tri 6291 18685 6389 18783 ne
rect 6389 18685 6743 18783
tri 6743 18685 6841 18783 sw
tri 6841 18685 6939 18783 ne
rect 6939 18685 7293 18783
tri 7293 18685 7391 18783 sw
tri 7391 18685 7489 18783 ne
rect 7489 18685 7843 18783
tri 7843 18685 7941 18783 sw
tri 7941 18685 8039 18783 ne
rect 8039 18685 8393 18783
tri 8393 18685 8491 18783 sw
tri 8491 18685 8589 18783 ne
rect 8589 18685 8943 18783
tri 8943 18685 9041 18783 sw
tri 9041 18685 9139 18783 ne
rect 9139 18685 9493 18783
tri 9493 18685 9591 18783 sw
tri 9591 18685 9689 18783 ne
rect 9689 18685 10043 18783
tri 10043 18685 10141 18783 sw
tri 10141 18685 10239 18783 ne
rect 10239 18685 10593 18783
tri 10593 18685 10691 18783 sw
tri 10691 18685 10789 18783 ne
rect 10789 18685 11143 18783
tri 11143 18685 11241 18783 sw
tri 11241 18685 11339 18783 ne
rect 11339 18685 11693 18783
tri 11693 18685 11791 18783 sw
tri 11791 18685 11889 18783 ne
rect 11889 18685 12243 18783
tri 12243 18685 12341 18783 sw
tri 12341 18685 12439 18783 ne
rect 12439 18685 12793 18783
tri 12793 18685 12891 18783 sw
tri 12891 18685 12989 18783 ne
rect 12989 18685 13343 18783
tri 13343 18685 13441 18783 sw
tri 13441 18685 13539 18783 ne
rect 13539 18685 13893 18783
tri 13893 18685 13991 18783 sw
tri 13991 18685 14089 18783 ne
rect 14089 18685 14443 18783
tri 14443 18685 14541 18783 sw
tri 14541 18685 14639 18783 ne
rect 14639 18685 14993 18783
tri 14993 18685 15091 18783 sw
tri 15091 18685 15189 18783 ne
rect 15189 18685 15543 18783
tri 15543 18685 15641 18783 sw
tri 15641 18685 15739 18783 ne
rect 15739 18685 16093 18783
tri 16093 18685 16191 18783 sw
tri 16191 18685 16289 18783 ne
rect 16289 18685 16643 18783
tri 16643 18685 16741 18783 sw
tri 16741 18685 16839 18783 ne
rect 16839 18685 17193 18783
tri 17193 18685 17291 18783 sw
tri 17291 18685 17389 18783 ne
rect 17389 18685 17743 18783
tri 17743 18685 17841 18783 sw
tri 17841 18685 17939 18783 ne
rect 17939 18685 18293 18783
tri 18293 18685 18391 18783 sw
tri 18391 18685 18489 18783 ne
rect 18489 18685 18843 18783
tri 18843 18685 18941 18783 sw
tri 18941 18685 19039 18783 ne
rect 19039 18685 19393 18783
tri 19393 18685 19491 18783 sw
tri 19491 18685 19589 18783 ne
rect 19589 18685 20300 18783
rect -2000 18587 241 18685
tri 241 18587 339 18685 sw
tri 339 18587 437 18685 ne
rect 437 18587 791 18685
tri 791 18587 889 18685 sw
tri 889 18587 987 18685 ne
rect 987 18587 1341 18685
tri 1341 18587 1439 18685 sw
tri 1439 18587 1537 18685 ne
rect 1537 18587 1891 18685
tri 1891 18587 1989 18685 sw
tri 1989 18587 2087 18685 ne
rect 2087 18587 2441 18685
tri 2441 18587 2539 18685 sw
tri 2539 18587 2637 18685 ne
rect 2637 18587 2991 18685
tri 2991 18587 3089 18685 sw
tri 3089 18587 3187 18685 ne
rect 3187 18587 3541 18685
tri 3541 18587 3639 18685 sw
tri 3639 18587 3737 18685 ne
rect 3737 18587 4091 18685
tri 4091 18587 4189 18685 sw
tri 4189 18587 4287 18685 ne
rect 4287 18587 4641 18685
tri 4641 18587 4739 18685 sw
tri 4739 18587 4837 18685 ne
rect 4837 18587 5191 18685
tri 5191 18587 5289 18685 sw
tri 5289 18587 5387 18685 ne
rect 5387 18587 5741 18685
tri 5741 18587 5839 18685 sw
tri 5839 18587 5937 18685 ne
rect 5937 18587 6291 18685
tri 6291 18587 6389 18685 sw
tri 6389 18587 6487 18685 ne
rect 6487 18587 6841 18685
tri 6841 18587 6939 18685 sw
tri 6939 18587 7037 18685 ne
rect 7037 18587 7391 18685
tri 7391 18587 7489 18685 sw
tri 7489 18587 7587 18685 ne
rect 7587 18587 7941 18685
tri 7941 18587 8039 18685 sw
tri 8039 18587 8137 18685 ne
rect 8137 18587 8491 18685
tri 8491 18587 8589 18685 sw
tri 8589 18587 8687 18685 ne
rect 8687 18587 9041 18685
tri 9041 18587 9139 18685 sw
tri 9139 18587 9237 18685 ne
rect 9237 18587 9591 18685
tri 9591 18587 9689 18685 sw
tri 9689 18587 9787 18685 ne
rect 9787 18587 10141 18685
tri 10141 18587 10239 18685 sw
tri 10239 18587 10337 18685 ne
rect 10337 18587 10691 18685
tri 10691 18587 10789 18685 sw
tri 10789 18587 10887 18685 ne
rect 10887 18587 11241 18685
tri 11241 18587 11339 18685 sw
tri 11339 18587 11437 18685 ne
rect 11437 18587 11791 18685
tri 11791 18587 11889 18685 sw
tri 11889 18587 11987 18685 ne
rect 11987 18587 12341 18685
tri 12341 18587 12439 18685 sw
tri 12439 18587 12537 18685 ne
rect 12537 18587 12891 18685
tri 12891 18587 12989 18685 sw
tri 12989 18587 13087 18685 ne
rect 13087 18587 13441 18685
tri 13441 18587 13539 18685 sw
tri 13539 18587 13637 18685 ne
rect 13637 18587 13991 18685
tri 13991 18587 14089 18685 sw
tri 14089 18587 14187 18685 ne
rect 14187 18587 14541 18685
tri 14541 18587 14639 18685 sw
tri 14639 18587 14737 18685 ne
rect 14737 18587 15091 18685
tri 15091 18587 15189 18685 sw
tri 15189 18587 15287 18685 ne
rect 15287 18587 15641 18685
tri 15641 18587 15739 18685 sw
tri 15739 18587 15837 18685 ne
rect 15837 18587 16191 18685
tri 16191 18587 16289 18685 sw
tri 16289 18587 16387 18685 ne
rect 16387 18587 16741 18685
tri 16741 18587 16839 18685 sw
tri 16839 18587 16937 18685 ne
rect 16937 18587 17291 18685
tri 17291 18587 17389 18685 sw
tri 17389 18587 17487 18685 ne
rect 17487 18587 17841 18685
tri 17841 18587 17939 18685 sw
tri 17939 18587 18037 18685 ne
rect 18037 18587 18391 18685
tri 18391 18587 18489 18685 sw
tri 18489 18587 18587 18685 ne
rect 18587 18587 18941 18685
tri 18941 18587 19039 18685 sw
tri 19039 18587 19137 18685 ne
rect 19137 18587 19491 18685
tri 19491 18587 19589 18685 sw
tri 19589 18587 19687 18685 ne
rect 19687 18587 20300 18685
rect -2000 18489 339 18587
tri 339 18489 437 18587 sw
tri 437 18489 535 18587 ne
rect 535 18489 889 18587
tri 889 18489 987 18587 sw
tri 987 18489 1085 18587 ne
rect 1085 18489 1439 18587
tri 1439 18489 1537 18587 sw
tri 1537 18489 1635 18587 ne
rect 1635 18489 1989 18587
tri 1989 18489 2087 18587 sw
tri 2087 18489 2185 18587 ne
rect 2185 18489 2539 18587
tri 2539 18489 2637 18587 sw
tri 2637 18489 2735 18587 ne
rect 2735 18489 3089 18587
tri 3089 18489 3187 18587 sw
tri 3187 18489 3285 18587 ne
rect 3285 18489 3639 18587
tri 3639 18489 3737 18587 sw
tri 3737 18489 3835 18587 ne
rect 3835 18489 4189 18587
tri 4189 18489 4287 18587 sw
tri 4287 18489 4385 18587 ne
rect 4385 18489 4739 18587
tri 4739 18489 4837 18587 sw
tri 4837 18489 4935 18587 ne
rect 4935 18489 5289 18587
tri 5289 18489 5387 18587 sw
tri 5387 18489 5485 18587 ne
rect 5485 18489 5839 18587
tri 5839 18489 5937 18587 sw
tri 5937 18489 6035 18587 ne
rect 6035 18489 6389 18587
tri 6389 18489 6487 18587 sw
tri 6487 18489 6585 18587 ne
rect 6585 18489 6939 18587
tri 6939 18489 7037 18587 sw
tri 7037 18489 7135 18587 ne
rect 7135 18489 7489 18587
tri 7489 18489 7587 18587 sw
tri 7587 18489 7685 18587 ne
rect 7685 18489 8039 18587
tri 8039 18489 8137 18587 sw
tri 8137 18489 8235 18587 ne
rect 8235 18489 8589 18587
tri 8589 18489 8687 18587 sw
tri 8687 18489 8785 18587 ne
rect 8785 18489 9139 18587
tri 9139 18489 9237 18587 sw
tri 9237 18489 9335 18587 ne
rect 9335 18489 9689 18587
tri 9689 18489 9787 18587 sw
tri 9787 18489 9885 18587 ne
rect 9885 18489 10239 18587
tri 10239 18489 10337 18587 sw
tri 10337 18489 10435 18587 ne
rect 10435 18489 10789 18587
tri 10789 18489 10887 18587 sw
tri 10887 18489 10985 18587 ne
rect 10985 18489 11339 18587
tri 11339 18489 11437 18587 sw
tri 11437 18489 11535 18587 ne
rect 11535 18489 11889 18587
tri 11889 18489 11987 18587 sw
tri 11987 18489 12085 18587 ne
rect 12085 18489 12439 18587
tri 12439 18489 12537 18587 sw
tri 12537 18489 12635 18587 ne
rect 12635 18489 12989 18587
tri 12989 18489 13087 18587 sw
tri 13087 18489 13185 18587 ne
rect 13185 18489 13539 18587
tri 13539 18489 13637 18587 sw
tri 13637 18489 13735 18587 ne
rect 13735 18489 14089 18587
tri 14089 18489 14187 18587 sw
tri 14187 18489 14285 18587 ne
rect 14285 18489 14639 18587
tri 14639 18489 14737 18587 sw
tri 14737 18489 14835 18587 ne
rect 14835 18489 15189 18587
tri 15189 18489 15287 18587 sw
tri 15287 18489 15385 18587 ne
rect 15385 18489 15739 18587
tri 15739 18489 15837 18587 sw
tri 15837 18489 15935 18587 ne
rect 15935 18489 16289 18587
tri 16289 18489 16387 18587 sw
tri 16387 18489 16485 18587 ne
rect 16485 18489 16839 18587
tri 16839 18489 16937 18587 sw
tri 16937 18489 17035 18587 ne
rect 17035 18489 17389 18587
tri 17389 18489 17487 18587 sw
tri 17487 18489 17585 18587 ne
rect 17585 18489 17939 18587
tri 17939 18489 18037 18587 sw
tri 18037 18489 18135 18587 ne
rect 18135 18489 18489 18587
tri 18489 18489 18587 18587 sw
tri 18587 18489 18685 18587 ne
rect 18685 18489 19039 18587
tri 19039 18489 19137 18587 sw
tri 19137 18489 19235 18587 ne
rect 19235 18489 19589 18587
tri 19589 18489 19687 18587 sw
rect 20800 18489 21800 19137
rect -2000 18485 437 18489
rect -2000 18365 215 18485
rect 335 18391 437 18485
tri 437 18391 535 18489 sw
tri 535 18391 633 18489 ne
rect 633 18485 987 18489
rect 633 18391 765 18485
rect 335 18365 535 18391
rect -2000 18361 535 18365
rect -2000 17713 -1000 18361
tri 113 18263 211 18361 ne
rect 211 18313 535 18361
tri 535 18313 613 18391 sw
tri 633 18313 711 18391 ne
rect 711 18365 765 18391
rect 885 18391 987 18485
tri 987 18391 1085 18489 sw
tri 1085 18391 1183 18489 ne
rect 1183 18485 1537 18489
rect 1183 18391 1315 18485
rect 885 18365 1085 18391
rect 711 18313 1085 18365
tri 1085 18313 1163 18391 sw
tri 1183 18313 1261 18391 ne
rect 1261 18365 1315 18391
rect 1435 18391 1537 18485
tri 1537 18391 1635 18489 sw
tri 1635 18391 1733 18489 ne
rect 1733 18485 2087 18489
rect 1733 18391 1865 18485
rect 1435 18365 1635 18391
rect 1261 18313 1635 18365
tri 1635 18313 1713 18391 sw
tri 1733 18313 1811 18391 ne
rect 1811 18365 1865 18391
rect 1985 18391 2087 18485
tri 2087 18391 2185 18489 sw
tri 2185 18391 2283 18489 ne
rect 2283 18485 2637 18489
rect 2283 18391 2415 18485
rect 1985 18365 2185 18391
rect 1811 18313 2185 18365
tri 2185 18313 2263 18391 sw
tri 2283 18313 2361 18391 ne
rect 2361 18365 2415 18391
rect 2535 18391 2637 18485
tri 2637 18391 2735 18489 sw
tri 2735 18391 2833 18489 ne
rect 2833 18485 3187 18489
rect 2833 18391 2965 18485
rect 2535 18365 2735 18391
rect 2361 18313 2735 18365
tri 2735 18313 2813 18391 sw
tri 2833 18313 2911 18391 ne
rect 2911 18365 2965 18391
rect 3085 18391 3187 18485
tri 3187 18391 3285 18489 sw
tri 3285 18391 3383 18489 ne
rect 3383 18485 3737 18489
rect 3383 18391 3515 18485
rect 3085 18365 3285 18391
rect 2911 18313 3285 18365
tri 3285 18313 3363 18391 sw
tri 3383 18313 3461 18391 ne
rect 3461 18365 3515 18391
rect 3635 18391 3737 18485
tri 3737 18391 3835 18489 sw
tri 3835 18391 3933 18489 ne
rect 3933 18485 4287 18489
rect 3933 18391 4065 18485
rect 3635 18365 3835 18391
rect 3461 18313 3835 18365
tri 3835 18313 3913 18391 sw
tri 3933 18313 4011 18391 ne
rect 4011 18365 4065 18391
rect 4185 18391 4287 18485
tri 4287 18391 4385 18489 sw
tri 4385 18391 4483 18489 ne
rect 4483 18485 4837 18489
rect 4483 18391 4615 18485
rect 4185 18365 4385 18391
rect 4011 18313 4385 18365
tri 4385 18313 4463 18391 sw
tri 4483 18313 4561 18391 ne
rect 4561 18365 4615 18391
rect 4735 18391 4837 18485
tri 4837 18391 4935 18489 sw
tri 4935 18391 5033 18489 ne
rect 5033 18485 5387 18489
rect 5033 18391 5165 18485
rect 4735 18365 4935 18391
rect 4561 18313 4935 18365
tri 4935 18313 5013 18391 sw
tri 5033 18313 5111 18391 ne
rect 5111 18365 5165 18391
rect 5285 18391 5387 18485
tri 5387 18391 5485 18489 sw
tri 5485 18391 5583 18489 ne
rect 5583 18485 5937 18489
rect 5583 18391 5715 18485
rect 5285 18365 5485 18391
rect 5111 18313 5485 18365
tri 5485 18313 5563 18391 sw
tri 5583 18313 5661 18391 ne
rect 5661 18365 5715 18391
rect 5835 18391 5937 18485
tri 5937 18391 6035 18489 sw
tri 6035 18391 6133 18489 ne
rect 6133 18485 6487 18489
rect 6133 18391 6265 18485
rect 5835 18365 6035 18391
rect 5661 18313 6035 18365
tri 6035 18313 6113 18391 sw
tri 6133 18313 6211 18391 ne
rect 6211 18365 6265 18391
rect 6385 18391 6487 18485
tri 6487 18391 6585 18489 sw
tri 6585 18391 6683 18489 ne
rect 6683 18485 7037 18489
rect 6683 18391 6815 18485
rect 6385 18365 6585 18391
rect 6211 18313 6585 18365
tri 6585 18313 6663 18391 sw
tri 6683 18313 6761 18391 ne
rect 6761 18365 6815 18391
rect 6935 18391 7037 18485
tri 7037 18391 7135 18489 sw
tri 7135 18391 7233 18489 ne
rect 7233 18485 7587 18489
rect 7233 18391 7365 18485
rect 6935 18365 7135 18391
rect 6761 18313 7135 18365
tri 7135 18313 7213 18391 sw
tri 7233 18313 7311 18391 ne
rect 7311 18365 7365 18391
rect 7485 18391 7587 18485
tri 7587 18391 7685 18489 sw
tri 7685 18391 7783 18489 ne
rect 7783 18485 8137 18489
rect 7783 18391 7915 18485
rect 7485 18365 7685 18391
rect 7311 18313 7685 18365
tri 7685 18313 7763 18391 sw
tri 7783 18313 7861 18391 ne
rect 7861 18365 7915 18391
rect 8035 18391 8137 18485
tri 8137 18391 8235 18489 sw
tri 8235 18391 8333 18489 ne
rect 8333 18485 8687 18489
rect 8333 18391 8465 18485
rect 8035 18365 8235 18391
rect 7861 18313 8235 18365
tri 8235 18313 8313 18391 sw
tri 8333 18313 8411 18391 ne
rect 8411 18365 8465 18391
rect 8585 18391 8687 18485
tri 8687 18391 8785 18489 sw
tri 8785 18391 8883 18489 ne
rect 8883 18485 9237 18489
rect 8883 18391 9015 18485
rect 8585 18365 8785 18391
rect 8411 18313 8785 18365
tri 8785 18313 8863 18391 sw
tri 8883 18313 8961 18391 ne
rect 8961 18365 9015 18391
rect 9135 18391 9237 18485
tri 9237 18391 9335 18489 sw
tri 9335 18391 9433 18489 ne
rect 9433 18485 9787 18489
rect 9433 18391 9565 18485
rect 9135 18365 9335 18391
rect 8961 18313 9335 18365
tri 9335 18313 9413 18391 sw
tri 9433 18313 9511 18391 ne
rect 9511 18365 9565 18391
rect 9685 18391 9787 18485
tri 9787 18391 9885 18489 sw
tri 9885 18391 9983 18489 ne
rect 9983 18485 10337 18489
rect 9983 18391 10115 18485
rect 9685 18365 9885 18391
rect 9511 18313 9885 18365
tri 9885 18313 9963 18391 sw
tri 9983 18313 10061 18391 ne
rect 10061 18365 10115 18391
rect 10235 18391 10337 18485
tri 10337 18391 10435 18489 sw
tri 10435 18391 10533 18489 ne
rect 10533 18485 10887 18489
rect 10533 18391 10665 18485
rect 10235 18365 10435 18391
rect 10061 18313 10435 18365
tri 10435 18313 10513 18391 sw
tri 10533 18313 10611 18391 ne
rect 10611 18365 10665 18391
rect 10785 18391 10887 18485
tri 10887 18391 10985 18489 sw
tri 10985 18391 11083 18489 ne
rect 11083 18485 11437 18489
rect 11083 18391 11215 18485
rect 10785 18365 10985 18391
rect 10611 18313 10985 18365
tri 10985 18313 11063 18391 sw
tri 11083 18313 11161 18391 ne
rect 11161 18365 11215 18391
rect 11335 18391 11437 18485
tri 11437 18391 11535 18489 sw
tri 11535 18391 11633 18489 ne
rect 11633 18485 11987 18489
rect 11633 18391 11765 18485
rect 11335 18365 11535 18391
rect 11161 18313 11535 18365
tri 11535 18313 11613 18391 sw
tri 11633 18313 11711 18391 ne
rect 11711 18365 11765 18391
rect 11885 18391 11987 18485
tri 11987 18391 12085 18489 sw
tri 12085 18391 12183 18489 ne
rect 12183 18485 12537 18489
rect 12183 18391 12315 18485
rect 11885 18365 12085 18391
rect 11711 18313 12085 18365
tri 12085 18313 12163 18391 sw
tri 12183 18313 12261 18391 ne
rect 12261 18365 12315 18391
rect 12435 18391 12537 18485
tri 12537 18391 12635 18489 sw
tri 12635 18391 12733 18489 ne
rect 12733 18485 13087 18489
rect 12733 18391 12865 18485
rect 12435 18365 12635 18391
rect 12261 18313 12635 18365
tri 12635 18313 12713 18391 sw
tri 12733 18313 12811 18391 ne
rect 12811 18365 12865 18391
rect 12985 18391 13087 18485
tri 13087 18391 13185 18489 sw
tri 13185 18391 13283 18489 ne
rect 13283 18485 13637 18489
rect 13283 18391 13415 18485
rect 12985 18365 13185 18391
rect 12811 18313 13185 18365
tri 13185 18313 13263 18391 sw
tri 13283 18313 13361 18391 ne
rect 13361 18365 13415 18391
rect 13535 18391 13637 18485
tri 13637 18391 13735 18489 sw
tri 13735 18391 13833 18489 ne
rect 13833 18485 14187 18489
rect 13833 18391 13965 18485
rect 13535 18365 13735 18391
rect 13361 18313 13735 18365
tri 13735 18313 13813 18391 sw
tri 13833 18313 13911 18391 ne
rect 13911 18365 13965 18391
rect 14085 18391 14187 18485
tri 14187 18391 14285 18489 sw
tri 14285 18391 14383 18489 ne
rect 14383 18485 14737 18489
rect 14383 18391 14515 18485
rect 14085 18365 14285 18391
rect 13911 18313 14285 18365
tri 14285 18313 14363 18391 sw
tri 14383 18313 14461 18391 ne
rect 14461 18365 14515 18391
rect 14635 18391 14737 18485
tri 14737 18391 14835 18489 sw
tri 14835 18391 14933 18489 ne
rect 14933 18485 15287 18489
rect 14933 18391 15065 18485
rect 14635 18365 14835 18391
rect 14461 18313 14835 18365
tri 14835 18313 14913 18391 sw
tri 14933 18313 15011 18391 ne
rect 15011 18365 15065 18391
rect 15185 18391 15287 18485
tri 15287 18391 15385 18489 sw
tri 15385 18391 15483 18489 ne
rect 15483 18485 15837 18489
rect 15483 18391 15615 18485
rect 15185 18365 15385 18391
rect 15011 18313 15385 18365
tri 15385 18313 15463 18391 sw
tri 15483 18313 15561 18391 ne
rect 15561 18365 15615 18391
rect 15735 18391 15837 18485
tri 15837 18391 15935 18489 sw
tri 15935 18391 16033 18489 ne
rect 16033 18485 16387 18489
rect 16033 18391 16165 18485
rect 15735 18365 15935 18391
rect 15561 18313 15935 18365
tri 15935 18313 16013 18391 sw
tri 16033 18313 16111 18391 ne
rect 16111 18365 16165 18391
rect 16285 18391 16387 18485
tri 16387 18391 16485 18489 sw
tri 16485 18391 16583 18489 ne
rect 16583 18485 16937 18489
rect 16583 18391 16715 18485
rect 16285 18365 16485 18391
rect 16111 18313 16485 18365
tri 16485 18313 16563 18391 sw
tri 16583 18313 16661 18391 ne
rect 16661 18365 16715 18391
rect 16835 18391 16937 18485
tri 16937 18391 17035 18489 sw
tri 17035 18391 17133 18489 ne
rect 17133 18485 17487 18489
rect 17133 18391 17265 18485
rect 16835 18365 17035 18391
rect 16661 18313 17035 18365
tri 17035 18313 17113 18391 sw
tri 17133 18313 17211 18391 ne
rect 17211 18365 17265 18391
rect 17385 18391 17487 18485
tri 17487 18391 17585 18489 sw
tri 17585 18391 17683 18489 ne
rect 17683 18485 18037 18489
rect 17683 18391 17815 18485
rect 17385 18365 17585 18391
rect 17211 18313 17585 18365
tri 17585 18313 17663 18391 sw
tri 17683 18313 17761 18391 ne
rect 17761 18365 17815 18391
rect 17935 18391 18037 18485
tri 18037 18391 18135 18489 sw
tri 18135 18391 18233 18489 ne
rect 18233 18485 18587 18489
rect 18233 18391 18365 18485
rect 17935 18365 18135 18391
rect 17761 18313 18135 18365
tri 18135 18313 18213 18391 sw
tri 18233 18313 18311 18391 ne
rect 18311 18365 18365 18391
rect 18485 18391 18587 18485
tri 18587 18391 18685 18489 sw
tri 18685 18391 18783 18489 ne
rect 18783 18485 19137 18489
rect 18783 18391 18915 18485
rect 18485 18365 18685 18391
rect 18311 18313 18685 18365
tri 18685 18313 18763 18391 sw
tri 18783 18313 18861 18391 ne
rect 18861 18365 18915 18391
rect 19035 18391 19137 18485
tri 19137 18391 19235 18489 sw
tri 19235 18391 19333 18489 ne
rect 19333 18485 21800 18489
rect 19333 18391 19465 18485
rect 19035 18365 19235 18391
rect 18861 18313 19235 18365
tri 19235 18313 19313 18391 sw
tri 19333 18313 19411 18391 ne
rect 19411 18365 19465 18391
rect 19585 18365 21800 18485
rect 19411 18313 21800 18365
rect 211 18263 613 18313
rect -500 18213 113 18263
tri 113 18213 163 18263 sw
tri 211 18213 261 18263 ne
rect 261 18233 613 18263
tri 613 18233 693 18313 sw
tri 711 18233 791 18313 ne
rect 791 18233 1163 18313
tri 1163 18233 1243 18313 sw
tri 1261 18233 1341 18313 ne
rect 1341 18233 1713 18313
tri 1713 18233 1793 18313 sw
tri 1811 18233 1891 18313 ne
rect 1891 18233 2263 18313
tri 2263 18233 2343 18313 sw
tri 2361 18233 2441 18313 ne
rect 2441 18233 2813 18313
tri 2813 18233 2893 18313 sw
tri 2911 18233 2991 18313 ne
rect 2991 18233 3363 18313
tri 3363 18233 3443 18313 sw
tri 3461 18233 3541 18313 ne
rect 3541 18233 3913 18313
tri 3913 18233 3993 18313 sw
tri 4011 18233 4091 18313 ne
rect 4091 18233 4463 18313
tri 4463 18233 4543 18313 sw
tri 4561 18233 4641 18313 ne
rect 4641 18233 5013 18313
tri 5013 18233 5093 18313 sw
tri 5111 18233 5191 18313 ne
rect 5191 18233 5563 18313
tri 5563 18233 5643 18313 sw
tri 5661 18233 5741 18313 ne
rect 5741 18233 6113 18313
tri 6113 18233 6193 18313 sw
tri 6211 18233 6291 18313 ne
rect 6291 18233 6663 18313
tri 6663 18233 6743 18313 sw
tri 6761 18233 6841 18313 ne
rect 6841 18233 7213 18313
tri 7213 18233 7293 18313 sw
tri 7311 18233 7391 18313 ne
rect 7391 18233 7763 18313
tri 7763 18233 7843 18313 sw
tri 7861 18233 7941 18313 ne
rect 7941 18233 8313 18313
tri 8313 18233 8393 18313 sw
tri 8411 18233 8491 18313 ne
rect 8491 18233 8863 18313
tri 8863 18233 8943 18313 sw
tri 8961 18233 9041 18313 ne
rect 9041 18233 9413 18313
tri 9413 18233 9493 18313 sw
tri 9511 18233 9591 18313 ne
rect 9591 18233 9963 18313
tri 9963 18233 10043 18313 sw
tri 10061 18233 10141 18313 ne
rect 10141 18233 10513 18313
tri 10513 18233 10593 18313 sw
tri 10611 18233 10691 18313 ne
rect 10691 18233 11063 18313
tri 11063 18233 11143 18313 sw
tri 11161 18233 11241 18313 ne
rect 11241 18233 11613 18313
tri 11613 18233 11693 18313 sw
tri 11711 18233 11791 18313 ne
rect 11791 18233 12163 18313
tri 12163 18233 12243 18313 sw
tri 12261 18233 12341 18313 ne
rect 12341 18233 12713 18313
tri 12713 18233 12793 18313 sw
tri 12811 18233 12891 18313 ne
rect 12891 18233 13263 18313
tri 13263 18233 13343 18313 sw
tri 13361 18233 13441 18313 ne
rect 13441 18233 13813 18313
tri 13813 18233 13893 18313 sw
tri 13911 18233 13991 18313 ne
rect 13991 18233 14363 18313
tri 14363 18233 14443 18313 sw
tri 14461 18233 14541 18313 ne
rect 14541 18233 14913 18313
tri 14913 18233 14993 18313 sw
tri 15011 18233 15091 18313 ne
rect 15091 18233 15463 18313
tri 15463 18233 15543 18313 sw
tri 15561 18233 15641 18313 ne
rect 15641 18233 16013 18313
tri 16013 18233 16093 18313 sw
tri 16111 18233 16191 18313 ne
rect 16191 18233 16563 18313
tri 16563 18233 16643 18313 sw
tri 16661 18233 16741 18313 ne
rect 16741 18233 17113 18313
tri 17113 18233 17193 18313 sw
tri 17211 18233 17291 18313 ne
rect 17291 18233 17663 18313
tri 17663 18233 17743 18313 sw
tri 17761 18233 17841 18313 ne
rect 17841 18233 18213 18313
tri 18213 18233 18293 18313 sw
tri 18311 18233 18391 18313 ne
rect 18391 18233 18763 18313
tri 18763 18233 18843 18313 sw
tri 18861 18233 18941 18313 ne
rect 18941 18233 19313 18313
tri 19313 18233 19393 18313 sw
tri 19411 18233 19491 18313 ne
rect 19491 18233 20100 18313
rect 261 18213 693 18233
rect -500 18135 163 18213
tri 163 18135 241 18213 sw
tri 261 18135 339 18213 ne
rect 339 18135 693 18213
tri 693 18135 791 18233 sw
tri 791 18135 889 18233 ne
rect 889 18135 1243 18233
tri 1243 18135 1341 18233 sw
tri 1341 18135 1439 18233 ne
rect 1439 18135 1793 18233
tri 1793 18135 1891 18233 sw
tri 1891 18135 1989 18233 ne
rect 1989 18135 2343 18233
tri 2343 18135 2441 18233 sw
tri 2441 18135 2539 18233 ne
rect 2539 18135 2893 18233
tri 2893 18135 2991 18233 sw
tri 2991 18135 3089 18233 ne
rect 3089 18135 3443 18233
tri 3443 18135 3541 18233 sw
tri 3541 18135 3639 18233 ne
rect 3639 18135 3993 18233
tri 3993 18135 4091 18233 sw
tri 4091 18135 4189 18233 ne
rect 4189 18135 4543 18233
tri 4543 18135 4641 18233 sw
tri 4641 18135 4739 18233 ne
rect 4739 18135 5093 18233
tri 5093 18135 5191 18233 sw
tri 5191 18135 5289 18233 ne
rect 5289 18135 5643 18233
tri 5643 18135 5741 18233 sw
tri 5741 18135 5839 18233 ne
rect 5839 18135 6193 18233
tri 6193 18135 6291 18233 sw
tri 6291 18135 6389 18233 ne
rect 6389 18135 6743 18233
tri 6743 18135 6841 18233 sw
tri 6841 18135 6939 18233 ne
rect 6939 18135 7293 18233
tri 7293 18135 7391 18233 sw
tri 7391 18135 7489 18233 ne
rect 7489 18135 7843 18233
tri 7843 18135 7941 18233 sw
tri 7941 18135 8039 18233 ne
rect 8039 18135 8393 18233
tri 8393 18135 8491 18233 sw
tri 8491 18135 8589 18233 ne
rect 8589 18135 8943 18233
tri 8943 18135 9041 18233 sw
tri 9041 18135 9139 18233 ne
rect 9139 18135 9493 18233
tri 9493 18135 9591 18233 sw
tri 9591 18135 9689 18233 ne
rect 9689 18135 10043 18233
tri 10043 18135 10141 18233 sw
tri 10141 18135 10239 18233 ne
rect 10239 18135 10593 18233
tri 10593 18135 10691 18233 sw
tri 10691 18135 10789 18233 ne
rect 10789 18135 11143 18233
tri 11143 18135 11241 18233 sw
tri 11241 18135 11339 18233 ne
rect 11339 18135 11693 18233
tri 11693 18135 11791 18233 sw
tri 11791 18135 11889 18233 ne
rect 11889 18135 12243 18233
tri 12243 18135 12341 18233 sw
tri 12341 18135 12439 18233 ne
rect 12439 18135 12793 18233
tri 12793 18135 12891 18233 sw
tri 12891 18135 12989 18233 ne
rect 12989 18135 13343 18233
tri 13343 18135 13441 18233 sw
tri 13441 18135 13539 18233 ne
rect 13539 18135 13893 18233
tri 13893 18135 13991 18233 sw
tri 13991 18135 14089 18233 ne
rect 14089 18135 14443 18233
tri 14443 18135 14541 18233 sw
tri 14541 18135 14639 18233 ne
rect 14639 18135 14993 18233
tri 14993 18135 15091 18233 sw
tri 15091 18135 15189 18233 ne
rect 15189 18135 15543 18233
tri 15543 18135 15641 18233 sw
tri 15641 18135 15739 18233 ne
rect 15739 18135 16093 18233
tri 16093 18135 16191 18233 sw
tri 16191 18135 16289 18233 ne
rect 16289 18135 16643 18233
tri 16643 18135 16741 18233 sw
tri 16741 18135 16839 18233 ne
rect 16839 18135 17193 18233
tri 17193 18135 17291 18233 sw
tri 17291 18135 17389 18233 ne
rect 17389 18135 17743 18233
tri 17743 18135 17841 18233 sw
tri 17841 18135 17939 18233 ne
rect 17939 18135 18293 18233
tri 18293 18135 18391 18233 sw
tri 18391 18135 18489 18233 ne
rect 18489 18135 18843 18233
tri 18843 18135 18941 18233 sw
tri 18941 18135 19039 18233 ne
rect 19039 18135 19393 18233
tri 19393 18135 19491 18233 sw
tri 19491 18135 19589 18233 ne
rect 19589 18213 20100 18233
rect 20200 18213 21800 18313
rect 19589 18135 21800 18213
rect -500 18087 241 18135
rect -500 17987 -400 18087
rect -300 18037 241 18087
tri 241 18037 339 18135 sw
tri 339 18037 437 18135 ne
rect 437 18037 791 18135
tri 791 18037 889 18135 sw
tri 889 18037 987 18135 ne
rect 987 18037 1341 18135
tri 1341 18037 1439 18135 sw
tri 1439 18037 1537 18135 ne
rect 1537 18037 1891 18135
tri 1891 18037 1989 18135 sw
tri 1989 18037 2087 18135 ne
rect 2087 18037 2441 18135
tri 2441 18037 2539 18135 sw
tri 2539 18037 2637 18135 ne
rect 2637 18037 2991 18135
tri 2991 18037 3089 18135 sw
tri 3089 18037 3187 18135 ne
rect 3187 18037 3541 18135
tri 3541 18037 3639 18135 sw
tri 3639 18037 3737 18135 ne
rect 3737 18037 4091 18135
tri 4091 18037 4189 18135 sw
tri 4189 18037 4287 18135 ne
rect 4287 18037 4641 18135
tri 4641 18037 4739 18135 sw
tri 4739 18037 4837 18135 ne
rect 4837 18037 5191 18135
tri 5191 18037 5289 18135 sw
tri 5289 18037 5387 18135 ne
rect 5387 18037 5741 18135
tri 5741 18037 5839 18135 sw
tri 5839 18037 5937 18135 ne
rect 5937 18037 6291 18135
tri 6291 18037 6389 18135 sw
tri 6389 18037 6487 18135 ne
rect 6487 18037 6841 18135
tri 6841 18037 6939 18135 sw
tri 6939 18037 7037 18135 ne
rect 7037 18037 7391 18135
tri 7391 18037 7489 18135 sw
tri 7489 18037 7587 18135 ne
rect 7587 18037 7941 18135
tri 7941 18037 8039 18135 sw
tri 8039 18037 8137 18135 ne
rect 8137 18037 8491 18135
tri 8491 18037 8589 18135 sw
tri 8589 18037 8687 18135 ne
rect 8687 18037 9041 18135
tri 9041 18037 9139 18135 sw
tri 9139 18037 9237 18135 ne
rect 9237 18037 9591 18135
tri 9591 18037 9689 18135 sw
tri 9689 18037 9787 18135 ne
rect 9787 18037 10141 18135
tri 10141 18037 10239 18135 sw
tri 10239 18037 10337 18135 ne
rect 10337 18037 10691 18135
tri 10691 18037 10789 18135 sw
tri 10789 18037 10887 18135 ne
rect 10887 18037 11241 18135
tri 11241 18037 11339 18135 sw
tri 11339 18037 11437 18135 ne
rect 11437 18037 11791 18135
tri 11791 18037 11889 18135 sw
tri 11889 18037 11987 18135 ne
rect 11987 18037 12341 18135
tri 12341 18037 12439 18135 sw
tri 12439 18037 12537 18135 ne
rect 12537 18037 12891 18135
tri 12891 18037 12989 18135 sw
tri 12989 18037 13087 18135 ne
rect 13087 18037 13441 18135
tri 13441 18037 13539 18135 sw
tri 13539 18037 13637 18135 ne
rect 13637 18037 13991 18135
tri 13991 18037 14089 18135 sw
tri 14089 18037 14187 18135 ne
rect 14187 18037 14541 18135
tri 14541 18037 14639 18135 sw
tri 14639 18037 14737 18135 ne
rect 14737 18037 15091 18135
tri 15091 18037 15189 18135 sw
tri 15189 18037 15287 18135 ne
rect 15287 18037 15641 18135
tri 15641 18037 15739 18135 sw
tri 15739 18037 15837 18135 ne
rect 15837 18037 16191 18135
tri 16191 18037 16289 18135 sw
tri 16289 18037 16387 18135 ne
rect 16387 18037 16741 18135
tri 16741 18037 16839 18135 sw
tri 16839 18037 16937 18135 ne
rect 16937 18037 17291 18135
tri 17291 18037 17389 18135 sw
tri 17389 18037 17487 18135 ne
rect 17487 18037 17841 18135
tri 17841 18037 17939 18135 sw
tri 17939 18037 18037 18135 ne
rect 18037 18037 18391 18135
tri 18391 18037 18489 18135 sw
tri 18489 18037 18587 18135 ne
rect 18587 18037 18941 18135
tri 18941 18037 19039 18135 sw
tri 19039 18037 19137 18135 ne
rect 19137 18037 19491 18135
tri 19491 18037 19589 18135 sw
tri 19589 18037 19687 18135 ne
rect 19687 18037 21800 18135
rect -300 17987 339 18037
rect -500 17939 339 17987
tri 339 17939 437 18037 sw
tri 437 17939 535 18037 ne
rect 535 17939 889 18037
tri 889 17939 987 18037 sw
tri 987 17939 1085 18037 ne
rect 1085 17939 1439 18037
tri 1439 17939 1537 18037 sw
tri 1537 17939 1635 18037 ne
rect 1635 17939 1989 18037
tri 1989 17939 2087 18037 sw
tri 2087 17939 2185 18037 ne
rect 2185 17939 2539 18037
tri 2539 17939 2637 18037 sw
tri 2637 17939 2735 18037 ne
rect 2735 17939 3089 18037
tri 3089 17939 3187 18037 sw
tri 3187 17939 3285 18037 ne
rect 3285 17939 3639 18037
tri 3639 17939 3737 18037 sw
tri 3737 17939 3835 18037 ne
rect 3835 17939 4189 18037
tri 4189 17939 4287 18037 sw
tri 4287 17939 4385 18037 ne
rect 4385 17939 4739 18037
tri 4739 17939 4837 18037 sw
tri 4837 17939 4935 18037 ne
rect 4935 17939 5289 18037
tri 5289 17939 5387 18037 sw
tri 5387 17939 5485 18037 ne
rect 5485 17939 5839 18037
tri 5839 17939 5937 18037 sw
tri 5937 17939 6035 18037 ne
rect 6035 17939 6389 18037
tri 6389 17939 6487 18037 sw
tri 6487 17939 6585 18037 ne
rect 6585 17939 6939 18037
tri 6939 17939 7037 18037 sw
tri 7037 17939 7135 18037 ne
rect 7135 17939 7489 18037
tri 7489 17939 7587 18037 sw
tri 7587 17939 7685 18037 ne
rect 7685 17939 8039 18037
tri 8039 17939 8137 18037 sw
tri 8137 17939 8235 18037 ne
rect 8235 17939 8589 18037
tri 8589 17939 8687 18037 sw
tri 8687 17939 8785 18037 ne
rect 8785 17939 9139 18037
tri 9139 17939 9237 18037 sw
tri 9237 17939 9335 18037 ne
rect 9335 17939 9689 18037
tri 9689 17939 9787 18037 sw
tri 9787 17939 9885 18037 ne
rect 9885 17939 10239 18037
tri 10239 17939 10337 18037 sw
tri 10337 17939 10435 18037 ne
rect 10435 17939 10789 18037
tri 10789 17939 10887 18037 sw
tri 10887 17939 10985 18037 ne
rect 10985 17939 11339 18037
tri 11339 17939 11437 18037 sw
tri 11437 17939 11535 18037 ne
rect 11535 17939 11889 18037
tri 11889 17939 11987 18037 sw
tri 11987 17939 12085 18037 ne
rect 12085 17939 12439 18037
tri 12439 17939 12537 18037 sw
tri 12537 17939 12635 18037 ne
rect 12635 17939 12989 18037
tri 12989 17939 13087 18037 sw
tri 13087 17939 13185 18037 ne
rect 13185 17939 13539 18037
tri 13539 17939 13637 18037 sw
tri 13637 17939 13735 18037 ne
rect 13735 17939 14089 18037
tri 14089 17939 14187 18037 sw
tri 14187 17939 14285 18037 ne
rect 14285 17939 14639 18037
tri 14639 17939 14737 18037 sw
tri 14737 17939 14835 18037 ne
rect 14835 17939 15189 18037
tri 15189 17939 15287 18037 sw
tri 15287 17939 15385 18037 ne
rect 15385 17939 15739 18037
tri 15739 17939 15837 18037 sw
tri 15837 17939 15935 18037 ne
rect 15935 17939 16289 18037
tri 16289 17939 16387 18037 sw
tri 16387 17939 16485 18037 ne
rect 16485 17939 16839 18037
tri 16839 17939 16937 18037 sw
tri 16937 17939 17035 18037 ne
rect 17035 17939 17389 18037
tri 17389 17939 17487 18037 sw
tri 17487 17939 17585 18037 ne
rect 17585 17939 17939 18037
tri 17939 17939 18037 18037 sw
tri 18037 17939 18135 18037 ne
rect 18135 17939 18489 18037
tri 18489 17939 18587 18037 sw
tri 18587 17939 18685 18037 ne
rect 18685 17939 19039 18037
tri 19039 17939 19137 18037 sw
tri 19137 17939 19235 18037 ne
rect 19235 17939 19589 18037
tri 19589 17939 19687 18037 sw
rect -500 17935 437 17939
rect -500 17815 215 17935
rect 335 17841 437 17935
tri 437 17841 535 17939 sw
tri 535 17841 633 17939 ne
rect 633 17935 987 17939
rect 633 17841 765 17935
rect 335 17815 535 17841
rect -500 17811 535 17815
tri 535 17811 565 17841 sw
tri 633 17811 663 17841 ne
rect 663 17815 765 17841
rect 885 17841 987 17935
tri 987 17841 1085 17939 sw
tri 1085 17841 1183 17939 ne
rect 1183 17935 1537 17939
rect 1183 17841 1315 17935
rect 885 17815 1085 17841
rect 663 17811 1085 17815
tri 1085 17811 1115 17841 sw
tri 1183 17811 1213 17841 ne
rect 1213 17815 1315 17841
rect 1435 17841 1537 17935
tri 1537 17841 1635 17939 sw
tri 1635 17841 1733 17939 ne
rect 1733 17935 2087 17939
rect 1733 17841 1865 17935
rect 1435 17815 1635 17841
rect 1213 17811 1635 17815
tri 1635 17811 1665 17841 sw
tri 1733 17811 1763 17841 ne
rect 1763 17815 1865 17841
rect 1985 17841 2087 17935
tri 2087 17841 2185 17939 sw
tri 2185 17841 2283 17939 ne
rect 2283 17935 2637 17939
rect 2283 17841 2415 17935
rect 1985 17815 2185 17841
rect 1763 17811 2185 17815
tri 2185 17811 2215 17841 sw
tri 2283 17811 2313 17841 ne
rect 2313 17815 2415 17841
rect 2535 17841 2637 17935
tri 2637 17841 2735 17939 sw
tri 2735 17841 2833 17939 ne
rect 2833 17935 3187 17939
rect 2833 17841 2965 17935
rect 2535 17815 2735 17841
rect 2313 17811 2735 17815
tri 2735 17811 2765 17841 sw
tri 2833 17811 2863 17841 ne
rect 2863 17815 2965 17841
rect 3085 17841 3187 17935
tri 3187 17841 3285 17939 sw
tri 3285 17841 3383 17939 ne
rect 3383 17935 3737 17939
rect 3383 17841 3515 17935
rect 3085 17815 3285 17841
rect 2863 17811 3285 17815
tri 3285 17811 3315 17841 sw
tri 3383 17811 3413 17841 ne
rect 3413 17815 3515 17841
rect 3635 17841 3737 17935
tri 3737 17841 3835 17939 sw
tri 3835 17841 3933 17939 ne
rect 3933 17935 4287 17939
rect 3933 17841 4065 17935
rect 3635 17815 3835 17841
rect 3413 17811 3835 17815
tri 3835 17811 3865 17841 sw
tri 3933 17811 3963 17841 ne
rect 3963 17815 4065 17841
rect 4185 17841 4287 17935
tri 4287 17841 4385 17939 sw
tri 4385 17841 4483 17939 ne
rect 4483 17935 4837 17939
rect 4483 17841 4615 17935
rect 4185 17815 4385 17841
rect 3963 17811 4385 17815
tri 4385 17811 4415 17841 sw
tri 4483 17811 4513 17841 ne
rect 4513 17815 4615 17841
rect 4735 17841 4837 17935
tri 4837 17841 4935 17939 sw
tri 4935 17841 5033 17939 ne
rect 5033 17935 5387 17939
rect 5033 17841 5165 17935
rect 4735 17815 4935 17841
rect 4513 17811 4935 17815
tri 4935 17811 4965 17841 sw
tri 5033 17811 5063 17841 ne
rect 5063 17815 5165 17841
rect 5285 17841 5387 17935
tri 5387 17841 5485 17939 sw
tri 5485 17841 5583 17939 ne
rect 5583 17935 5937 17939
rect 5583 17841 5715 17935
rect 5285 17815 5485 17841
rect 5063 17811 5485 17815
tri 5485 17811 5515 17841 sw
tri 5583 17811 5613 17841 ne
rect 5613 17815 5715 17841
rect 5835 17841 5937 17935
tri 5937 17841 6035 17939 sw
tri 6035 17841 6133 17939 ne
rect 6133 17935 6487 17939
rect 6133 17841 6265 17935
rect 5835 17815 6035 17841
rect 5613 17811 6035 17815
tri 6035 17811 6065 17841 sw
tri 6133 17811 6163 17841 ne
rect 6163 17815 6265 17841
rect 6385 17841 6487 17935
tri 6487 17841 6585 17939 sw
tri 6585 17841 6683 17939 ne
rect 6683 17935 7037 17939
rect 6683 17841 6815 17935
rect 6385 17815 6585 17841
rect 6163 17811 6585 17815
tri 6585 17811 6615 17841 sw
tri 6683 17811 6713 17841 ne
rect 6713 17815 6815 17841
rect 6935 17841 7037 17935
tri 7037 17841 7135 17939 sw
tri 7135 17841 7233 17939 ne
rect 7233 17935 7587 17939
rect 7233 17841 7365 17935
rect 6935 17815 7135 17841
rect 6713 17811 7135 17815
tri 7135 17811 7165 17841 sw
tri 7233 17811 7263 17841 ne
rect 7263 17815 7365 17841
rect 7485 17841 7587 17935
tri 7587 17841 7685 17939 sw
tri 7685 17841 7783 17939 ne
rect 7783 17935 8137 17939
rect 7783 17841 7915 17935
rect 7485 17815 7685 17841
rect 7263 17811 7685 17815
tri 7685 17811 7715 17841 sw
tri 7783 17811 7813 17841 ne
rect 7813 17815 7915 17841
rect 8035 17841 8137 17935
tri 8137 17841 8235 17939 sw
tri 8235 17841 8333 17939 ne
rect 8333 17935 8687 17939
rect 8333 17841 8465 17935
rect 8035 17815 8235 17841
rect 7813 17811 8235 17815
tri 8235 17811 8265 17841 sw
tri 8333 17811 8363 17841 ne
rect 8363 17815 8465 17841
rect 8585 17841 8687 17935
tri 8687 17841 8785 17939 sw
tri 8785 17841 8883 17939 ne
rect 8883 17935 9237 17939
rect 8883 17841 9015 17935
rect 8585 17815 8785 17841
rect 8363 17811 8785 17815
tri 8785 17811 8815 17841 sw
tri 8883 17811 8913 17841 ne
rect 8913 17815 9015 17841
rect 9135 17841 9237 17935
tri 9237 17841 9335 17939 sw
tri 9335 17841 9433 17939 ne
rect 9433 17935 9787 17939
rect 9433 17841 9565 17935
rect 9135 17815 9335 17841
rect 8913 17811 9335 17815
tri 9335 17811 9365 17841 sw
tri 9433 17811 9463 17841 ne
rect 9463 17815 9565 17841
rect 9685 17841 9787 17935
tri 9787 17841 9885 17939 sw
tri 9885 17841 9983 17939 ne
rect 9983 17935 10337 17939
rect 9983 17841 10115 17935
rect 9685 17815 9885 17841
rect 9463 17811 9885 17815
tri 9885 17811 9915 17841 sw
tri 9983 17811 10013 17841 ne
rect 10013 17815 10115 17841
rect 10235 17841 10337 17935
tri 10337 17841 10435 17939 sw
tri 10435 17841 10533 17939 ne
rect 10533 17935 10887 17939
rect 10533 17841 10665 17935
rect 10235 17815 10435 17841
rect 10013 17811 10435 17815
tri 10435 17811 10465 17841 sw
tri 10533 17811 10563 17841 ne
rect 10563 17815 10665 17841
rect 10785 17841 10887 17935
tri 10887 17841 10985 17939 sw
tri 10985 17841 11083 17939 ne
rect 11083 17935 11437 17939
rect 11083 17841 11215 17935
rect 10785 17815 10985 17841
rect 10563 17811 10985 17815
tri 10985 17811 11015 17841 sw
tri 11083 17811 11113 17841 ne
rect 11113 17815 11215 17841
rect 11335 17841 11437 17935
tri 11437 17841 11535 17939 sw
tri 11535 17841 11633 17939 ne
rect 11633 17935 11987 17939
rect 11633 17841 11765 17935
rect 11335 17815 11535 17841
rect 11113 17811 11535 17815
tri 11535 17811 11565 17841 sw
tri 11633 17811 11663 17841 ne
rect 11663 17815 11765 17841
rect 11885 17841 11987 17935
tri 11987 17841 12085 17939 sw
tri 12085 17841 12183 17939 ne
rect 12183 17935 12537 17939
rect 12183 17841 12315 17935
rect 11885 17815 12085 17841
rect 11663 17811 12085 17815
tri 12085 17811 12115 17841 sw
tri 12183 17811 12213 17841 ne
rect 12213 17815 12315 17841
rect 12435 17841 12537 17935
tri 12537 17841 12635 17939 sw
tri 12635 17841 12733 17939 ne
rect 12733 17935 13087 17939
rect 12733 17841 12865 17935
rect 12435 17815 12635 17841
rect 12213 17811 12635 17815
tri 12635 17811 12665 17841 sw
tri 12733 17811 12763 17841 ne
rect 12763 17815 12865 17841
rect 12985 17841 13087 17935
tri 13087 17841 13185 17939 sw
tri 13185 17841 13283 17939 ne
rect 13283 17935 13637 17939
rect 13283 17841 13415 17935
rect 12985 17815 13185 17841
rect 12763 17811 13185 17815
tri 13185 17811 13215 17841 sw
tri 13283 17811 13313 17841 ne
rect 13313 17815 13415 17841
rect 13535 17841 13637 17935
tri 13637 17841 13735 17939 sw
tri 13735 17841 13833 17939 ne
rect 13833 17935 14187 17939
rect 13833 17841 13965 17935
rect 13535 17815 13735 17841
rect 13313 17811 13735 17815
tri 13735 17811 13765 17841 sw
tri 13833 17811 13863 17841 ne
rect 13863 17815 13965 17841
rect 14085 17841 14187 17935
tri 14187 17841 14285 17939 sw
tri 14285 17841 14383 17939 ne
rect 14383 17935 14737 17939
rect 14383 17841 14515 17935
rect 14085 17815 14285 17841
rect 13863 17811 14285 17815
tri 14285 17811 14315 17841 sw
tri 14383 17811 14413 17841 ne
rect 14413 17815 14515 17841
rect 14635 17841 14737 17935
tri 14737 17841 14835 17939 sw
tri 14835 17841 14933 17939 ne
rect 14933 17935 15287 17939
rect 14933 17841 15065 17935
rect 14635 17815 14835 17841
rect 14413 17811 14835 17815
tri 14835 17811 14865 17841 sw
tri 14933 17811 14963 17841 ne
rect 14963 17815 15065 17841
rect 15185 17841 15287 17935
tri 15287 17841 15385 17939 sw
tri 15385 17841 15483 17939 ne
rect 15483 17935 15837 17939
rect 15483 17841 15615 17935
rect 15185 17815 15385 17841
rect 14963 17811 15385 17815
tri 15385 17811 15415 17841 sw
tri 15483 17811 15513 17841 ne
rect 15513 17815 15615 17841
rect 15735 17841 15837 17935
tri 15837 17841 15935 17939 sw
tri 15935 17841 16033 17939 ne
rect 16033 17935 16387 17939
rect 16033 17841 16165 17935
rect 15735 17815 15935 17841
rect 15513 17811 15935 17815
tri 15935 17811 15965 17841 sw
tri 16033 17811 16063 17841 ne
rect 16063 17815 16165 17841
rect 16285 17841 16387 17935
tri 16387 17841 16485 17939 sw
tri 16485 17841 16583 17939 ne
rect 16583 17935 16937 17939
rect 16583 17841 16715 17935
rect 16285 17815 16485 17841
rect 16063 17811 16485 17815
tri 16485 17811 16515 17841 sw
tri 16583 17811 16613 17841 ne
rect 16613 17815 16715 17841
rect 16835 17841 16937 17935
tri 16937 17841 17035 17939 sw
tri 17035 17841 17133 17939 ne
rect 17133 17935 17487 17939
rect 17133 17841 17265 17935
rect 16835 17815 17035 17841
rect 16613 17811 17035 17815
tri 17035 17811 17065 17841 sw
tri 17133 17811 17163 17841 ne
rect 17163 17815 17265 17841
rect 17385 17841 17487 17935
tri 17487 17841 17585 17939 sw
tri 17585 17841 17683 17939 ne
rect 17683 17935 18037 17939
rect 17683 17841 17815 17935
rect 17385 17815 17585 17841
rect 17163 17811 17585 17815
tri 17585 17811 17615 17841 sw
tri 17683 17811 17713 17841 ne
rect 17713 17815 17815 17841
rect 17935 17841 18037 17935
tri 18037 17841 18135 17939 sw
tri 18135 17841 18233 17939 ne
rect 18233 17935 18587 17939
rect 18233 17841 18365 17935
rect 17935 17815 18135 17841
rect 17713 17811 18135 17815
tri 18135 17811 18165 17841 sw
tri 18233 17811 18263 17841 ne
rect 18263 17815 18365 17841
rect 18485 17841 18587 17935
tri 18587 17841 18685 17939 sw
tri 18685 17841 18783 17939 ne
rect 18783 17935 19137 17939
rect 18783 17841 18915 17935
rect 18485 17815 18685 17841
rect 18263 17811 18685 17815
tri 18685 17811 18715 17841 sw
tri 18783 17811 18813 17841 ne
rect 18813 17815 18915 17841
rect 19035 17841 19137 17935
tri 19137 17841 19235 17939 sw
tri 19235 17841 19333 17939 ne
rect 19333 17935 20300 17939
rect 19333 17841 19465 17935
rect 19035 17815 19235 17841
rect 18813 17811 19235 17815
tri 19235 17811 19265 17841 sw
tri 19333 17811 19363 17841 ne
rect 19363 17815 19465 17841
rect 19585 17815 20300 17935
rect 19363 17811 20300 17815
tri 113 17713 211 17811 ne
rect 211 17713 565 17811
tri 565 17713 663 17811 sw
tri 663 17713 761 17811 ne
rect 761 17713 1115 17811
tri 1115 17713 1213 17811 sw
tri 1213 17713 1311 17811 ne
rect 1311 17713 1665 17811
tri 1665 17713 1763 17811 sw
tri 1763 17713 1861 17811 ne
rect 1861 17713 2215 17811
tri 2215 17713 2313 17811 sw
tri 2313 17713 2411 17811 ne
rect 2411 17713 2765 17811
tri 2765 17713 2863 17811 sw
tri 2863 17713 2961 17811 ne
rect 2961 17713 3315 17811
tri 3315 17713 3413 17811 sw
tri 3413 17713 3511 17811 ne
rect 3511 17713 3865 17811
tri 3865 17713 3963 17811 sw
tri 3963 17713 4061 17811 ne
rect 4061 17713 4415 17811
tri 4415 17713 4513 17811 sw
tri 4513 17713 4611 17811 ne
rect 4611 17713 4965 17811
tri 4965 17713 5063 17811 sw
tri 5063 17713 5161 17811 ne
rect 5161 17713 5515 17811
tri 5515 17713 5613 17811 sw
tri 5613 17713 5711 17811 ne
rect 5711 17713 6065 17811
tri 6065 17713 6163 17811 sw
tri 6163 17713 6261 17811 ne
rect 6261 17713 6615 17811
tri 6615 17713 6713 17811 sw
tri 6713 17713 6811 17811 ne
rect 6811 17713 7165 17811
tri 7165 17713 7263 17811 sw
tri 7263 17713 7361 17811 ne
rect 7361 17713 7715 17811
tri 7715 17713 7813 17811 sw
tri 7813 17713 7911 17811 ne
rect 7911 17713 8265 17811
tri 8265 17713 8363 17811 sw
tri 8363 17713 8461 17811 ne
rect 8461 17713 8815 17811
tri 8815 17713 8913 17811 sw
tri 8913 17713 9011 17811 ne
rect 9011 17713 9365 17811
tri 9365 17713 9463 17811 sw
tri 9463 17713 9561 17811 ne
rect 9561 17713 9915 17811
tri 9915 17713 10013 17811 sw
tri 10013 17713 10111 17811 ne
rect 10111 17713 10465 17811
tri 10465 17713 10563 17811 sw
tri 10563 17713 10661 17811 ne
rect 10661 17713 11015 17811
tri 11015 17713 11113 17811 sw
tri 11113 17713 11211 17811 ne
rect 11211 17713 11565 17811
tri 11565 17713 11663 17811 sw
tri 11663 17713 11761 17811 ne
rect 11761 17713 12115 17811
tri 12115 17713 12213 17811 sw
tri 12213 17713 12311 17811 ne
rect 12311 17713 12665 17811
tri 12665 17713 12763 17811 sw
tri 12763 17713 12861 17811 ne
rect 12861 17713 13215 17811
tri 13215 17713 13313 17811 sw
tri 13313 17713 13411 17811 ne
rect 13411 17713 13765 17811
tri 13765 17713 13863 17811 sw
tri 13863 17713 13961 17811 ne
rect 13961 17713 14315 17811
tri 14315 17713 14413 17811 sw
tri 14413 17713 14511 17811 ne
rect 14511 17713 14865 17811
tri 14865 17713 14963 17811 sw
tri 14963 17713 15061 17811 ne
rect 15061 17713 15415 17811
tri 15415 17713 15513 17811 sw
tri 15513 17713 15611 17811 ne
rect 15611 17713 15965 17811
tri 15965 17713 16063 17811 sw
tri 16063 17713 16161 17811 ne
rect 16161 17713 16515 17811
tri 16515 17713 16613 17811 sw
tri 16613 17713 16711 17811 ne
rect 16711 17713 17065 17811
tri 17065 17713 17163 17811 sw
tri 17163 17713 17261 17811 ne
rect 17261 17713 17615 17811
tri 17615 17713 17713 17811 sw
tri 17713 17713 17811 17811 ne
rect 17811 17713 18165 17811
tri 18165 17713 18263 17811 sw
tri 18263 17713 18361 17811 ne
rect 18361 17713 18715 17811
tri 18715 17713 18813 17811 sw
tri 18813 17713 18911 17811 ne
rect 18911 17713 19265 17811
tri 19265 17713 19363 17811 sw
tri 19363 17713 19461 17811 ne
rect 19461 17713 20300 17811
rect -2000 17683 113 17713
tri 113 17683 143 17713 sw
tri 211 17683 241 17713 ne
rect 241 17683 663 17713
tri 663 17683 693 17713 sw
tri 761 17683 791 17713 ne
rect 791 17683 1213 17713
tri 1213 17683 1243 17713 sw
tri 1311 17683 1341 17713 ne
rect 1341 17683 1763 17713
tri 1763 17683 1793 17713 sw
tri 1861 17683 1891 17713 ne
rect 1891 17683 2313 17713
tri 2313 17683 2343 17713 sw
tri 2411 17683 2441 17713 ne
rect 2441 17683 2863 17713
tri 2863 17683 2893 17713 sw
tri 2961 17683 2991 17713 ne
rect 2991 17683 3413 17713
tri 3413 17683 3443 17713 sw
tri 3511 17683 3541 17713 ne
rect 3541 17683 3963 17713
tri 3963 17683 3993 17713 sw
tri 4061 17683 4091 17713 ne
rect 4091 17683 4513 17713
tri 4513 17683 4543 17713 sw
tri 4611 17683 4641 17713 ne
rect 4641 17683 5063 17713
tri 5063 17683 5093 17713 sw
tri 5161 17683 5191 17713 ne
rect 5191 17683 5613 17713
tri 5613 17683 5643 17713 sw
tri 5711 17683 5741 17713 ne
rect 5741 17683 6163 17713
tri 6163 17683 6193 17713 sw
tri 6261 17683 6291 17713 ne
rect 6291 17683 6713 17713
tri 6713 17683 6743 17713 sw
tri 6811 17683 6841 17713 ne
rect 6841 17683 7263 17713
tri 7263 17683 7293 17713 sw
tri 7361 17683 7391 17713 ne
rect 7391 17683 7813 17713
tri 7813 17683 7843 17713 sw
tri 7911 17683 7941 17713 ne
rect 7941 17683 8363 17713
tri 8363 17683 8393 17713 sw
tri 8461 17683 8491 17713 ne
rect 8491 17683 8913 17713
tri 8913 17683 8943 17713 sw
tri 9011 17683 9041 17713 ne
rect 9041 17683 9463 17713
tri 9463 17683 9493 17713 sw
tri 9561 17683 9591 17713 ne
rect 9591 17683 10013 17713
tri 10013 17683 10043 17713 sw
tri 10111 17683 10141 17713 ne
rect 10141 17683 10563 17713
tri 10563 17683 10593 17713 sw
tri 10661 17683 10691 17713 ne
rect 10691 17683 11113 17713
tri 11113 17683 11143 17713 sw
tri 11211 17683 11241 17713 ne
rect 11241 17683 11663 17713
tri 11663 17683 11693 17713 sw
tri 11761 17683 11791 17713 ne
rect 11791 17683 12213 17713
tri 12213 17683 12243 17713 sw
tri 12311 17683 12341 17713 ne
rect 12341 17683 12763 17713
tri 12763 17683 12793 17713 sw
tri 12861 17683 12891 17713 ne
rect 12891 17683 13313 17713
tri 13313 17683 13343 17713 sw
tri 13411 17683 13441 17713 ne
rect 13441 17683 13863 17713
tri 13863 17683 13893 17713 sw
tri 13961 17683 13991 17713 ne
rect 13991 17683 14413 17713
tri 14413 17683 14443 17713 sw
tri 14511 17683 14541 17713 ne
rect 14541 17683 14963 17713
tri 14963 17683 14993 17713 sw
tri 15061 17683 15091 17713 ne
rect 15091 17683 15513 17713
tri 15513 17683 15543 17713 sw
tri 15611 17683 15641 17713 ne
rect 15641 17683 16063 17713
tri 16063 17683 16093 17713 sw
tri 16161 17683 16191 17713 ne
rect 16191 17683 16613 17713
tri 16613 17683 16643 17713 sw
tri 16711 17683 16741 17713 ne
rect 16741 17683 17163 17713
tri 17163 17683 17193 17713 sw
tri 17261 17683 17291 17713 ne
rect 17291 17683 17713 17713
tri 17713 17683 17743 17713 sw
tri 17811 17683 17841 17713 ne
rect 17841 17683 18263 17713
tri 18263 17683 18293 17713 sw
tri 18361 17683 18391 17713 ne
rect 18391 17683 18813 17713
tri 18813 17683 18843 17713 sw
tri 18911 17683 18941 17713 ne
rect 18941 17683 19363 17713
tri 19363 17683 19393 17713 sw
tri 19461 17683 19491 17713 ne
rect 19491 17683 20300 17713
rect -2000 17585 143 17683
tri 143 17585 241 17683 sw
tri 241 17585 339 17683 ne
rect 339 17585 693 17683
tri 693 17585 791 17683 sw
tri 791 17585 889 17683 ne
rect 889 17585 1243 17683
tri 1243 17585 1341 17683 sw
tri 1341 17585 1439 17683 ne
rect 1439 17585 1793 17683
tri 1793 17585 1891 17683 sw
tri 1891 17585 1989 17683 ne
rect 1989 17585 2343 17683
tri 2343 17585 2441 17683 sw
tri 2441 17585 2539 17683 ne
rect 2539 17585 2893 17683
tri 2893 17585 2991 17683 sw
tri 2991 17585 3089 17683 ne
rect 3089 17585 3443 17683
tri 3443 17585 3541 17683 sw
tri 3541 17585 3639 17683 ne
rect 3639 17585 3993 17683
tri 3993 17585 4091 17683 sw
tri 4091 17585 4189 17683 ne
rect 4189 17585 4543 17683
tri 4543 17585 4641 17683 sw
tri 4641 17585 4739 17683 ne
rect 4739 17585 5093 17683
tri 5093 17585 5191 17683 sw
tri 5191 17585 5289 17683 ne
rect 5289 17585 5643 17683
tri 5643 17585 5741 17683 sw
tri 5741 17585 5839 17683 ne
rect 5839 17585 6193 17683
tri 6193 17585 6291 17683 sw
tri 6291 17585 6389 17683 ne
rect 6389 17585 6743 17683
tri 6743 17585 6841 17683 sw
tri 6841 17585 6939 17683 ne
rect 6939 17585 7293 17683
tri 7293 17585 7391 17683 sw
tri 7391 17585 7489 17683 ne
rect 7489 17585 7843 17683
tri 7843 17585 7941 17683 sw
tri 7941 17585 8039 17683 ne
rect 8039 17585 8393 17683
tri 8393 17585 8491 17683 sw
tri 8491 17585 8589 17683 ne
rect 8589 17585 8943 17683
tri 8943 17585 9041 17683 sw
tri 9041 17585 9139 17683 ne
rect 9139 17585 9493 17683
tri 9493 17585 9591 17683 sw
tri 9591 17585 9689 17683 ne
rect 9689 17585 10043 17683
tri 10043 17585 10141 17683 sw
tri 10141 17585 10239 17683 ne
rect 10239 17585 10593 17683
tri 10593 17585 10691 17683 sw
tri 10691 17585 10789 17683 ne
rect 10789 17585 11143 17683
tri 11143 17585 11241 17683 sw
tri 11241 17585 11339 17683 ne
rect 11339 17585 11693 17683
tri 11693 17585 11791 17683 sw
tri 11791 17585 11889 17683 ne
rect 11889 17585 12243 17683
tri 12243 17585 12341 17683 sw
tri 12341 17585 12439 17683 ne
rect 12439 17585 12793 17683
tri 12793 17585 12891 17683 sw
tri 12891 17585 12989 17683 ne
rect 12989 17585 13343 17683
tri 13343 17585 13441 17683 sw
tri 13441 17585 13539 17683 ne
rect 13539 17585 13893 17683
tri 13893 17585 13991 17683 sw
tri 13991 17585 14089 17683 ne
rect 14089 17585 14443 17683
tri 14443 17585 14541 17683 sw
tri 14541 17585 14639 17683 ne
rect 14639 17585 14993 17683
tri 14993 17585 15091 17683 sw
tri 15091 17585 15189 17683 ne
rect 15189 17585 15543 17683
tri 15543 17585 15641 17683 sw
tri 15641 17585 15739 17683 ne
rect 15739 17585 16093 17683
tri 16093 17585 16191 17683 sw
tri 16191 17585 16289 17683 ne
rect 16289 17585 16643 17683
tri 16643 17585 16741 17683 sw
tri 16741 17585 16839 17683 ne
rect 16839 17585 17193 17683
tri 17193 17585 17291 17683 sw
tri 17291 17585 17389 17683 ne
rect 17389 17585 17743 17683
tri 17743 17585 17841 17683 sw
tri 17841 17585 17939 17683 ne
rect 17939 17585 18293 17683
tri 18293 17585 18391 17683 sw
tri 18391 17585 18489 17683 ne
rect 18489 17585 18843 17683
tri 18843 17585 18941 17683 sw
tri 18941 17585 19039 17683 ne
rect 19039 17585 19393 17683
tri 19393 17585 19491 17683 sw
tri 19491 17585 19589 17683 ne
rect 19589 17585 20300 17683
rect -2000 17487 241 17585
tri 241 17487 339 17585 sw
tri 339 17487 437 17585 ne
rect 437 17487 791 17585
tri 791 17487 889 17585 sw
tri 889 17487 987 17585 ne
rect 987 17487 1341 17585
tri 1341 17487 1439 17585 sw
tri 1439 17487 1537 17585 ne
rect 1537 17487 1891 17585
tri 1891 17487 1989 17585 sw
tri 1989 17487 2087 17585 ne
rect 2087 17487 2441 17585
tri 2441 17487 2539 17585 sw
tri 2539 17487 2637 17585 ne
rect 2637 17487 2991 17585
tri 2991 17487 3089 17585 sw
tri 3089 17487 3187 17585 ne
rect 3187 17487 3541 17585
tri 3541 17487 3639 17585 sw
tri 3639 17487 3737 17585 ne
rect 3737 17487 4091 17585
tri 4091 17487 4189 17585 sw
tri 4189 17487 4287 17585 ne
rect 4287 17487 4641 17585
tri 4641 17487 4739 17585 sw
tri 4739 17487 4837 17585 ne
rect 4837 17487 5191 17585
tri 5191 17487 5289 17585 sw
tri 5289 17487 5387 17585 ne
rect 5387 17487 5741 17585
tri 5741 17487 5839 17585 sw
tri 5839 17487 5937 17585 ne
rect 5937 17487 6291 17585
tri 6291 17487 6389 17585 sw
tri 6389 17487 6487 17585 ne
rect 6487 17487 6841 17585
tri 6841 17487 6939 17585 sw
tri 6939 17487 7037 17585 ne
rect 7037 17487 7391 17585
tri 7391 17487 7489 17585 sw
tri 7489 17487 7587 17585 ne
rect 7587 17487 7941 17585
tri 7941 17487 8039 17585 sw
tri 8039 17487 8137 17585 ne
rect 8137 17487 8491 17585
tri 8491 17487 8589 17585 sw
tri 8589 17487 8687 17585 ne
rect 8687 17487 9041 17585
tri 9041 17487 9139 17585 sw
tri 9139 17487 9237 17585 ne
rect 9237 17487 9591 17585
tri 9591 17487 9689 17585 sw
tri 9689 17487 9787 17585 ne
rect 9787 17487 10141 17585
tri 10141 17487 10239 17585 sw
tri 10239 17487 10337 17585 ne
rect 10337 17487 10691 17585
tri 10691 17487 10789 17585 sw
tri 10789 17487 10887 17585 ne
rect 10887 17487 11241 17585
tri 11241 17487 11339 17585 sw
tri 11339 17487 11437 17585 ne
rect 11437 17487 11791 17585
tri 11791 17487 11889 17585 sw
tri 11889 17487 11987 17585 ne
rect 11987 17487 12341 17585
tri 12341 17487 12439 17585 sw
tri 12439 17487 12537 17585 ne
rect 12537 17487 12891 17585
tri 12891 17487 12989 17585 sw
tri 12989 17487 13087 17585 ne
rect 13087 17487 13441 17585
tri 13441 17487 13539 17585 sw
tri 13539 17487 13637 17585 ne
rect 13637 17487 13991 17585
tri 13991 17487 14089 17585 sw
tri 14089 17487 14187 17585 ne
rect 14187 17487 14541 17585
tri 14541 17487 14639 17585 sw
tri 14639 17487 14737 17585 ne
rect 14737 17487 15091 17585
tri 15091 17487 15189 17585 sw
tri 15189 17487 15287 17585 ne
rect 15287 17487 15641 17585
tri 15641 17487 15739 17585 sw
tri 15739 17487 15837 17585 ne
rect 15837 17487 16191 17585
tri 16191 17487 16289 17585 sw
tri 16289 17487 16387 17585 ne
rect 16387 17487 16741 17585
tri 16741 17487 16839 17585 sw
tri 16839 17487 16937 17585 ne
rect 16937 17487 17291 17585
tri 17291 17487 17389 17585 sw
tri 17389 17487 17487 17585 ne
rect 17487 17487 17841 17585
tri 17841 17487 17939 17585 sw
tri 17939 17487 18037 17585 ne
rect 18037 17487 18391 17585
tri 18391 17487 18489 17585 sw
tri 18489 17487 18587 17585 ne
rect 18587 17487 18941 17585
tri 18941 17487 19039 17585 sw
tri 19039 17487 19137 17585 ne
rect 19137 17487 19491 17585
tri 19491 17487 19589 17585 sw
tri 19589 17487 19687 17585 ne
rect 19687 17487 20300 17585
rect -2000 17389 339 17487
tri 339 17389 437 17487 sw
tri 437 17389 535 17487 ne
rect 535 17389 889 17487
tri 889 17389 987 17487 sw
tri 987 17389 1085 17487 ne
rect 1085 17389 1439 17487
tri 1439 17389 1537 17487 sw
tri 1537 17389 1635 17487 ne
rect 1635 17389 1989 17487
tri 1989 17389 2087 17487 sw
tri 2087 17389 2185 17487 ne
rect 2185 17389 2539 17487
tri 2539 17389 2637 17487 sw
tri 2637 17389 2735 17487 ne
rect 2735 17389 3089 17487
tri 3089 17389 3187 17487 sw
tri 3187 17389 3285 17487 ne
rect 3285 17389 3639 17487
tri 3639 17389 3737 17487 sw
tri 3737 17389 3835 17487 ne
rect 3835 17389 4189 17487
tri 4189 17389 4287 17487 sw
tri 4287 17389 4385 17487 ne
rect 4385 17389 4739 17487
tri 4739 17389 4837 17487 sw
tri 4837 17389 4935 17487 ne
rect 4935 17389 5289 17487
tri 5289 17389 5387 17487 sw
tri 5387 17389 5485 17487 ne
rect 5485 17389 5839 17487
tri 5839 17389 5937 17487 sw
tri 5937 17389 6035 17487 ne
rect 6035 17389 6389 17487
tri 6389 17389 6487 17487 sw
tri 6487 17389 6585 17487 ne
rect 6585 17389 6939 17487
tri 6939 17389 7037 17487 sw
tri 7037 17389 7135 17487 ne
rect 7135 17389 7489 17487
tri 7489 17389 7587 17487 sw
tri 7587 17389 7685 17487 ne
rect 7685 17389 8039 17487
tri 8039 17389 8137 17487 sw
tri 8137 17389 8235 17487 ne
rect 8235 17389 8589 17487
tri 8589 17389 8687 17487 sw
tri 8687 17389 8785 17487 ne
rect 8785 17389 9139 17487
tri 9139 17389 9237 17487 sw
tri 9237 17389 9335 17487 ne
rect 9335 17389 9689 17487
tri 9689 17389 9787 17487 sw
tri 9787 17389 9885 17487 ne
rect 9885 17389 10239 17487
tri 10239 17389 10337 17487 sw
tri 10337 17389 10435 17487 ne
rect 10435 17389 10789 17487
tri 10789 17389 10887 17487 sw
tri 10887 17389 10985 17487 ne
rect 10985 17389 11339 17487
tri 11339 17389 11437 17487 sw
tri 11437 17389 11535 17487 ne
rect 11535 17389 11889 17487
tri 11889 17389 11987 17487 sw
tri 11987 17389 12085 17487 ne
rect 12085 17389 12439 17487
tri 12439 17389 12537 17487 sw
tri 12537 17389 12635 17487 ne
rect 12635 17389 12989 17487
tri 12989 17389 13087 17487 sw
tri 13087 17389 13185 17487 ne
rect 13185 17389 13539 17487
tri 13539 17389 13637 17487 sw
tri 13637 17389 13735 17487 ne
rect 13735 17389 14089 17487
tri 14089 17389 14187 17487 sw
tri 14187 17389 14285 17487 ne
rect 14285 17389 14639 17487
tri 14639 17389 14737 17487 sw
tri 14737 17389 14835 17487 ne
rect 14835 17389 15189 17487
tri 15189 17389 15287 17487 sw
tri 15287 17389 15385 17487 ne
rect 15385 17389 15739 17487
tri 15739 17389 15837 17487 sw
tri 15837 17389 15935 17487 ne
rect 15935 17389 16289 17487
tri 16289 17389 16387 17487 sw
tri 16387 17389 16485 17487 ne
rect 16485 17389 16839 17487
tri 16839 17389 16937 17487 sw
tri 16937 17389 17035 17487 ne
rect 17035 17389 17389 17487
tri 17389 17389 17487 17487 sw
tri 17487 17389 17585 17487 ne
rect 17585 17389 17939 17487
tri 17939 17389 18037 17487 sw
tri 18037 17389 18135 17487 ne
rect 18135 17389 18489 17487
tri 18489 17389 18587 17487 sw
tri 18587 17389 18685 17487 ne
rect 18685 17389 19039 17487
tri 19039 17389 19137 17487 sw
tri 19137 17389 19235 17487 ne
rect 19235 17389 19589 17487
tri 19589 17389 19687 17487 sw
rect 20800 17389 21800 18037
rect -2000 17385 437 17389
rect -2000 17265 215 17385
rect 335 17291 437 17385
tri 437 17291 535 17389 sw
tri 535 17291 633 17389 ne
rect 633 17385 987 17389
rect 633 17291 765 17385
rect 335 17265 535 17291
rect -2000 17261 535 17265
rect -2000 16613 -1000 17261
tri 113 17163 211 17261 ne
rect 211 17213 535 17261
tri 535 17213 613 17291 sw
tri 633 17213 711 17291 ne
rect 711 17265 765 17291
rect 885 17291 987 17385
tri 987 17291 1085 17389 sw
tri 1085 17291 1183 17389 ne
rect 1183 17385 1537 17389
rect 1183 17291 1315 17385
rect 885 17265 1085 17291
rect 711 17213 1085 17265
tri 1085 17213 1163 17291 sw
tri 1183 17213 1261 17291 ne
rect 1261 17265 1315 17291
rect 1435 17291 1537 17385
tri 1537 17291 1635 17389 sw
tri 1635 17291 1733 17389 ne
rect 1733 17385 2087 17389
rect 1733 17291 1865 17385
rect 1435 17265 1635 17291
rect 1261 17213 1635 17265
tri 1635 17213 1713 17291 sw
tri 1733 17213 1811 17291 ne
rect 1811 17265 1865 17291
rect 1985 17291 2087 17385
tri 2087 17291 2185 17389 sw
tri 2185 17291 2283 17389 ne
rect 2283 17385 2637 17389
rect 2283 17291 2415 17385
rect 1985 17265 2185 17291
rect 1811 17213 2185 17265
tri 2185 17213 2263 17291 sw
tri 2283 17213 2361 17291 ne
rect 2361 17265 2415 17291
rect 2535 17291 2637 17385
tri 2637 17291 2735 17389 sw
tri 2735 17291 2833 17389 ne
rect 2833 17385 3187 17389
rect 2833 17291 2965 17385
rect 2535 17265 2735 17291
rect 2361 17213 2735 17265
tri 2735 17213 2813 17291 sw
tri 2833 17213 2911 17291 ne
rect 2911 17265 2965 17291
rect 3085 17291 3187 17385
tri 3187 17291 3285 17389 sw
tri 3285 17291 3383 17389 ne
rect 3383 17385 3737 17389
rect 3383 17291 3515 17385
rect 3085 17265 3285 17291
rect 2911 17213 3285 17265
tri 3285 17213 3363 17291 sw
tri 3383 17213 3461 17291 ne
rect 3461 17265 3515 17291
rect 3635 17291 3737 17385
tri 3737 17291 3835 17389 sw
tri 3835 17291 3933 17389 ne
rect 3933 17385 4287 17389
rect 3933 17291 4065 17385
rect 3635 17265 3835 17291
rect 3461 17213 3835 17265
tri 3835 17213 3913 17291 sw
tri 3933 17213 4011 17291 ne
rect 4011 17265 4065 17291
rect 4185 17291 4287 17385
tri 4287 17291 4385 17389 sw
tri 4385 17291 4483 17389 ne
rect 4483 17385 4837 17389
rect 4483 17291 4615 17385
rect 4185 17265 4385 17291
rect 4011 17213 4385 17265
tri 4385 17213 4463 17291 sw
tri 4483 17213 4561 17291 ne
rect 4561 17265 4615 17291
rect 4735 17291 4837 17385
tri 4837 17291 4935 17389 sw
tri 4935 17291 5033 17389 ne
rect 5033 17385 5387 17389
rect 5033 17291 5165 17385
rect 4735 17265 4935 17291
rect 4561 17213 4935 17265
tri 4935 17213 5013 17291 sw
tri 5033 17213 5111 17291 ne
rect 5111 17265 5165 17291
rect 5285 17291 5387 17385
tri 5387 17291 5485 17389 sw
tri 5485 17291 5583 17389 ne
rect 5583 17385 5937 17389
rect 5583 17291 5715 17385
rect 5285 17265 5485 17291
rect 5111 17213 5485 17265
tri 5485 17213 5563 17291 sw
tri 5583 17213 5661 17291 ne
rect 5661 17265 5715 17291
rect 5835 17291 5937 17385
tri 5937 17291 6035 17389 sw
tri 6035 17291 6133 17389 ne
rect 6133 17385 6487 17389
rect 6133 17291 6265 17385
rect 5835 17265 6035 17291
rect 5661 17213 6035 17265
tri 6035 17213 6113 17291 sw
tri 6133 17213 6211 17291 ne
rect 6211 17265 6265 17291
rect 6385 17291 6487 17385
tri 6487 17291 6585 17389 sw
tri 6585 17291 6683 17389 ne
rect 6683 17385 7037 17389
rect 6683 17291 6815 17385
rect 6385 17265 6585 17291
rect 6211 17213 6585 17265
tri 6585 17213 6663 17291 sw
tri 6683 17213 6761 17291 ne
rect 6761 17265 6815 17291
rect 6935 17291 7037 17385
tri 7037 17291 7135 17389 sw
tri 7135 17291 7233 17389 ne
rect 7233 17385 7587 17389
rect 7233 17291 7365 17385
rect 6935 17265 7135 17291
rect 6761 17213 7135 17265
tri 7135 17213 7213 17291 sw
tri 7233 17213 7311 17291 ne
rect 7311 17265 7365 17291
rect 7485 17291 7587 17385
tri 7587 17291 7685 17389 sw
tri 7685 17291 7783 17389 ne
rect 7783 17385 8137 17389
rect 7783 17291 7915 17385
rect 7485 17265 7685 17291
rect 7311 17213 7685 17265
tri 7685 17213 7763 17291 sw
tri 7783 17213 7861 17291 ne
rect 7861 17265 7915 17291
rect 8035 17291 8137 17385
tri 8137 17291 8235 17389 sw
tri 8235 17291 8333 17389 ne
rect 8333 17385 8687 17389
rect 8333 17291 8465 17385
rect 8035 17265 8235 17291
rect 7861 17213 8235 17265
tri 8235 17213 8313 17291 sw
tri 8333 17213 8411 17291 ne
rect 8411 17265 8465 17291
rect 8585 17291 8687 17385
tri 8687 17291 8785 17389 sw
tri 8785 17291 8883 17389 ne
rect 8883 17385 9237 17389
rect 8883 17291 9015 17385
rect 8585 17265 8785 17291
rect 8411 17213 8785 17265
tri 8785 17213 8863 17291 sw
tri 8883 17213 8961 17291 ne
rect 8961 17265 9015 17291
rect 9135 17291 9237 17385
tri 9237 17291 9335 17389 sw
tri 9335 17291 9433 17389 ne
rect 9433 17385 9787 17389
rect 9433 17291 9565 17385
rect 9135 17265 9335 17291
rect 8961 17213 9335 17265
tri 9335 17213 9413 17291 sw
tri 9433 17213 9511 17291 ne
rect 9511 17265 9565 17291
rect 9685 17291 9787 17385
tri 9787 17291 9885 17389 sw
tri 9885 17291 9983 17389 ne
rect 9983 17385 10337 17389
rect 9983 17291 10115 17385
rect 9685 17265 9885 17291
rect 9511 17213 9885 17265
tri 9885 17213 9963 17291 sw
tri 9983 17213 10061 17291 ne
rect 10061 17265 10115 17291
rect 10235 17291 10337 17385
tri 10337 17291 10435 17389 sw
tri 10435 17291 10533 17389 ne
rect 10533 17385 10887 17389
rect 10533 17291 10665 17385
rect 10235 17265 10435 17291
rect 10061 17213 10435 17265
tri 10435 17213 10513 17291 sw
tri 10533 17213 10611 17291 ne
rect 10611 17265 10665 17291
rect 10785 17291 10887 17385
tri 10887 17291 10985 17389 sw
tri 10985 17291 11083 17389 ne
rect 11083 17385 11437 17389
rect 11083 17291 11215 17385
rect 10785 17265 10985 17291
rect 10611 17213 10985 17265
tri 10985 17213 11063 17291 sw
tri 11083 17213 11161 17291 ne
rect 11161 17265 11215 17291
rect 11335 17291 11437 17385
tri 11437 17291 11535 17389 sw
tri 11535 17291 11633 17389 ne
rect 11633 17385 11987 17389
rect 11633 17291 11765 17385
rect 11335 17265 11535 17291
rect 11161 17213 11535 17265
tri 11535 17213 11613 17291 sw
tri 11633 17213 11711 17291 ne
rect 11711 17265 11765 17291
rect 11885 17291 11987 17385
tri 11987 17291 12085 17389 sw
tri 12085 17291 12183 17389 ne
rect 12183 17385 12537 17389
rect 12183 17291 12315 17385
rect 11885 17265 12085 17291
rect 11711 17213 12085 17265
tri 12085 17213 12163 17291 sw
tri 12183 17213 12261 17291 ne
rect 12261 17265 12315 17291
rect 12435 17291 12537 17385
tri 12537 17291 12635 17389 sw
tri 12635 17291 12733 17389 ne
rect 12733 17385 13087 17389
rect 12733 17291 12865 17385
rect 12435 17265 12635 17291
rect 12261 17213 12635 17265
tri 12635 17213 12713 17291 sw
tri 12733 17213 12811 17291 ne
rect 12811 17265 12865 17291
rect 12985 17291 13087 17385
tri 13087 17291 13185 17389 sw
tri 13185 17291 13283 17389 ne
rect 13283 17385 13637 17389
rect 13283 17291 13415 17385
rect 12985 17265 13185 17291
rect 12811 17213 13185 17265
tri 13185 17213 13263 17291 sw
tri 13283 17213 13361 17291 ne
rect 13361 17265 13415 17291
rect 13535 17291 13637 17385
tri 13637 17291 13735 17389 sw
tri 13735 17291 13833 17389 ne
rect 13833 17385 14187 17389
rect 13833 17291 13965 17385
rect 13535 17265 13735 17291
rect 13361 17213 13735 17265
tri 13735 17213 13813 17291 sw
tri 13833 17213 13911 17291 ne
rect 13911 17265 13965 17291
rect 14085 17291 14187 17385
tri 14187 17291 14285 17389 sw
tri 14285 17291 14383 17389 ne
rect 14383 17385 14737 17389
rect 14383 17291 14515 17385
rect 14085 17265 14285 17291
rect 13911 17213 14285 17265
tri 14285 17213 14363 17291 sw
tri 14383 17213 14461 17291 ne
rect 14461 17265 14515 17291
rect 14635 17291 14737 17385
tri 14737 17291 14835 17389 sw
tri 14835 17291 14933 17389 ne
rect 14933 17385 15287 17389
rect 14933 17291 15065 17385
rect 14635 17265 14835 17291
rect 14461 17213 14835 17265
tri 14835 17213 14913 17291 sw
tri 14933 17213 15011 17291 ne
rect 15011 17265 15065 17291
rect 15185 17291 15287 17385
tri 15287 17291 15385 17389 sw
tri 15385 17291 15483 17389 ne
rect 15483 17385 15837 17389
rect 15483 17291 15615 17385
rect 15185 17265 15385 17291
rect 15011 17213 15385 17265
tri 15385 17213 15463 17291 sw
tri 15483 17213 15561 17291 ne
rect 15561 17265 15615 17291
rect 15735 17291 15837 17385
tri 15837 17291 15935 17389 sw
tri 15935 17291 16033 17389 ne
rect 16033 17385 16387 17389
rect 16033 17291 16165 17385
rect 15735 17265 15935 17291
rect 15561 17213 15935 17265
tri 15935 17213 16013 17291 sw
tri 16033 17213 16111 17291 ne
rect 16111 17265 16165 17291
rect 16285 17291 16387 17385
tri 16387 17291 16485 17389 sw
tri 16485 17291 16583 17389 ne
rect 16583 17385 16937 17389
rect 16583 17291 16715 17385
rect 16285 17265 16485 17291
rect 16111 17213 16485 17265
tri 16485 17213 16563 17291 sw
tri 16583 17213 16661 17291 ne
rect 16661 17265 16715 17291
rect 16835 17291 16937 17385
tri 16937 17291 17035 17389 sw
tri 17035 17291 17133 17389 ne
rect 17133 17385 17487 17389
rect 17133 17291 17265 17385
rect 16835 17265 17035 17291
rect 16661 17213 17035 17265
tri 17035 17213 17113 17291 sw
tri 17133 17213 17211 17291 ne
rect 17211 17265 17265 17291
rect 17385 17291 17487 17385
tri 17487 17291 17585 17389 sw
tri 17585 17291 17683 17389 ne
rect 17683 17385 18037 17389
rect 17683 17291 17815 17385
rect 17385 17265 17585 17291
rect 17211 17213 17585 17265
tri 17585 17213 17663 17291 sw
tri 17683 17213 17761 17291 ne
rect 17761 17265 17815 17291
rect 17935 17291 18037 17385
tri 18037 17291 18135 17389 sw
tri 18135 17291 18233 17389 ne
rect 18233 17385 18587 17389
rect 18233 17291 18365 17385
rect 17935 17265 18135 17291
rect 17761 17213 18135 17265
tri 18135 17213 18213 17291 sw
tri 18233 17213 18311 17291 ne
rect 18311 17265 18365 17291
rect 18485 17291 18587 17385
tri 18587 17291 18685 17389 sw
tri 18685 17291 18783 17389 ne
rect 18783 17385 19137 17389
rect 18783 17291 18915 17385
rect 18485 17265 18685 17291
rect 18311 17213 18685 17265
tri 18685 17213 18763 17291 sw
tri 18783 17213 18861 17291 ne
rect 18861 17265 18915 17291
rect 19035 17291 19137 17385
tri 19137 17291 19235 17389 sw
tri 19235 17291 19333 17389 ne
rect 19333 17385 21800 17389
rect 19333 17291 19465 17385
rect 19035 17265 19235 17291
rect 18861 17213 19235 17265
tri 19235 17213 19313 17291 sw
tri 19333 17213 19411 17291 ne
rect 19411 17265 19465 17291
rect 19585 17265 21800 17385
rect 19411 17213 21800 17265
rect 211 17163 613 17213
rect -500 17113 113 17163
tri 113 17113 163 17163 sw
tri 211 17113 261 17163 ne
rect 261 17133 613 17163
tri 613 17133 693 17213 sw
tri 711 17133 791 17213 ne
rect 791 17133 1163 17213
tri 1163 17133 1243 17213 sw
tri 1261 17133 1341 17213 ne
rect 1341 17133 1713 17213
tri 1713 17133 1793 17213 sw
tri 1811 17133 1891 17213 ne
rect 1891 17133 2263 17213
tri 2263 17133 2343 17213 sw
tri 2361 17133 2441 17213 ne
rect 2441 17133 2813 17213
tri 2813 17133 2893 17213 sw
tri 2911 17133 2991 17213 ne
rect 2991 17133 3363 17213
tri 3363 17133 3443 17213 sw
tri 3461 17133 3541 17213 ne
rect 3541 17133 3913 17213
tri 3913 17133 3993 17213 sw
tri 4011 17133 4091 17213 ne
rect 4091 17133 4463 17213
tri 4463 17133 4543 17213 sw
tri 4561 17133 4641 17213 ne
rect 4641 17133 5013 17213
tri 5013 17133 5093 17213 sw
tri 5111 17133 5191 17213 ne
rect 5191 17133 5563 17213
tri 5563 17133 5643 17213 sw
tri 5661 17133 5741 17213 ne
rect 5741 17133 6113 17213
tri 6113 17133 6193 17213 sw
tri 6211 17133 6291 17213 ne
rect 6291 17133 6663 17213
tri 6663 17133 6743 17213 sw
tri 6761 17133 6841 17213 ne
rect 6841 17133 7213 17213
tri 7213 17133 7293 17213 sw
tri 7311 17133 7391 17213 ne
rect 7391 17133 7763 17213
tri 7763 17133 7843 17213 sw
tri 7861 17133 7941 17213 ne
rect 7941 17133 8313 17213
tri 8313 17133 8393 17213 sw
tri 8411 17133 8491 17213 ne
rect 8491 17133 8863 17213
tri 8863 17133 8943 17213 sw
tri 8961 17133 9041 17213 ne
rect 9041 17133 9413 17213
tri 9413 17133 9493 17213 sw
tri 9511 17133 9591 17213 ne
rect 9591 17133 9963 17213
tri 9963 17133 10043 17213 sw
tri 10061 17133 10141 17213 ne
rect 10141 17133 10513 17213
tri 10513 17133 10593 17213 sw
tri 10611 17133 10691 17213 ne
rect 10691 17133 11063 17213
tri 11063 17133 11143 17213 sw
tri 11161 17133 11241 17213 ne
rect 11241 17133 11613 17213
tri 11613 17133 11693 17213 sw
tri 11711 17133 11791 17213 ne
rect 11791 17133 12163 17213
tri 12163 17133 12243 17213 sw
tri 12261 17133 12341 17213 ne
rect 12341 17133 12713 17213
tri 12713 17133 12793 17213 sw
tri 12811 17133 12891 17213 ne
rect 12891 17133 13263 17213
tri 13263 17133 13343 17213 sw
tri 13361 17133 13441 17213 ne
rect 13441 17133 13813 17213
tri 13813 17133 13893 17213 sw
tri 13911 17133 13991 17213 ne
rect 13991 17133 14363 17213
tri 14363 17133 14443 17213 sw
tri 14461 17133 14541 17213 ne
rect 14541 17133 14913 17213
tri 14913 17133 14993 17213 sw
tri 15011 17133 15091 17213 ne
rect 15091 17133 15463 17213
tri 15463 17133 15543 17213 sw
tri 15561 17133 15641 17213 ne
rect 15641 17133 16013 17213
tri 16013 17133 16093 17213 sw
tri 16111 17133 16191 17213 ne
rect 16191 17133 16563 17213
tri 16563 17133 16643 17213 sw
tri 16661 17133 16741 17213 ne
rect 16741 17133 17113 17213
tri 17113 17133 17193 17213 sw
tri 17211 17133 17291 17213 ne
rect 17291 17133 17663 17213
tri 17663 17133 17743 17213 sw
tri 17761 17133 17841 17213 ne
rect 17841 17133 18213 17213
tri 18213 17133 18293 17213 sw
tri 18311 17133 18391 17213 ne
rect 18391 17133 18763 17213
tri 18763 17133 18843 17213 sw
tri 18861 17133 18941 17213 ne
rect 18941 17133 19313 17213
tri 19313 17133 19393 17213 sw
tri 19411 17133 19491 17213 ne
rect 19491 17133 20100 17213
rect 261 17113 693 17133
rect -500 17035 163 17113
tri 163 17035 241 17113 sw
tri 261 17035 339 17113 ne
rect 339 17035 693 17113
tri 693 17035 791 17133 sw
tri 791 17035 889 17133 ne
rect 889 17035 1243 17133
tri 1243 17035 1341 17133 sw
tri 1341 17035 1439 17133 ne
rect 1439 17035 1793 17133
tri 1793 17035 1891 17133 sw
tri 1891 17035 1989 17133 ne
rect 1989 17035 2343 17133
tri 2343 17035 2441 17133 sw
tri 2441 17035 2539 17133 ne
rect 2539 17035 2893 17133
tri 2893 17035 2991 17133 sw
tri 2991 17035 3089 17133 ne
rect 3089 17035 3443 17133
tri 3443 17035 3541 17133 sw
tri 3541 17035 3639 17133 ne
rect 3639 17035 3993 17133
tri 3993 17035 4091 17133 sw
tri 4091 17035 4189 17133 ne
rect 4189 17035 4543 17133
tri 4543 17035 4641 17133 sw
tri 4641 17035 4739 17133 ne
rect 4739 17035 5093 17133
tri 5093 17035 5191 17133 sw
tri 5191 17035 5289 17133 ne
rect 5289 17035 5643 17133
tri 5643 17035 5741 17133 sw
tri 5741 17035 5839 17133 ne
rect 5839 17035 6193 17133
tri 6193 17035 6291 17133 sw
tri 6291 17035 6389 17133 ne
rect 6389 17035 6743 17133
tri 6743 17035 6841 17133 sw
tri 6841 17035 6939 17133 ne
rect 6939 17035 7293 17133
tri 7293 17035 7391 17133 sw
tri 7391 17035 7489 17133 ne
rect 7489 17035 7843 17133
tri 7843 17035 7941 17133 sw
tri 7941 17035 8039 17133 ne
rect 8039 17035 8393 17133
tri 8393 17035 8491 17133 sw
tri 8491 17035 8589 17133 ne
rect 8589 17035 8943 17133
tri 8943 17035 9041 17133 sw
tri 9041 17035 9139 17133 ne
rect 9139 17035 9493 17133
tri 9493 17035 9591 17133 sw
tri 9591 17035 9689 17133 ne
rect 9689 17035 10043 17133
tri 10043 17035 10141 17133 sw
tri 10141 17035 10239 17133 ne
rect 10239 17035 10593 17133
tri 10593 17035 10691 17133 sw
tri 10691 17035 10789 17133 ne
rect 10789 17035 11143 17133
tri 11143 17035 11241 17133 sw
tri 11241 17035 11339 17133 ne
rect 11339 17035 11693 17133
tri 11693 17035 11791 17133 sw
tri 11791 17035 11889 17133 ne
rect 11889 17035 12243 17133
tri 12243 17035 12341 17133 sw
tri 12341 17035 12439 17133 ne
rect 12439 17035 12793 17133
tri 12793 17035 12891 17133 sw
tri 12891 17035 12989 17133 ne
rect 12989 17035 13343 17133
tri 13343 17035 13441 17133 sw
tri 13441 17035 13539 17133 ne
rect 13539 17035 13893 17133
tri 13893 17035 13991 17133 sw
tri 13991 17035 14089 17133 ne
rect 14089 17035 14443 17133
tri 14443 17035 14541 17133 sw
tri 14541 17035 14639 17133 ne
rect 14639 17035 14993 17133
tri 14993 17035 15091 17133 sw
tri 15091 17035 15189 17133 ne
rect 15189 17035 15543 17133
tri 15543 17035 15641 17133 sw
tri 15641 17035 15739 17133 ne
rect 15739 17035 16093 17133
tri 16093 17035 16191 17133 sw
tri 16191 17035 16289 17133 ne
rect 16289 17035 16643 17133
tri 16643 17035 16741 17133 sw
tri 16741 17035 16839 17133 ne
rect 16839 17035 17193 17133
tri 17193 17035 17291 17133 sw
tri 17291 17035 17389 17133 ne
rect 17389 17035 17743 17133
tri 17743 17035 17841 17133 sw
tri 17841 17035 17939 17133 ne
rect 17939 17035 18293 17133
tri 18293 17035 18391 17133 sw
tri 18391 17035 18489 17133 ne
rect 18489 17035 18843 17133
tri 18843 17035 18941 17133 sw
tri 18941 17035 19039 17133 ne
rect 19039 17035 19393 17133
tri 19393 17035 19491 17133 sw
tri 19491 17035 19589 17133 ne
rect 19589 17113 20100 17133
rect 20200 17113 21800 17213
rect 19589 17035 21800 17113
rect -500 16987 241 17035
rect -500 16887 -400 16987
rect -300 16937 241 16987
tri 241 16937 339 17035 sw
tri 339 16937 437 17035 ne
rect 437 16937 791 17035
tri 791 16937 889 17035 sw
tri 889 16937 987 17035 ne
rect 987 16937 1341 17035
tri 1341 16937 1439 17035 sw
tri 1439 16937 1537 17035 ne
rect 1537 16937 1891 17035
tri 1891 16937 1989 17035 sw
tri 1989 16937 2087 17035 ne
rect 2087 16937 2441 17035
tri 2441 16937 2539 17035 sw
tri 2539 16937 2637 17035 ne
rect 2637 16937 2991 17035
tri 2991 16937 3089 17035 sw
tri 3089 16937 3187 17035 ne
rect 3187 16937 3541 17035
tri 3541 16937 3639 17035 sw
tri 3639 16937 3737 17035 ne
rect 3737 16937 4091 17035
tri 4091 16937 4189 17035 sw
tri 4189 16937 4287 17035 ne
rect 4287 16937 4641 17035
tri 4641 16937 4739 17035 sw
tri 4739 16937 4837 17035 ne
rect 4837 16937 5191 17035
tri 5191 16937 5289 17035 sw
tri 5289 16937 5387 17035 ne
rect 5387 16937 5741 17035
tri 5741 16937 5839 17035 sw
tri 5839 16937 5937 17035 ne
rect 5937 16937 6291 17035
tri 6291 16937 6389 17035 sw
tri 6389 16937 6487 17035 ne
rect 6487 16937 6841 17035
tri 6841 16937 6939 17035 sw
tri 6939 16937 7037 17035 ne
rect 7037 16937 7391 17035
tri 7391 16937 7489 17035 sw
tri 7489 16937 7587 17035 ne
rect 7587 16937 7941 17035
tri 7941 16937 8039 17035 sw
tri 8039 16937 8137 17035 ne
rect 8137 16937 8491 17035
tri 8491 16937 8589 17035 sw
tri 8589 16937 8687 17035 ne
rect 8687 16937 9041 17035
tri 9041 16937 9139 17035 sw
tri 9139 16937 9237 17035 ne
rect 9237 16937 9591 17035
tri 9591 16937 9689 17035 sw
tri 9689 16937 9787 17035 ne
rect 9787 16937 10141 17035
tri 10141 16937 10239 17035 sw
tri 10239 16937 10337 17035 ne
rect 10337 16937 10691 17035
tri 10691 16937 10789 17035 sw
tri 10789 16937 10887 17035 ne
rect 10887 16937 11241 17035
tri 11241 16937 11339 17035 sw
tri 11339 16937 11437 17035 ne
rect 11437 16937 11791 17035
tri 11791 16937 11889 17035 sw
tri 11889 16937 11987 17035 ne
rect 11987 16937 12341 17035
tri 12341 16937 12439 17035 sw
tri 12439 16937 12537 17035 ne
rect 12537 16937 12891 17035
tri 12891 16937 12989 17035 sw
tri 12989 16937 13087 17035 ne
rect 13087 16937 13441 17035
tri 13441 16937 13539 17035 sw
tri 13539 16937 13637 17035 ne
rect 13637 16937 13991 17035
tri 13991 16937 14089 17035 sw
tri 14089 16937 14187 17035 ne
rect 14187 16937 14541 17035
tri 14541 16937 14639 17035 sw
tri 14639 16937 14737 17035 ne
rect 14737 16937 15091 17035
tri 15091 16937 15189 17035 sw
tri 15189 16937 15287 17035 ne
rect 15287 16937 15641 17035
tri 15641 16937 15739 17035 sw
tri 15739 16937 15837 17035 ne
rect 15837 16937 16191 17035
tri 16191 16937 16289 17035 sw
tri 16289 16937 16387 17035 ne
rect 16387 16937 16741 17035
tri 16741 16937 16839 17035 sw
tri 16839 16937 16937 17035 ne
rect 16937 16937 17291 17035
tri 17291 16937 17389 17035 sw
tri 17389 16937 17487 17035 ne
rect 17487 16937 17841 17035
tri 17841 16937 17939 17035 sw
tri 17939 16937 18037 17035 ne
rect 18037 16937 18391 17035
tri 18391 16937 18489 17035 sw
tri 18489 16937 18587 17035 ne
rect 18587 16937 18941 17035
tri 18941 16937 19039 17035 sw
tri 19039 16937 19137 17035 ne
rect 19137 16937 19491 17035
tri 19491 16937 19589 17035 sw
tri 19589 16937 19687 17035 ne
rect 19687 16937 21800 17035
rect -300 16887 339 16937
rect -500 16839 339 16887
tri 339 16839 437 16937 sw
tri 437 16839 535 16937 ne
rect 535 16839 889 16937
tri 889 16839 987 16937 sw
tri 987 16839 1085 16937 ne
rect 1085 16839 1439 16937
tri 1439 16839 1537 16937 sw
tri 1537 16839 1635 16937 ne
rect 1635 16839 1989 16937
tri 1989 16839 2087 16937 sw
tri 2087 16839 2185 16937 ne
rect 2185 16839 2539 16937
tri 2539 16839 2637 16937 sw
tri 2637 16839 2735 16937 ne
rect 2735 16839 3089 16937
tri 3089 16839 3187 16937 sw
tri 3187 16839 3285 16937 ne
rect 3285 16839 3639 16937
tri 3639 16839 3737 16937 sw
tri 3737 16839 3835 16937 ne
rect 3835 16839 4189 16937
tri 4189 16839 4287 16937 sw
tri 4287 16839 4385 16937 ne
rect 4385 16839 4739 16937
tri 4739 16839 4837 16937 sw
tri 4837 16839 4935 16937 ne
rect 4935 16839 5289 16937
tri 5289 16839 5387 16937 sw
tri 5387 16839 5485 16937 ne
rect 5485 16839 5839 16937
tri 5839 16839 5937 16937 sw
tri 5937 16839 6035 16937 ne
rect 6035 16839 6389 16937
tri 6389 16839 6487 16937 sw
tri 6487 16839 6585 16937 ne
rect 6585 16839 6939 16937
tri 6939 16839 7037 16937 sw
tri 7037 16839 7135 16937 ne
rect 7135 16839 7489 16937
tri 7489 16839 7587 16937 sw
tri 7587 16839 7685 16937 ne
rect 7685 16839 8039 16937
tri 8039 16839 8137 16937 sw
tri 8137 16839 8235 16937 ne
rect 8235 16839 8589 16937
tri 8589 16839 8687 16937 sw
tri 8687 16839 8785 16937 ne
rect 8785 16839 9139 16937
tri 9139 16839 9237 16937 sw
tri 9237 16839 9335 16937 ne
rect 9335 16839 9689 16937
tri 9689 16839 9787 16937 sw
tri 9787 16839 9885 16937 ne
rect 9885 16839 10239 16937
tri 10239 16839 10337 16937 sw
tri 10337 16839 10435 16937 ne
rect 10435 16839 10789 16937
tri 10789 16839 10887 16937 sw
tri 10887 16839 10985 16937 ne
rect 10985 16839 11339 16937
tri 11339 16839 11437 16937 sw
tri 11437 16839 11535 16937 ne
rect 11535 16839 11889 16937
tri 11889 16839 11987 16937 sw
tri 11987 16839 12085 16937 ne
rect 12085 16839 12439 16937
tri 12439 16839 12537 16937 sw
tri 12537 16839 12635 16937 ne
rect 12635 16839 12989 16937
tri 12989 16839 13087 16937 sw
tri 13087 16839 13185 16937 ne
rect 13185 16839 13539 16937
tri 13539 16839 13637 16937 sw
tri 13637 16839 13735 16937 ne
rect 13735 16839 14089 16937
tri 14089 16839 14187 16937 sw
tri 14187 16839 14285 16937 ne
rect 14285 16839 14639 16937
tri 14639 16839 14737 16937 sw
tri 14737 16839 14835 16937 ne
rect 14835 16839 15189 16937
tri 15189 16839 15287 16937 sw
tri 15287 16839 15385 16937 ne
rect 15385 16839 15739 16937
tri 15739 16839 15837 16937 sw
tri 15837 16839 15935 16937 ne
rect 15935 16839 16289 16937
tri 16289 16839 16387 16937 sw
tri 16387 16839 16485 16937 ne
rect 16485 16839 16839 16937
tri 16839 16839 16937 16937 sw
tri 16937 16839 17035 16937 ne
rect 17035 16839 17389 16937
tri 17389 16839 17487 16937 sw
tri 17487 16839 17585 16937 ne
rect 17585 16839 17939 16937
tri 17939 16839 18037 16937 sw
tri 18037 16839 18135 16937 ne
rect 18135 16839 18489 16937
tri 18489 16839 18587 16937 sw
tri 18587 16839 18685 16937 ne
rect 18685 16839 19039 16937
tri 19039 16839 19137 16937 sw
tri 19137 16839 19235 16937 ne
rect 19235 16839 19589 16937
tri 19589 16839 19687 16937 sw
rect -500 16835 437 16839
rect -500 16715 215 16835
rect 335 16741 437 16835
tri 437 16741 535 16839 sw
tri 535 16741 633 16839 ne
rect 633 16835 987 16839
rect 633 16741 765 16835
rect 335 16715 535 16741
rect -500 16711 535 16715
tri 535 16711 565 16741 sw
tri 633 16711 663 16741 ne
rect 663 16715 765 16741
rect 885 16741 987 16835
tri 987 16741 1085 16839 sw
tri 1085 16741 1183 16839 ne
rect 1183 16835 1537 16839
rect 1183 16741 1315 16835
rect 885 16715 1085 16741
rect 663 16711 1085 16715
tri 1085 16711 1115 16741 sw
tri 1183 16711 1213 16741 ne
rect 1213 16715 1315 16741
rect 1435 16741 1537 16835
tri 1537 16741 1635 16839 sw
tri 1635 16741 1733 16839 ne
rect 1733 16835 2087 16839
rect 1733 16741 1865 16835
rect 1435 16715 1635 16741
rect 1213 16711 1635 16715
tri 1635 16711 1665 16741 sw
tri 1733 16711 1763 16741 ne
rect 1763 16715 1865 16741
rect 1985 16741 2087 16835
tri 2087 16741 2185 16839 sw
tri 2185 16741 2283 16839 ne
rect 2283 16835 2637 16839
rect 2283 16741 2415 16835
rect 1985 16715 2185 16741
rect 1763 16711 2185 16715
tri 2185 16711 2215 16741 sw
tri 2283 16711 2313 16741 ne
rect 2313 16715 2415 16741
rect 2535 16741 2637 16835
tri 2637 16741 2735 16839 sw
tri 2735 16741 2833 16839 ne
rect 2833 16835 3187 16839
rect 2833 16741 2965 16835
rect 2535 16715 2735 16741
rect 2313 16711 2735 16715
tri 2735 16711 2765 16741 sw
tri 2833 16711 2863 16741 ne
rect 2863 16715 2965 16741
rect 3085 16741 3187 16835
tri 3187 16741 3285 16839 sw
tri 3285 16741 3383 16839 ne
rect 3383 16835 3737 16839
rect 3383 16741 3515 16835
rect 3085 16715 3285 16741
rect 2863 16711 3285 16715
tri 3285 16711 3315 16741 sw
tri 3383 16711 3413 16741 ne
rect 3413 16715 3515 16741
rect 3635 16741 3737 16835
tri 3737 16741 3835 16839 sw
tri 3835 16741 3933 16839 ne
rect 3933 16835 4287 16839
rect 3933 16741 4065 16835
rect 3635 16715 3835 16741
rect 3413 16711 3835 16715
tri 3835 16711 3865 16741 sw
tri 3933 16711 3963 16741 ne
rect 3963 16715 4065 16741
rect 4185 16741 4287 16835
tri 4287 16741 4385 16839 sw
tri 4385 16741 4483 16839 ne
rect 4483 16835 4837 16839
rect 4483 16741 4615 16835
rect 4185 16715 4385 16741
rect 3963 16711 4385 16715
tri 4385 16711 4415 16741 sw
tri 4483 16711 4513 16741 ne
rect 4513 16715 4615 16741
rect 4735 16741 4837 16835
tri 4837 16741 4935 16839 sw
tri 4935 16741 5033 16839 ne
rect 5033 16835 5387 16839
rect 5033 16741 5165 16835
rect 4735 16715 4935 16741
rect 4513 16711 4935 16715
tri 4935 16711 4965 16741 sw
tri 5033 16711 5063 16741 ne
rect 5063 16715 5165 16741
rect 5285 16741 5387 16835
tri 5387 16741 5485 16839 sw
tri 5485 16741 5583 16839 ne
rect 5583 16835 5937 16839
rect 5583 16741 5715 16835
rect 5285 16715 5485 16741
rect 5063 16711 5485 16715
tri 5485 16711 5515 16741 sw
tri 5583 16711 5613 16741 ne
rect 5613 16715 5715 16741
rect 5835 16741 5937 16835
tri 5937 16741 6035 16839 sw
tri 6035 16741 6133 16839 ne
rect 6133 16835 6487 16839
rect 6133 16741 6265 16835
rect 5835 16715 6035 16741
rect 5613 16711 6035 16715
tri 6035 16711 6065 16741 sw
tri 6133 16711 6163 16741 ne
rect 6163 16715 6265 16741
rect 6385 16741 6487 16835
tri 6487 16741 6585 16839 sw
tri 6585 16741 6683 16839 ne
rect 6683 16835 7037 16839
rect 6683 16741 6815 16835
rect 6385 16715 6585 16741
rect 6163 16711 6585 16715
tri 6585 16711 6615 16741 sw
tri 6683 16711 6713 16741 ne
rect 6713 16715 6815 16741
rect 6935 16741 7037 16835
tri 7037 16741 7135 16839 sw
tri 7135 16741 7233 16839 ne
rect 7233 16835 7587 16839
rect 7233 16741 7365 16835
rect 6935 16715 7135 16741
rect 6713 16711 7135 16715
tri 7135 16711 7165 16741 sw
tri 7233 16711 7263 16741 ne
rect 7263 16715 7365 16741
rect 7485 16741 7587 16835
tri 7587 16741 7685 16839 sw
tri 7685 16741 7783 16839 ne
rect 7783 16835 8137 16839
rect 7783 16741 7915 16835
rect 7485 16715 7685 16741
rect 7263 16711 7685 16715
tri 7685 16711 7715 16741 sw
tri 7783 16711 7813 16741 ne
rect 7813 16715 7915 16741
rect 8035 16741 8137 16835
tri 8137 16741 8235 16839 sw
tri 8235 16741 8333 16839 ne
rect 8333 16835 8687 16839
rect 8333 16741 8465 16835
rect 8035 16715 8235 16741
rect 7813 16711 8235 16715
tri 8235 16711 8265 16741 sw
tri 8333 16711 8363 16741 ne
rect 8363 16715 8465 16741
rect 8585 16741 8687 16835
tri 8687 16741 8785 16839 sw
tri 8785 16741 8883 16839 ne
rect 8883 16835 9237 16839
rect 8883 16741 9015 16835
rect 8585 16715 8785 16741
rect 8363 16711 8785 16715
tri 8785 16711 8815 16741 sw
tri 8883 16711 8913 16741 ne
rect 8913 16715 9015 16741
rect 9135 16741 9237 16835
tri 9237 16741 9335 16839 sw
tri 9335 16741 9433 16839 ne
rect 9433 16835 9787 16839
rect 9433 16741 9565 16835
rect 9135 16715 9335 16741
rect 8913 16711 9335 16715
tri 9335 16711 9365 16741 sw
tri 9433 16711 9463 16741 ne
rect 9463 16715 9565 16741
rect 9685 16741 9787 16835
tri 9787 16741 9885 16839 sw
tri 9885 16741 9983 16839 ne
rect 9983 16835 10337 16839
rect 9983 16741 10115 16835
rect 9685 16715 9885 16741
rect 9463 16711 9885 16715
tri 9885 16711 9915 16741 sw
tri 9983 16711 10013 16741 ne
rect 10013 16715 10115 16741
rect 10235 16741 10337 16835
tri 10337 16741 10435 16839 sw
tri 10435 16741 10533 16839 ne
rect 10533 16835 10887 16839
rect 10533 16741 10665 16835
rect 10235 16715 10435 16741
rect 10013 16711 10435 16715
tri 10435 16711 10465 16741 sw
tri 10533 16711 10563 16741 ne
rect 10563 16715 10665 16741
rect 10785 16741 10887 16835
tri 10887 16741 10985 16839 sw
tri 10985 16741 11083 16839 ne
rect 11083 16835 11437 16839
rect 11083 16741 11215 16835
rect 10785 16715 10985 16741
rect 10563 16711 10985 16715
tri 10985 16711 11015 16741 sw
tri 11083 16711 11113 16741 ne
rect 11113 16715 11215 16741
rect 11335 16741 11437 16835
tri 11437 16741 11535 16839 sw
tri 11535 16741 11633 16839 ne
rect 11633 16835 11987 16839
rect 11633 16741 11765 16835
rect 11335 16715 11535 16741
rect 11113 16711 11535 16715
tri 11535 16711 11565 16741 sw
tri 11633 16711 11663 16741 ne
rect 11663 16715 11765 16741
rect 11885 16741 11987 16835
tri 11987 16741 12085 16839 sw
tri 12085 16741 12183 16839 ne
rect 12183 16835 12537 16839
rect 12183 16741 12315 16835
rect 11885 16715 12085 16741
rect 11663 16711 12085 16715
tri 12085 16711 12115 16741 sw
tri 12183 16711 12213 16741 ne
rect 12213 16715 12315 16741
rect 12435 16741 12537 16835
tri 12537 16741 12635 16839 sw
tri 12635 16741 12733 16839 ne
rect 12733 16835 13087 16839
rect 12733 16741 12865 16835
rect 12435 16715 12635 16741
rect 12213 16711 12635 16715
tri 12635 16711 12665 16741 sw
tri 12733 16711 12763 16741 ne
rect 12763 16715 12865 16741
rect 12985 16741 13087 16835
tri 13087 16741 13185 16839 sw
tri 13185 16741 13283 16839 ne
rect 13283 16835 13637 16839
rect 13283 16741 13415 16835
rect 12985 16715 13185 16741
rect 12763 16711 13185 16715
tri 13185 16711 13215 16741 sw
tri 13283 16711 13313 16741 ne
rect 13313 16715 13415 16741
rect 13535 16741 13637 16835
tri 13637 16741 13735 16839 sw
tri 13735 16741 13833 16839 ne
rect 13833 16835 14187 16839
rect 13833 16741 13965 16835
rect 13535 16715 13735 16741
rect 13313 16711 13735 16715
tri 13735 16711 13765 16741 sw
tri 13833 16711 13863 16741 ne
rect 13863 16715 13965 16741
rect 14085 16741 14187 16835
tri 14187 16741 14285 16839 sw
tri 14285 16741 14383 16839 ne
rect 14383 16835 14737 16839
rect 14383 16741 14515 16835
rect 14085 16715 14285 16741
rect 13863 16711 14285 16715
tri 14285 16711 14315 16741 sw
tri 14383 16711 14413 16741 ne
rect 14413 16715 14515 16741
rect 14635 16741 14737 16835
tri 14737 16741 14835 16839 sw
tri 14835 16741 14933 16839 ne
rect 14933 16835 15287 16839
rect 14933 16741 15065 16835
rect 14635 16715 14835 16741
rect 14413 16711 14835 16715
tri 14835 16711 14865 16741 sw
tri 14933 16711 14963 16741 ne
rect 14963 16715 15065 16741
rect 15185 16741 15287 16835
tri 15287 16741 15385 16839 sw
tri 15385 16741 15483 16839 ne
rect 15483 16835 15837 16839
rect 15483 16741 15615 16835
rect 15185 16715 15385 16741
rect 14963 16711 15385 16715
tri 15385 16711 15415 16741 sw
tri 15483 16711 15513 16741 ne
rect 15513 16715 15615 16741
rect 15735 16741 15837 16835
tri 15837 16741 15935 16839 sw
tri 15935 16741 16033 16839 ne
rect 16033 16835 16387 16839
rect 16033 16741 16165 16835
rect 15735 16715 15935 16741
rect 15513 16711 15935 16715
tri 15935 16711 15965 16741 sw
tri 16033 16711 16063 16741 ne
rect 16063 16715 16165 16741
rect 16285 16741 16387 16835
tri 16387 16741 16485 16839 sw
tri 16485 16741 16583 16839 ne
rect 16583 16835 16937 16839
rect 16583 16741 16715 16835
rect 16285 16715 16485 16741
rect 16063 16711 16485 16715
tri 16485 16711 16515 16741 sw
tri 16583 16711 16613 16741 ne
rect 16613 16715 16715 16741
rect 16835 16741 16937 16835
tri 16937 16741 17035 16839 sw
tri 17035 16741 17133 16839 ne
rect 17133 16835 17487 16839
rect 17133 16741 17265 16835
rect 16835 16715 17035 16741
rect 16613 16711 17035 16715
tri 17035 16711 17065 16741 sw
tri 17133 16711 17163 16741 ne
rect 17163 16715 17265 16741
rect 17385 16741 17487 16835
tri 17487 16741 17585 16839 sw
tri 17585 16741 17683 16839 ne
rect 17683 16835 18037 16839
rect 17683 16741 17815 16835
rect 17385 16715 17585 16741
rect 17163 16711 17585 16715
tri 17585 16711 17615 16741 sw
tri 17683 16711 17713 16741 ne
rect 17713 16715 17815 16741
rect 17935 16741 18037 16835
tri 18037 16741 18135 16839 sw
tri 18135 16741 18233 16839 ne
rect 18233 16835 18587 16839
rect 18233 16741 18365 16835
rect 17935 16715 18135 16741
rect 17713 16711 18135 16715
tri 18135 16711 18165 16741 sw
tri 18233 16711 18263 16741 ne
rect 18263 16715 18365 16741
rect 18485 16741 18587 16835
tri 18587 16741 18685 16839 sw
tri 18685 16741 18783 16839 ne
rect 18783 16835 19137 16839
rect 18783 16741 18915 16835
rect 18485 16715 18685 16741
rect 18263 16711 18685 16715
tri 18685 16711 18715 16741 sw
tri 18783 16711 18813 16741 ne
rect 18813 16715 18915 16741
rect 19035 16741 19137 16835
tri 19137 16741 19235 16839 sw
tri 19235 16741 19333 16839 ne
rect 19333 16835 20300 16839
rect 19333 16741 19465 16835
rect 19035 16715 19235 16741
rect 18813 16711 19235 16715
tri 19235 16711 19265 16741 sw
tri 19333 16711 19363 16741 ne
rect 19363 16715 19465 16741
rect 19585 16715 20300 16835
rect 19363 16711 20300 16715
tri 113 16613 211 16711 ne
rect 211 16613 565 16711
tri 565 16613 663 16711 sw
tri 663 16613 761 16711 ne
rect 761 16613 1115 16711
tri 1115 16613 1213 16711 sw
tri 1213 16613 1311 16711 ne
rect 1311 16613 1665 16711
tri 1665 16613 1763 16711 sw
tri 1763 16613 1861 16711 ne
rect 1861 16613 2215 16711
tri 2215 16613 2313 16711 sw
tri 2313 16613 2411 16711 ne
rect 2411 16613 2765 16711
tri 2765 16613 2863 16711 sw
tri 2863 16613 2961 16711 ne
rect 2961 16613 3315 16711
tri 3315 16613 3413 16711 sw
tri 3413 16613 3511 16711 ne
rect 3511 16613 3865 16711
tri 3865 16613 3963 16711 sw
tri 3963 16613 4061 16711 ne
rect 4061 16613 4415 16711
tri 4415 16613 4513 16711 sw
tri 4513 16613 4611 16711 ne
rect 4611 16613 4965 16711
tri 4965 16613 5063 16711 sw
tri 5063 16613 5161 16711 ne
rect 5161 16613 5515 16711
tri 5515 16613 5613 16711 sw
tri 5613 16613 5711 16711 ne
rect 5711 16613 6065 16711
tri 6065 16613 6163 16711 sw
tri 6163 16613 6261 16711 ne
rect 6261 16613 6615 16711
tri 6615 16613 6713 16711 sw
tri 6713 16613 6811 16711 ne
rect 6811 16613 7165 16711
tri 7165 16613 7263 16711 sw
tri 7263 16613 7361 16711 ne
rect 7361 16613 7715 16711
tri 7715 16613 7813 16711 sw
tri 7813 16613 7911 16711 ne
rect 7911 16613 8265 16711
tri 8265 16613 8363 16711 sw
tri 8363 16613 8461 16711 ne
rect 8461 16613 8815 16711
tri 8815 16613 8913 16711 sw
tri 8913 16613 9011 16711 ne
rect 9011 16613 9365 16711
tri 9365 16613 9463 16711 sw
tri 9463 16613 9561 16711 ne
rect 9561 16613 9915 16711
tri 9915 16613 10013 16711 sw
tri 10013 16613 10111 16711 ne
rect 10111 16613 10465 16711
tri 10465 16613 10563 16711 sw
tri 10563 16613 10661 16711 ne
rect 10661 16613 11015 16711
tri 11015 16613 11113 16711 sw
tri 11113 16613 11211 16711 ne
rect 11211 16613 11565 16711
tri 11565 16613 11663 16711 sw
tri 11663 16613 11761 16711 ne
rect 11761 16613 12115 16711
tri 12115 16613 12213 16711 sw
tri 12213 16613 12311 16711 ne
rect 12311 16613 12665 16711
tri 12665 16613 12763 16711 sw
tri 12763 16613 12861 16711 ne
rect 12861 16613 13215 16711
tri 13215 16613 13313 16711 sw
tri 13313 16613 13411 16711 ne
rect 13411 16613 13765 16711
tri 13765 16613 13863 16711 sw
tri 13863 16613 13961 16711 ne
rect 13961 16613 14315 16711
tri 14315 16613 14413 16711 sw
tri 14413 16613 14511 16711 ne
rect 14511 16613 14865 16711
tri 14865 16613 14963 16711 sw
tri 14963 16613 15061 16711 ne
rect 15061 16613 15415 16711
tri 15415 16613 15513 16711 sw
tri 15513 16613 15611 16711 ne
rect 15611 16613 15965 16711
tri 15965 16613 16063 16711 sw
tri 16063 16613 16161 16711 ne
rect 16161 16613 16515 16711
tri 16515 16613 16613 16711 sw
tri 16613 16613 16711 16711 ne
rect 16711 16613 17065 16711
tri 17065 16613 17163 16711 sw
tri 17163 16613 17261 16711 ne
rect 17261 16613 17615 16711
tri 17615 16613 17713 16711 sw
tri 17713 16613 17811 16711 ne
rect 17811 16613 18165 16711
tri 18165 16613 18263 16711 sw
tri 18263 16613 18361 16711 ne
rect 18361 16613 18715 16711
tri 18715 16613 18813 16711 sw
tri 18813 16613 18911 16711 ne
rect 18911 16613 19265 16711
tri 19265 16613 19363 16711 sw
tri 19363 16613 19461 16711 ne
rect 19461 16613 20300 16711
rect -2000 16583 113 16613
tri 113 16583 143 16613 sw
tri 211 16583 241 16613 ne
rect 241 16583 663 16613
tri 663 16583 693 16613 sw
tri 761 16583 791 16613 ne
rect 791 16583 1213 16613
tri 1213 16583 1243 16613 sw
tri 1311 16583 1341 16613 ne
rect 1341 16583 1763 16613
tri 1763 16583 1793 16613 sw
tri 1861 16583 1891 16613 ne
rect 1891 16583 2313 16613
tri 2313 16583 2343 16613 sw
tri 2411 16583 2441 16613 ne
rect 2441 16583 2863 16613
tri 2863 16583 2893 16613 sw
tri 2961 16583 2991 16613 ne
rect 2991 16583 3413 16613
tri 3413 16583 3443 16613 sw
tri 3511 16583 3541 16613 ne
rect 3541 16583 3963 16613
tri 3963 16583 3993 16613 sw
tri 4061 16583 4091 16613 ne
rect 4091 16583 4513 16613
tri 4513 16583 4543 16613 sw
tri 4611 16583 4641 16613 ne
rect 4641 16583 5063 16613
tri 5063 16583 5093 16613 sw
tri 5161 16583 5191 16613 ne
rect 5191 16583 5613 16613
tri 5613 16583 5643 16613 sw
tri 5711 16583 5741 16613 ne
rect 5741 16583 6163 16613
tri 6163 16583 6193 16613 sw
tri 6261 16583 6291 16613 ne
rect 6291 16583 6713 16613
tri 6713 16583 6743 16613 sw
tri 6811 16583 6841 16613 ne
rect 6841 16583 7263 16613
tri 7263 16583 7293 16613 sw
tri 7361 16583 7391 16613 ne
rect 7391 16583 7813 16613
tri 7813 16583 7843 16613 sw
tri 7911 16583 7941 16613 ne
rect 7941 16583 8363 16613
tri 8363 16583 8393 16613 sw
tri 8461 16583 8491 16613 ne
rect 8491 16583 8913 16613
tri 8913 16583 8943 16613 sw
tri 9011 16583 9041 16613 ne
rect 9041 16583 9463 16613
tri 9463 16583 9493 16613 sw
tri 9561 16583 9591 16613 ne
rect 9591 16583 10013 16613
tri 10013 16583 10043 16613 sw
tri 10111 16583 10141 16613 ne
rect 10141 16583 10563 16613
tri 10563 16583 10593 16613 sw
tri 10661 16583 10691 16613 ne
rect 10691 16583 11113 16613
tri 11113 16583 11143 16613 sw
tri 11211 16583 11241 16613 ne
rect 11241 16583 11663 16613
tri 11663 16583 11693 16613 sw
tri 11761 16583 11791 16613 ne
rect 11791 16583 12213 16613
tri 12213 16583 12243 16613 sw
tri 12311 16583 12341 16613 ne
rect 12341 16583 12763 16613
tri 12763 16583 12793 16613 sw
tri 12861 16583 12891 16613 ne
rect 12891 16583 13313 16613
tri 13313 16583 13343 16613 sw
tri 13411 16583 13441 16613 ne
rect 13441 16583 13863 16613
tri 13863 16583 13893 16613 sw
tri 13961 16583 13991 16613 ne
rect 13991 16583 14413 16613
tri 14413 16583 14443 16613 sw
tri 14511 16583 14541 16613 ne
rect 14541 16583 14963 16613
tri 14963 16583 14993 16613 sw
tri 15061 16583 15091 16613 ne
rect 15091 16583 15513 16613
tri 15513 16583 15543 16613 sw
tri 15611 16583 15641 16613 ne
rect 15641 16583 16063 16613
tri 16063 16583 16093 16613 sw
tri 16161 16583 16191 16613 ne
rect 16191 16583 16613 16613
tri 16613 16583 16643 16613 sw
tri 16711 16583 16741 16613 ne
rect 16741 16583 17163 16613
tri 17163 16583 17193 16613 sw
tri 17261 16583 17291 16613 ne
rect 17291 16583 17713 16613
tri 17713 16583 17743 16613 sw
tri 17811 16583 17841 16613 ne
rect 17841 16583 18263 16613
tri 18263 16583 18293 16613 sw
tri 18361 16583 18391 16613 ne
rect 18391 16583 18813 16613
tri 18813 16583 18843 16613 sw
tri 18911 16583 18941 16613 ne
rect 18941 16583 19363 16613
tri 19363 16583 19393 16613 sw
tri 19461 16583 19491 16613 ne
rect 19491 16583 20300 16613
rect -2000 16485 143 16583
tri 143 16485 241 16583 sw
tri 241 16485 339 16583 ne
rect 339 16485 693 16583
tri 693 16485 791 16583 sw
tri 791 16485 889 16583 ne
rect 889 16485 1243 16583
tri 1243 16485 1341 16583 sw
tri 1341 16485 1439 16583 ne
rect 1439 16485 1793 16583
tri 1793 16485 1891 16583 sw
tri 1891 16485 1989 16583 ne
rect 1989 16485 2343 16583
tri 2343 16485 2441 16583 sw
tri 2441 16485 2539 16583 ne
rect 2539 16485 2893 16583
tri 2893 16485 2991 16583 sw
tri 2991 16485 3089 16583 ne
rect 3089 16485 3443 16583
tri 3443 16485 3541 16583 sw
tri 3541 16485 3639 16583 ne
rect 3639 16485 3993 16583
tri 3993 16485 4091 16583 sw
tri 4091 16485 4189 16583 ne
rect 4189 16485 4543 16583
tri 4543 16485 4641 16583 sw
tri 4641 16485 4739 16583 ne
rect 4739 16485 5093 16583
tri 5093 16485 5191 16583 sw
tri 5191 16485 5289 16583 ne
rect 5289 16485 5643 16583
tri 5643 16485 5741 16583 sw
tri 5741 16485 5839 16583 ne
rect 5839 16485 6193 16583
tri 6193 16485 6291 16583 sw
tri 6291 16485 6389 16583 ne
rect 6389 16485 6743 16583
tri 6743 16485 6841 16583 sw
tri 6841 16485 6939 16583 ne
rect 6939 16485 7293 16583
tri 7293 16485 7391 16583 sw
tri 7391 16485 7489 16583 ne
rect 7489 16485 7843 16583
tri 7843 16485 7941 16583 sw
tri 7941 16485 8039 16583 ne
rect 8039 16485 8393 16583
tri 8393 16485 8491 16583 sw
tri 8491 16485 8589 16583 ne
rect 8589 16485 8943 16583
tri 8943 16485 9041 16583 sw
tri 9041 16485 9139 16583 ne
rect 9139 16485 9493 16583
tri 9493 16485 9591 16583 sw
tri 9591 16485 9689 16583 ne
rect 9689 16485 10043 16583
tri 10043 16485 10141 16583 sw
tri 10141 16485 10239 16583 ne
rect 10239 16485 10593 16583
tri 10593 16485 10691 16583 sw
tri 10691 16485 10789 16583 ne
rect 10789 16485 11143 16583
tri 11143 16485 11241 16583 sw
tri 11241 16485 11339 16583 ne
rect 11339 16485 11693 16583
tri 11693 16485 11791 16583 sw
tri 11791 16485 11889 16583 ne
rect 11889 16485 12243 16583
tri 12243 16485 12341 16583 sw
tri 12341 16485 12439 16583 ne
rect 12439 16485 12793 16583
tri 12793 16485 12891 16583 sw
tri 12891 16485 12989 16583 ne
rect 12989 16485 13343 16583
tri 13343 16485 13441 16583 sw
tri 13441 16485 13539 16583 ne
rect 13539 16485 13893 16583
tri 13893 16485 13991 16583 sw
tri 13991 16485 14089 16583 ne
rect 14089 16485 14443 16583
tri 14443 16485 14541 16583 sw
tri 14541 16485 14639 16583 ne
rect 14639 16485 14993 16583
tri 14993 16485 15091 16583 sw
tri 15091 16485 15189 16583 ne
rect 15189 16485 15543 16583
tri 15543 16485 15641 16583 sw
tri 15641 16485 15739 16583 ne
rect 15739 16485 16093 16583
tri 16093 16485 16191 16583 sw
tri 16191 16485 16289 16583 ne
rect 16289 16485 16643 16583
tri 16643 16485 16741 16583 sw
tri 16741 16485 16839 16583 ne
rect 16839 16485 17193 16583
tri 17193 16485 17291 16583 sw
tri 17291 16485 17389 16583 ne
rect 17389 16485 17743 16583
tri 17743 16485 17841 16583 sw
tri 17841 16485 17939 16583 ne
rect 17939 16485 18293 16583
tri 18293 16485 18391 16583 sw
tri 18391 16485 18489 16583 ne
rect 18489 16485 18843 16583
tri 18843 16485 18941 16583 sw
tri 18941 16485 19039 16583 ne
rect 19039 16485 19393 16583
tri 19393 16485 19491 16583 sw
tri 19491 16485 19589 16583 ne
rect 19589 16485 20300 16583
rect -2000 16387 241 16485
tri 241 16387 339 16485 sw
tri 339 16387 437 16485 ne
rect 437 16387 791 16485
tri 791 16387 889 16485 sw
tri 889 16387 987 16485 ne
rect 987 16387 1341 16485
tri 1341 16387 1439 16485 sw
tri 1439 16387 1537 16485 ne
rect 1537 16387 1891 16485
tri 1891 16387 1989 16485 sw
tri 1989 16387 2087 16485 ne
rect 2087 16387 2441 16485
tri 2441 16387 2539 16485 sw
tri 2539 16387 2637 16485 ne
rect 2637 16387 2991 16485
tri 2991 16387 3089 16485 sw
tri 3089 16387 3187 16485 ne
rect 3187 16387 3541 16485
tri 3541 16387 3639 16485 sw
tri 3639 16387 3737 16485 ne
rect 3737 16387 4091 16485
tri 4091 16387 4189 16485 sw
tri 4189 16387 4287 16485 ne
rect 4287 16387 4641 16485
tri 4641 16387 4739 16485 sw
tri 4739 16387 4837 16485 ne
rect 4837 16387 5191 16485
tri 5191 16387 5289 16485 sw
tri 5289 16387 5387 16485 ne
rect 5387 16387 5741 16485
tri 5741 16387 5839 16485 sw
tri 5839 16387 5937 16485 ne
rect 5937 16387 6291 16485
tri 6291 16387 6389 16485 sw
tri 6389 16387 6487 16485 ne
rect 6487 16387 6841 16485
tri 6841 16387 6939 16485 sw
tri 6939 16387 7037 16485 ne
rect 7037 16387 7391 16485
tri 7391 16387 7489 16485 sw
tri 7489 16387 7587 16485 ne
rect 7587 16387 7941 16485
tri 7941 16387 8039 16485 sw
tri 8039 16387 8137 16485 ne
rect 8137 16387 8491 16485
tri 8491 16387 8589 16485 sw
tri 8589 16387 8687 16485 ne
rect 8687 16387 9041 16485
tri 9041 16387 9139 16485 sw
tri 9139 16387 9237 16485 ne
rect 9237 16387 9591 16485
tri 9591 16387 9689 16485 sw
tri 9689 16387 9787 16485 ne
rect 9787 16387 10141 16485
tri 10141 16387 10239 16485 sw
tri 10239 16387 10337 16485 ne
rect 10337 16387 10691 16485
tri 10691 16387 10789 16485 sw
tri 10789 16387 10887 16485 ne
rect 10887 16387 11241 16485
tri 11241 16387 11339 16485 sw
tri 11339 16387 11437 16485 ne
rect 11437 16387 11791 16485
tri 11791 16387 11889 16485 sw
tri 11889 16387 11987 16485 ne
rect 11987 16387 12341 16485
tri 12341 16387 12439 16485 sw
tri 12439 16387 12537 16485 ne
rect 12537 16387 12891 16485
tri 12891 16387 12989 16485 sw
tri 12989 16387 13087 16485 ne
rect 13087 16387 13441 16485
tri 13441 16387 13539 16485 sw
tri 13539 16387 13637 16485 ne
rect 13637 16387 13991 16485
tri 13991 16387 14089 16485 sw
tri 14089 16387 14187 16485 ne
rect 14187 16387 14541 16485
tri 14541 16387 14639 16485 sw
tri 14639 16387 14737 16485 ne
rect 14737 16387 15091 16485
tri 15091 16387 15189 16485 sw
tri 15189 16387 15287 16485 ne
rect 15287 16387 15641 16485
tri 15641 16387 15739 16485 sw
tri 15739 16387 15837 16485 ne
rect 15837 16387 16191 16485
tri 16191 16387 16289 16485 sw
tri 16289 16387 16387 16485 ne
rect 16387 16387 16741 16485
tri 16741 16387 16839 16485 sw
tri 16839 16387 16937 16485 ne
rect 16937 16387 17291 16485
tri 17291 16387 17389 16485 sw
tri 17389 16387 17487 16485 ne
rect 17487 16387 17841 16485
tri 17841 16387 17939 16485 sw
tri 17939 16387 18037 16485 ne
rect 18037 16387 18391 16485
tri 18391 16387 18489 16485 sw
tri 18489 16387 18587 16485 ne
rect 18587 16387 18941 16485
tri 18941 16387 19039 16485 sw
tri 19039 16387 19137 16485 ne
rect 19137 16387 19491 16485
tri 19491 16387 19589 16485 sw
tri 19589 16387 19687 16485 ne
rect 19687 16387 20300 16485
rect -2000 16289 339 16387
tri 339 16289 437 16387 sw
tri 437 16289 535 16387 ne
rect 535 16289 889 16387
tri 889 16289 987 16387 sw
tri 987 16289 1085 16387 ne
rect 1085 16289 1439 16387
tri 1439 16289 1537 16387 sw
tri 1537 16289 1635 16387 ne
rect 1635 16289 1989 16387
tri 1989 16289 2087 16387 sw
tri 2087 16289 2185 16387 ne
rect 2185 16289 2539 16387
tri 2539 16289 2637 16387 sw
tri 2637 16289 2735 16387 ne
rect 2735 16289 3089 16387
tri 3089 16289 3187 16387 sw
tri 3187 16289 3285 16387 ne
rect 3285 16289 3639 16387
tri 3639 16289 3737 16387 sw
tri 3737 16289 3835 16387 ne
rect 3835 16289 4189 16387
tri 4189 16289 4287 16387 sw
tri 4287 16289 4385 16387 ne
rect 4385 16289 4739 16387
tri 4739 16289 4837 16387 sw
tri 4837 16289 4935 16387 ne
rect 4935 16289 5289 16387
tri 5289 16289 5387 16387 sw
tri 5387 16289 5485 16387 ne
rect 5485 16289 5839 16387
tri 5839 16289 5937 16387 sw
tri 5937 16289 6035 16387 ne
rect 6035 16289 6389 16387
tri 6389 16289 6487 16387 sw
tri 6487 16289 6585 16387 ne
rect 6585 16289 6939 16387
tri 6939 16289 7037 16387 sw
tri 7037 16289 7135 16387 ne
rect 7135 16289 7489 16387
tri 7489 16289 7587 16387 sw
tri 7587 16289 7685 16387 ne
rect 7685 16289 8039 16387
tri 8039 16289 8137 16387 sw
tri 8137 16289 8235 16387 ne
rect 8235 16289 8589 16387
tri 8589 16289 8687 16387 sw
tri 8687 16289 8785 16387 ne
rect 8785 16289 9139 16387
tri 9139 16289 9237 16387 sw
tri 9237 16289 9335 16387 ne
rect 9335 16289 9689 16387
tri 9689 16289 9787 16387 sw
tri 9787 16289 9885 16387 ne
rect 9885 16289 10239 16387
tri 10239 16289 10337 16387 sw
tri 10337 16289 10435 16387 ne
rect 10435 16289 10789 16387
tri 10789 16289 10887 16387 sw
tri 10887 16289 10985 16387 ne
rect 10985 16289 11339 16387
tri 11339 16289 11437 16387 sw
tri 11437 16289 11535 16387 ne
rect 11535 16289 11889 16387
tri 11889 16289 11987 16387 sw
tri 11987 16289 12085 16387 ne
rect 12085 16289 12439 16387
tri 12439 16289 12537 16387 sw
tri 12537 16289 12635 16387 ne
rect 12635 16289 12989 16387
tri 12989 16289 13087 16387 sw
tri 13087 16289 13185 16387 ne
rect 13185 16289 13539 16387
tri 13539 16289 13637 16387 sw
tri 13637 16289 13735 16387 ne
rect 13735 16289 14089 16387
tri 14089 16289 14187 16387 sw
tri 14187 16289 14285 16387 ne
rect 14285 16289 14639 16387
tri 14639 16289 14737 16387 sw
tri 14737 16289 14835 16387 ne
rect 14835 16289 15189 16387
tri 15189 16289 15287 16387 sw
tri 15287 16289 15385 16387 ne
rect 15385 16289 15739 16387
tri 15739 16289 15837 16387 sw
tri 15837 16289 15935 16387 ne
rect 15935 16289 16289 16387
tri 16289 16289 16387 16387 sw
tri 16387 16289 16485 16387 ne
rect 16485 16289 16839 16387
tri 16839 16289 16937 16387 sw
tri 16937 16289 17035 16387 ne
rect 17035 16289 17389 16387
tri 17389 16289 17487 16387 sw
tri 17487 16289 17585 16387 ne
rect 17585 16289 17939 16387
tri 17939 16289 18037 16387 sw
tri 18037 16289 18135 16387 ne
rect 18135 16289 18489 16387
tri 18489 16289 18587 16387 sw
tri 18587 16289 18685 16387 ne
rect 18685 16289 19039 16387
tri 19039 16289 19137 16387 sw
tri 19137 16289 19235 16387 ne
rect 19235 16289 19589 16387
tri 19589 16289 19687 16387 sw
rect 20800 16289 21800 16937
rect -2000 16285 437 16289
rect -2000 16165 215 16285
rect 335 16191 437 16285
tri 437 16191 535 16289 sw
tri 535 16191 633 16289 ne
rect 633 16285 987 16289
rect 633 16191 765 16285
rect 335 16165 535 16191
rect -2000 16161 535 16165
rect -2000 15513 -1000 16161
tri 113 16063 211 16161 ne
rect 211 16113 535 16161
tri 535 16113 613 16191 sw
tri 633 16113 711 16191 ne
rect 711 16165 765 16191
rect 885 16191 987 16285
tri 987 16191 1085 16289 sw
tri 1085 16191 1183 16289 ne
rect 1183 16285 1537 16289
rect 1183 16191 1315 16285
rect 885 16165 1085 16191
rect 711 16113 1085 16165
tri 1085 16113 1163 16191 sw
tri 1183 16113 1261 16191 ne
rect 1261 16165 1315 16191
rect 1435 16191 1537 16285
tri 1537 16191 1635 16289 sw
tri 1635 16191 1733 16289 ne
rect 1733 16285 2087 16289
rect 1733 16191 1865 16285
rect 1435 16165 1635 16191
rect 1261 16113 1635 16165
tri 1635 16113 1713 16191 sw
tri 1733 16113 1811 16191 ne
rect 1811 16165 1865 16191
rect 1985 16191 2087 16285
tri 2087 16191 2185 16289 sw
tri 2185 16191 2283 16289 ne
rect 2283 16285 2637 16289
rect 2283 16191 2415 16285
rect 1985 16165 2185 16191
rect 1811 16113 2185 16165
tri 2185 16113 2263 16191 sw
tri 2283 16113 2361 16191 ne
rect 2361 16165 2415 16191
rect 2535 16191 2637 16285
tri 2637 16191 2735 16289 sw
tri 2735 16191 2833 16289 ne
rect 2833 16285 3187 16289
rect 2833 16191 2965 16285
rect 2535 16165 2735 16191
rect 2361 16113 2735 16165
tri 2735 16113 2813 16191 sw
tri 2833 16113 2911 16191 ne
rect 2911 16165 2965 16191
rect 3085 16191 3187 16285
tri 3187 16191 3285 16289 sw
tri 3285 16191 3383 16289 ne
rect 3383 16285 3737 16289
rect 3383 16191 3515 16285
rect 3085 16165 3285 16191
rect 2911 16113 3285 16165
tri 3285 16113 3363 16191 sw
tri 3383 16113 3461 16191 ne
rect 3461 16165 3515 16191
rect 3635 16191 3737 16285
tri 3737 16191 3835 16289 sw
tri 3835 16191 3933 16289 ne
rect 3933 16285 4287 16289
rect 3933 16191 4065 16285
rect 3635 16165 3835 16191
rect 3461 16113 3835 16165
tri 3835 16113 3913 16191 sw
tri 3933 16113 4011 16191 ne
rect 4011 16165 4065 16191
rect 4185 16191 4287 16285
tri 4287 16191 4385 16289 sw
tri 4385 16191 4483 16289 ne
rect 4483 16285 4837 16289
rect 4483 16191 4615 16285
rect 4185 16165 4385 16191
rect 4011 16113 4385 16165
tri 4385 16113 4463 16191 sw
tri 4483 16113 4561 16191 ne
rect 4561 16165 4615 16191
rect 4735 16191 4837 16285
tri 4837 16191 4935 16289 sw
tri 4935 16191 5033 16289 ne
rect 5033 16285 5387 16289
rect 5033 16191 5165 16285
rect 4735 16165 4935 16191
rect 4561 16113 4935 16165
tri 4935 16113 5013 16191 sw
tri 5033 16113 5111 16191 ne
rect 5111 16165 5165 16191
rect 5285 16191 5387 16285
tri 5387 16191 5485 16289 sw
tri 5485 16191 5583 16289 ne
rect 5583 16285 5937 16289
rect 5583 16191 5715 16285
rect 5285 16165 5485 16191
rect 5111 16113 5485 16165
tri 5485 16113 5563 16191 sw
tri 5583 16113 5661 16191 ne
rect 5661 16165 5715 16191
rect 5835 16191 5937 16285
tri 5937 16191 6035 16289 sw
tri 6035 16191 6133 16289 ne
rect 6133 16285 6487 16289
rect 6133 16191 6265 16285
rect 5835 16165 6035 16191
rect 5661 16113 6035 16165
tri 6035 16113 6113 16191 sw
tri 6133 16113 6211 16191 ne
rect 6211 16165 6265 16191
rect 6385 16191 6487 16285
tri 6487 16191 6585 16289 sw
tri 6585 16191 6683 16289 ne
rect 6683 16285 7037 16289
rect 6683 16191 6815 16285
rect 6385 16165 6585 16191
rect 6211 16113 6585 16165
tri 6585 16113 6663 16191 sw
tri 6683 16113 6761 16191 ne
rect 6761 16165 6815 16191
rect 6935 16191 7037 16285
tri 7037 16191 7135 16289 sw
tri 7135 16191 7233 16289 ne
rect 7233 16285 7587 16289
rect 7233 16191 7365 16285
rect 6935 16165 7135 16191
rect 6761 16113 7135 16165
tri 7135 16113 7213 16191 sw
tri 7233 16113 7311 16191 ne
rect 7311 16165 7365 16191
rect 7485 16191 7587 16285
tri 7587 16191 7685 16289 sw
tri 7685 16191 7783 16289 ne
rect 7783 16285 8137 16289
rect 7783 16191 7915 16285
rect 7485 16165 7685 16191
rect 7311 16113 7685 16165
tri 7685 16113 7763 16191 sw
tri 7783 16113 7861 16191 ne
rect 7861 16165 7915 16191
rect 8035 16191 8137 16285
tri 8137 16191 8235 16289 sw
tri 8235 16191 8333 16289 ne
rect 8333 16285 8687 16289
rect 8333 16191 8465 16285
rect 8035 16165 8235 16191
rect 7861 16113 8235 16165
tri 8235 16113 8313 16191 sw
tri 8333 16113 8411 16191 ne
rect 8411 16165 8465 16191
rect 8585 16191 8687 16285
tri 8687 16191 8785 16289 sw
tri 8785 16191 8883 16289 ne
rect 8883 16285 9237 16289
rect 8883 16191 9015 16285
rect 8585 16165 8785 16191
rect 8411 16113 8785 16165
tri 8785 16113 8863 16191 sw
tri 8883 16113 8961 16191 ne
rect 8961 16165 9015 16191
rect 9135 16191 9237 16285
tri 9237 16191 9335 16289 sw
tri 9335 16191 9433 16289 ne
rect 9433 16285 9787 16289
rect 9433 16191 9565 16285
rect 9135 16165 9335 16191
rect 8961 16113 9335 16165
tri 9335 16113 9413 16191 sw
tri 9433 16113 9511 16191 ne
rect 9511 16165 9565 16191
rect 9685 16191 9787 16285
tri 9787 16191 9885 16289 sw
tri 9885 16191 9983 16289 ne
rect 9983 16285 10337 16289
rect 9983 16191 10115 16285
rect 9685 16165 9885 16191
rect 9511 16113 9885 16165
tri 9885 16113 9963 16191 sw
tri 9983 16113 10061 16191 ne
rect 10061 16165 10115 16191
rect 10235 16191 10337 16285
tri 10337 16191 10435 16289 sw
tri 10435 16191 10533 16289 ne
rect 10533 16285 10887 16289
rect 10533 16191 10665 16285
rect 10235 16165 10435 16191
rect 10061 16113 10435 16165
tri 10435 16113 10513 16191 sw
tri 10533 16113 10611 16191 ne
rect 10611 16165 10665 16191
rect 10785 16191 10887 16285
tri 10887 16191 10985 16289 sw
tri 10985 16191 11083 16289 ne
rect 11083 16285 11437 16289
rect 11083 16191 11215 16285
rect 10785 16165 10985 16191
rect 10611 16113 10985 16165
tri 10985 16113 11063 16191 sw
tri 11083 16113 11161 16191 ne
rect 11161 16165 11215 16191
rect 11335 16191 11437 16285
tri 11437 16191 11535 16289 sw
tri 11535 16191 11633 16289 ne
rect 11633 16285 11987 16289
rect 11633 16191 11765 16285
rect 11335 16165 11535 16191
rect 11161 16113 11535 16165
tri 11535 16113 11613 16191 sw
tri 11633 16113 11711 16191 ne
rect 11711 16165 11765 16191
rect 11885 16191 11987 16285
tri 11987 16191 12085 16289 sw
tri 12085 16191 12183 16289 ne
rect 12183 16285 12537 16289
rect 12183 16191 12315 16285
rect 11885 16165 12085 16191
rect 11711 16113 12085 16165
tri 12085 16113 12163 16191 sw
tri 12183 16113 12261 16191 ne
rect 12261 16165 12315 16191
rect 12435 16191 12537 16285
tri 12537 16191 12635 16289 sw
tri 12635 16191 12733 16289 ne
rect 12733 16285 13087 16289
rect 12733 16191 12865 16285
rect 12435 16165 12635 16191
rect 12261 16113 12635 16165
tri 12635 16113 12713 16191 sw
tri 12733 16113 12811 16191 ne
rect 12811 16165 12865 16191
rect 12985 16191 13087 16285
tri 13087 16191 13185 16289 sw
tri 13185 16191 13283 16289 ne
rect 13283 16285 13637 16289
rect 13283 16191 13415 16285
rect 12985 16165 13185 16191
rect 12811 16113 13185 16165
tri 13185 16113 13263 16191 sw
tri 13283 16113 13361 16191 ne
rect 13361 16165 13415 16191
rect 13535 16191 13637 16285
tri 13637 16191 13735 16289 sw
tri 13735 16191 13833 16289 ne
rect 13833 16285 14187 16289
rect 13833 16191 13965 16285
rect 13535 16165 13735 16191
rect 13361 16113 13735 16165
tri 13735 16113 13813 16191 sw
tri 13833 16113 13911 16191 ne
rect 13911 16165 13965 16191
rect 14085 16191 14187 16285
tri 14187 16191 14285 16289 sw
tri 14285 16191 14383 16289 ne
rect 14383 16285 14737 16289
rect 14383 16191 14515 16285
rect 14085 16165 14285 16191
rect 13911 16113 14285 16165
tri 14285 16113 14363 16191 sw
tri 14383 16113 14461 16191 ne
rect 14461 16165 14515 16191
rect 14635 16191 14737 16285
tri 14737 16191 14835 16289 sw
tri 14835 16191 14933 16289 ne
rect 14933 16285 15287 16289
rect 14933 16191 15065 16285
rect 14635 16165 14835 16191
rect 14461 16113 14835 16165
tri 14835 16113 14913 16191 sw
tri 14933 16113 15011 16191 ne
rect 15011 16165 15065 16191
rect 15185 16191 15287 16285
tri 15287 16191 15385 16289 sw
tri 15385 16191 15483 16289 ne
rect 15483 16285 15837 16289
rect 15483 16191 15615 16285
rect 15185 16165 15385 16191
rect 15011 16113 15385 16165
tri 15385 16113 15463 16191 sw
tri 15483 16113 15561 16191 ne
rect 15561 16165 15615 16191
rect 15735 16191 15837 16285
tri 15837 16191 15935 16289 sw
tri 15935 16191 16033 16289 ne
rect 16033 16285 16387 16289
rect 16033 16191 16165 16285
rect 15735 16165 15935 16191
rect 15561 16113 15935 16165
tri 15935 16113 16013 16191 sw
tri 16033 16113 16111 16191 ne
rect 16111 16165 16165 16191
rect 16285 16191 16387 16285
tri 16387 16191 16485 16289 sw
tri 16485 16191 16583 16289 ne
rect 16583 16285 16937 16289
rect 16583 16191 16715 16285
rect 16285 16165 16485 16191
rect 16111 16113 16485 16165
tri 16485 16113 16563 16191 sw
tri 16583 16113 16661 16191 ne
rect 16661 16165 16715 16191
rect 16835 16191 16937 16285
tri 16937 16191 17035 16289 sw
tri 17035 16191 17133 16289 ne
rect 17133 16285 17487 16289
rect 17133 16191 17265 16285
rect 16835 16165 17035 16191
rect 16661 16113 17035 16165
tri 17035 16113 17113 16191 sw
tri 17133 16113 17211 16191 ne
rect 17211 16165 17265 16191
rect 17385 16191 17487 16285
tri 17487 16191 17585 16289 sw
tri 17585 16191 17683 16289 ne
rect 17683 16285 18037 16289
rect 17683 16191 17815 16285
rect 17385 16165 17585 16191
rect 17211 16113 17585 16165
tri 17585 16113 17663 16191 sw
tri 17683 16113 17761 16191 ne
rect 17761 16165 17815 16191
rect 17935 16191 18037 16285
tri 18037 16191 18135 16289 sw
tri 18135 16191 18233 16289 ne
rect 18233 16285 18587 16289
rect 18233 16191 18365 16285
rect 17935 16165 18135 16191
rect 17761 16113 18135 16165
tri 18135 16113 18213 16191 sw
tri 18233 16113 18311 16191 ne
rect 18311 16165 18365 16191
rect 18485 16191 18587 16285
tri 18587 16191 18685 16289 sw
tri 18685 16191 18783 16289 ne
rect 18783 16285 19137 16289
rect 18783 16191 18915 16285
rect 18485 16165 18685 16191
rect 18311 16113 18685 16165
tri 18685 16113 18763 16191 sw
tri 18783 16113 18861 16191 ne
rect 18861 16165 18915 16191
rect 19035 16191 19137 16285
tri 19137 16191 19235 16289 sw
tri 19235 16191 19333 16289 ne
rect 19333 16285 21800 16289
rect 19333 16191 19465 16285
rect 19035 16165 19235 16191
rect 18861 16113 19235 16165
tri 19235 16113 19313 16191 sw
tri 19333 16113 19411 16191 ne
rect 19411 16165 19465 16191
rect 19585 16165 21800 16285
rect 19411 16113 21800 16165
rect 211 16063 613 16113
rect -500 16013 113 16063
tri 113 16013 163 16063 sw
tri 211 16013 261 16063 ne
rect 261 16033 613 16063
tri 613 16033 693 16113 sw
tri 711 16033 791 16113 ne
rect 791 16033 1163 16113
tri 1163 16033 1243 16113 sw
tri 1261 16033 1341 16113 ne
rect 1341 16033 1713 16113
tri 1713 16033 1793 16113 sw
tri 1811 16033 1891 16113 ne
rect 1891 16033 2263 16113
tri 2263 16033 2343 16113 sw
tri 2361 16033 2441 16113 ne
rect 2441 16033 2813 16113
tri 2813 16033 2893 16113 sw
tri 2911 16033 2991 16113 ne
rect 2991 16033 3363 16113
tri 3363 16033 3443 16113 sw
tri 3461 16033 3541 16113 ne
rect 3541 16033 3913 16113
tri 3913 16033 3993 16113 sw
tri 4011 16033 4091 16113 ne
rect 4091 16033 4463 16113
tri 4463 16033 4543 16113 sw
tri 4561 16033 4641 16113 ne
rect 4641 16033 5013 16113
tri 5013 16033 5093 16113 sw
tri 5111 16033 5191 16113 ne
rect 5191 16033 5563 16113
tri 5563 16033 5643 16113 sw
tri 5661 16033 5741 16113 ne
rect 5741 16033 6113 16113
tri 6113 16033 6193 16113 sw
tri 6211 16033 6291 16113 ne
rect 6291 16033 6663 16113
tri 6663 16033 6743 16113 sw
tri 6761 16033 6841 16113 ne
rect 6841 16033 7213 16113
tri 7213 16033 7293 16113 sw
tri 7311 16033 7391 16113 ne
rect 7391 16033 7763 16113
tri 7763 16033 7843 16113 sw
tri 7861 16033 7941 16113 ne
rect 7941 16033 8313 16113
tri 8313 16033 8393 16113 sw
tri 8411 16033 8491 16113 ne
rect 8491 16033 8863 16113
tri 8863 16033 8943 16113 sw
tri 8961 16033 9041 16113 ne
rect 9041 16033 9413 16113
tri 9413 16033 9493 16113 sw
tri 9511 16033 9591 16113 ne
rect 9591 16033 9963 16113
tri 9963 16033 10043 16113 sw
tri 10061 16033 10141 16113 ne
rect 10141 16033 10513 16113
tri 10513 16033 10593 16113 sw
tri 10611 16033 10691 16113 ne
rect 10691 16033 11063 16113
tri 11063 16033 11143 16113 sw
tri 11161 16033 11241 16113 ne
rect 11241 16033 11613 16113
tri 11613 16033 11693 16113 sw
tri 11711 16033 11791 16113 ne
rect 11791 16033 12163 16113
tri 12163 16033 12243 16113 sw
tri 12261 16033 12341 16113 ne
rect 12341 16033 12713 16113
tri 12713 16033 12793 16113 sw
tri 12811 16033 12891 16113 ne
rect 12891 16033 13263 16113
tri 13263 16033 13343 16113 sw
tri 13361 16033 13441 16113 ne
rect 13441 16033 13813 16113
tri 13813 16033 13893 16113 sw
tri 13911 16033 13991 16113 ne
rect 13991 16033 14363 16113
tri 14363 16033 14443 16113 sw
tri 14461 16033 14541 16113 ne
rect 14541 16033 14913 16113
tri 14913 16033 14993 16113 sw
tri 15011 16033 15091 16113 ne
rect 15091 16033 15463 16113
tri 15463 16033 15543 16113 sw
tri 15561 16033 15641 16113 ne
rect 15641 16033 16013 16113
tri 16013 16033 16093 16113 sw
tri 16111 16033 16191 16113 ne
rect 16191 16033 16563 16113
tri 16563 16033 16643 16113 sw
tri 16661 16033 16741 16113 ne
rect 16741 16033 17113 16113
tri 17113 16033 17193 16113 sw
tri 17211 16033 17291 16113 ne
rect 17291 16033 17663 16113
tri 17663 16033 17743 16113 sw
tri 17761 16033 17841 16113 ne
rect 17841 16033 18213 16113
tri 18213 16033 18293 16113 sw
tri 18311 16033 18391 16113 ne
rect 18391 16033 18763 16113
tri 18763 16033 18843 16113 sw
tri 18861 16033 18941 16113 ne
rect 18941 16033 19313 16113
tri 19313 16033 19393 16113 sw
tri 19411 16033 19491 16113 ne
rect 19491 16033 20100 16113
rect 261 16013 693 16033
rect -500 15935 163 16013
tri 163 15935 241 16013 sw
tri 261 15935 339 16013 ne
rect 339 15935 693 16013
tri 693 15935 791 16033 sw
tri 791 15935 889 16033 ne
rect 889 15935 1243 16033
tri 1243 15935 1341 16033 sw
tri 1341 15935 1439 16033 ne
rect 1439 15935 1793 16033
tri 1793 15935 1891 16033 sw
tri 1891 15935 1989 16033 ne
rect 1989 15935 2343 16033
tri 2343 15935 2441 16033 sw
tri 2441 15935 2539 16033 ne
rect 2539 15935 2893 16033
tri 2893 15935 2991 16033 sw
tri 2991 15935 3089 16033 ne
rect 3089 15935 3443 16033
tri 3443 15935 3541 16033 sw
tri 3541 15935 3639 16033 ne
rect 3639 15935 3993 16033
tri 3993 15935 4091 16033 sw
tri 4091 15935 4189 16033 ne
rect 4189 15935 4543 16033
tri 4543 15935 4641 16033 sw
tri 4641 15935 4739 16033 ne
rect 4739 15935 5093 16033
tri 5093 15935 5191 16033 sw
tri 5191 15935 5289 16033 ne
rect 5289 15935 5643 16033
tri 5643 15935 5741 16033 sw
tri 5741 15935 5839 16033 ne
rect 5839 15935 6193 16033
tri 6193 15935 6291 16033 sw
tri 6291 15935 6389 16033 ne
rect 6389 15935 6743 16033
tri 6743 15935 6841 16033 sw
tri 6841 15935 6939 16033 ne
rect 6939 15935 7293 16033
tri 7293 15935 7391 16033 sw
tri 7391 15935 7489 16033 ne
rect 7489 15935 7843 16033
tri 7843 15935 7941 16033 sw
tri 7941 15935 8039 16033 ne
rect 8039 15935 8393 16033
tri 8393 15935 8491 16033 sw
tri 8491 15935 8589 16033 ne
rect 8589 15935 8943 16033
tri 8943 15935 9041 16033 sw
tri 9041 15935 9139 16033 ne
rect 9139 15935 9493 16033
tri 9493 15935 9591 16033 sw
tri 9591 15935 9689 16033 ne
rect 9689 15935 10043 16033
tri 10043 15935 10141 16033 sw
tri 10141 15935 10239 16033 ne
rect 10239 15935 10593 16033
tri 10593 15935 10691 16033 sw
tri 10691 15935 10789 16033 ne
rect 10789 15935 11143 16033
tri 11143 15935 11241 16033 sw
tri 11241 15935 11339 16033 ne
rect 11339 15935 11693 16033
tri 11693 15935 11791 16033 sw
tri 11791 15935 11889 16033 ne
rect 11889 15935 12243 16033
tri 12243 15935 12341 16033 sw
tri 12341 15935 12439 16033 ne
rect 12439 15935 12793 16033
tri 12793 15935 12891 16033 sw
tri 12891 15935 12989 16033 ne
rect 12989 15935 13343 16033
tri 13343 15935 13441 16033 sw
tri 13441 15935 13539 16033 ne
rect 13539 15935 13893 16033
tri 13893 15935 13991 16033 sw
tri 13991 15935 14089 16033 ne
rect 14089 15935 14443 16033
tri 14443 15935 14541 16033 sw
tri 14541 15935 14639 16033 ne
rect 14639 15935 14993 16033
tri 14993 15935 15091 16033 sw
tri 15091 15935 15189 16033 ne
rect 15189 15935 15543 16033
tri 15543 15935 15641 16033 sw
tri 15641 15935 15739 16033 ne
rect 15739 15935 16093 16033
tri 16093 15935 16191 16033 sw
tri 16191 15935 16289 16033 ne
rect 16289 15935 16643 16033
tri 16643 15935 16741 16033 sw
tri 16741 15935 16839 16033 ne
rect 16839 15935 17193 16033
tri 17193 15935 17291 16033 sw
tri 17291 15935 17389 16033 ne
rect 17389 15935 17743 16033
tri 17743 15935 17841 16033 sw
tri 17841 15935 17939 16033 ne
rect 17939 15935 18293 16033
tri 18293 15935 18391 16033 sw
tri 18391 15935 18489 16033 ne
rect 18489 15935 18843 16033
tri 18843 15935 18941 16033 sw
tri 18941 15935 19039 16033 ne
rect 19039 15935 19393 16033
tri 19393 15935 19491 16033 sw
tri 19491 15935 19589 16033 ne
rect 19589 16013 20100 16033
rect 20200 16013 21800 16113
rect 19589 15935 21800 16013
rect -500 15887 241 15935
rect -500 15787 -400 15887
rect -300 15837 241 15887
tri 241 15837 339 15935 sw
tri 339 15837 437 15935 ne
rect 437 15837 791 15935
tri 791 15837 889 15935 sw
tri 889 15837 987 15935 ne
rect 987 15837 1341 15935
tri 1341 15837 1439 15935 sw
tri 1439 15837 1537 15935 ne
rect 1537 15837 1891 15935
tri 1891 15837 1989 15935 sw
tri 1989 15837 2087 15935 ne
rect 2087 15837 2441 15935
tri 2441 15837 2539 15935 sw
tri 2539 15837 2637 15935 ne
rect 2637 15837 2991 15935
tri 2991 15837 3089 15935 sw
tri 3089 15837 3187 15935 ne
rect 3187 15837 3541 15935
tri 3541 15837 3639 15935 sw
tri 3639 15837 3737 15935 ne
rect 3737 15837 4091 15935
tri 4091 15837 4189 15935 sw
tri 4189 15837 4287 15935 ne
rect 4287 15837 4641 15935
tri 4641 15837 4739 15935 sw
tri 4739 15837 4837 15935 ne
rect 4837 15837 5191 15935
tri 5191 15837 5289 15935 sw
tri 5289 15837 5387 15935 ne
rect 5387 15837 5741 15935
tri 5741 15837 5839 15935 sw
tri 5839 15837 5937 15935 ne
rect 5937 15837 6291 15935
tri 6291 15837 6389 15935 sw
tri 6389 15837 6487 15935 ne
rect 6487 15837 6841 15935
tri 6841 15837 6939 15935 sw
tri 6939 15837 7037 15935 ne
rect 7037 15837 7391 15935
tri 7391 15837 7489 15935 sw
tri 7489 15837 7587 15935 ne
rect 7587 15837 7941 15935
tri 7941 15837 8039 15935 sw
tri 8039 15837 8137 15935 ne
rect 8137 15837 8491 15935
tri 8491 15837 8589 15935 sw
tri 8589 15837 8687 15935 ne
rect 8687 15837 9041 15935
tri 9041 15837 9139 15935 sw
tri 9139 15837 9237 15935 ne
rect 9237 15837 9591 15935
tri 9591 15837 9689 15935 sw
tri 9689 15837 9787 15935 ne
rect 9787 15837 10141 15935
tri 10141 15837 10239 15935 sw
tri 10239 15837 10337 15935 ne
rect 10337 15837 10691 15935
tri 10691 15837 10789 15935 sw
tri 10789 15837 10887 15935 ne
rect 10887 15837 11241 15935
tri 11241 15837 11339 15935 sw
tri 11339 15837 11437 15935 ne
rect 11437 15837 11791 15935
tri 11791 15837 11889 15935 sw
tri 11889 15837 11987 15935 ne
rect 11987 15837 12341 15935
tri 12341 15837 12439 15935 sw
tri 12439 15837 12537 15935 ne
rect 12537 15837 12891 15935
tri 12891 15837 12989 15935 sw
tri 12989 15837 13087 15935 ne
rect 13087 15837 13441 15935
tri 13441 15837 13539 15935 sw
tri 13539 15837 13637 15935 ne
rect 13637 15837 13991 15935
tri 13991 15837 14089 15935 sw
tri 14089 15837 14187 15935 ne
rect 14187 15837 14541 15935
tri 14541 15837 14639 15935 sw
tri 14639 15837 14737 15935 ne
rect 14737 15837 15091 15935
tri 15091 15837 15189 15935 sw
tri 15189 15837 15287 15935 ne
rect 15287 15837 15641 15935
tri 15641 15837 15739 15935 sw
tri 15739 15837 15837 15935 ne
rect 15837 15837 16191 15935
tri 16191 15837 16289 15935 sw
tri 16289 15837 16387 15935 ne
rect 16387 15837 16741 15935
tri 16741 15837 16839 15935 sw
tri 16839 15837 16937 15935 ne
rect 16937 15837 17291 15935
tri 17291 15837 17389 15935 sw
tri 17389 15837 17487 15935 ne
rect 17487 15837 17841 15935
tri 17841 15837 17939 15935 sw
tri 17939 15837 18037 15935 ne
rect 18037 15837 18391 15935
tri 18391 15837 18489 15935 sw
tri 18489 15837 18587 15935 ne
rect 18587 15837 18941 15935
tri 18941 15837 19039 15935 sw
tri 19039 15837 19137 15935 ne
rect 19137 15837 19491 15935
tri 19491 15837 19589 15935 sw
tri 19589 15837 19687 15935 ne
rect 19687 15837 21800 15935
rect -300 15787 339 15837
rect -500 15739 339 15787
tri 339 15739 437 15837 sw
tri 437 15739 535 15837 ne
rect 535 15739 889 15837
tri 889 15739 987 15837 sw
tri 987 15739 1085 15837 ne
rect 1085 15739 1439 15837
tri 1439 15739 1537 15837 sw
tri 1537 15739 1635 15837 ne
rect 1635 15739 1989 15837
tri 1989 15739 2087 15837 sw
tri 2087 15739 2185 15837 ne
rect 2185 15739 2539 15837
tri 2539 15739 2637 15837 sw
tri 2637 15739 2735 15837 ne
rect 2735 15739 3089 15837
tri 3089 15739 3187 15837 sw
tri 3187 15739 3285 15837 ne
rect 3285 15739 3639 15837
tri 3639 15739 3737 15837 sw
tri 3737 15739 3835 15837 ne
rect 3835 15739 4189 15837
tri 4189 15739 4287 15837 sw
tri 4287 15739 4385 15837 ne
rect 4385 15739 4739 15837
tri 4739 15739 4837 15837 sw
tri 4837 15739 4935 15837 ne
rect 4935 15739 5289 15837
tri 5289 15739 5387 15837 sw
tri 5387 15739 5485 15837 ne
rect 5485 15739 5839 15837
tri 5839 15739 5937 15837 sw
tri 5937 15739 6035 15837 ne
rect 6035 15739 6389 15837
tri 6389 15739 6487 15837 sw
tri 6487 15739 6585 15837 ne
rect 6585 15739 6939 15837
tri 6939 15739 7037 15837 sw
tri 7037 15739 7135 15837 ne
rect 7135 15739 7489 15837
tri 7489 15739 7587 15837 sw
tri 7587 15739 7685 15837 ne
rect 7685 15739 8039 15837
tri 8039 15739 8137 15837 sw
tri 8137 15739 8235 15837 ne
rect 8235 15739 8589 15837
tri 8589 15739 8687 15837 sw
tri 8687 15739 8785 15837 ne
rect 8785 15739 9139 15837
tri 9139 15739 9237 15837 sw
tri 9237 15739 9335 15837 ne
rect 9335 15739 9689 15837
tri 9689 15739 9787 15837 sw
tri 9787 15739 9885 15837 ne
rect 9885 15739 10239 15837
tri 10239 15739 10337 15837 sw
tri 10337 15739 10435 15837 ne
rect 10435 15739 10789 15837
tri 10789 15739 10887 15837 sw
tri 10887 15739 10985 15837 ne
rect 10985 15739 11339 15837
tri 11339 15739 11437 15837 sw
tri 11437 15739 11535 15837 ne
rect 11535 15739 11889 15837
tri 11889 15739 11987 15837 sw
tri 11987 15739 12085 15837 ne
rect 12085 15739 12439 15837
tri 12439 15739 12537 15837 sw
tri 12537 15739 12635 15837 ne
rect 12635 15739 12989 15837
tri 12989 15739 13087 15837 sw
tri 13087 15739 13185 15837 ne
rect 13185 15739 13539 15837
tri 13539 15739 13637 15837 sw
tri 13637 15739 13735 15837 ne
rect 13735 15739 14089 15837
tri 14089 15739 14187 15837 sw
tri 14187 15739 14285 15837 ne
rect 14285 15739 14639 15837
tri 14639 15739 14737 15837 sw
tri 14737 15739 14835 15837 ne
rect 14835 15739 15189 15837
tri 15189 15739 15287 15837 sw
tri 15287 15739 15385 15837 ne
rect 15385 15739 15739 15837
tri 15739 15739 15837 15837 sw
tri 15837 15739 15935 15837 ne
rect 15935 15739 16289 15837
tri 16289 15739 16387 15837 sw
tri 16387 15739 16485 15837 ne
rect 16485 15739 16839 15837
tri 16839 15739 16937 15837 sw
tri 16937 15739 17035 15837 ne
rect 17035 15739 17389 15837
tri 17389 15739 17487 15837 sw
tri 17487 15739 17585 15837 ne
rect 17585 15739 17939 15837
tri 17939 15739 18037 15837 sw
tri 18037 15739 18135 15837 ne
rect 18135 15739 18489 15837
tri 18489 15739 18587 15837 sw
tri 18587 15739 18685 15837 ne
rect 18685 15739 19039 15837
tri 19039 15739 19137 15837 sw
tri 19137 15739 19235 15837 ne
rect 19235 15739 19589 15837
tri 19589 15739 19687 15837 sw
rect -500 15735 437 15739
rect -500 15615 215 15735
rect 335 15641 437 15735
tri 437 15641 535 15739 sw
tri 535 15641 633 15739 ne
rect 633 15735 987 15739
rect 633 15641 765 15735
rect 335 15615 535 15641
rect -500 15611 535 15615
tri 535 15611 565 15641 sw
tri 633 15611 663 15641 ne
rect 663 15615 765 15641
rect 885 15641 987 15735
tri 987 15641 1085 15739 sw
tri 1085 15641 1183 15739 ne
rect 1183 15735 1537 15739
rect 1183 15641 1315 15735
rect 885 15615 1085 15641
rect 663 15611 1085 15615
tri 1085 15611 1115 15641 sw
tri 1183 15611 1213 15641 ne
rect 1213 15615 1315 15641
rect 1435 15641 1537 15735
tri 1537 15641 1635 15739 sw
tri 1635 15641 1733 15739 ne
rect 1733 15735 2087 15739
rect 1733 15641 1865 15735
rect 1435 15615 1635 15641
rect 1213 15611 1635 15615
tri 1635 15611 1665 15641 sw
tri 1733 15611 1763 15641 ne
rect 1763 15615 1865 15641
rect 1985 15641 2087 15735
tri 2087 15641 2185 15739 sw
tri 2185 15641 2283 15739 ne
rect 2283 15735 2637 15739
rect 2283 15641 2415 15735
rect 1985 15615 2185 15641
rect 1763 15611 2185 15615
tri 2185 15611 2215 15641 sw
tri 2283 15611 2313 15641 ne
rect 2313 15615 2415 15641
rect 2535 15641 2637 15735
tri 2637 15641 2735 15739 sw
tri 2735 15641 2833 15739 ne
rect 2833 15735 3187 15739
rect 2833 15641 2965 15735
rect 2535 15615 2735 15641
rect 2313 15611 2735 15615
tri 2735 15611 2765 15641 sw
tri 2833 15611 2863 15641 ne
rect 2863 15615 2965 15641
rect 3085 15641 3187 15735
tri 3187 15641 3285 15739 sw
tri 3285 15641 3383 15739 ne
rect 3383 15735 3737 15739
rect 3383 15641 3515 15735
rect 3085 15615 3285 15641
rect 2863 15611 3285 15615
tri 3285 15611 3315 15641 sw
tri 3383 15611 3413 15641 ne
rect 3413 15615 3515 15641
rect 3635 15641 3737 15735
tri 3737 15641 3835 15739 sw
tri 3835 15641 3933 15739 ne
rect 3933 15735 4287 15739
rect 3933 15641 4065 15735
rect 3635 15615 3835 15641
rect 3413 15611 3835 15615
tri 3835 15611 3865 15641 sw
tri 3933 15611 3963 15641 ne
rect 3963 15615 4065 15641
rect 4185 15641 4287 15735
tri 4287 15641 4385 15739 sw
tri 4385 15641 4483 15739 ne
rect 4483 15735 4837 15739
rect 4483 15641 4615 15735
rect 4185 15615 4385 15641
rect 3963 15611 4385 15615
tri 4385 15611 4415 15641 sw
tri 4483 15611 4513 15641 ne
rect 4513 15615 4615 15641
rect 4735 15641 4837 15735
tri 4837 15641 4935 15739 sw
tri 4935 15641 5033 15739 ne
rect 5033 15735 5387 15739
rect 5033 15641 5165 15735
rect 4735 15615 4935 15641
rect 4513 15611 4935 15615
tri 4935 15611 4965 15641 sw
tri 5033 15611 5063 15641 ne
rect 5063 15615 5165 15641
rect 5285 15641 5387 15735
tri 5387 15641 5485 15739 sw
tri 5485 15641 5583 15739 ne
rect 5583 15735 5937 15739
rect 5583 15641 5715 15735
rect 5285 15615 5485 15641
rect 5063 15611 5485 15615
tri 5485 15611 5515 15641 sw
tri 5583 15611 5613 15641 ne
rect 5613 15615 5715 15641
rect 5835 15641 5937 15735
tri 5937 15641 6035 15739 sw
tri 6035 15641 6133 15739 ne
rect 6133 15735 6487 15739
rect 6133 15641 6265 15735
rect 5835 15615 6035 15641
rect 5613 15611 6035 15615
tri 6035 15611 6065 15641 sw
tri 6133 15611 6163 15641 ne
rect 6163 15615 6265 15641
rect 6385 15641 6487 15735
tri 6487 15641 6585 15739 sw
tri 6585 15641 6683 15739 ne
rect 6683 15735 7037 15739
rect 6683 15641 6815 15735
rect 6385 15615 6585 15641
rect 6163 15611 6585 15615
tri 6585 15611 6615 15641 sw
tri 6683 15611 6713 15641 ne
rect 6713 15615 6815 15641
rect 6935 15641 7037 15735
tri 7037 15641 7135 15739 sw
tri 7135 15641 7233 15739 ne
rect 7233 15735 7587 15739
rect 7233 15641 7365 15735
rect 6935 15615 7135 15641
rect 6713 15611 7135 15615
tri 7135 15611 7165 15641 sw
tri 7233 15611 7263 15641 ne
rect 7263 15615 7365 15641
rect 7485 15641 7587 15735
tri 7587 15641 7685 15739 sw
tri 7685 15641 7783 15739 ne
rect 7783 15735 8137 15739
rect 7783 15641 7915 15735
rect 7485 15615 7685 15641
rect 7263 15611 7685 15615
tri 7685 15611 7715 15641 sw
tri 7783 15611 7813 15641 ne
rect 7813 15615 7915 15641
rect 8035 15641 8137 15735
tri 8137 15641 8235 15739 sw
tri 8235 15641 8333 15739 ne
rect 8333 15735 8687 15739
rect 8333 15641 8465 15735
rect 8035 15615 8235 15641
rect 7813 15611 8235 15615
tri 8235 15611 8265 15641 sw
tri 8333 15611 8363 15641 ne
rect 8363 15615 8465 15641
rect 8585 15641 8687 15735
tri 8687 15641 8785 15739 sw
tri 8785 15641 8883 15739 ne
rect 8883 15735 9237 15739
rect 8883 15641 9015 15735
rect 8585 15615 8785 15641
rect 8363 15611 8785 15615
tri 8785 15611 8815 15641 sw
tri 8883 15611 8913 15641 ne
rect 8913 15615 9015 15641
rect 9135 15641 9237 15735
tri 9237 15641 9335 15739 sw
tri 9335 15641 9433 15739 ne
rect 9433 15735 9787 15739
rect 9433 15641 9565 15735
rect 9135 15615 9335 15641
rect 8913 15611 9335 15615
tri 9335 15611 9365 15641 sw
tri 9433 15611 9463 15641 ne
rect 9463 15615 9565 15641
rect 9685 15641 9787 15735
tri 9787 15641 9885 15739 sw
tri 9885 15641 9983 15739 ne
rect 9983 15735 10337 15739
rect 9983 15641 10115 15735
rect 9685 15615 9885 15641
rect 9463 15611 9885 15615
tri 9885 15611 9915 15641 sw
tri 9983 15611 10013 15641 ne
rect 10013 15615 10115 15641
rect 10235 15641 10337 15735
tri 10337 15641 10435 15739 sw
tri 10435 15641 10533 15739 ne
rect 10533 15735 10887 15739
rect 10533 15641 10665 15735
rect 10235 15615 10435 15641
rect 10013 15611 10435 15615
tri 10435 15611 10465 15641 sw
tri 10533 15611 10563 15641 ne
rect 10563 15615 10665 15641
rect 10785 15641 10887 15735
tri 10887 15641 10985 15739 sw
tri 10985 15641 11083 15739 ne
rect 11083 15735 11437 15739
rect 11083 15641 11215 15735
rect 10785 15615 10985 15641
rect 10563 15611 10985 15615
tri 10985 15611 11015 15641 sw
tri 11083 15611 11113 15641 ne
rect 11113 15615 11215 15641
rect 11335 15641 11437 15735
tri 11437 15641 11535 15739 sw
tri 11535 15641 11633 15739 ne
rect 11633 15735 11987 15739
rect 11633 15641 11765 15735
rect 11335 15615 11535 15641
rect 11113 15611 11535 15615
tri 11535 15611 11565 15641 sw
tri 11633 15611 11663 15641 ne
rect 11663 15615 11765 15641
rect 11885 15641 11987 15735
tri 11987 15641 12085 15739 sw
tri 12085 15641 12183 15739 ne
rect 12183 15735 12537 15739
rect 12183 15641 12315 15735
rect 11885 15615 12085 15641
rect 11663 15611 12085 15615
tri 12085 15611 12115 15641 sw
tri 12183 15611 12213 15641 ne
rect 12213 15615 12315 15641
rect 12435 15641 12537 15735
tri 12537 15641 12635 15739 sw
tri 12635 15641 12733 15739 ne
rect 12733 15735 13087 15739
rect 12733 15641 12865 15735
rect 12435 15615 12635 15641
rect 12213 15611 12635 15615
tri 12635 15611 12665 15641 sw
tri 12733 15611 12763 15641 ne
rect 12763 15615 12865 15641
rect 12985 15641 13087 15735
tri 13087 15641 13185 15739 sw
tri 13185 15641 13283 15739 ne
rect 13283 15735 13637 15739
rect 13283 15641 13415 15735
rect 12985 15615 13185 15641
rect 12763 15611 13185 15615
tri 13185 15611 13215 15641 sw
tri 13283 15611 13313 15641 ne
rect 13313 15615 13415 15641
rect 13535 15641 13637 15735
tri 13637 15641 13735 15739 sw
tri 13735 15641 13833 15739 ne
rect 13833 15735 14187 15739
rect 13833 15641 13965 15735
rect 13535 15615 13735 15641
rect 13313 15611 13735 15615
tri 13735 15611 13765 15641 sw
tri 13833 15611 13863 15641 ne
rect 13863 15615 13965 15641
rect 14085 15641 14187 15735
tri 14187 15641 14285 15739 sw
tri 14285 15641 14383 15739 ne
rect 14383 15735 14737 15739
rect 14383 15641 14515 15735
rect 14085 15615 14285 15641
rect 13863 15611 14285 15615
tri 14285 15611 14315 15641 sw
tri 14383 15611 14413 15641 ne
rect 14413 15615 14515 15641
rect 14635 15641 14737 15735
tri 14737 15641 14835 15739 sw
tri 14835 15641 14933 15739 ne
rect 14933 15735 15287 15739
rect 14933 15641 15065 15735
rect 14635 15615 14835 15641
rect 14413 15611 14835 15615
tri 14835 15611 14865 15641 sw
tri 14933 15611 14963 15641 ne
rect 14963 15615 15065 15641
rect 15185 15641 15287 15735
tri 15287 15641 15385 15739 sw
tri 15385 15641 15483 15739 ne
rect 15483 15735 15837 15739
rect 15483 15641 15615 15735
rect 15185 15615 15385 15641
rect 14963 15611 15385 15615
tri 15385 15611 15415 15641 sw
tri 15483 15611 15513 15641 ne
rect 15513 15615 15615 15641
rect 15735 15641 15837 15735
tri 15837 15641 15935 15739 sw
tri 15935 15641 16033 15739 ne
rect 16033 15735 16387 15739
rect 16033 15641 16165 15735
rect 15735 15615 15935 15641
rect 15513 15611 15935 15615
tri 15935 15611 15965 15641 sw
tri 16033 15611 16063 15641 ne
rect 16063 15615 16165 15641
rect 16285 15641 16387 15735
tri 16387 15641 16485 15739 sw
tri 16485 15641 16583 15739 ne
rect 16583 15735 16937 15739
rect 16583 15641 16715 15735
rect 16285 15615 16485 15641
rect 16063 15611 16485 15615
tri 16485 15611 16515 15641 sw
tri 16583 15611 16613 15641 ne
rect 16613 15615 16715 15641
rect 16835 15641 16937 15735
tri 16937 15641 17035 15739 sw
tri 17035 15641 17133 15739 ne
rect 17133 15735 17487 15739
rect 17133 15641 17265 15735
rect 16835 15615 17035 15641
rect 16613 15611 17035 15615
tri 17035 15611 17065 15641 sw
tri 17133 15611 17163 15641 ne
rect 17163 15615 17265 15641
rect 17385 15641 17487 15735
tri 17487 15641 17585 15739 sw
tri 17585 15641 17683 15739 ne
rect 17683 15735 18037 15739
rect 17683 15641 17815 15735
rect 17385 15615 17585 15641
rect 17163 15611 17585 15615
tri 17585 15611 17615 15641 sw
tri 17683 15611 17713 15641 ne
rect 17713 15615 17815 15641
rect 17935 15641 18037 15735
tri 18037 15641 18135 15739 sw
tri 18135 15641 18233 15739 ne
rect 18233 15735 18587 15739
rect 18233 15641 18365 15735
rect 17935 15615 18135 15641
rect 17713 15611 18135 15615
tri 18135 15611 18165 15641 sw
tri 18233 15611 18263 15641 ne
rect 18263 15615 18365 15641
rect 18485 15641 18587 15735
tri 18587 15641 18685 15739 sw
tri 18685 15641 18783 15739 ne
rect 18783 15735 19137 15739
rect 18783 15641 18915 15735
rect 18485 15615 18685 15641
rect 18263 15611 18685 15615
tri 18685 15611 18715 15641 sw
tri 18783 15611 18813 15641 ne
rect 18813 15615 18915 15641
rect 19035 15641 19137 15735
tri 19137 15641 19235 15739 sw
tri 19235 15641 19333 15739 ne
rect 19333 15735 20300 15739
rect 19333 15641 19465 15735
rect 19035 15615 19235 15641
rect 18813 15611 19235 15615
tri 19235 15611 19265 15641 sw
tri 19333 15611 19363 15641 ne
rect 19363 15615 19465 15641
rect 19585 15615 20300 15735
rect 19363 15611 20300 15615
tri 113 15513 211 15611 ne
rect 211 15513 565 15611
tri 565 15513 663 15611 sw
tri 663 15513 761 15611 ne
rect 761 15513 1115 15611
tri 1115 15513 1213 15611 sw
tri 1213 15513 1311 15611 ne
rect 1311 15513 1665 15611
tri 1665 15513 1763 15611 sw
tri 1763 15513 1861 15611 ne
rect 1861 15513 2215 15611
tri 2215 15513 2313 15611 sw
tri 2313 15513 2411 15611 ne
rect 2411 15513 2765 15611
tri 2765 15513 2863 15611 sw
tri 2863 15513 2961 15611 ne
rect 2961 15513 3315 15611
tri 3315 15513 3413 15611 sw
tri 3413 15513 3511 15611 ne
rect 3511 15513 3865 15611
tri 3865 15513 3963 15611 sw
tri 3963 15513 4061 15611 ne
rect 4061 15513 4415 15611
tri 4415 15513 4513 15611 sw
tri 4513 15513 4611 15611 ne
rect 4611 15513 4965 15611
tri 4965 15513 5063 15611 sw
tri 5063 15513 5161 15611 ne
rect 5161 15513 5515 15611
tri 5515 15513 5613 15611 sw
tri 5613 15513 5711 15611 ne
rect 5711 15513 6065 15611
tri 6065 15513 6163 15611 sw
tri 6163 15513 6261 15611 ne
rect 6261 15513 6615 15611
tri 6615 15513 6713 15611 sw
tri 6713 15513 6811 15611 ne
rect 6811 15513 7165 15611
tri 7165 15513 7263 15611 sw
tri 7263 15513 7361 15611 ne
rect 7361 15513 7715 15611
tri 7715 15513 7813 15611 sw
tri 7813 15513 7911 15611 ne
rect 7911 15513 8265 15611
tri 8265 15513 8363 15611 sw
tri 8363 15513 8461 15611 ne
rect 8461 15513 8815 15611
tri 8815 15513 8913 15611 sw
tri 8913 15513 9011 15611 ne
rect 9011 15513 9365 15611
tri 9365 15513 9463 15611 sw
tri 9463 15513 9561 15611 ne
rect 9561 15513 9915 15611
tri 9915 15513 10013 15611 sw
tri 10013 15513 10111 15611 ne
rect 10111 15513 10465 15611
tri 10465 15513 10563 15611 sw
tri 10563 15513 10661 15611 ne
rect 10661 15513 11015 15611
tri 11015 15513 11113 15611 sw
tri 11113 15513 11211 15611 ne
rect 11211 15513 11565 15611
tri 11565 15513 11663 15611 sw
tri 11663 15513 11761 15611 ne
rect 11761 15513 12115 15611
tri 12115 15513 12213 15611 sw
tri 12213 15513 12311 15611 ne
rect 12311 15513 12665 15611
tri 12665 15513 12763 15611 sw
tri 12763 15513 12861 15611 ne
rect 12861 15513 13215 15611
tri 13215 15513 13313 15611 sw
tri 13313 15513 13411 15611 ne
rect 13411 15513 13765 15611
tri 13765 15513 13863 15611 sw
tri 13863 15513 13961 15611 ne
rect 13961 15513 14315 15611
tri 14315 15513 14413 15611 sw
tri 14413 15513 14511 15611 ne
rect 14511 15513 14865 15611
tri 14865 15513 14963 15611 sw
tri 14963 15513 15061 15611 ne
rect 15061 15513 15415 15611
tri 15415 15513 15513 15611 sw
tri 15513 15513 15611 15611 ne
rect 15611 15513 15965 15611
tri 15965 15513 16063 15611 sw
tri 16063 15513 16161 15611 ne
rect 16161 15513 16515 15611
tri 16515 15513 16613 15611 sw
tri 16613 15513 16711 15611 ne
rect 16711 15513 17065 15611
tri 17065 15513 17163 15611 sw
tri 17163 15513 17261 15611 ne
rect 17261 15513 17615 15611
tri 17615 15513 17713 15611 sw
tri 17713 15513 17811 15611 ne
rect 17811 15513 18165 15611
tri 18165 15513 18263 15611 sw
tri 18263 15513 18361 15611 ne
rect 18361 15513 18715 15611
tri 18715 15513 18813 15611 sw
tri 18813 15513 18911 15611 ne
rect 18911 15513 19265 15611
tri 19265 15513 19363 15611 sw
tri 19363 15513 19461 15611 ne
rect 19461 15513 20300 15611
rect -2000 15483 113 15513
tri 113 15483 143 15513 sw
tri 211 15483 241 15513 ne
rect 241 15483 663 15513
tri 663 15483 693 15513 sw
tri 761 15483 791 15513 ne
rect 791 15483 1213 15513
tri 1213 15483 1243 15513 sw
tri 1311 15483 1341 15513 ne
rect 1341 15483 1763 15513
tri 1763 15483 1793 15513 sw
tri 1861 15483 1891 15513 ne
rect 1891 15483 2313 15513
tri 2313 15483 2343 15513 sw
tri 2411 15483 2441 15513 ne
rect 2441 15483 2863 15513
tri 2863 15483 2893 15513 sw
tri 2961 15483 2991 15513 ne
rect 2991 15483 3413 15513
tri 3413 15483 3443 15513 sw
tri 3511 15483 3541 15513 ne
rect 3541 15483 3963 15513
tri 3963 15483 3993 15513 sw
tri 4061 15483 4091 15513 ne
rect 4091 15483 4513 15513
tri 4513 15483 4543 15513 sw
tri 4611 15483 4641 15513 ne
rect 4641 15483 5063 15513
tri 5063 15483 5093 15513 sw
tri 5161 15483 5191 15513 ne
rect 5191 15483 5613 15513
tri 5613 15483 5643 15513 sw
tri 5711 15483 5741 15513 ne
rect 5741 15483 6163 15513
tri 6163 15483 6193 15513 sw
tri 6261 15483 6291 15513 ne
rect 6291 15483 6713 15513
tri 6713 15483 6743 15513 sw
tri 6811 15483 6841 15513 ne
rect 6841 15483 7263 15513
tri 7263 15483 7293 15513 sw
tri 7361 15483 7391 15513 ne
rect 7391 15483 7813 15513
tri 7813 15483 7843 15513 sw
tri 7911 15483 7941 15513 ne
rect 7941 15483 8363 15513
tri 8363 15483 8393 15513 sw
tri 8461 15483 8491 15513 ne
rect 8491 15483 8913 15513
tri 8913 15483 8943 15513 sw
tri 9011 15483 9041 15513 ne
rect 9041 15483 9463 15513
tri 9463 15483 9493 15513 sw
tri 9561 15483 9591 15513 ne
rect 9591 15483 10013 15513
tri 10013 15483 10043 15513 sw
tri 10111 15483 10141 15513 ne
rect 10141 15483 10563 15513
tri 10563 15483 10593 15513 sw
tri 10661 15483 10691 15513 ne
rect 10691 15483 11113 15513
tri 11113 15483 11143 15513 sw
tri 11211 15483 11241 15513 ne
rect 11241 15483 11663 15513
tri 11663 15483 11693 15513 sw
tri 11761 15483 11791 15513 ne
rect 11791 15483 12213 15513
tri 12213 15483 12243 15513 sw
tri 12311 15483 12341 15513 ne
rect 12341 15483 12763 15513
tri 12763 15483 12793 15513 sw
tri 12861 15483 12891 15513 ne
rect 12891 15483 13313 15513
tri 13313 15483 13343 15513 sw
tri 13411 15483 13441 15513 ne
rect 13441 15483 13863 15513
tri 13863 15483 13893 15513 sw
tri 13961 15483 13991 15513 ne
rect 13991 15483 14413 15513
tri 14413 15483 14443 15513 sw
tri 14511 15483 14541 15513 ne
rect 14541 15483 14963 15513
tri 14963 15483 14993 15513 sw
tri 15061 15483 15091 15513 ne
rect 15091 15483 15513 15513
tri 15513 15483 15543 15513 sw
tri 15611 15483 15641 15513 ne
rect 15641 15483 16063 15513
tri 16063 15483 16093 15513 sw
tri 16161 15483 16191 15513 ne
rect 16191 15483 16613 15513
tri 16613 15483 16643 15513 sw
tri 16711 15483 16741 15513 ne
rect 16741 15483 17163 15513
tri 17163 15483 17193 15513 sw
tri 17261 15483 17291 15513 ne
rect 17291 15483 17713 15513
tri 17713 15483 17743 15513 sw
tri 17811 15483 17841 15513 ne
rect 17841 15483 18263 15513
tri 18263 15483 18293 15513 sw
tri 18361 15483 18391 15513 ne
rect 18391 15483 18813 15513
tri 18813 15483 18843 15513 sw
tri 18911 15483 18941 15513 ne
rect 18941 15483 19363 15513
tri 19363 15483 19393 15513 sw
tri 19461 15483 19491 15513 ne
rect 19491 15483 20300 15513
rect -2000 15385 143 15483
tri 143 15385 241 15483 sw
tri 241 15385 339 15483 ne
rect 339 15385 693 15483
tri 693 15385 791 15483 sw
tri 791 15385 889 15483 ne
rect 889 15385 1243 15483
tri 1243 15385 1341 15483 sw
tri 1341 15385 1439 15483 ne
rect 1439 15385 1793 15483
tri 1793 15385 1891 15483 sw
tri 1891 15385 1989 15483 ne
rect 1989 15385 2343 15483
tri 2343 15385 2441 15483 sw
tri 2441 15385 2539 15483 ne
rect 2539 15385 2893 15483
tri 2893 15385 2991 15483 sw
tri 2991 15385 3089 15483 ne
rect 3089 15385 3443 15483
tri 3443 15385 3541 15483 sw
tri 3541 15385 3639 15483 ne
rect 3639 15385 3993 15483
tri 3993 15385 4091 15483 sw
tri 4091 15385 4189 15483 ne
rect 4189 15385 4543 15483
tri 4543 15385 4641 15483 sw
tri 4641 15385 4739 15483 ne
rect 4739 15385 5093 15483
tri 5093 15385 5191 15483 sw
tri 5191 15385 5289 15483 ne
rect 5289 15385 5643 15483
tri 5643 15385 5741 15483 sw
tri 5741 15385 5839 15483 ne
rect 5839 15385 6193 15483
tri 6193 15385 6291 15483 sw
tri 6291 15385 6389 15483 ne
rect 6389 15385 6743 15483
tri 6743 15385 6841 15483 sw
tri 6841 15385 6939 15483 ne
rect 6939 15385 7293 15483
tri 7293 15385 7391 15483 sw
tri 7391 15385 7489 15483 ne
rect 7489 15385 7843 15483
tri 7843 15385 7941 15483 sw
tri 7941 15385 8039 15483 ne
rect 8039 15385 8393 15483
tri 8393 15385 8491 15483 sw
tri 8491 15385 8589 15483 ne
rect 8589 15385 8943 15483
tri 8943 15385 9041 15483 sw
tri 9041 15385 9139 15483 ne
rect 9139 15385 9493 15483
tri 9493 15385 9591 15483 sw
tri 9591 15385 9689 15483 ne
rect 9689 15385 10043 15483
tri 10043 15385 10141 15483 sw
tri 10141 15385 10239 15483 ne
rect 10239 15385 10593 15483
tri 10593 15385 10691 15483 sw
tri 10691 15385 10789 15483 ne
rect 10789 15385 11143 15483
tri 11143 15385 11241 15483 sw
tri 11241 15385 11339 15483 ne
rect 11339 15385 11693 15483
tri 11693 15385 11791 15483 sw
tri 11791 15385 11889 15483 ne
rect 11889 15385 12243 15483
tri 12243 15385 12341 15483 sw
tri 12341 15385 12439 15483 ne
rect 12439 15385 12793 15483
tri 12793 15385 12891 15483 sw
tri 12891 15385 12989 15483 ne
rect 12989 15385 13343 15483
tri 13343 15385 13441 15483 sw
tri 13441 15385 13539 15483 ne
rect 13539 15385 13893 15483
tri 13893 15385 13991 15483 sw
tri 13991 15385 14089 15483 ne
rect 14089 15385 14443 15483
tri 14443 15385 14541 15483 sw
tri 14541 15385 14639 15483 ne
rect 14639 15385 14993 15483
tri 14993 15385 15091 15483 sw
tri 15091 15385 15189 15483 ne
rect 15189 15385 15543 15483
tri 15543 15385 15641 15483 sw
tri 15641 15385 15739 15483 ne
rect 15739 15385 16093 15483
tri 16093 15385 16191 15483 sw
tri 16191 15385 16289 15483 ne
rect 16289 15385 16643 15483
tri 16643 15385 16741 15483 sw
tri 16741 15385 16839 15483 ne
rect 16839 15385 17193 15483
tri 17193 15385 17291 15483 sw
tri 17291 15385 17389 15483 ne
rect 17389 15385 17743 15483
tri 17743 15385 17841 15483 sw
tri 17841 15385 17939 15483 ne
rect 17939 15385 18293 15483
tri 18293 15385 18391 15483 sw
tri 18391 15385 18489 15483 ne
rect 18489 15385 18843 15483
tri 18843 15385 18941 15483 sw
tri 18941 15385 19039 15483 ne
rect 19039 15385 19393 15483
tri 19393 15385 19491 15483 sw
tri 19491 15385 19589 15483 ne
rect 19589 15385 20300 15483
rect -2000 15287 241 15385
tri 241 15287 339 15385 sw
tri 339 15287 437 15385 ne
rect 437 15287 791 15385
tri 791 15287 889 15385 sw
tri 889 15287 987 15385 ne
rect 987 15287 1341 15385
tri 1341 15287 1439 15385 sw
tri 1439 15287 1537 15385 ne
rect 1537 15287 1891 15385
tri 1891 15287 1989 15385 sw
tri 1989 15287 2087 15385 ne
rect 2087 15287 2441 15385
tri 2441 15287 2539 15385 sw
tri 2539 15287 2637 15385 ne
rect 2637 15287 2991 15385
tri 2991 15287 3089 15385 sw
tri 3089 15287 3187 15385 ne
rect 3187 15287 3541 15385
tri 3541 15287 3639 15385 sw
tri 3639 15287 3737 15385 ne
rect 3737 15287 4091 15385
tri 4091 15287 4189 15385 sw
tri 4189 15287 4287 15385 ne
rect 4287 15287 4641 15385
tri 4641 15287 4739 15385 sw
tri 4739 15287 4837 15385 ne
rect 4837 15287 5191 15385
tri 5191 15287 5289 15385 sw
tri 5289 15287 5387 15385 ne
rect 5387 15287 5741 15385
tri 5741 15287 5839 15385 sw
tri 5839 15287 5937 15385 ne
rect 5937 15287 6291 15385
tri 6291 15287 6389 15385 sw
tri 6389 15287 6487 15385 ne
rect 6487 15287 6841 15385
tri 6841 15287 6939 15385 sw
tri 6939 15287 7037 15385 ne
rect 7037 15287 7391 15385
tri 7391 15287 7489 15385 sw
tri 7489 15287 7587 15385 ne
rect 7587 15287 7941 15385
tri 7941 15287 8039 15385 sw
tri 8039 15287 8137 15385 ne
rect 8137 15287 8491 15385
tri 8491 15287 8589 15385 sw
tri 8589 15287 8687 15385 ne
rect 8687 15287 9041 15385
tri 9041 15287 9139 15385 sw
tri 9139 15287 9237 15385 ne
rect 9237 15287 9591 15385
tri 9591 15287 9689 15385 sw
tri 9689 15287 9787 15385 ne
rect 9787 15287 10141 15385
tri 10141 15287 10239 15385 sw
tri 10239 15287 10337 15385 ne
rect 10337 15287 10691 15385
tri 10691 15287 10789 15385 sw
tri 10789 15287 10887 15385 ne
rect 10887 15287 11241 15385
tri 11241 15287 11339 15385 sw
tri 11339 15287 11437 15385 ne
rect 11437 15287 11791 15385
tri 11791 15287 11889 15385 sw
tri 11889 15287 11987 15385 ne
rect 11987 15287 12341 15385
tri 12341 15287 12439 15385 sw
tri 12439 15287 12537 15385 ne
rect 12537 15287 12891 15385
tri 12891 15287 12989 15385 sw
tri 12989 15287 13087 15385 ne
rect 13087 15287 13441 15385
tri 13441 15287 13539 15385 sw
tri 13539 15287 13637 15385 ne
rect 13637 15287 13991 15385
tri 13991 15287 14089 15385 sw
tri 14089 15287 14187 15385 ne
rect 14187 15287 14541 15385
tri 14541 15287 14639 15385 sw
tri 14639 15287 14737 15385 ne
rect 14737 15287 15091 15385
tri 15091 15287 15189 15385 sw
tri 15189 15287 15287 15385 ne
rect 15287 15287 15641 15385
tri 15641 15287 15739 15385 sw
tri 15739 15287 15837 15385 ne
rect 15837 15287 16191 15385
tri 16191 15287 16289 15385 sw
tri 16289 15287 16387 15385 ne
rect 16387 15287 16741 15385
tri 16741 15287 16839 15385 sw
tri 16839 15287 16937 15385 ne
rect 16937 15287 17291 15385
tri 17291 15287 17389 15385 sw
tri 17389 15287 17487 15385 ne
rect 17487 15287 17841 15385
tri 17841 15287 17939 15385 sw
tri 17939 15287 18037 15385 ne
rect 18037 15287 18391 15385
tri 18391 15287 18489 15385 sw
tri 18489 15287 18587 15385 ne
rect 18587 15287 18941 15385
tri 18941 15287 19039 15385 sw
tri 19039 15287 19137 15385 ne
rect 19137 15287 19491 15385
tri 19491 15287 19589 15385 sw
tri 19589 15287 19687 15385 ne
rect 19687 15287 20300 15385
rect -2000 15189 339 15287
tri 339 15189 437 15287 sw
tri 437 15189 535 15287 ne
rect 535 15189 889 15287
tri 889 15189 987 15287 sw
tri 987 15189 1085 15287 ne
rect 1085 15189 1439 15287
tri 1439 15189 1537 15287 sw
tri 1537 15189 1635 15287 ne
rect 1635 15189 1989 15287
tri 1989 15189 2087 15287 sw
tri 2087 15189 2185 15287 ne
rect 2185 15189 2539 15287
tri 2539 15189 2637 15287 sw
tri 2637 15189 2735 15287 ne
rect 2735 15189 3089 15287
tri 3089 15189 3187 15287 sw
tri 3187 15189 3285 15287 ne
rect 3285 15189 3639 15287
tri 3639 15189 3737 15287 sw
tri 3737 15189 3835 15287 ne
rect 3835 15189 4189 15287
tri 4189 15189 4287 15287 sw
tri 4287 15189 4385 15287 ne
rect 4385 15189 4739 15287
tri 4739 15189 4837 15287 sw
tri 4837 15189 4935 15287 ne
rect 4935 15189 5289 15287
tri 5289 15189 5387 15287 sw
tri 5387 15189 5485 15287 ne
rect 5485 15189 5839 15287
tri 5839 15189 5937 15287 sw
tri 5937 15189 6035 15287 ne
rect 6035 15189 6389 15287
tri 6389 15189 6487 15287 sw
tri 6487 15189 6585 15287 ne
rect 6585 15189 6939 15287
tri 6939 15189 7037 15287 sw
tri 7037 15189 7135 15287 ne
rect 7135 15189 7489 15287
tri 7489 15189 7587 15287 sw
tri 7587 15189 7685 15287 ne
rect 7685 15189 8039 15287
tri 8039 15189 8137 15287 sw
tri 8137 15189 8235 15287 ne
rect 8235 15189 8589 15287
tri 8589 15189 8687 15287 sw
tri 8687 15189 8785 15287 ne
rect 8785 15189 9139 15287
tri 9139 15189 9237 15287 sw
tri 9237 15189 9335 15287 ne
rect 9335 15189 9689 15287
tri 9689 15189 9787 15287 sw
tri 9787 15189 9885 15287 ne
rect 9885 15189 10239 15287
tri 10239 15189 10337 15287 sw
tri 10337 15189 10435 15287 ne
rect 10435 15189 10789 15287
tri 10789 15189 10887 15287 sw
tri 10887 15189 10985 15287 ne
rect 10985 15189 11339 15287
tri 11339 15189 11437 15287 sw
tri 11437 15189 11535 15287 ne
rect 11535 15189 11889 15287
tri 11889 15189 11987 15287 sw
tri 11987 15189 12085 15287 ne
rect 12085 15189 12439 15287
tri 12439 15189 12537 15287 sw
tri 12537 15189 12635 15287 ne
rect 12635 15189 12989 15287
tri 12989 15189 13087 15287 sw
tri 13087 15189 13185 15287 ne
rect 13185 15189 13539 15287
tri 13539 15189 13637 15287 sw
tri 13637 15189 13735 15287 ne
rect 13735 15189 14089 15287
tri 14089 15189 14187 15287 sw
tri 14187 15189 14285 15287 ne
rect 14285 15189 14639 15287
tri 14639 15189 14737 15287 sw
tri 14737 15189 14835 15287 ne
rect 14835 15189 15189 15287
tri 15189 15189 15287 15287 sw
tri 15287 15189 15385 15287 ne
rect 15385 15189 15739 15287
tri 15739 15189 15837 15287 sw
tri 15837 15189 15935 15287 ne
rect 15935 15189 16289 15287
tri 16289 15189 16387 15287 sw
tri 16387 15189 16485 15287 ne
rect 16485 15189 16839 15287
tri 16839 15189 16937 15287 sw
tri 16937 15189 17035 15287 ne
rect 17035 15189 17389 15287
tri 17389 15189 17487 15287 sw
tri 17487 15189 17585 15287 ne
rect 17585 15189 17939 15287
tri 17939 15189 18037 15287 sw
tri 18037 15189 18135 15287 ne
rect 18135 15189 18489 15287
tri 18489 15189 18587 15287 sw
tri 18587 15189 18685 15287 ne
rect 18685 15189 19039 15287
tri 19039 15189 19137 15287 sw
tri 19137 15189 19235 15287 ne
rect 19235 15189 19589 15287
tri 19589 15189 19687 15287 sw
rect 20800 15189 21800 15837
rect -2000 15185 437 15189
rect -2000 15065 215 15185
rect 335 15091 437 15185
tri 437 15091 535 15189 sw
tri 535 15091 633 15189 ne
rect 633 15185 987 15189
rect 633 15091 765 15185
rect 335 15065 535 15091
rect -2000 15061 535 15065
rect -2000 14413 -1000 15061
tri 113 14963 211 15061 ne
rect 211 15013 535 15061
tri 535 15013 613 15091 sw
tri 633 15013 711 15091 ne
rect 711 15065 765 15091
rect 885 15091 987 15185
tri 987 15091 1085 15189 sw
tri 1085 15091 1183 15189 ne
rect 1183 15185 1537 15189
rect 1183 15091 1315 15185
rect 885 15065 1085 15091
rect 711 15013 1085 15065
tri 1085 15013 1163 15091 sw
tri 1183 15013 1261 15091 ne
rect 1261 15065 1315 15091
rect 1435 15091 1537 15185
tri 1537 15091 1635 15189 sw
tri 1635 15091 1733 15189 ne
rect 1733 15185 2087 15189
rect 1733 15091 1865 15185
rect 1435 15065 1635 15091
rect 1261 15013 1635 15065
tri 1635 15013 1713 15091 sw
tri 1733 15013 1811 15091 ne
rect 1811 15065 1865 15091
rect 1985 15091 2087 15185
tri 2087 15091 2185 15189 sw
tri 2185 15091 2283 15189 ne
rect 2283 15185 2637 15189
rect 2283 15091 2415 15185
rect 1985 15065 2185 15091
rect 1811 15013 2185 15065
tri 2185 15013 2263 15091 sw
tri 2283 15013 2361 15091 ne
rect 2361 15065 2415 15091
rect 2535 15091 2637 15185
tri 2637 15091 2735 15189 sw
tri 2735 15091 2833 15189 ne
rect 2833 15185 3187 15189
rect 2833 15091 2965 15185
rect 2535 15065 2735 15091
rect 2361 15013 2735 15065
tri 2735 15013 2813 15091 sw
tri 2833 15013 2911 15091 ne
rect 2911 15065 2965 15091
rect 3085 15091 3187 15185
tri 3187 15091 3285 15189 sw
tri 3285 15091 3383 15189 ne
rect 3383 15185 3737 15189
rect 3383 15091 3515 15185
rect 3085 15065 3285 15091
rect 2911 15013 3285 15065
tri 3285 15013 3363 15091 sw
tri 3383 15013 3461 15091 ne
rect 3461 15065 3515 15091
rect 3635 15091 3737 15185
tri 3737 15091 3835 15189 sw
tri 3835 15091 3933 15189 ne
rect 3933 15185 4287 15189
rect 3933 15091 4065 15185
rect 3635 15065 3835 15091
rect 3461 15013 3835 15065
tri 3835 15013 3913 15091 sw
tri 3933 15013 4011 15091 ne
rect 4011 15065 4065 15091
rect 4185 15091 4287 15185
tri 4287 15091 4385 15189 sw
tri 4385 15091 4483 15189 ne
rect 4483 15185 4837 15189
rect 4483 15091 4615 15185
rect 4185 15065 4385 15091
rect 4011 15013 4385 15065
tri 4385 15013 4463 15091 sw
tri 4483 15013 4561 15091 ne
rect 4561 15065 4615 15091
rect 4735 15091 4837 15185
tri 4837 15091 4935 15189 sw
tri 4935 15091 5033 15189 ne
rect 5033 15185 5387 15189
rect 5033 15091 5165 15185
rect 4735 15065 4935 15091
rect 4561 15013 4935 15065
tri 4935 15013 5013 15091 sw
tri 5033 15013 5111 15091 ne
rect 5111 15065 5165 15091
rect 5285 15091 5387 15185
tri 5387 15091 5485 15189 sw
tri 5485 15091 5583 15189 ne
rect 5583 15185 5937 15189
rect 5583 15091 5715 15185
rect 5285 15065 5485 15091
rect 5111 15013 5485 15065
tri 5485 15013 5563 15091 sw
tri 5583 15013 5661 15091 ne
rect 5661 15065 5715 15091
rect 5835 15091 5937 15185
tri 5937 15091 6035 15189 sw
tri 6035 15091 6133 15189 ne
rect 6133 15185 6487 15189
rect 6133 15091 6265 15185
rect 5835 15065 6035 15091
rect 5661 15013 6035 15065
tri 6035 15013 6113 15091 sw
tri 6133 15013 6211 15091 ne
rect 6211 15065 6265 15091
rect 6385 15091 6487 15185
tri 6487 15091 6585 15189 sw
tri 6585 15091 6683 15189 ne
rect 6683 15185 7037 15189
rect 6683 15091 6815 15185
rect 6385 15065 6585 15091
rect 6211 15013 6585 15065
tri 6585 15013 6663 15091 sw
tri 6683 15013 6761 15091 ne
rect 6761 15065 6815 15091
rect 6935 15091 7037 15185
tri 7037 15091 7135 15189 sw
tri 7135 15091 7233 15189 ne
rect 7233 15185 7587 15189
rect 7233 15091 7365 15185
rect 6935 15065 7135 15091
rect 6761 15013 7135 15065
tri 7135 15013 7213 15091 sw
tri 7233 15013 7311 15091 ne
rect 7311 15065 7365 15091
rect 7485 15091 7587 15185
tri 7587 15091 7685 15189 sw
tri 7685 15091 7783 15189 ne
rect 7783 15185 8137 15189
rect 7783 15091 7915 15185
rect 7485 15065 7685 15091
rect 7311 15013 7685 15065
tri 7685 15013 7763 15091 sw
tri 7783 15013 7861 15091 ne
rect 7861 15065 7915 15091
rect 8035 15091 8137 15185
tri 8137 15091 8235 15189 sw
tri 8235 15091 8333 15189 ne
rect 8333 15185 8687 15189
rect 8333 15091 8465 15185
rect 8035 15065 8235 15091
rect 7861 15013 8235 15065
tri 8235 15013 8313 15091 sw
tri 8333 15013 8411 15091 ne
rect 8411 15065 8465 15091
rect 8585 15091 8687 15185
tri 8687 15091 8785 15189 sw
tri 8785 15091 8883 15189 ne
rect 8883 15185 9237 15189
rect 8883 15091 9015 15185
rect 8585 15065 8785 15091
rect 8411 15013 8785 15065
tri 8785 15013 8863 15091 sw
tri 8883 15013 8961 15091 ne
rect 8961 15065 9015 15091
rect 9135 15091 9237 15185
tri 9237 15091 9335 15189 sw
tri 9335 15091 9433 15189 ne
rect 9433 15185 9787 15189
rect 9433 15091 9565 15185
rect 9135 15065 9335 15091
rect 8961 15013 9335 15065
tri 9335 15013 9413 15091 sw
tri 9433 15013 9511 15091 ne
rect 9511 15065 9565 15091
rect 9685 15091 9787 15185
tri 9787 15091 9885 15189 sw
tri 9885 15091 9983 15189 ne
rect 9983 15185 10337 15189
rect 9983 15091 10115 15185
rect 9685 15065 9885 15091
rect 9511 15013 9885 15065
tri 9885 15013 9963 15091 sw
tri 9983 15013 10061 15091 ne
rect 10061 15065 10115 15091
rect 10235 15091 10337 15185
tri 10337 15091 10435 15189 sw
tri 10435 15091 10533 15189 ne
rect 10533 15185 10887 15189
rect 10533 15091 10665 15185
rect 10235 15065 10435 15091
rect 10061 15013 10435 15065
tri 10435 15013 10513 15091 sw
tri 10533 15013 10611 15091 ne
rect 10611 15065 10665 15091
rect 10785 15091 10887 15185
tri 10887 15091 10985 15189 sw
tri 10985 15091 11083 15189 ne
rect 11083 15185 11437 15189
rect 11083 15091 11215 15185
rect 10785 15065 10985 15091
rect 10611 15013 10985 15065
tri 10985 15013 11063 15091 sw
tri 11083 15013 11161 15091 ne
rect 11161 15065 11215 15091
rect 11335 15091 11437 15185
tri 11437 15091 11535 15189 sw
tri 11535 15091 11633 15189 ne
rect 11633 15185 11987 15189
rect 11633 15091 11765 15185
rect 11335 15065 11535 15091
rect 11161 15013 11535 15065
tri 11535 15013 11613 15091 sw
tri 11633 15013 11711 15091 ne
rect 11711 15065 11765 15091
rect 11885 15091 11987 15185
tri 11987 15091 12085 15189 sw
tri 12085 15091 12183 15189 ne
rect 12183 15185 12537 15189
rect 12183 15091 12315 15185
rect 11885 15065 12085 15091
rect 11711 15013 12085 15065
tri 12085 15013 12163 15091 sw
tri 12183 15013 12261 15091 ne
rect 12261 15065 12315 15091
rect 12435 15091 12537 15185
tri 12537 15091 12635 15189 sw
tri 12635 15091 12733 15189 ne
rect 12733 15185 13087 15189
rect 12733 15091 12865 15185
rect 12435 15065 12635 15091
rect 12261 15013 12635 15065
tri 12635 15013 12713 15091 sw
tri 12733 15013 12811 15091 ne
rect 12811 15065 12865 15091
rect 12985 15091 13087 15185
tri 13087 15091 13185 15189 sw
tri 13185 15091 13283 15189 ne
rect 13283 15185 13637 15189
rect 13283 15091 13415 15185
rect 12985 15065 13185 15091
rect 12811 15013 13185 15065
tri 13185 15013 13263 15091 sw
tri 13283 15013 13361 15091 ne
rect 13361 15065 13415 15091
rect 13535 15091 13637 15185
tri 13637 15091 13735 15189 sw
tri 13735 15091 13833 15189 ne
rect 13833 15185 14187 15189
rect 13833 15091 13965 15185
rect 13535 15065 13735 15091
rect 13361 15013 13735 15065
tri 13735 15013 13813 15091 sw
tri 13833 15013 13911 15091 ne
rect 13911 15065 13965 15091
rect 14085 15091 14187 15185
tri 14187 15091 14285 15189 sw
tri 14285 15091 14383 15189 ne
rect 14383 15185 14737 15189
rect 14383 15091 14515 15185
rect 14085 15065 14285 15091
rect 13911 15013 14285 15065
tri 14285 15013 14363 15091 sw
tri 14383 15013 14461 15091 ne
rect 14461 15065 14515 15091
rect 14635 15091 14737 15185
tri 14737 15091 14835 15189 sw
tri 14835 15091 14933 15189 ne
rect 14933 15185 15287 15189
rect 14933 15091 15065 15185
rect 14635 15065 14835 15091
rect 14461 15013 14835 15065
tri 14835 15013 14913 15091 sw
tri 14933 15013 15011 15091 ne
rect 15011 15065 15065 15091
rect 15185 15091 15287 15185
tri 15287 15091 15385 15189 sw
tri 15385 15091 15483 15189 ne
rect 15483 15185 15837 15189
rect 15483 15091 15615 15185
rect 15185 15065 15385 15091
rect 15011 15013 15385 15065
tri 15385 15013 15463 15091 sw
tri 15483 15013 15561 15091 ne
rect 15561 15065 15615 15091
rect 15735 15091 15837 15185
tri 15837 15091 15935 15189 sw
tri 15935 15091 16033 15189 ne
rect 16033 15185 16387 15189
rect 16033 15091 16165 15185
rect 15735 15065 15935 15091
rect 15561 15013 15935 15065
tri 15935 15013 16013 15091 sw
tri 16033 15013 16111 15091 ne
rect 16111 15065 16165 15091
rect 16285 15091 16387 15185
tri 16387 15091 16485 15189 sw
tri 16485 15091 16583 15189 ne
rect 16583 15185 16937 15189
rect 16583 15091 16715 15185
rect 16285 15065 16485 15091
rect 16111 15013 16485 15065
tri 16485 15013 16563 15091 sw
tri 16583 15013 16661 15091 ne
rect 16661 15065 16715 15091
rect 16835 15091 16937 15185
tri 16937 15091 17035 15189 sw
tri 17035 15091 17133 15189 ne
rect 17133 15185 17487 15189
rect 17133 15091 17265 15185
rect 16835 15065 17035 15091
rect 16661 15013 17035 15065
tri 17035 15013 17113 15091 sw
tri 17133 15013 17211 15091 ne
rect 17211 15065 17265 15091
rect 17385 15091 17487 15185
tri 17487 15091 17585 15189 sw
tri 17585 15091 17683 15189 ne
rect 17683 15185 18037 15189
rect 17683 15091 17815 15185
rect 17385 15065 17585 15091
rect 17211 15013 17585 15065
tri 17585 15013 17663 15091 sw
tri 17683 15013 17761 15091 ne
rect 17761 15065 17815 15091
rect 17935 15091 18037 15185
tri 18037 15091 18135 15189 sw
tri 18135 15091 18233 15189 ne
rect 18233 15185 18587 15189
rect 18233 15091 18365 15185
rect 17935 15065 18135 15091
rect 17761 15013 18135 15065
tri 18135 15013 18213 15091 sw
tri 18233 15013 18311 15091 ne
rect 18311 15065 18365 15091
rect 18485 15091 18587 15185
tri 18587 15091 18685 15189 sw
tri 18685 15091 18783 15189 ne
rect 18783 15185 19137 15189
rect 18783 15091 18915 15185
rect 18485 15065 18685 15091
rect 18311 15013 18685 15065
tri 18685 15013 18763 15091 sw
tri 18783 15013 18861 15091 ne
rect 18861 15065 18915 15091
rect 19035 15091 19137 15185
tri 19137 15091 19235 15189 sw
tri 19235 15091 19333 15189 ne
rect 19333 15185 21800 15189
rect 19333 15091 19465 15185
rect 19035 15065 19235 15091
rect 18861 15013 19235 15065
tri 19235 15013 19313 15091 sw
tri 19333 15013 19411 15091 ne
rect 19411 15065 19465 15091
rect 19585 15065 21800 15185
rect 19411 15013 21800 15065
rect 211 14963 613 15013
rect -500 14913 113 14963
tri 113 14913 163 14963 sw
tri 211 14913 261 14963 ne
rect 261 14933 613 14963
tri 613 14933 693 15013 sw
tri 711 14933 791 15013 ne
rect 791 14933 1163 15013
tri 1163 14933 1243 15013 sw
tri 1261 14933 1341 15013 ne
rect 1341 14933 1713 15013
tri 1713 14933 1793 15013 sw
tri 1811 14933 1891 15013 ne
rect 1891 14933 2263 15013
tri 2263 14933 2343 15013 sw
tri 2361 14933 2441 15013 ne
rect 2441 14933 2813 15013
tri 2813 14933 2893 15013 sw
tri 2911 14933 2991 15013 ne
rect 2991 14933 3363 15013
tri 3363 14933 3443 15013 sw
tri 3461 14933 3541 15013 ne
rect 3541 14933 3913 15013
tri 3913 14933 3993 15013 sw
tri 4011 14933 4091 15013 ne
rect 4091 14933 4463 15013
tri 4463 14933 4543 15013 sw
tri 4561 14933 4641 15013 ne
rect 4641 14933 5013 15013
tri 5013 14933 5093 15013 sw
tri 5111 14933 5191 15013 ne
rect 5191 14933 5563 15013
tri 5563 14933 5643 15013 sw
tri 5661 14933 5741 15013 ne
rect 5741 14933 6113 15013
tri 6113 14933 6193 15013 sw
tri 6211 14933 6291 15013 ne
rect 6291 14933 6663 15013
tri 6663 14933 6743 15013 sw
tri 6761 14933 6841 15013 ne
rect 6841 14933 7213 15013
tri 7213 14933 7293 15013 sw
tri 7311 14933 7391 15013 ne
rect 7391 14933 7763 15013
tri 7763 14933 7843 15013 sw
tri 7861 14933 7941 15013 ne
rect 7941 14933 8313 15013
tri 8313 14933 8393 15013 sw
tri 8411 14933 8491 15013 ne
rect 8491 14933 8863 15013
tri 8863 14933 8943 15013 sw
tri 8961 14933 9041 15013 ne
rect 9041 14933 9413 15013
tri 9413 14933 9493 15013 sw
tri 9511 14933 9591 15013 ne
rect 9591 14933 9963 15013
tri 9963 14933 10043 15013 sw
tri 10061 14933 10141 15013 ne
rect 10141 14933 10513 15013
tri 10513 14933 10593 15013 sw
tri 10611 14933 10691 15013 ne
rect 10691 14933 11063 15013
tri 11063 14933 11143 15013 sw
tri 11161 14933 11241 15013 ne
rect 11241 14933 11613 15013
tri 11613 14933 11693 15013 sw
tri 11711 14933 11791 15013 ne
rect 11791 14933 12163 15013
tri 12163 14933 12243 15013 sw
tri 12261 14933 12341 15013 ne
rect 12341 14933 12713 15013
tri 12713 14933 12793 15013 sw
tri 12811 14933 12891 15013 ne
rect 12891 14933 13263 15013
tri 13263 14933 13343 15013 sw
tri 13361 14933 13441 15013 ne
rect 13441 14933 13813 15013
tri 13813 14933 13893 15013 sw
tri 13911 14933 13991 15013 ne
rect 13991 14933 14363 15013
tri 14363 14933 14443 15013 sw
tri 14461 14933 14541 15013 ne
rect 14541 14933 14913 15013
tri 14913 14933 14993 15013 sw
tri 15011 14933 15091 15013 ne
rect 15091 14933 15463 15013
tri 15463 14933 15543 15013 sw
tri 15561 14933 15641 15013 ne
rect 15641 14933 16013 15013
tri 16013 14933 16093 15013 sw
tri 16111 14933 16191 15013 ne
rect 16191 14933 16563 15013
tri 16563 14933 16643 15013 sw
tri 16661 14933 16741 15013 ne
rect 16741 14933 17113 15013
tri 17113 14933 17193 15013 sw
tri 17211 14933 17291 15013 ne
rect 17291 14933 17663 15013
tri 17663 14933 17743 15013 sw
tri 17761 14933 17841 15013 ne
rect 17841 14933 18213 15013
tri 18213 14933 18293 15013 sw
tri 18311 14933 18391 15013 ne
rect 18391 14933 18763 15013
tri 18763 14933 18843 15013 sw
tri 18861 14933 18941 15013 ne
rect 18941 14933 19313 15013
tri 19313 14933 19393 15013 sw
tri 19411 14933 19491 15013 ne
rect 19491 14933 20100 15013
rect 261 14913 693 14933
rect -500 14835 163 14913
tri 163 14835 241 14913 sw
tri 261 14835 339 14913 ne
rect 339 14835 693 14913
tri 693 14835 791 14933 sw
tri 791 14835 889 14933 ne
rect 889 14835 1243 14933
tri 1243 14835 1341 14933 sw
tri 1341 14835 1439 14933 ne
rect 1439 14835 1793 14933
tri 1793 14835 1891 14933 sw
tri 1891 14835 1989 14933 ne
rect 1989 14835 2343 14933
tri 2343 14835 2441 14933 sw
tri 2441 14835 2539 14933 ne
rect 2539 14835 2893 14933
tri 2893 14835 2991 14933 sw
tri 2991 14835 3089 14933 ne
rect 3089 14835 3443 14933
tri 3443 14835 3541 14933 sw
tri 3541 14835 3639 14933 ne
rect 3639 14835 3993 14933
tri 3993 14835 4091 14933 sw
tri 4091 14835 4189 14933 ne
rect 4189 14835 4543 14933
tri 4543 14835 4641 14933 sw
tri 4641 14835 4739 14933 ne
rect 4739 14835 5093 14933
tri 5093 14835 5191 14933 sw
tri 5191 14835 5289 14933 ne
rect 5289 14835 5643 14933
tri 5643 14835 5741 14933 sw
tri 5741 14835 5839 14933 ne
rect 5839 14835 6193 14933
tri 6193 14835 6291 14933 sw
tri 6291 14835 6389 14933 ne
rect 6389 14835 6743 14933
tri 6743 14835 6841 14933 sw
tri 6841 14835 6939 14933 ne
rect 6939 14835 7293 14933
tri 7293 14835 7391 14933 sw
tri 7391 14835 7489 14933 ne
rect 7489 14835 7843 14933
tri 7843 14835 7941 14933 sw
tri 7941 14835 8039 14933 ne
rect 8039 14835 8393 14933
tri 8393 14835 8491 14933 sw
tri 8491 14835 8589 14933 ne
rect 8589 14835 8943 14933
tri 8943 14835 9041 14933 sw
tri 9041 14835 9139 14933 ne
rect 9139 14835 9493 14933
tri 9493 14835 9591 14933 sw
tri 9591 14835 9689 14933 ne
rect 9689 14835 10043 14933
tri 10043 14835 10141 14933 sw
tri 10141 14835 10239 14933 ne
rect 10239 14835 10593 14933
tri 10593 14835 10691 14933 sw
tri 10691 14835 10789 14933 ne
rect 10789 14835 11143 14933
tri 11143 14835 11241 14933 sw
tri 11241 14835 11339 14933 ne
rect 11339 14835 11693 14933
tri 11693 14835 11791 14933 sw
tri 11791 14835 11889 14933 ne
rect 11889 14835 12243 14933
tri 12243 14835 12341 14933 sw
tri 12341 14835 12439 14933 ne
rect 12439 14835 12793 14933
tri 12793 14835 12891 14933 sw
tri 12891 14835 12989 14933 ne
rect 12989 14835 13343 14933
tri 13343 14835 13441 14933 sw
tri 13441 14835 13539 14933 ne
rect 13539 14835 13893 14933
tri 13893 14835 13991 14933 sw
tri 13991 14835 14089 14933 ne
rect 14089 14835 14443 14933
tri 14443 14835 14541 14933 sw
tri 14541 14835 14639 14933 ne
rect 14639 14835 14993 14933
tri 14993 14835 15091 14933 sw
tri 15091 14835 15189 14933 ne
rect 15189 14835 15543 14933
tri 15543 14835 15641 14933 sw
tri 15641 14835 15739 14933 ne
rect 15739 14835 16093 14933
tri 16093 14835 16191 14933 sw
tri 16191 14835 16289 14933 ne
rect 16289 14835 16643 14933
tri 16643 14835 16741 14933 sw
tri 16741 14835 16839 14933 ne
rect 16839 14835 17193 14933
tri 17193 14835 17291 14933 sw
tri 17291 14835 17389 14933 ne
rect 17389 14835 17743 14933
tri 17743 14835 17841 14933 sw
tri 17841 14835 17939 14933 ne
rect 17939 14835 18293 14933
tri 18293 14835 18391 14933 sw
tri 18391 14835 18489 14933 ne
rect 18489 14835 18843 14933
tri 18843 14835 18941 14933 sw
tri 18941 14835 19039 14933 ne
rect 19039 14835 19393 14933
tri 19393 14835 19491 14933 sw
tri 19491 14835 19589 14933 ne
rect 19589 14913 20100 14933
rect 20200 14913 21800 15013
rect 19589 14835 21800 14913
rect -500 14787 241 14835
rect -500 14687 -400 14787
rect -300 14737 241 14787
tri 241 14737 339 14835 sw
tri 339 14737 437 14835 ne
rect 437 14737 791 14835
tri 791 14737 889 14835 sw
tri 889 14737 987 14835 ne
rect 987 14737 1341 14835
tri 1341 14737 1439 14835 sw
tri 1439 14737 1537 14835 ne
rect 1537 14737 1891 14835
tri 1891 14737 1989 14835 sw
tri 1989 14737 2087 14835 ne
rect 2087 14737 2441 14835
tri 2441 14737 2539 14835 sw
tri 2539 14737 2637 14835 ne
rect 2637 14737 2991 14835
tri 2991 14737 3089 14835 sw
tri 3089 14737 3187 14835 ne
rect 3187 14737 3541 14835
tri 3541 14737 3639 14835 sw
tri 3639 14737 3737 14835 ne
rect 3737 14737 4091 14835
tri 4091 14737 4189 14835 sw
tri 4189 14737 4287 14835 ne
rect 4287 14737 4641 14835
tri 4641 14737 4739 14835 sw
tri 4739 14737 4837 14835 ne
rect 4837 14737 5191 14835
tri 5191 14737 5289 14835 sw
tri 5289 14737 5387 14835 ne
rect 5387 14737 5741 14835
tri 5741 14737 5839 14835 sw
tri 5839 14737 5937 14835 ne
rect 5937 14737 6291 14835
tri 6291 14737 6389 14835 sw
tri 6389 14737 6487 14835 ne
rect 6487 14737 6841 14835
tri 6841 14737 6939 14835 sw
tri 6939 14737 7037 14835 ne
rect 7037 14737 7391 14835
tri 7391 14737 7489 14835 sw
tri 7489 14737 7587 14835 ne
rect 7587 14737 7941 14835
tri 7941 14737 8039 14835 sw
tri 8039 14737 8137 14835 ne
rect 8137 14737 8491 14835
tri 8491 14737 8589 14835 sw
tri 8589 14737 8687 14835 ne
rect 8687 14737 9041 14835
tri 9041 14737 9139 14835 sw
tri 9139 14737 9237 14835 ne
rect 9237 14737 9591 14835
tri 9591 14737 9689 14835 sw
tri 9689 14737 9787 14835 ne
rect 9787 14737 10141 14835
tri 10141 14737 10239 14835 sw
tri 10239 14737 10337 14835 ne
rect 10337 14737 10691 14835
tri 10691 14737 10789 14835 sw
tri 10789 14737 10887 14835 ne
rect 10887 14737 11241 14835
tri 11241 14737 11339 14835 sw
tri 11339 14737 11437 14835 ne
rect 11437 14737 11791 14835
tri 11791 14737 11889 14835 sw
tri 11889 14737 11987 14835 ne
rect 11987 14737 12341 14835
tri 12341 14737 12439 14835 sw
tri 12439 14737 12537 14835 ne
rect 12537 14737 12891 14835
tri 12891 14737 12989 14835 sw
tri 12989 14737 13087 14835 ne
rect 13087 14737 13441 14835
tri 13441 14737 13539 14835 sw
tri 13539 14737 13637 14835 ne
rect 13637 14737 13991 14835
tri 13991 14737 14089 14835 sw
tri 14089 14737 14187 14835 ne
rect 14187 14737 14541 14835
tri 14541 14737 14639 14835 sw
tri 14639 14737 14737 14835 ne
rect 14737 14737 15091 14835
tri 15091 14737 15189 14835 sw
tri 15189 14737 15287 14835 ne
rect 15287 14737 15641 14835
tri 15641 14737 15739 14835 sw
tri 15739 14737 15837 14835 ne
rect 15837 14737 16191 14835
tri 16191 14737 16289 14835 sw
tri 16289 14737 16387 14835 ne
rect 16387 14737 16741 14835
tri 16741 14737 16839 14835 sw
tri 16839 14737 16937 14835 ne
rect 16937 14737 17291 14835
tri 17291 14737 17389 14835 sw
tri 17389 14737 17487 14835 ne
rect 17487 14737 17841 14835
tri 17841 14737 17939 14835 sw
tri 17939 14737 18037 14835 ne
rect 18037 14737 18391 14835
tri 18391 14737 18489 14835 sw
tri 18489 14737 18587 14835 ne
rect 18587 14737 18941 14835
tri 18941 14737 19039 14835 sw
tri 19039 14737 19137 14835 ne
rect 19137 14737 19491 14835
tri 19491 14737 19589 14835 sw
tri 19589 14737 19687 14835 ne
rect 19687 14737 21800 14835
rect -300 14687 339 14737
rect -500 14639 339 14687
tri 339 14639 437 14737 sw
tri 437 14639 535 14737 ne
rect 535 14639 889 14737
tri 889 14639 987 14737 sw
tri 987 14639 1085 14737 ne
rect 1085 14639 1439 14737
tri 1439 14639 1537 14737 sw
tri 1537 14639 1635 14737 ne
rect 1635 14639 1989 14737
tri 1989 14639 2087 14737 sw
tri 2087 14639 2185 14737 ne
rect 2185 14639 2539 14737
tri 2539 14639 2637 14737 sw
tri 2637 14639 2735 14737 ne
rect 2735 14639 3089 14737
tri 3089 14639 3187 14737 sw
tri 3187 14639 3285 14737 ne
rect 3285 14639 3639 14737
tri 3639 14639 3737 14737 sw
tri 3737 14639 3835 14737 ne
rect 3835 14639 4189 14737
tri 4189 14639 4287 14737 sw
tri 4287 14639 4385 14737 ne
rect 4385 14639 4739 14737
tri 4739 14639 4837 14737 sw
tri 4837 14639 4935 14737 ne
rect 4935 14639 5289 14737
tri 5289 14639 5387 14737 sw
tri 5387 14639 5485 14737 ne
rect 5485 14639 5839 14737
tri 5839 14639 5937 14737 sw
tri 5937 14639 6035 14737 ne
rect 6035 14639 6389 14737
tri 6389 14639 6487 14737 sw
tri 6487 14639 6585 14737 ne
rect 6585 14639 6939 14737
tri 6939 14639 7037 14737 sw
tri 7037 14639 7135 14737 ne
rect 7135 14639 7489 14737
tri 7489 14639 7587 14737 sw
tri 7587 14639 7685 14737 ne
rect 7685 14639 8039 14737
tri 8039 14639 8137 14737 sw
tri 8137 14639 8235 14737 ne
rect 8235 14639 8589 14737
tri 8589 14639 8687 14737 sw
tri 8687 14639 8785 14737 ne
rect 8785 14639 9139 14737
tri 9139 14639 9237 14737 sw
tri 9237 14639 9335 14737 ne
rect 9335 14639 9689 14737
tri 9689 14639 9787 14737 sw
tri 9787 14639 9885 14737 ne
rect 9885 14639 10239 14737
tri 10239 14639 10337 14737 sw
tri 10337 14639 10435 14737 ne
rect 10435 14639 10789 14737
tri 10789 14639 10887 14737 sw
tri 10887 14639 10985 14737 ne
rect 10985 14639 11339 14737
tri 11339 14639 11437 14737 sw
tri 11437 14639 11535 14737 ne
rect 11535 14639 11889 14737
tri 11889 14639 11987 14737 sw
tri 11987 14639 12085 14737 ne
rect 12085 14639 12439 14737
tri 12439 14639 12537 14737 sw
tri 12537 14639 12635 14737 ne
rect 12635 14639 12989 14737
tri 12989 14639 13087 14737 sw
tri 13087 14639 13185 14737 ne
rect 13185 14639 13539 14737
tri 13539 14639 13637 14737 sw
tri 13637 14639 13735 14737 ne
rect 13735 14639 14089 14737
tri 14089 14639 14187 14737 sw
tri 14187 14639 14285 14737 ne
rect 14285 14639 14639 14737
tri 14639 14639 14737 14737 sw
tri 14737 14639 14835 14737 ne
rect 14835 14639 15189 14737
tri 15189 14639 15287 14737 sw
tri 15287 14639 15385 14737 ne
rect 15385 14639 15739 14737
tri 15739 14639 15837 14737 sw
tri 15837 14639 15935 14737 ne
rect 15935 14639 16289 14737
tri 16289 14639 16387 14737 sw
tri 16387 14639 16485 14737 ne
rect 16485 14639 16839 14737
tri 16839 14639 16937 14737 sw
tri 16937 14639 17035 14737 ne
rect 17035 14639 17389 14737
tri 17389 14639 17487 14737 sw
tri 17487 14639 17585 14737 ne
rect 17585 14639 17939 14737
tri 17939 14639 18037 14737 sw
tri 18037 14639 18135 14737 ne
rect 18135 14639 18489 14737
tri 18489 14639 18587 14737 sw
tri 18587 14639 18685 14737 ne
rect 18685 14639 19039 14737
tri 19039 14639 19137 14737 sw
tri 19137 14639 19235 14737 ne
rect 19235 14639 19589 14737
tri 19589 14639 19687 14737 sw
rect -500 14635 437 14639
rect -500 14515 215 14635
rect 335 14541 437 14635
tri 437 14541 535 14639 sw
tri 535 14541 633 14639 ne
rect 633 14635 987 14639
rect 633 14541 765 14635
rect 335 14515 535 14541
rect -500 14511 535 14515
tri 535 14511 565 14541 sw
tri 633 14511 663 14541 ne
rect 663 14515 765 14541
rect 885 14541 987 14635
tri 987 14541 1085 14639 sw
tri 1085 14541 1183 14639 ne
rect 1183 14635 1537 14639
rect 1183 14541 1315 14635
rect 885 14515 1085 14541
rect 663 14511 1085 14515
tri 1085 14511 1115 14541 sw
tri 1183 14511 1213 14541 ne
rect 1213 14515 1315 14541
rect 1435 14541 1537 14635
tri 1537 14541 1635 14639 sw
tri 1635 14541 1733 14639 ne
rect 1733 14635 2087 14639
rect 1733 14541 1865 14635
rect 1435 14515 1635 14541
rect 1213 14511 1635 14515
tri 1635 14511 1665 14541 sw
tri 1733 14511 1763 14541 ne
rect 1763 14515 1865 14541
rect 1985 14541 2087 14635
tri 2087 14541 2185 14639 sw
tri 2185 14541 2283 14639 ne
rect 2283 14635 2637 14639
rect 2283 14541 2415 14635
rect 1985 14515 2185 14541
rect 1763 14511 2185 14515
tri 2185 14511 2215 14541 sw
tri 2283 14511 2313 14541 ne
rect 2313 14515 2415 14541
rect 2535 14541 2637 14635
tri 2637 14541 2735 14639 sw
tri 2735 14541 2833 14639 ne
rect 2833 14635 3187 14639
rect 2833 14541 2965 14635
rect 2535 14515 2735 14541
rect 2313 14511 2735 14515
tri 2735 14511 2765 14541 sw
tri 2833 14511 2863 14541 ne
rect 2863 14515 2965 14541
rect 3085 14541 3187 14635
tri 3187 14541 3285 14639 sw
tri 3285 14541 3383 14639 ne
rect 3383 14635 3737 14639
rect 3383 14541 3515 14635
rect 3085 14515 3285 14541
rect 2863 14511 3285 14515
tri 3285 14511 3315 14541 sw
tri 3383 14511 3413 14541 ne
rect 3413 14515 3515 14541
rect 3635 14541 3737 14635
tri 3737 14541 3835 14639 sw
tri 3835 14541 3933 14639 ne
rect 3933 14635 4287 14639
rect 3933 14541 4065 14635
rect 3635 14515 3835 14541
rect 3413 14511 3835 14515
tri 3835 14511 3865 14541 sw
tri 3933 14511 3963 14541 ne
rect 3963 14515 4065 14541
rect 4185 14541 4287 14635
tri 4287 14541 4385 14639 sw
tri 4385 14541 4483 14639 ne
rect 4483 14635 4837 14639
rect 4483 14541 4615 14635
rect 4185 14515 4385 14541
rect 3963 14511 4385 14515
tri 4385 14511 4415 14541 sw
tri 4483 14511 4513 14541 ne
rect 4513 14515 4615 14541
rect 4735 14541 4837 14635
tri 4837 14541 4935 14639 sw
tri 4935 14541 5033 14639 ne
rect 5033 14635 5387 14639
rect 5033 14541 5165 14635
rect 4735 14515 4935 14541
rect 4513 14511 4935 14515
tri 4935 14511 4965 14541 sw
tri 5033 14511 5063 14541 ne
rect 5063 14515 5165 14541
rect 5285 14541 5387 14635
tri 5387 14541 5485 14639 sw
tri 5485 14541 5583 14639 ne
rect 5583 14635 5937 14639
rect 5583 14541 5715 14635
rect 5285 14515 5485 14541
rect 5063 14511 5485 14515
tri 5485 14511 5515 14541 sw
tri 5583 14511 5613 14541 ne
rect 5613 14515 5715 14541
rect 5835 14541 5937 14635
tri 5937 14541 6035 14639 sw
tri 6035 14541 6133 14639 ne
rect 6133 14635 6487 14639
rect 6133 14541 6265 14635
rect 5835 14515 6035 14541
rect 5613 14511 6035 14515
tri 6035 14511 6065 14541 sw
tri 6133 14511 6163 14541 ne
rect 6163 14515 6265 14541
rect 6385 14541 6487 14635
tri 6487 14541 6585 14639 sw
tri 6585 14541 6683 14639 ne
rect 6683 14635 7037 14639
rect 6683 14541 6815 14635
rect 6385 14515 6585 14541
rect 6163 14511 6585 14515
tri 6585 14511 6615 14541 sw
tri 6683 14511 6713 14541 ne
rect 6713 14515 6815 14541
rect 6935 14541 7037 14635
tri 7037 14541 7135 14639 sw
tri 7135 14541 7233 14639 ne
rect 7233 14635 7587 14639
rect 7233 14541 7365 14635
rect 6935 14515 7135 14541
rect 6713 14511 7135 14515
tri 7135 14511 7165 14541 sw
tri 7233 14511 7263 14541 ne
rect 7263 14515 7365 14541
rect 7485 14541 7587 14635
tri 7587 14541 7685 14639 sw
tri 7685 14541 7783 14639 ne
rect 7783 14635 8137 14639
rect 7783 14541 7915 14635
rect 7485 14515 7685 14541
rect 7263 14511 7685 14515
tri 7685 14511 7715 14541 sw
tri 7783 14511 7813 14541 ne
rect 7813 14515 7915 14541
rect 8035 14541 8137 14635
tri 8137 14541 8235 14639 sw
tri 8235 14541 8333 14639 ne
rect 8333 14635 8687 14639
rect 8333 14541 8465 14635
rect 8035 14515 8235 14541
rect 7813 14511 8235 14515
tri 8235 14511 8265 14541 sw
tri 8333 14511 8363 14541 ne
rect 8363 14515 8465 14541
rect 8585 14541 8687 14635
tri 8687 14541 8785 14639 sw
tri 8785 14541 8883 14639 ne
rect 8883 14635 9237 14639
rect 8883 14541 9015 14635
rect 8585 14515 8785 14541
rect 8363 14511 8785 14515
tri 8785 14511 8815 14541 sw
tri 8883 14511 8913 14541 ne
rect 8913 14515 9015 14541
rect 9135 14541 9237 14635
tri 9237 14541 9335 14639 sw
tri 9335 14541 9433 14639 ne
rect 9433 14635 9787 14639
rect 9433 14541 9565 14635
rect 9135 14515 9335 14541
rect 8913 14511 9335 14515
tri 9335 14511 9365 14541 sw
tri 9433 14511 9463 14541 ne
rect 9463 14515 9565 14541
rect 9685 14541 9787 14635
tri 9787 14541 9885 14639 sw
tri 9885 14541 9983 14639 ne
rect 9983 14635 10337 14639
rect 9983 14541 10115 14635
rect 9685 14515 9885 14541
rect 9463 14511 9885 14515
tri 9885 14511 9915 14541 sw
tri 9983 14511 10013 14541 ne
rect 10013 14515 10115 14541
rect 10235 14541 10337 14635
tri 10337 14541 10435 14639 sw
tri 10435 14541 10533 14639 ne
rect 10533 14635 10887 14639
rect 10533 14541 10665 14635
rect 10235 14515 10435 14541
rect 10013 14511 10435 14515
tri 10435 14511 10465 14541 sw
tri 10533 14511 10563 14541 ne
rect 10563 14515 10665 14541
rect 10785 14541 10887 14635
tri 10887 14541 10985 14639 sw
tri 10985 14541 11083 14639 ne
rect 11083 14635 11437 14639
rect 11083 14541 11215 14635
rect 10785 14515 10985 14541
rect 10563 14511 10985 14515
tri 10985 14511 11015 14541 sw
tri 11083 14511 11113 14541 ne
rect 11113 14515 11215 14541
rect 11335 14541 11437 14635
tri 11437 14541 11535 14639 sw
tri 11535 14541 11633 14639 ne
rect 11633 14635 11987 14639
rect 11633 14541 11765 14635
rect 11335 14515 11535 14541
rect 11113 14511 11535 14515
tri 11535 14511 11565 14541 sw
tri 11633 14511 11663 14541 ne
rect 11663 14515 11765 14541
rect 11885 14541 11987 14635
tri 11987 14541 12085 14639 sw
tri 12085 14541 12183 14639 ne
rect 12183 14635 12537 14639
rect 12183 14541 12315 14635
rect 11885 14515 12085 14541
rect 11663 14511 12085 14515
tri 12085 14511 12115 14541 sw
tri 12183 14511 12213 14541 ne
rect 12213 14515 12315 14541
rect 12435 14541 12537 14635
tri 12537 14541 12635 14639 sw
tri 12635 14541 12733 14639 ne
rect 12733 14635 13087 14639
rect 12733 14541 12865 14635
rect 12435 14515 12635 14541
rect 12213 14511 12635 14515
tri 12635 14511 12665 14541 sw
tri 12733 14511 12763 14541 ne
rect 12763 14515 12865 14541
rect 12985 14541 13087 14635
tri 13087 14541 13185 14639 sw
tri 13185 14541 13283 14639 ne
rect 13283 14635 13637 14639
rect 13283 14541 13415 14635
rect 12985 14515 13185 14541
rect 12763 14511 13185 14515
tri 13185 14511 13215 14541 sw
tri 13283 14511 13313 14541 ne
rect 13313 14515 13415 14541
rect 13535 14541 13637 14635
tri 13637 14541 13735 14639 sw
tri 13735 14541 13833 14639 ne
rect 13833 14635 14187 14639
rect 13833 14541 13965 14635
rect 13535 14515 13735 14541
rect 13313 14511 13735 14515
tri 13735 14511 13765 14541 sw
tri 13833 14511 13863 14541 ne
rect 13863 14515 13965 14541
rect 14085 14541 14187 14635
tri 14187 14541 14285 14639 sw
tri 14285 14541 14383 14639 ne
rect 14383 14635 14737 14639
rect 14383 14541 14515 14635
rect 14085 14515 14285 14541
rect 13863 14511 14285 14515
tri 14285 14511 14315 14541 sw
tri 14383 14511 14413 14541 ne
rect 14413 14515 14515 14541
rect 14635 14541 14737 14635
tri 14737 14541 14835 14639 sw
tri 14835 14541 14933 14639 ne
rect 14933 14635 15287 14639
rect 14933 14541 15065 14635
rect 14635 14515 14835 14541
rect 14413 14511 14835 14515
tri 14835 14511 14865 14541 sw
tri 14933 14511 14963 14541 ne
rect 14963 14515 15065 14541
rect 15185 14541 15287 14635
tri 15287 14541 15385 14639 sw
tri 15385 14541 15483 14639 ne
rect 15483 14635 15837 14639
rect 15483 14541 15615 14635
rect 15185 14515 15385 14541
rect 14963 14511 15385 14515
tri 15385 14511 15415 14541 sw
tri 15483 14511 15513 14541 ne
rect 15513 14515 15615 14541
rect 15735 14541 15837 14635
tri 15837 14541 15935 14639 sw
tri 15935 14541 16033 14639 ne
rect 16033 14635 16387 14639
rect 16033 14541 16165 14635
rect 15735 14515 15935 14541
rect 15513 14511 15935 14515
tri 15935 14511 15965 14541 sw
tri 16033 14511 16063 14541 ne
rect 16063 14515 16165 14541
rect 16285 14541 16387 14635
tri 16387 14541 16485 14639 sw
tri 16485 14541 16583 14639 ne
rect 16583 14635 16937 14639
rect 16583 14541 16715 14635
rect 16285 14515 16485 14541
rect 16063 14511 16485 14515
tri 16485 14511 16515 14541 sw
tri 16583 14511 16613 14541 ne
rect 16613 14515 16715 14541
rect 16835 14541 16937 14635
tri 16937 14541 17035 14639 sw
tri 17035 14541 17133 14639 ne
rect 17133 14635 17487 14639
rect 17133 14541 17265 14635
rect 16835 14515 17035 14541
rect 16613 14511 17035 14515
tri 17035 14511 17065 14541 sw
tri 17133 14511 17163 14541 ne
rect 17163 14515 17265 14541
rect 17385 14541 17487 14635
tri 17487 14541 17585 14639 sw
tri 17585 14541 17683 14639 ne
rect 17683 14635 18037 14639
rect 17683 14541 17815 14635
rect 17385 14515 17585 14541
rect 17163 14511 17585 14515
tri 17585 14511 17615 14541 sw
tri 17683 14511 17713 14541 ne
rect 17713 14515 17815 14541
rect 17935 14541 18037 14635
tri 18037 14541 18135 14639 sw
tri 18135 14541 18233 14639 ne
rect 18233 14635 18587 14639
rect 18233 14541 18365 14635
rect 17935 14515 18135 14541
rect 17713 14511 18135 14515
tri 18135 14511 18165 14541 sw
tri 18233 14511 18263 14541 ne
rect 18263 14515 18365 14541
rect 18485 14541 18587 14635
tri 18587 14541 18685 14639 sw
tri 18685 14541 18783 14639 ne
rect 18783 14635 19137 14639
rect 18783 14541 18915 14635
rect 18485 14515 18685 14541
rect 18263 14511 18685 14515
tri 18685 14511 18715 14541 sw
tri 18783 14511 18813 14541 ne
rect 18813 14515 18915 14541
rect 19035 14541 19137 14635
tri 19137 14541 19235 14639 sw
tri 19235 14541 19333 14639 ne
rect 19333 14635 20300 14639
rect 19333 14541 19465 14635
rect 19035 14515 19235 14541
rect 18813 14511 19235 14515
tri 19235 14511 19265 14541 sw
tri 19333 14511 19363 14541 ne
rect 19363 14515 19465 14541
rect 19585 14515 20300 14635
rect 19363 14511 20300 14515
tri 113 14413 211 14511 ne
rect 211 14413 565 14511
tri 565 14413 663 14511 sw
tri 663 14413 761 14511 ne
rect 761 14413 1115 14511
tri 1115 14413 1213 14511 sw
tri 1213 14413 1311 14511 ne
rect 1311 14413 1665 14511
tri 1665 14413 1763 14511 sw
tri 1763 14413 1861 14511 ne
rect 1861 14413 2215 14511
tri 2215 14413 2313 14511 sw
tri 2313 14413 2411 14511 ne
rect 2411 14413 2765 14511
tri 2765 14413 2863 14511 sw
tri 2863 14413 2961 14511 ne
rect 2961 14413 3315 14511
tri 3315 14413 3413 14511 sw
tri 3413 14413 3511 14511 ne
rect 3511 14413 3865 14511
tri 3865 14413 3963 14511 sw
tri 3963 14413 4061 14511 ne
rect 4061 14413 4415 14511
tri 4415 14413 4513 14511 sw
tri 4513 14413 4611 14511 ne
rect 4611 14413 4965 14511
tri 4965 14413 5063 14511 sw
tri 5063 14413 5161 14511 ne
rect 5161 14413 5515 14511
tri 5515 14413 5613 14511 sw
tri 5613 14413 5711 14511 ne
rect 5711 14413 6065 14511
tri 6065 14413 6163 14511 sw
tri 6163 14413 6261 14511 ne
rect 6261 14413 6615 14511
tri 6615 14413 6713 14511 sw
tri 6713 14413 6811 14511 ne
rect 6811 14413 7165 14511
tri 7165 14413 7263 14511 sw
tri 7263 14413 7361 14511 ne
rect 7361 14413 7715 14511
tri 7715 14413 7813 14511 sw
tri 7813 14413 7911 14511 ne
rect 7911 14413 8265 14511
tri 8265 14413 8363 14511 sw
tri 8363 14413 8461 14511 ne
rect 8461 14413 8815 14511
tri 8815 14413 8913 14511 sw
tri 8913 14413 9011 14511 ne
rect 9011 14413 9365 14511
tri 9365 14413 9463 14511 sw
tri 9463 14413 9561 14511 ne
rect 9561 14413 9915 14511
tri 9915 14413 10013 14511 sw
tri 10013 14413 10111 14511 ne
rect 10111 14413 10465 14511
tri 10465 14413 10563 14511 sw
tri 10563 14413 10661 14511 ne
rect 10661 14413 11015 14511
tri 11015 14413 11113 14511 sw
tri 11113 14413 11211 14511 ne
rect 11211 14413 11565 14511
tri 11565 14413 11663 14511 sw
tri 11663 14413 11761 14511 ne
rect 11761 14413 12115 14511
tri 12115 14413 12213 14511 sw
tri 12213 14413 12311 14511 ne
rect 12311 14413 12665 14511
tri 12665 14413 12763 14511 sw
tri 12763 14413 12861 14511 ne
rect 12861 14413 13215 14511
tri 13215 14413 13313 14511 sw
tri 13313 14413 13411 14511 ne
rect 13411 14413 13765 14511
tri 13765 14413 13863 14511 sw
tri 13863 14413 13961 14511 ne
rect 13961 14413 14315 14511
tri 14315 14413 14413 14511 sw
tri 14413 14413 14511 14511 ne
rect 14511 14413 14865 14511
tri 14865 14413 14963 14511 sw
tri 14963 14413 15061 14511 ne
rect 15061 14413 15415 14511
tri 15415 14413 15513 14511 sw
tri 15513 14413 15611 14511 ne
rect 15611 14413 15965 14511
tri 15965 14413 16063 14511 sw
tri 16063 14413 16161 14511 ne
rect 16161 14413 16515 14511
tri 16515 14413 16613 14511 sw
tri 16613 14413 16711 14511 ne
rect 16711 14413 17065 14511
tri 17065 14413 17163 14511 sw
tri 17163 14413 17261 14511 ne
rect 17261 14413 17615 14511
tri 17615 14413 17713 14511 sw
tri 17713 14413 17811 14511 ne
rect 17811 14413 18165 14511
tri 18165 14413 18263 14511 sw
tri 18263 14413 18361 14511 ne
rect 18361 14413 18715 14511
tri 18715 14413 18813 14511 sw
tri 18813 14413 18911 14511 ne
rect 18911 14413 19265 14511
tri 19265 14413 19363 14511 sw
tri 19363 14413 19461 14511 ne
rect 19461 14413 20300 14511
rect -2000 14383 113 14413
tri 113 14383 143 14413 sw
tri 211 14383 241 14413 ne
rect 241 14383 663 14413
tri 663 14383 693 14413 sw
tri 761 14383 791 14413 ne
rect 791 14383 1213 14413
tri 1213 14383 1243 14413 sw
tri 1311 14383 1341 14413 ne
rect 1341 14383 1763 14413
tri 1763 14383 1793 14413 sw
tri 1861 14383 1891 14413 ne
rect 1891 14383 2313 14413
tri 2313 14383 2343 14413 sw
tri 2411 14383 2441 14413 ne
rect 2441 14383 2863 14413
tri 2863 14383 2893 14413 sw
tri 2961 14383 2991 14413 ne
rect 2991 14383 3413 14413
tri 3413 14383 3443 14413 sw
tri 3511 14383 3541 14413 ne
rect 3541 14383 3963 14413
tri 3963 14383 3993 14413 sw
tri 4061 14383 4091 14413 ne
rect 4091 14383 4513 14413
tri 4513 14383 4543 14413 sw
tri 4611 14383 4641 14413 ne
rect 4641 14383 5063 14413
tri 5063 14383 5093 14413 sw
tri 5161 14383 5191 14413 ne
rect 5191 14383 5613 14413
tri 5613 14383 5643 14413 sw
tri 5711 14383 5741 14413 ne
rect 5741 14383 6163 14413
tri 6163 14383 6193 14413 sw
tri 6261 14383 6291 14413 ne
rect 6291 14383 6713 14413
tri 6713 14383 6743 14413 sw
tri 6811 14383 6841 14413 ne
rect 6841 14383 7263 14413
tri 7263 14383 7293 14413 sw
tri 7361 14383 7391 14413 ne
rect 7391 14383 7813 14413
tri 7813 14383 7843 14413 sw
tri 7911 14383 7941 14413 ne
rect 7941 14383 8363 14413
tri 8363 14383 8393 14413 sw
tri 8461 14383 8491 14413 ne
rect 8491 14383 8913 14413
tri 8913 14383 8943 14413 sw
tri 9011 14383 9041 14413 ne
rect 9041 14383 9463 14413
tri 9463 14383 9493 14413 sw
tri 9561 14383 9591 14413 ne
rect 9591 14383 10013 14413
tri 10013 14383 10043 14413 sw
tri 10111 14383 10141 14413 ne
rect 10141 14383 10563 14413
tri 10563 14383 10593 14413 sw
tri 10661 14383 10691 14413 ne
rect 10691 14383 11113 14413
tri 11113 14383 11143 14413 sw
tri 11211 14383 11241 14413 ne
rect 11241 14383 11663 14413
tri 11663 14383 11693 14413 sw
tri 11761 14383 11791 14413 ne
rect 11791 14383 12213 14413
tri 12213 14383 12243 14413 sw
tri 12311 14383 12341 14413 ne
rect 12341 14383 12763 14413
tri 12763 14383 12793 14413 sw
tri 12861 14383 12891 14413 ne
rect 12891 14383 13313 14413
tri 13313 14383 13343 14413 sw
tri 13411 14383 13441 14413 ne
rect 13441 14383 13863 14413
tri 13863 14383 13893 14413 sw
tri 13961 14383 13991 14413 ne
rect 13991 14383 14413 14413
tri 14413 14383 14443 14413 sw
tri 14511 14383 14541 14413 ne
rect 14541 14383 14963 14413
tri 14963 14383 14993 14413 sw
tri 15061 14383 15091 14413 ne
rect 15091 14383 15513 14413
tri 15513 14383 15543 14413 sw
tri 15611 14383 15641 14413 ne
rect 15641 14383 16063 14413
tri 16063 14383 16093 14413 sw
tri 16161 14383 16191 14413 ne
rect 16191 14383 16613 14413
tri 16613 14383 16643 14413 sw
tri 16711 14383 16741 14413 ne
rect 16741 14383 17163 14413
tri 17163 14383 17193 14413 sw
tri 17261 14383 17291 14413 ne
rect 17291 14383 17713 14413
tri 17713 14383 17743 14413 sw
tri 17811 14383 17841 14413 ne
rect 17841 14383 18263 14413
tri 18263 14383 18293 14413 sw
tri 18361 14383 18391 14413 ne
rect 18391 14383 18813 14413
tri 18813 14383 18843 14413 sw
tri 18911 14383 18941 14413 ne
rect 18941 14383 19363 14413
tri 19363 14383 19393 14413 sw
tri 19461 14383 19491 14413 ne
rect 19491 14383 20300 14413
rect -2000 14285 143 14383
tri 143 14285 241 14383 sw
tri 241 14285 339 14383 ne
rect 339 14285 693 14383
tri 693 14285 791 14383 sw
tri 791 14285 889 14383 ne
rect 889 14285 1243 14383
tri 1243 14285 1341 14383 sw
tri 1341 14285 1439 14383 ne
rect 1439 14285 1793 14383
tri 1793 14285 1891 14383 sw
tri 1891 14285 1989 14383 ne
rect 1989 14285 2343 14383
tri 2343 14285 2441 14383 sw
tri 2441 14285 2539 14383 ne
rect 2539 14285 2893 14383
tri 2893 14285 2991 14383 sw
tri 2991 14285 3089 14383 ne
rect 3089 14285 3443 14383
tri 3443 14285 3541 14383 sw
tri 3541 14285 3639 14383 ne
rect 3639 14285 3993 14383
tri 3993 14285 4091 14383 sw
tri 4091 14285 4189 14383 ne
rect 4189 14285 4543 14383
tri 4543 14285 4641 14383 sw
tri 4641 14285 4739 14383 ne
rect 4739 14285 5093 14383
tri 5093 14285 5191 14383 sw
tri 5191 14285 5289 14383 ne
rect 5289 14285 5643 14383
tri 5643 14285 5741 14383 sw
tri 5741 14285 5839 14383 ne
rect 5839 14285 6193 14383
tri 6193 14285 6291 14383 sw
tri 6291 14285 6389 14383 ne
rect 6389 14285 6743 14383
tri 6743 14285 6841 14383 sw
tri 6841 14285 6939 14383 ne
rect 6939 14285 7293 14383
tri 7293 14285 7391 14383 sw
tri 7391 14285 7489 14383 ne
rect 7489 14285 7843 14383
tri 7843 14285 7941 14383 sw
tri 7941 14285 8039 14383 ne
rect 8039 14285 8393 14383
tri 8393 14285 8491 14383 sw
tri 8491 14285 8589 14383 ne
rect 8589 14285 8943 14383
tri 8943 14285 9041 14383 sw
tri 9041 14285 9139 14383 ne
rect 9139 14285 9493 14383
tri 9493 14285 9591 14383 sw
tri 9591 14285 9689 14383 ne
rect 9689 14285 10043 14383
tri 10043 14285 10141 14383 sw
tri 10141 14285 10239 14383 ne
rect 10239 14285 10593 14383
tri 10593 14285 10691 14383 sw
tri 10691 14285 10789 14383 ne
rect 10789 14285 11143 14383
tri 11143 14285 11241 14383 sw
tri 11241 14285 11339 14383 ne
rect 11339 14285 11693 14383
tri 11693 14285 11791 14383 sw
tri 11791 14285 11889 14383 ne
rect 11889 14285 12243 14383
tri 12243 14285 12341 14383 sw
tri 12341 14285 12439 14383 ne
rect 12439 14285 12793 14383
tri 12793 14285 12891 14383 sw
tri 12891 14285 12989 14383 ne
rect 12989 14285 13343 14383
tri 13343 14285 13441 14383 sw
tri 13441 14285 13539 14383 ne
rect 13539 14285 13893 14383
tri 13893 14285 13991 14383 sw
tri 13991 14285 14089 14383 ne
rect 14089 14285 14443 14383
tri 14443 14285 14541 14383 sw
tri 14541 14285 14639 14383 ne
rect 14639 14285 14993 14383
tri 14993 14285 15091 14383 sw
tri 15091 14285 15189 14383 ne
rect 15189 14285 15543 14383
tri 15543 14285 15641 14383 sw
tri 15641 14285 15739 14383 ne
rect 15739 14285 16093 14383
tri 16093 14285 16191 14383 sw
tri 16191 14285 16289 14383 ne
rect 16289 14285 16643 14383
tri 16643 14285 16741 14383 sw
tri 16741 14285 16839 14383 ne
rect 16839 14285 17193 14383
tri 17193 14285 17291 14383 sw
tri 17291 14285 17389 14383 ne
rect 17389 14285 17743 14383
tri 17743 14285 17841 14383 sw
tri 17841 14285 17939 14383 ne
rect 17939 14285 18293 14383
tri 18293 14285 18391 14383 sw
tri 18391 14285 18489 14383 ne
rect 18489 14285 18843 14383
tri 18843 14285 18941 14383 sw
tri 18941 14285 19039 14383 ne
rect 19039 14285 19393 14383
tri 19393 14285 19491 14383 sw
tri 19491 14285 19589 14383 ne
rect 19589 14285 20300 14383
rect -2000 14187 241 14285
tri 241 14187 339 14285 sw
tri 339 14187 437 14285 ne
rect 437 14187 791 14285
tri 791 14187 889 14285 sw
tri 889 14187 987 14285 ne
rect 987 14187 1341 14285
tri 1341 14187 1439 14285 sw
tri 1439 14187 1537 14285 ne
rect 1537 14187 1891 14285
tri 1891 14187 1989 14285 sw
tri 1989 14187 2087 14285 ne
rect 2087 14187 2441 14285
tri 2441 14187 2539 14285 sw
tri 2539 14187 2637 14285 ne
rect 2637 14187 2991 14285
tri 2991 14187 3089 14285 sw
tri 3089 14187 3187 14285 ne
rect 3187 14187 3541 14285
tri 3541 14187 3639 14285 sw
tri 3639 14187 3737 14285 ne
rect 3737 14187 4091 14285
tri 4091 14187 4189 14285 sw
tri 4189 14187 4287 14285 ne
rect 4287 14187 4641 14285
tri 4641 14187 4739 14285 sw
tri 4739 14187 4837 14285 ne
rect 4837 14187 5191 14285
tri 5191 14187 5289 14285 sw
tri 5289 14187 5387 14285 ne
rect 5387 14187 5741 14285
tri 5741 14187 5839 14285 sw
tri 5839 14187 5937 14285 ne
rect 5937 14187 6291 14285
tri 6291 14187 6389 14285 sw
tri 6389 14187 6487 14285 ne
rect 6487 14187 6841 14285
tri 6841 14187 6939 14285 sw
tri 6939 14187 7037 14285 ne
rect 7037 14187 7391 14285
tri 7391 14187 7489 14285 sw
tri 7489 14187 7587 14285 ne
rect 7587 14187 7941 14285
tri 7941 14187 8039 14285 sw
tri 8039 14187 8137 14285 ne
rect 8137 14187 8491 14285
tri 8491 14187 8589 14285 sw
tri 8589 14187 8687 14285 ne
rect 8687 14187 9041 14285
tri 9041 14187 9139 14285 sw
tri 9139 14187 9237 14285 ne
rect 9237 14187 9591 14285
tri 9591 14187 9689 14285 sw
tri 9689 14187 9787 14285 ne
rect 9787 14187 10141 14285
tri 10141 14187 10239 14285 sw
tri 10239 14187 10337 14285 ne
rect 10337 14187 10691 14285
tri 10691 14187 10789 14285 sw
tri 10789 14187 10887 14285 ne
rect 10887 14187 11241 14285
tri 11241 14187 11339 14285 sw
tri 11339 14187 11437 14285 ne
rect 11437 14187 11791 14285
tri 11791 14187 11889 14285 sw
tri 11889 14187 11987 14285 ne
rect 11987 14187 12341 14285
tri 12341 14187 12439 14285 sw
tri 12439 14187 12537 14285 ne
rect 12537 14187 12891 14285
tri 12891 14187 12989 14285 sw
tri 12989 14187 13087 14285 ne
rect 13087 14187 13441 14285
tri 13441 14187 13539 14285 sw
tri 13539 14187 13637 14285 ne
rect 13637 14187 13991 14285
tri 13991 14187 14089 14285 sw
tri 14089 14187 14187 14285 ne
rect 14187 14187 14541 14285
tri 14541 14187 14639 14285 sw
tri 14639 14187 14737 14285 ne
rect 14737 14187 15091 14285
tri 15091 14187 15189 14285 sw
tri 15189 14187 15287 14285 ne
rect 15287 14187 15641 14285
tri 15641 14187 15739 14285 sw
tri 15739 14187 15837 14285 ne
rect 15837 14187 16191 14285
tri 16191 14187 16289 14285 sw
tri 16289 14187 16387 14285 ne
rect 16387 14187 16741 14285
tri 16741 14187 16839 14285 sw
tri 16839 14187 16937 14285 ne
rect 16937 14187 17291 14285
tri 17291 14187 17389 14285 sw
tri 17389 14187 17487 14285 ne
rect 17487 14187 17841 14285
tri 17841 14187 17939 14285 sw
tri 17939 14187 18037 14285 ne
rect 18037 14187 18391 14285
tri 18391 14187 18489 14285 sw
tri 18489 14187 18587 14285 ne
rect 18587 14187 18941 14285
tri 18941 14187 19039 14285 sw
tri 19039 14187 19137 14285 ne
rect 19137 14187 19491 14285
tri 19491 14187 19589 14285 sw
tri 19589 14187 19687 14285 ne
rect 19687 14187 20300 14285
rect -2000 14089 339 14187
tri 339 14089 437 14187 sw
tri 437 14089 535 14187 ne
rect 535 14089 889 14187
tri 889 14089 987 14187 sw
tri 987 14089 1085 14187 ne
rect 1085 14089 1439 14187
tri 1439 14089 1537 14187 sw
tri 1537 14089 1635 14187 ne
rect 1635 14089 1989 14187
tri 1989 14089 2087 14187 sw
tri 2087 14089 2185 14187 ne
rect 2185 14089 2539 14187
tri 2539 14089 2637 14187 sw
tri 2637 14089 2735 14187 ne
rect 2735 14089 3089 14187
tri 3089 14089 3187 14187 sw
tri 3187 14089 3285 14187 ne
rect 3285 14089 3639 14187
tri 3639 14089 3737 14187 sw
tri 3737 14089 3835 14187 ne
rect 3835 14089 4189 14187
tri 4189 14089 4287 14187 sw
tri 4287 14089 4385 14187 ne
rect 4385 14089 4739 14187
tri 4739 14089 4837 14187 sw
tri 4837 14089 4935 14187 ne
rect 4935 14089 5289 14187
tri 5289 14089 5387 14187 sw
tri 5387 14089 5485 14187 ne
rect 5485 14089 5839 14187
tri 5839 14089 5937 14187 sw
tri 5937 14089 6035 14187 ne
rect 6035 14089 6389 14187
tri 6389 14089 6487 14187 sw
tri 6487 14089 6585 14187 ne
rect 6585 14089 6939 14187
tri 6939 14089 7037 14187 sw
tri 7037 14089 7135 14187 ne
rect 7135 14089 7489 14187
tri 7489 14089 7587 14187 sw
tri 7587 14089 7685 14187 ne
rect 7685 14089 8039 14187
tri 8039 14089 8137 14187 sw
tri 8137 14089 8235 14187 ne
rect 8235 14089 8589 14187
tri 8589 14089 8687 14187 sw
tri 8687 14089 8785 14187 ne
rect 8785 14089 9139 14187
tri 9139 14089 9237 14187 sw
tri 9237 14089 9335 14187 ne
rect 9335 14089 9689 14187
tri 9689 14089 9787 14187 sw
tri 9787 14089 9885 14187 ne
rect 9885 14089 10239 14187
tri 10239 14089 10337 14187 sw
tri 10337 14089 10435 14187 ne
rect 10435 14089 10789 14187
tri 10789 14089 10887 14187 sw
tri 10887 14089 10985 14187 ne
rect 10985 14089 11339 14187
tri 11339 14089 11437 14187 sw
tri 11437 14089 11535 14187 ne
rect 11535 14089 11889 14187
tri 11889 14089 11987 14187 sw
tri 11987 14089 12085 14187 ne
rect 12085 14089 12439 14187
tri 12439 14089 12537 14187 sw
tri 12537 14089 12635 14187 ne
rect 12635 14089 12989 14187
tri 12989 14089 13087 14187 sw
tri 13087 14089 13185 14187 ne
rect 13185 14089 13539 14187
tri 13539 14089 13637 14187 sw
tri 13637 14089 13735 14187 ne
rect 13735 14089 14089 14187
tri 14089 14089 14187 14187 sw
tri 14187 14089 14285 14187 ne
rect 14285 14089 14639 14187
tri 14639 14089 14737 14187 sw
tri 14737 14089 14835 14187 ne
rect 14835 14089 15189 14187
tri 15189 14089 15287 14187 sw
tri 15287 14089 15385 14187 ne
rect 15385 14089 15739 14187
tri 15739 14089 15837 14187 sw
tri 15837 14089 15935 14187 ne
rect 15935 14089 16289 14187
tri 16289 14089 16387 14187 sw
tri 16387 14089 16485 14187 ne
rect 16485 14089 16839 14187
tri 16839 14089 16937 14187 sw
tri 16937 14089 17035 14187 ne
rect 17035 14089 17389 14187
tri 17389 14089 17487 14187 sw
tri 17487 14089 17585 14187 ne
rect 17585 14089 17939 14187
tri 17939 14089 18037 14187 sw
tri 18037 14089 18135 14187 ne
rect 18135 14089 18489 14187
tri 18489 14089 18587 14187 sw
tri 18587 14089 18685 14187 ne
rect 18685 14089 19039 14187
tri 19039 14089 19137 14187 sw
tri 19137 14089 19235 14187 ne
rect 19235 14089 19589 14187
tri 19589 14089 19687 14187 sw
rect 20800 14089 21800 14737
rect -2000 14085 437 14089
rect -2000 13965 215 14085
rect 335 13991 437 14085
tri 437 13991 535 14089 sw
tri 535 13991 633 14089 ne
rect 633 14085 987 14089
rect 633 13991 765 14085
rect 335 13965 535 13991
rect -2000 13961 535 13965
rect -2000 13313 -1000 13961
tri 113 13863 211 13961 ne
rect 211 13913 535 13961
tri 535 13913 613 13991 sw
tri 633 13913 711 13991 ne
rect 711 13965 765 13991
rect 885 13991 987 14085
tri 987 13991 1085 14089 sw
tri 1085 13991 1183 14089 ne
rect 1183 14085 1537 14089
rect 1183 13991 1315 14085
rect 885 13965 1085 13991
rect 711 13913 1085 13965
tri 1085 13913 1163 13991 sw
tri 1183 13913 1261 13991 ne
rect 1261 13965 1315 13991
rect 1435 13991 1537 14085
tri 1537 13991 1635 14089 sw
tri 1635 13991 1733 14089 ne
rect 1733 14085 2087 14089
rect 1733 13991 1865 14085
rect 1435 13965 1635 13991
rect 1261 13913 1635 13965
tri 1635 13913 1713 13991 sw
tri 1733 13913 1811 13991 ne
rect 1811 13965 1865 13991
rect 1985 13991 2087 14085
tri 2087 13991 2185 14089 sw
tri 2185 13991 2283 14089 ne
rect 2283 14085 2637 14089
rect 2283 13991 2415 14085
rect 1985 13965 2185 13991
rect 1811 13913 2185 13965
tri 2185 13913 2263 13991 sw
tri 2283 13913 2361 13991 ne
rect 2361 13965 2415 13991
rect 2535 13991 2637 14085
tri 2637 13991 2735 14089 sw
tri 2735 13991 2833 14089 ne
rect 2833 14085 3187 14089
rect 2833 13991 2965 14085
rect 2535 13965 2735 13991
rect 2361 13913 2735 13965
tri 2735 13913 2813 13991 sw
tri 2833 13913 2911 13991 ne
rect 2911 13965 2965 13991
rect 3085 13991 3187 14085
tri 3187 13991 3285 14089 sw
tri 3285 13991 3383 14089 ne
rect 3383 14085 3737 14089
rect 3383 13991 3515 14085
rect 3085 13965 3285 13991
rect 2911 13913 3285 13965
tri 3285 13913 3363 13991 sw
tri 3383 13913 3461 13991 ne
rect 3461 13965 3515 13991
rect 3635 13991 3737 14085
tri 3737 13991 3835 14089 sw
tri 3835 13991 3933 14089 ne
rect 3933 14085 4287 14089
rect 3933 13991 4065 14085
rect 3635 13965 3835 13991
rect 3461 13913 3835 13965
tri 3835 13913 3913 13991 sw
tri 3933 13913 4011 13991 ne
rect 4011 13965 4065 13991
rect 4185 13991 4287 14085
tri 4287 13991 4385 14089 sw
tri 4385 13991 4483 14089 ne
rect 4483 14085 4837 14089
rect 4483 13991 4615 14085
rect 4185 13965 4385 13991
rect 4011 13913 4385 13965
tri 4385 13913 4463 13991 sw
tri 4483 13913 4561 13991 ne
rect 4561 13965 4615 13991
rect 4735 13991 4837 14085
tri 4837 13991 4935 14089 sw
tri 4935 13991 5033 14089 ne
rect 5033 14085 5387 14089
rect 5033 13991 5165 14085
rect 4735 13965 4935 13991
rect 4561 13913 4935 13965
tri 4935 13913 5013 13991 sw
tri 5033 13913 5111 13991 ne
rect 5111 13965 5165 13991
rect 5285 13991 5387 14085
tri 5387 13991 5485 14089 sw
tri 5485 13991 5583 14089 ne
rect 5583 14085 5937 14089
rect 5583 13991 5715 14085
rect 5285 13965 5485 13991
rect 5111 13913 5485 13965
tri 5485 13913 5563 13991 sw
tri 5583 13913 5661 13991 ne
rect 5661 13965 5715 13991
rect 5835 13991 5937 14085
tri 5937 13991 6035 14089 sw
tri 6035 13991 6133 14089 ne
rect 6133 14085 6487 14089
rect 6133 13991 6265 14085
rect 5835 13965 6035 13991
rect 5661 13913 6035 13965
tri 6035 13913 6113 13991 sw
tri 6133 13913 6211 13991 ne
rect 6211 13965 6265 13991
rect 6385 13991 6487 14085
tri 6487 13991 6585 14089 sw
tri 6585 13991 6683 14089 ne
rect 6683 14085 7037 14089
rect 6683 13991 6815 14085
rect 6385 13965 6585 13991
rect 6211 13913 6585 13965
tri 6585 13913 6663 13991 sw
tri 6683 13913 6761 13991 ne
rect 6761 13965 6815 13991
rect 6935 13991 7037 14085
tri 7037 13991 7135 14089 sw
tri 7135 13991 7233 14089 ne
rect 7233 14085 7587 14089
rect 7233 13991 7365 14085
rect 6935 13965 7135 13991
rect 6761 13913 7135 13965
tri 7135 13913 7213 13991 sw
tri 7233 13913 7311 13991 ne
rect 7311 13965 7365 13991
rect 7485 13991 7587 14085
tri 7587 13991 7685 14089 sw
tri 7685 13991 7783 14089 ne
rect 7783 14085 8137 14089
rect 7783 13991 7915 14085
rect 7485 13965 7685 13991
rect 7311 13913 7685 13965
tri 7685 13913 7763 13991 sw
tri 7783 13913 7861 13991 ne
rect 7861 13965 7915 13991
rect 8035 13991 8137 14085
tri 8137 13991 8235 14089 sw
tri 8235 13991 8333 14089 ne
rect 8333 14085 8687 14089
rect 8333 13991 8465 14085
rect 8035 13965 8235 13991
rect 7861 13913 8235 13965
tri 8235 13913 8313 13991 sw
tri 8333 13913 8411 13991 ne
rect 8411 13965 8465 13991
rect 8585 13991 8687 14085
tri 8687 13991 8785 14089 sw
tri 8785 13991 8883 14089 ne
rect 8883 14085 9237 14089
rect 8883 13991 9015 14085
rect 8585 13965 8785 13991
rect 8411 13913 8785 13965
tri 8785 13913 8863 13991 sw
tri 8883 13913 8961 13991 ne
rect 8961 13965 9015 13991
rect 9135 13991 9237 14085
tri 9237 13991 9335 14089 sw
tri 9335 13991 9433 14089 ne
rect 9433 14085 9787 14089
rect 9433 13991 9565 14085
rect 9135 13965 9335 13991
rect 8961 13913 9335 13965
tri 9335 13913 9413 13991 sw
tri 9433 13913 9511 13991 ne
rect 9511 13965 9565 13991
rect 9685 13991 9787 14085
tri 9787 13991 9885 14089 sw
tri 9885 13991 9983 14089 ne
rect 9983 14085 10337 14089
rect 9983 13991 10115 14085
rect 9685 13965 9885 13991
rect 9511 13913 9885 13965
tri 9885 13913 9963 13991 sw
tri 9983 13913 10061 13991 ne
rect 10061 13965 10115 13991
rect 10235 13991 10337 14085
tri 10337 13991 10435 14089 sw
tri 10435 13991 10533 14089 ne
rect 10533 14085 10887 14089
rect 10533 13991 10665 14085
rect 10235 13965 10435 13991
rect 10061 13913 10435 13965
tri 10435 13913 10513 13991 sw
tri 10533 13913 10611 13991 ne
rect 10611 13965 10665 13991
rect 10785 13991 10887 14085
tri 10887 13991 10985 14089 sw
tri 10985 13991 11083 14089 ne
rect 11083 14085 11437 14089
rect 11083 13991 11215 14085
rect 10785 13965 10985 13991
rect 10611 13913 10985 13965
tri 10985 13913 11063 13991 sw
tri 11083 13913 11161 13991 ne
rect 11161 13965 11215 13991
rect 11335 13991 11437 14085
tri 11437 13991 11535 14089 sw
tri 11535 13991 11633 14089 ne
rect 11633 14085 11987 14089
rect 11633 13991 11765 14085
rect 11335 13965 11535 13991
rect 11161 13913 11535 13965
tri 11535 13913 11613 13991 sw
tri 11633 13913 11711 13991 ne
rect 11711 13965 11765 13991
rect 11885 13991 11987 14085
tri 11987 13991 12085 14089 sw
tri 12085 13991 12183 14089 ne
rect 12183 14085 12537 14089
rect 12183 13991 12315 14085
rect 11885 13965 12085 13991
rect 11711 13913 12085 13965
tri 12085 13913 12163 13991 sw
tri 12183 13913 12261 13991 ne
rect 12261 13965 12315 13991
rect 12435 13991 12537 14085
tri 12537 13991 12635 14089 sw
tri 12635 13991 12733 14089 ne
rect 12733 14085 13087 14089
rect 12733 13991 12865 14085
rect 12435 13965 12635 13991
rect 12261 13913 12635 13965
tri 12635 13913 12713 13991 sw
tri 12733 13913 12811 13991 ne
rect 12811 13965 12865 13991
rect 12985 13991 13087 14085
tri 13087 13991 13185 14089 sw
tri 13185 13991 13283 14089 ne
rect 13283 14085 13637 14089
rect 13283 13991 13415 14085
rect 12985 13965 13185 13991
rect 12811 13913 13185 13965
tri 13185 13913 13263 13991 sw
tri 13283 13913 13361 13991 ne
rect 13361 13965 13415 13991
rect 13535 13991 13637 14085
tri 13637 13991 13735 14089 sw
tri 13735 13991 13833 14089 ne
rect 13833 14085 14187 14089
rect 13833 13991 13965 14085
rect 13535 13965 13735 13991
rect 13361 13913 13735 13965
tri 13735 13913 13813 13991 sw
tri 13833 13913 13911 13991 ne
rect 13911 13965 13965 13991
rect 14085 13991 14187 14085
tri 14187 13991 14285 14089 sw
tri 14285 13991 14383 14089 ne
rect 14383 14085 14737 14089
rect 14383 13991 14515 14085
rect 14085 13965 14285 13991
rect 13911 13913 14285 13965
tri 14285 13913 14363 13991 sw
tri 14383 13913 14461 13991 ne
rect 14461 13965 14515 13991
rect 14635 13991 14737 14085
tri 14737 13991 14835 14089 sw
tri 14835 13991 14933 14089 ne
rect 14933 14085 15287 14089
rect 14933 13991 15065 14085
rect 14635 13965 14835 13991
rect 14461 13913 14835 13965
tri 14835 13913 14913 13991 sw
tri 14933 13913 15011 13991 ne
rect 15011 13965 15065 13991
rect 15185 13991 15287 14085
tri 15287 13991 15385 14089 sw
tri 15385 13991 15483 14089 ne
rect 15483 14085 15837 14089
rect 15483 13991 15615 14085
rect 15185 13965 15385 13991
rect 15011 13913 15385 13965
tri 15385 13913 15463 13991 sw
tri 15483 13913 15561 13991 ne
rect 15561 13965 15615 13991
rect 15735 13991 15837 14085
tri 15837 13991 15935 14089 sw
tri 15935 13991 16033 14089 ne
rect 16033 14085 16387 14089
rect 16033 13991 16165 14085
rect 15735 13965 15935 13991
rect 15561 13913 15935 13965
tri 15935 13913 16013 13991 sw
tri 16033 13913 16111 13991 ne
rect 16111 13965 16165 13991
rect 16285 13991 16387 14085
tri 16387 13991 16485 14089 sw
tri 16485 13991 16583 14089 ne
rect 16583 14085 16937 14089
rect 16583 13991 16715 14085
rect 16285 13965 16485 13991
rect 16111 13913 16485 13965
tri 16485 13913 16563 13991 sw
tri 16583 13913 16661 13991 ne
rect 16661 13965 16715 13991
rect 16835 13991 16937 14085
tri 16937 13991 17035 14089 sw
tri 17035 13991 17133 14089 ne
rect 17133 14085 17487 14089
rect 17133 13991 17265 14085
rect 16835 13965 17035 13991
rect 16661 13913 17035 13965
tri 17035 13913 17113 13991 sw
tri 17133 13913 17211 13991 ne
rect 17211 13965 17265 13991
rect 17385 13991 17487 14085
tri 17487 13991 17585 14089 sw
tri 17585 13991 17683 14089 ne
rect 17683 14085 18037 14089
rect 17683 13991 17815 14085
rect 17385 13965 17585 13991
rect 17211 13913 17585 13965
tri 17585 13913 17663 13991 sw
tri 17683 13913 17761 13991 ne
rect 17761 13965 17815 13991
rect 17935 13991 18037 14085
tri 18037 13991 18135 14089 sw
tri 18135 13991 18233 14089 ne
rect 18233 14085 18587 14089
rect 18233 13991 18365 14085
rect 17935 13965 18135 13991
rect 17761 13913 18135 13965
tri 18135 13913 18213 13991 sw
tri 18233 13913 18311 13991 ne
rect 18311 13965 18365 13991
rect 18485 13991 18587 14085
tri 18587 13991 18685 14089 sw
tri 18685 13991 18783 14089 ne
rect 18783 14085 19137 14089
rect 18783 13991 18915 14085
rect 18485 13965 18685 13991
rect 18311 13913 18685 13965
tri 18685 13913 18763 13991 sw
tri 18783 13913 18861 13991 ne
rect 18861 13965 18915 13991
rect 19035 13991 19137 14085
tri 19137 13991 19235 14089 sw
tri 19235 13991 19333 14089 ne
rect 19333 14085 21800 14089
rect 19333 13991 19465 14085
rect 19035 13965 19235 13991
rect 18861 13913 19235 13965
tri 19235 13913 19313 13991 sw
tri 19333 13913 19411 13991 ne
rect 19411 13965 19465 13991
rect 19585 13965 21800 14085
rect 19411 13913 21800 13965
rect 211 13863 613 13913
rect -500 13813 113 13863
tri 113 13813 163 13863 sw
tri 211 13813 261 13863 ne
rect 261 13833 613 13863
tri 613 13833 693 13913 sw
tri 711 13833 791 13913 ne
rect 791 13833 1163 13913
tri 1163 13833 1243 13913 sw
tri 1261 13833 1341 13913 ne
rect 1341 13833 1713 13913
tri 1713 13833 1793 13913 sw
tri 1811 13833 1891 13913 ne
rect 1891 13833 2263 13913
tri 2263 13833 2343 13913 sw
tri 2361 13833 2441 13913 ne
rect 2441 13833 2813 13913
tri 2813 13833 2893 13913 sw
tri 2911 13833 2991 13913 ne
rect 2991 13833 3363 13913
tri 3363 13833 3443 13913 sw
tri 3461 13833 3541 13913 ne
rect 3541 13833 3913 13913
tri 3913 13833 3993 13913 sw
tri 4011 13833 4091 13913 ne
rect 4091 13833 4463 13913
tri 4463 13833 4543 13913 sw
tri 4561 13833 4641 13913 ne
rect 4641 13833 5013 13913
tri 5013 13833 5093 13913 sw
tri 5111 13833 5191 13913 ne
rect 5191 13833 5563 13913
tri 5563 13833 5643 13913 sw
tri 5661 13833 5741 13913 ne
rect 5741 13833 6113 13913
tri 6113 13833 6193 13913 sw
tri 6211 13833 6291 13913 ne
rect 6291 13833 6663 13913
tri 6663 13833 6743 13913 sw
tri 6761 13833 6841 13913 ne
rect 6841 13833 7213 13913
tri 7213 13833 7293 13913 sw
tri 7311 13833 7391 13913 ne
rect 7391 13833 7763 13913
tri 7763 13833 7843 13913 sw
tri 7861 13833 7941 13913 ne
rect 7941 13833 8313 13913
tri 8313 13833 8393 13913 sw
tri 8411 13833 8491 13913 ne
rect 8491 13833 8863 13913
tri 8863 13833 8943 13913 sw
tri 8961 13833 9041 13913 ne
rect 9041 13833 9413 13913
tri 9413 13833 9493 13913 sw
tri 9511 13833 9591 13913 ne
rect 9591 13833 9963 13913
tri 9963 13833 10043 13913 sw
tri 10061 13833 10141 13913 ne
rect 10141 13833 10513 13913
tri 10513 13833 10593 13913 sw
tri 10611 13833 10691 13913 ne
rect 10691 13833 11063 13913
tri 11063 13833 11143 13913 sw
tri 11161 13833 11241 13913 ne
rect 11241 13833 11613 13913
tri 11613 13833 11693 13913 sw
tri 11711 13833 11791 13913 ne
rect 11791 13833 12163 13913
tri 12163 13833 12243 13913 sw
tri 12261 13833 12341 13913 ne
rect 12341 13833 12713 13913
tri 12713 13833 12793 13913 sw
tri 12811 13833 12891 13913 ne
rect 12891 13833 13263 13913
tri 13263 13833 13343 13913 sw
tri 13361 13833 13441 13913 ne
rect 13441 13833 13813 13913
tri 13813 13833 13893 13913 sw
tri 13911 13833 13991 13913 ne
rect 13991 13833 14363 13913
tri 14363 13833 14443 13913 sw
tri 14461 13833 14541 13913 ne
rect 14541 13833 14913 13913
tri 14913 13833 14993 13913 sw
tri 15011 13833 15091 13913 ne
rect 15091 13833 15463 13913
tri 15463 13833 15543 13913 sw
tri 15561 13833 15641 13913 ne
rect 15641 13833 16013 13913
tri 16013 13833 16093 13913 sw
tri 16111 13833 16191 13913 ne
rect 16191 13833 16563 13913
tri 16563 13833 16643 13913 sw
tri 16661 13833 16741 13913 ne
rect 16741 13833 17113 13913
tri 17113 13833 17193 13913 sw
tri 17211 13833 17291 13913 ne
rect 17291 13833 17663 13913
tri 17663 13833 17743 13913 sw
tri 17761 13833 17841 13913 ne
rect 17841 13833 18213 13913
tri 18213 13833 18293 13913 sw
tri 18311 13833 18391 13913 ne
rect 18391 13833 18763 13913
tri 18763 13833 18843 13913 sw
tri 18861 13833 18941 13913 ne
rect 18941 13833 19313 13913
tri 19313 13833 19393 13913 sw
tri 19411 13833 19491 13913 ne
rect 19491 13833 20100 13913
rect 261 13813 693 13833
rect -500 13735 163 13813
tri 163 13735 241 13813 sw
tri 261 13735 339 13813 ne
rect 339 13735 693 13813
tri 693 13735 791 13833 sw
tri 791 13735 889 13833 ne
rect 889 13735 1243 13833
tri 1243 13735 1341 13833 sw
tri 1341 13735 1439 13833 ne
rect 1439 13735 1793 13833
tri 1793 13735 1891 13833 sw
tri 1891 13735 1989 13833 ne
rect 1989 13735 2343 13833
tri 2343 13735 2441 13833 sw
tri 2441 13735 2539 13833 ne
rect 2539 13735 2893 13833
tri 2893 13735 2991 13833 sw
tri 2991 13735 3089 13833 ne
rect 3089 13735 3443 13833
tri 3443 13735 3541 13833 sw
tri 3541 13735 3639 13833 ne
rect 3639 13735 3993 13833
tri 3993 13735 4091 13833 sw
tri 4091 13735 4189 13833 ne
rect 4189 13735 4543 13833
tri 4543 13735 4641 13833 sw
tri 4641 13735 4739 13833 ne
rect 4739 13735 5093 13833
tri 5093 13735 5191 13833 sw
tri 5191 13735 5289 13833 ne
rect 5289 13735 5643 13833
tri 5643 13735 5741 13833 sw
tri 5741 13735 5839 13833 ne
rect 5839 13735 6193 13833
tri 6193 13735 6291 13833 sw
tri 6291 13735 6389 13833 ne
rect 6389 13735 6743 13833
tri 6743 13735 6841 13833 sw
tri 6841 13735 6939 13833 ne
rect 6939 13735 7293 13833
tri 7293 13735 7391 13833 sw
tri 7391 13735 7489 13833 ne
rect 7489 13735 7843 13833
tri 7843 13735 7941 13833 sw
tri 7941 13735 8039 13833 ne
rect 8039 13735 8393 13833
tri 8393 13735 8491 13833 sw
tri 8491 13735 8589 13833 ne
rect 8589 13735 8943 13833
tri 8943 13735 9041 13833 sw
tri 9041 13735 9139 13833 ne
rect 9139 13735 9493 13833
tri 9493 13735 9591 13833 sw
tri 9591 13735 9689 13833 ne
rect 9689 13735 10043 13833
tri 10043 13735 10141 13833 sw
tri 10141 13735 10239 13833 ne
rect 10239 13735 10593 13833
tri 10593 13735 10691 13833 sw
tri 10691 13735 10789 13833 ne
rect 10789 13735 11143 13833
tri 11143 13735 11241 13833 sw
tri 11241 13735 11339 13833 ne
rect 11339 13735 11693 13833
tri 11693 13735 11791 13833 sw
tri 11791 13735 11889 13833 ne
rect 11889 13735 12243 13833
tri 12243 13735 12341 13833 sw
tri 12341 13735 12439 13833 ne
rect 12439 13735 12793 13833
tri 12793 13735 12891 13833 sw
tri 12891 13735 12989 13833 ne
rect 12989 13735 13343 13833
tri 13343 13735 13441 13833 sw
tri 13441 13735 13539 13833 ne
rect 13539 13735 13893 13833
tri 13893 13735 13991 13833 sw
tri 13991 13735 14089 13833 ne
rect 14089 13735 14443 13833
tri 14443 13735 14541 13833 sw
tri 14541 13735 14639 13833 ne
rect 14639 13735 14993 13833
tri 14993 13735 15091 13833 sw
tri 15091 13735 15189 13833 ne
rect 15189 13735 15543 13833
tri 15543 13735 15641 13833 sw
tri 15641 13735 15739 13833 ne
rect 15739 13735 16093 13833
tri 16093 13735 16191 13833 sw
tri 16191 13735 16289 13833 ne
rect 16289 13735 16643 13833
tri 16643 13735 16741 13833 sw
tri 16741 13735 16839 13833 ne
rect 16839 13735 17193 13833
tri 17193 13735 17291 13833 sw
tri 17291 13735 17389 13833 ne
rect 17389 13735 17743 13833
tri 17743 13735 17841 13833 sw
tri 17841 13735 17939 13833 ne
rect 17939 13735 18293 13833
tri 18293 13735 18391 13833 sw
tri 18391 13735 18489 13833 ne
rect 18489 13735 18843 13833
tri 18843 13735 18941 13833 sw
tri 18941 13735 19039 13833 ne
rect 19039 13735 19393 13833
tri 19393 13735 19491 13833 sw
tri 19491 13735 19589 13833 ne
rect 19589 13813 20100 13833
rect 20200 13813 21800 13913
rect 19589 13735 21800 13813
rect -500 13687 241 13735
rect -500 13587 -400 13687
rect -300 13637 241 13687
tri 241 13637 339 13735 sw
tri 339 13637 437 13735 ne
rect 437 13637 791 13735
tri 791 13637 889 13735 sw
tri 889 13637 987 13735 ne
rect 987 13637 1341 13735
tri 1341 13637 1439 13735 sw
tri 1439 13637 1537 13735 ne
rect 1537 13637 1891 13735
tri 1891 13637 1989 13735 sw
tri 1989 13637 2087 13735 ne
rect 2087 13637 2441 13735
tri 2441 13637 2539 13735 sw
tri 2539 13637 2637 13735 ne
rect 2637 13637 2991 13735
tri 2991 13637 3089 13735 sw
tri 3089 13637 3187 13735 ne
rect 3187 13637 3541 13735
tri 3541 13637 3639 13735 sw
tri 3639 13637 3737 13735 ne
rect 3737 13637 4091 13735
tri 4091 13637 4189 13735 sw
tri 4189 13637 4287 13735 ne
rect 4287 13637 4641 13735
tri 4641 13637 4739 13735 sw
tri 4739 13637 4837 13735 ne
rect 4837 13637 5191 13735
tri 5191 13637 5289 13735 sw
tri 5289 13637 5387 13735 ne
rect 5387 13637 5741 13735
tri 5741 13637 5839 13735 sw
tri 5839 13637 5937 13735 ne
rect 5937 13637 6291 13735
tri 6291 13637 6389 13735 sw
tri 6389 13637 6487 13735 ne
rect 6487 13637 6841 13735
tri 6841 13637 6939 13735 sw
tri 6939 13637 7037 13735 ne
rect 7037 13637 7391 13735
tri 7391 13637 7489 13735 sw
tri 7489 13637 7587 13735 ne
rect 7587 13637 7941 13735
tri 7941 13637 8039 13735 sw
tri 8039 13637 8137 13735 ne
rect 8137 13637 8491 13735
tri 8491 13637 8589 13735 sw
tri 8589 13637 8687 13735 ne
rect 8687 13637 9041 13735
tri 9041 13637 9139 13735 sw
tri 9139 13637 9237 13735 ne
rect 9237 13637 9591 13735
tri 9591 13637 9689 13735 sw
tri 9689 13637 9787 13735 ne
rect 9787 13637 10141 13735
tri 10141 13637 10239 13735 sw
tri 10239 13637 10337 13735 ne
rect 10337 13637 10691 13735
tri 10691 13637 10789 13735 sw
tri 10789 13637 10887 13735 ne
rect 10887 13637 11241 13735
tri 11241 13637 11339 13735 sw
tri 11339 13637 11437 13735 ne
rect 11437 13637 11791 13735
tri 11791 13637 11889 13735 sw
tri 11889 13637 11987 13735 ne
rect 11987 13637 12341 13735
tri 12341 13637 12439 13735 sw
tri 12439 13637 12537 13735 ne
rect 12537 13637 12891 13735
tri 12891 13637 12989 13735 sw
tri 12989 13637 13087 13735 ne
rect 13087 13637 13441 13735
tri 13441 13637 13539 13735 sw
tri 13539 13637 13637 13735 ne
rect 13637 13637 13991 13735
tri 13991 13637 14089 13735 sw
tri 14089 13637 14187 13735 ne
rect 14187 13637 14541 13735
tri 14541 13637 14639 13735 sw
tri 14639 13637 14737 13735 ne
rect 14737 13637 15091 13735
tri 15091 13637 15189 13735 sw
tri 15189 13637 15287 13735 ne
rect 15287 13637 15641 13735
tri 15641 13637 15739 13735 sw
tri 15739 13637 15837 13735 ne
rect 15837 13637 16191 13735
tri 16191 13637 16289 13735 sw
tri 16289 13637 16387 13735 ne
rect 16387 13637 16741 13735
tri 16741 13637 16839 13735 sw
tri 16839 13637 16937 13735 ne
rect 16937 13637 17291 13735
tri 17291 13637 17389 13735 sw
tri 17389 13637 17487 13735 ne
rect 17487 13637 17841 13735
tri 17841 13637 17939 13735 sw
tri 17939 13637 18037 13735 ne
rect 18037 13637 18391 13735
tri 18391 13637 18489 13735 sw
tri 18489 13637 18587 13735 ne
rect 18587 13637 18941 13735
tri 18941 13637 19039 13735 sw
tri 19039 13637 19137 13735 ne
rect 19137 13637 19491 13735
tri 19491 13637 19589 13735 sw
tri 19589 13637 19687 13735 ne
rect 19687 13637 21800 13735
rect -300 13587 339 13637
rect -500 13539 339 13587
tri 339 13539 437 13637 sw
tri 437 13539 535 13637 ne
rect 535 13539 889 13637
tri 889 13539 987 13637 sw
tri 987 13539 1085 13637 ne
rect 1085 13539 1439 13637
tri 1439 13539 1537 13637 sw
tri 1537 13539 1635 13637 ne
rect 1635 13539 1989 13637
tri 1989 13539 2087 13637 sw
tri 2087 13539 2185 13637 ne
rect 2185 13539 2539 13637
tri 2539 13539 2637 13637 sw
tri 2637 13539 2735 13637 ne
rect 2735 13539 3089 13637
tri 3089 13539 3187 13637 sw
tri 3187 13539 3285 13637 ne
rect 3285 13539 3639 13637
tri 3639 13539 3737 13637 sw
tri 3737 13539 3835 13637 ne
rect 3835 13539 4189 13637
tri 4189 13539 4287 13637 sw
tri 4287 13539 4385 13637 ne
rect 4385 13539 4739 13637
tri 4739 13539 4837 13637 sw
tri 4837 13539 4935 13637 ne
rect 4935 13539 5289 13637
tri 5289 13539 5387 13637 sw
tri 5387 13539 5485 13637 ne
rect 5485 13539 5839 13637
tri 5839 13539 5937 13637 sw
tri 5937 13539 6035 13637 ne
rect 6035 13539 6389 13637
tri 6389 13539 6487 13637 sw
tri 6487 13539 6585 13637 ne
rect 6585 13539 6939 13637
tri 6939 13539 7037 13637 sw
tri 7037 13539 7135 13637 ne
rect 7135 13539 7489 13637
tri 7489 13539 7587 13637 sw
tri 7587 13539 7685 13637 ne
rect 7685 13539 8039 13637
tri 8039 13539 8137 13637 sw
tri 8137 13539 8235 13637 ne
rect 8235 13539 8589 13637
tri 8589 13539 8687 13637 sw
tri 8687 13539 8785 13637 ne
rect 8785 13539 9139 13637
tri 9139 13539 9237 13637 sw
tri 9237 13539 9335 13637 ne
rect 9335 13539 9689 13637
tri 9689 13539 9787 13637 sw
tri 9787 13539 9885 13637 ne
rect 9885 13539 10239 13637
tri 10239 13539 10337 13637 sw
tri 10337 13539 10435 13637 ne
rect 10435 13539 10789 13637
tri 10789 13539 10887 13637 sw
tri 10887 13539 10985 13637 ne
rect 10985 13539 11339 13637
tri 11339 13539 11437 13637 sw
tri 11437 13539 11535 13637 ne
rect 11535 13539 11889 13637
tri 11889 13539 11987 13637 sw
tri 11987 13539 12085 13637 ne
rect 12085 13539 12439 13637
tri 12439 13539 12537 13637 sw
tri 12537 13539 12635 13637 ne
rect 12635 13539 12989 13637
tri 12989 13539 13087 13637 sw
tri 13087 13539 13185 13637 ne
rect 13185 13539 13539 13637
tri 13539 13539 13637 13637 sw
tri 13637 13539 13735 13637 ne
rect 13735 13539 14089 13637
tri 14089 13539 14187 13637 sw
tri 14187 13539 14285 13637 ne
rect 14285 13539 14639 13637
tri 14639 13539 14737 13637 sw
tri 14737 13539 14835 13637 ne
rect 14835 13539 15189 13637
tri 15189 13539 15287 13637 sw
tri 15287 13539 15385 13637 ne
rect 15385 13539 15739 13637
tri 15739 13539 15837 13637 sw
tri 15837 13539 15935 13637 ne
rect 15935 13539 16289 13637
tri 16289 13539 16387 13637 sw
tri 16387 13539 16485 13637 ne
rect 16485 13539 16839 13637
tri 16839 13539 16937 13637 sw
tri 16937 13539 17035 13637 ne
rect 17035 13539 17389 13637
tri 17389 13539 17487 13637 sw
tri 17487 13539 17585 13637 ne
rect 17585 13539 17939 13637
tri 17939 13539 18037 13637 sw
tri 18037 13539 18135 13637 ne
rect 18135 13539 18489 13637
tri 18489 13539 18587 13637 sw
tri 18587 13539 18685 13637 ne
rect 18685 13539 19039 13637
tri 19039 13539 19137 13637 sw
tri 19137 13539 19235 13637 ne
rect 19235 13539 19589 13637
tri 19589 13539 19687 13637 sw
rect -500 13535 437 13539
rect -500 13415 215 13535
rect 335 13441 437 13535
tri 437 13441 535 13539 sw
tri 535 13441 633 13539 ne
rect 633 13535 987 13539
rect 633 13441 765 13535
rect 335 13415 535 13441
rect -500 13411 535 13415
tri 535 13411 565 13441 sw
tri 633 13411 663 13441 ne
rect 663 13415 765 13441
rect 885 13441 987 13535
tri 987 13441 1085 13539 sw
tri 1085 13441 1183 13539 ne
rect 1183 13535 1537 13539
rect 1183 13441 1315 13535
rect 885 13415 1085 13441
rect 663 13411 1085 13415
tri 1085 13411 1115 13441 sw
tri 1183 13411 1213 13441 ne
rect 1213 13415 1315 13441
rect 1435 13441 1537 13535
tri 1537 13441 1635 13539 sw
tri 1635 13441 1733 13539 ne
rect 1733 13535 2087 13539
rect 1733 13441 1865 13535
rect 1435 13415 1635 13441
rect 1213 13411 1635 13415
tri 1635 13411 1665 13441 sw
tri 1733 13411 1763 13441 ne
rect 1763 13415 1865 13441
rect 1985 13441 2087 13535
tri 2087 13441 2185 13539 sw
tri 2185 13441 2283 13539 ne
rect 2283 13535 2637 13539
rect 2283 13441 2415 13535
rect 1985 13415 2185 13441
rect 1763 13411 2185 13415
tri 2185 13411 2215 13441 sw
tri 2283 13411 2313 13441 ne
rect 2313 13415 2415 13441
rect 2535 13441 2637 13535
tri 2637 13441 2735 13539 sw
tri 2735 13441 2833 13539 ne
rect 2833 13535 3187 13539
rect 2833 13441 2965 13535
rect 2535 13415 2735 13441
rect 2313 13411 2735 13415
tri 2735 13411 2765 13441 sw
tri 2833 13411 2863 13441 ne
rect 2863 13415 2965 13441
rect 3085 13441 3187 13535
tri 3187 13441 3285 13539 sw
tri 3285 13441 3383 13539 ne
rect 3383 13535 3737 13539
rect 3383 13441 3515 13535
rect 3085 13415 3285 13441
rect 2863 13411 3285 13415
tri 3285 13411 3315 13441 sw
tri 3383 13411 3413 13441 ne
rect 3413 13415 3515 13441
rect 3635 13441 3737 13535
tri 3737 13441 3835 13539 sw
tri 3835 13441 3933 13539 ne
rect 3933 13535 4287 13539
rect 3933 13441 4065 13535
rect 3635 13415 3835 13441
rect 3413 13411 3835 13415
tri 3835 13411 3865 13441 sw
tri 3933 13411 3963 13441 ne
rect 3963 13415 4065 13441
rect 4185 13441 4287 13535
tri 4287 13441 4385 13539 sw
tri 4385 13441 4483 13539 ne
rect 4483 13535 4837 13539
rect 4483 13441 4615 13535
rect 4185 13415 4385 13441
rect 3963 13411 4385 13415
tri 4385 13411 4415 13441 sw
tri 4483 13411 4513 13441 ne
rect 4513 13415 4615 13441
rect 4735 13441 4837 13535
tri 4837 13441 4935 13539 sw
tri 4935 13441 5033 13539 ne
rect 5033 13535 5387 13539
rect 5033 13441 5165 13535
rect 4735 13415 4935 13441
rect 4513 13411 4935 13415
tri 4935 13411 4965 13441 sw
tri 5033 13411 5063 13441 ne
rect 5063 13415 5165 13441
rect 5285 13441 5387 13535
tri 5387 13441 5485 13539 sw
tri 5485 13441 5583 13539 ne
rect 5583 13535 5937 13539
rect 5583 13441 5715 13535
rect 5285 13415 5485 13441
rect 5063 13411 5485 13415
tri 5485 13411 5515 13441 sw
tri 5583 13411 5613 13441 ne
rect 5613 13415 5715 13441
rect 5835 13441 5937 13535
tri 5937 13441 6035 13539 sw
tri 6035 13441 6133 13539 ne
rect 6133 13535 6487 13539
rect 6133 13441 6265 13535
rect 5835 13415 6035 13441
rect 5613 13411 6035 13415
tri 6035 13411 6065 13441 sw
tri 6133 13411 6163 13441 ne
rect 6163 13415 6265 13441
rect 6385 13441 6487 13535
tri 6487 13441 6585 13539 sw
tri 6585 13441 6683 13539 ne
rect 6683 13535 7037 13539
rect 6683 13441 6815 13535
rect 6385 13415 6585 13441
rect 6163 13411 6585 13415
tri 6585 13411 6615 13441 sw
tri 6683 13411 6713 13441 ne
rect 6713 13415 6815 13441
rect 6935 13441 7037 13535
tri 7037 13441 7135 13539 sw
tri 7135 13441 7233 13539 ne
rect 7233 13535 7587 13539
rect 7233 13441 7365 13535
rect 6935 13415 7135 13441
rect 6713 13411 7135 13415
tri 7135 13411 7165 13441 sw
tri 7233 13411 7263 13441 ne
rect 7263 13415 7365 13441
rect 7485 13441 7587 13535
tri 7587 13441 7685 13539 sw
tri 7685 13441 7783 13539 ne
rect 7783 13535 8137 13539
rect 7783 13441 7915 13535
rect 7485 13415 7685 13441
rect 7263 13411 7685 13415
tri 7685 13411 7715 13441 sw
tri 7783 13411 7813 13441 ne
rect 7813 13415 7915 13441
rect 8035 13441 8137 13535
tri 8137 13441 8235 13539 sw
tri 8235 13441 8333 13539 ne
rect 8333 13535 8687 13539
rect 8333 13441 8465 13535
rect 8035 13415 8235 13441
rect 7813 13411 8235 13415
tri 8235 13411 8265 13441 sw
tri 8333 13411 8363 13441 ne
rect 8363 13415 8465 13441
rect 8585 13441 8687 13535
tri 8687 13441 8785 13539 sw
tri 8785 13441 8883 13539 ne
rect 8883 13535 9237 13539
rect 8883 13441 9015 13535
rect 8585 13415 8785 13441
rect 8363 13411 8785 13415
tri 8785 13411 8815 13441 sw
tri 8883 13411 8913 13441 ne
rect 8913 13415 9015 13441
rect 9135 13441 9237 13535
tri 9237 13441 9335 13539 sw
tri 9335 13441 9433 13539 ne
rect 9433 13535 9787 13539
rect 9433 13441 9565 13535
rect 9135 13415 9335 13441
rect 8913 13411 9335 13415
tri 9335 13411 9365 13441 sw
tri 9433 13411 9463 13441 ne
rect 9463 13415 9565 13441
rect 9685 13441 9787 13535
tri 9787 13441 9885 13539 sw
tri 9885 13441 9983 13539 ne
rect 9983 13535 10337 13539
rect 9983 13441 10115 13535
rect 9685 13415 9885 13441
rect 9463 13411 9885 13415
tri 9885 13411 9915 13441 sw
tri 9983 13411 10013 13441 ne
rect 10013 13415 10115 13441
rect 10235 13441 10337 13535
tri 10337 13441 10435 13539 sw
tri 10435 13441 10533 13539 ne
rect 10533 13535 10887 13539
rect 10533 13441 10665 13535
rect 10235 13415 10435 13441
rect 10013 13411 10435 13415
tri 10435 13411 10465 13441 sw
tri 10533 13411 10563 13441 ne
rect 10563 13415 10665 13441
rect 10785 13441 10887 13535
tri 10887 13441 10985 13539 sw
tri 10985 13441 11083 13539 ne
rect 11083 13535 11437 13539
rect 11083 13441 11215 13535
rect 10785 13415 10985 13441
rect 10563 13411 10985 13415
tri 10985 13411 11015 13441 sw
tri 11083 13411 11113 13441 ne
rect 11113 13415 11215 13441
rect 11335 13441 11437 13535
tri 11437 13441 11535 13539 sw
tri 11535 13441 11633 13539 ne
rect 11633 13535 11987 13539
rect 11633 13441 11765 13535
rect 11335 13415 11535 13441
rect 11113 13411 11535 13415
tri 11535 13411 11565 13441 sw
tri 11633 13411 11663 13441 ne
rect 11663 13415 11765 13441
rect 11885 13441 11987 13535
tri 11987 13441 12085 13539 sw
tri 12085 13441 12183 13539 ne
rect 12183 13535 12537 13539
rect 12183 13441 12315 13535
rect 11885 13415 12085 13441
rect 11663 13411 12085 13415
tri 12085 13411 12115 13441 sw
tri 12183 13411 12213 13441 ne
rect 12213 13415 12315 13441
rect 12435 13441 12537 13535
tri 12537 13441 12635 13539 sw
tri 12635 13441 12733 13539 ne
rect 12733 13535 13087 13539
rect 12733 13441 12865 13535
rect 12435 13415 12635 13441
rect 12213 13411 12635 13415
tri 12635 13411 12665 13441 sw
tri 12733 13411 12763 13441 ne
rect 12763 13415 12865 13441
rect 12985 13441 13087 13535
tri 13087 13441 13185 13539 sw
tri 13185 13441 13283 13539 ne
rect 13283 13535 13637 13539
rect 13283 13441 13415 13535
rect 12985 13415 13185 13441
rect 12763 13411 13185 13415
tri 13185 13411 13215 13441 sw
tri 13283 13411 13313 13441 ne
rect 13313 13415 13415 13441
rect 13535 13441 13637 13535
tri 13637 13441 13735 13539 sw
tri 13735 13441 13833 13539 ne
rect 13833 13535 14187 13539
rect 13833 13441 13965 13535
rect 13535 13415 13735 13441
rect 13313 13411 13735 13415
tri 13735 13411 13765 13441 sw
tri 13833 13411 13863 13441 ne
rect 13863 13415 13965 13441
rect 14085 13441 14187 13535
tri 14187 13441 14285 13539 sw
tri 14285 13441 14383 13539 ne
rect 14383 13535 14737 13539
rect 14383 13441 14515 13535
rect 14085 13415 14285 13441
rect 13863 13411 14285 13415
tri 14285 13411 14315 13441 sw
tri 14383 13411 14413 13441 ne
rect 14413 13415 14515 13441
rect 14635 13441 14737 13535
tri 14737 13441 14835 13539 sw
tri 14835 13441 14933 13539 ne
rect 14933 13535 15287 13539
rect 14933 13441 15065 13535
rect 14635 13415 14835 13441
rect 14413 13411 14835 13415
tri 14835 13411 14865 13441 sw
tri 14933 13411 14963 13441 ne
rect 14963 13415 15065 13441
rect 15185 13441 15287 13535
tri 15287 13441 15385 13539 sw
tri 15385 13441 15483 13539 ne
rect 15483 13535 15837 13539
rect 15483 13441 15615 13535
rect 15185 13415 15385 13441
rect 14963 13411 15385 13415
tri 15385 13411 15415 13441 sw
tri 15483 13411 15513 13441 ne
rect 15513 13415 15615 13441
rect 15735 13441 15837 13535
tri 15837 13441 15935 13539 sw
tri 15935 13441 16033 13539 ne
rect 16033 13535 16387 13539
rect 16033 13441 16165 13535
rect 15735 13415 15935 13441
rect 15513 13411 15935 13415
tri 15935 13411 15965 13441 sw
tri 16033 13411 16063 13441 ne
rect 16063 13415 16165 13441
rect 16285 13441 16387 13535
tri 16387 13441 16485 13539 sw
tri 16485 13441 16583 13539 ne
rect 16583 13535 16937 13539
rect 16583 13441 16715 13535
rect 16285 13415 16485 13441
rect 16063 13411 16485 13415
tri 16485 13411 16515 13441 sw
tri 16583 13411 16613 13441 ne
rect 16613 13415 16715 13441
rect 16835 13441 16937 13535
tri 16937 13441 17035 13539 sw
tri 17035 13441 17133 13539 ne
rect 17133 13535 17487 13539
rect 17133 13441 17265 13535
rect 16835 13415 17035 13441
rect 16613 13411 17035 13415
tri 17035 13411 17065 13441 sw
tri 17133 13411 17163 13441 ne
rect 17163 13415 17265 13441
rect 17385 13441 17487 13535
tri 17487 13441 17585 13539 sw
tri 17585 13441 17683 13539 ne
rect 17683 13535 18037 13539
rect 17683 13441 17815 13535
rect 17385 13415 17585 13441
rect 17163 13411 17585 13415
tri 17585 13411 17615 13441 sw
tri 17683 13411 17713 13441 ne
rect 17713 13415 17815 13441
rect 17935 13441 18037 13535
tri 18037 13441 18135 13539 sw
tri 18135 13441 18233 13539 ne
rect 18233 13535 18587 13539
rect 18233 13441 18365 13535
rect 17935 13415 18135 13441
rect 17713 13411 18135 13415
tri 18135 13411 18165 13441 sw
tri 18233 13411 18263 13441 ne
rect 18263 13415 18365 13441
rect 18485 13441 18587 13535
tri 18587 13441 18685 13539 sw
tri 18685 13441 18783 13539 ne
rect 18783 13535 19137 13539
rect 18783 13441 18915 13535
rect 18485 13415 18685 13441
rect 18263 13411 18685 13415
tri 18685 13411 18715 13441 sw
tri 18783 13411 18813 13441 ne
rect 18813 13415 18915 13441
rect 19035 13441 19137 13535
tri 19137 13441 19235 13539 sw
tri 19235 13441 19333 13539 ne
rect 19333 13535 20300 13539
rect 19333 13441 19465 13535
rect 19035 13415 19235 13441
rect 18813 13411 19235 13415
tri 19235 13411 19265 13441 sw
tri 19333 13411 19363 13441 ne
rect 19363 13415 19465 13441
rect 19585 13415 20300 13535
rect 19363 13411 20300 13415
tri 113 13313 211 13411 ne
rect 211 13313 565 13411
tri 565 13313 663 13411 sw
tri 663 13313 761 13411 ne
rect 761 13313 1115 13411
tri 1115 13313 1213 13411 sw
tri 1213 13313 1311 13411 ne
rect 1311 13313 1665 13411
tri 1665 13313 1763 13411 sw
tri 1763 13313 1861 13411 ne
rect 1861 13313 2215 13411
tri 2215 13313 2313 13411 sw
tri 2313 13313 2411 13411 ne
rect 2411 13313 2765 13411
tri 2765 13313 2863 13411 sw
tri 2863 13313 2961 13411 ne
rect 2961 13313 3315 13411
tri 3315 13313 3413 13411 sw
tri 3413 13313 3511 13411 ne
rect 3511 13313 3865 13411
tri 3865 13313 3963 13411 sw
tri 3963 13313 4061 13411 ne
rect 4061 13313 4415 13411
tri 4415 13313 4513 13411 sw
tri 4513 13313 4611 13411 ne
rect 4611 13313 4965 13411
tri 4965 13313 5063 13411 sw
tri 5063 13313 5161 13411 ne
rect 5161 13313 5515 13411
tri 5515 13313 5613 13411 sw
tri 5613 13313 5711 13411 ne
rect 5711 13313 6065 13411
tri 6065 13313 6163 13411 sw
tri 6163 13313 6261 13411 ne
rect 6261 13313 6615 13411
tri 6615 13313 6713 13411 sw
tri 6713 13313 6811 13411 ne
rect 6811 13313 7165 13411
tri 7165 13313 7263 13411 sw
tri 7263 13313 7361 13411 ne
rect 7361 13313 7715 13411
tri 7715 13313 7813 13411 sw
tri 7813 13313 7911 13411 ne
rect 7911 13313 8265 13411
tri 8265 13313 8363 13411 sw
tri 8363 13313 8461 13411 ne
rect 8461 13313 8815 13411
tri 8815 13313 8913 13411 sw
tri 8913 13313 9011 13411 ne
rect 9011 13313 9365 13411
tri 9365 13313 9463 13411 sw
tri 9463 13313 9561 13411 ne
rect 9561 13313 9915 13411
tri 9915 13313 10013 13411 sw
tri 10013 13313 10111 13411 ne
rect 10111 13313 10465 13411
tri 10465 13313 10563 13411 sw
tri 10563 13313 10661 13411 ne
rect 10661 13313 11015 13411
tri 11015 13313 11113 13411 sw
tri 11113 13313 11211 13411 ne
rect 11211 13313 11565 13411
tri 11565 13313 11663 13411 sw
tri 11663 13313 11761 13411 ne
rect 11761 13313 12115 13411
tri 12115 13313 12213 13411 sw
tri 12213 13313 12311 13411 ne
rect 12311 13313 12665 13411
tri 12665 13313 12763 13411 sw
tri 12763 13313 12861 13411 ne
rect 12861 13313 13215 13411
tri 13215 13313 13313 13411 sw
tri 13313 13313 13411 13411 ne
rect 13411 13313 13765 13411
tri 13765 13313 13863 13411 sw
tri 13863 13313 13961 13411 ne
rect 13961 13313 14315 13411
tri 14315 13313 14413 13411 sw
tri 14413 13313 14511 13411 ne
rect 14511 13313 14865 13411
tri 14865 13313 14963 13411 sw
tri 14963 13313 15061 13411 ne
rect 15061 13313 15415 13411
tri 15415 13313 15513 13411 sw
tri 15513 13313 15611 13411 ne
rect 15611 13313 15965 13411
tri 15965 13313 16063 13411 sw
tri 16063 13313 16161 13411 ne
rect 16161 13313 16515 13411
tri 16515 13313 16613 13411 sw
tri 16613 13313 16711 13411 ne
rect 16711 13313 17065 13411
tri 17065 13313 17163 13411 sw
tri 17163 13313 17261 13411 ne
rect 17261 13313 17615 13411
tri 17615 13313 17713 13411 sw
tri 17713 13313 17811 13411 ne
rect 17811 13313 18165 13411
tri 18165 13313 18263 13411 sw
tri 18263 13313 18361 13411 ne
rect 18361 13313 18715 13411
tri 18715 13313 18813 13411 sw
tri 18813 13313 18911 13411 ne
rect 18911 13313 19265 13411
tri 19265 13313 19363 13411 sw
tri 19363 13313 19461 13411 ne
rect 19461 13313 20300 13411
rect -2000 13283 113 13313
tri 113 13283 143 13313 sw
tri 211 13283 241 13313 ne
rect 241 13283 663 13313
tri 663 13283 693 13313 sw
tri 761 13283 791 13313 ne
rect 791 13283 1213 13313
tri 1213 13283 1243 13313 sw
tri 1311 13283 1341 13313 ne
rect 1341 13283 1763 13313
tri 1763 13283 1793 13313 sw
tri 1861 13283 1891 13313 ne
rect 1891 13283 2313 13313
tri 2313 13283 2343 13313 sw
tri 2411 13283 2441 13313 ne
rect 2441 13283 2863 13313
tri 2863 13283 2893 13313 sw
tri 2961 13283 2991 13313 ne
rect 2991 13283 3413 13313
tri 3413 13283 3443 13313 sw
tri 3511 13283 3541 13313 ne
rect 3541 13283 3963 13313
tri 3963 13283 3993 13313 sw
tri 4061 13283 4091 13313 ne
rect 4091 13283 4513 13313
tri 4513 13283 4543 13313 sw
tri 4611 13283 4641 13313 ne
rect 4641 13283 5063 13313
tri 5063 13283 5093 13313 sw
tri 5161 13283 5191 13313 ne
rect 5191 13283 5613 13313
tri 5613 13283 5643 13313 sw
tri 5711 13283 5741 13313 ne
rect 5741 13283 6163 13313
tri 6163 13283 6193 13313 sw
tri 6261 13283 6291 13313 ne
rect 6291 13283 6713 13313
tri 6713 13283 6743 13313 sw
tri 6811 13283 6841 13313 ne
rect 6841 13283 7263 13313
tri 7263 13283 7293 13313 sw
tri 7361 13283 7391 13313 ne
rect 7391 13283 7813 13313
tri 7813 13283 7843 13313 sw
tri 7911 13283 7941 13313 ne
rect 7941 13283 8363 13313
tri 8363 13283 8393 13313 sw
tri 8461 13283 8491 13313 ne
rect 8491 13283 8913 13313
tri 8913 13283 8943 13313 sw
tri 9011 13283 9041 13313 ne
rect 9041 13283 9463 13313
tri 9463 13283 9493 13313 sw
tri 9561 13283 9591 13313 ne
rect 9591 13283 10013 13313
tri 10013 13283 10043 13313 sw
tri 10111 13283 10141 13313 ne
rect 10141 13283 10563 13313
tri 10563 13283 10593 13313 sw
tri 10661 13283 10691 13313 ne
rect 10691 13283 11113 13313
tri 11113 13283 11143 13313 sw
tri 11211 13283 11241 13313 ne
rect 11241 13283 11663 13313
tri 11663 13283 11693 13313 sw
tri 11761 13283 11791 13313 ne
rect 11791 13283 12213 13313
tri 12213 13283 12243 13313 sw
tri 12311 13283 12341 13313 ne
rect 12341 13283 12763 13313
tri 12763 13283 12793 13313 sw
tri 12861 13283 12891 13313 ne
rect 12891 13283 13313 13313
tri 13313 13283 13343 13313 sw
tri 13411 13283 13441 13313 ne
rect 13441 13283 13863 13313
tri 13863 13283 13893 13313 sw
tri 13961 13283 13991 13313 ne
rect 13991 13283 14413 13313
tri 14413 13283 14443 13313 sw
tri 14511 13283 14541 13313 ne
rect 14541 13283 14963 13313
tri 14963 13283 14993 13313 sw
tri 15061 13283 15091 13313 ne
rect 15091 13283 15513 13313
tri 15513 13283 15543 13313 sw
tri 15611 13283 15641 13313 ne
rect 15641 13283 16063 13313
tri 16063 13283 16093 13313 sw
tri 16161 13283 16191 13313 ne
rect 16191 13283 16613 13313
tri 16613 13283 16643 13313 sw
tri 16711 13283 16741 13313 ne
rect 16741 13283 17163 13313
tri 17163 13283 17193 13313 sw
tri 17261 13283 17291 13313 ne
rect 17291 13283 17713 13313
tri 17713 13283 17743 13313 sw
tri 17811 13283 17841 13313 ne
rect 17841 13283 18263 13313
tri 18263 13283 18293 13313 sw
tri 18361 13283 18391 13313 ne
rect 18391 13283 18813 13313
tri 18813 13283 18843 13313 sw
tri 18911 13283 18941 13313 ne
rect 18941 13283 19363 13313
tri 19363 13283 19393 13313 sw
tri 19461 13283 19491 13313 ne
rect 19491 13283 20300 13313
rect -2000 13185 143 13283
tri 143 13185 241 13283 sw
tri 241 13185 339 13283 ne
rect 339 13185 693 13283
tri 693 13185 791 13283 sw
tri 791 13185 889 13283 ne
rect 889 13185 1243 13283
tri 1243 13185 1341 13283 sw
tri 1341 13185 1439 13283 ne
rect 1439 13185 1793 13283
tri 1793 13185 1891 13283 sw
tri 1891 13185 1989 13283 ne
rect 1989 13185 2343 13283
tri 2343 13185 2441 13283 sw
tri 2441 13185 2539 13283 ne
rect 2539 13185 2893 13283
tri 2893 13185 2991 13283 sw
tri 2991 13185 3089 13283 ne
rect 3089 13185 3443 13283
tri 3443 13185 3541 13283 sw
tri 3541 13185 3639 13283 ne
rect 3639 13185 3993 13283
tri 3993 13185 4091 13283 sw
tri 4091 13185 4189 13283 ne
rect 4189 13185 4543 13283
tri 4543 13185 4641 13283 sw
tri 4641 13185 4739 13283 ne
rect 4739 13185 5093 13283
tri 5093 13185 5191 13283 sw
tri 5191 13185 5289 13283 ne
rect 5289 13185 5643 13283
tri 5643 13185 5741 13283 sw
tri 5741 13185 5839 13283 ne
rect 5839 13185 6193 13283
tri 6193 13185 6291 13283 sw
tri 6291 13185 6389 13283 ne
rect 6389 13185 6743 13283
tri 6743 13185 6841 13283 sw
tri 6841 13185 6939 13283 ne
rect 6939 13185 7293 13283
tri 7293 13185 7391 13283 sw
tri 7391 13185 7489 13283 ne
rect 7489 13185 7843 13283
tri 7843 13185 7941 13283 sw
tri 7941 13185 8039 13283 ne
rect 8039 13185 8393 13283
tri 8393 13185 8491 13283 sw
tri 8491 13185 8589 13283 ne
rect 8589 13185 8943 13283
tri 8943 13185 9041 13283 sw
tri 9041 13185 9139 13283 ne
rect 9139 13185 9493 13283
tri 9493 13185 9591 13283 sw
tri 9591 13185 9689 13283 ne
rect 9689 13185 10043 13283
tri 10043 13185 10141 13283 sw
tri 10141 13185 10239 13283 ne
rect 10239 13185 10593 13283
tri 10593 13185 10691 13283 sw
tri 10691 13185 10789 13283 ne
rect 10789 13185 11143 13283
tri 11143 13185 11241 13283 sw
tri 11241 13185 11339 13283 ne
rect 11339 13185 11693 13283
tri 11693 13185 11791 13283 sw
tri 11791 13185 11889 13283 ne
rect 11889 13185 12243 13283
tri 12243 13185 12341 13283 sw
tri 12341 13185 12439 13283 ne
rect 12439 13185 12793 13283
tri 12793 13185 12891 13283 sw
tri 12891 13185 12989 13283 ne
rect 12989 13185 13343 13283
tri 13343 13185 13441 13283 sw
tri 13441 13185 13539 13283 ne
rect 13539 13185 13893 13283
tri 13893 13185 13991 13283 sw
tri 13991 13185 14089 13283 ne
rect 14089 13185 14443 13283
tri 14443 13185 14541 13283 sw
tri 14541 13185 14639 13283 ne
rect 14639 13185 14993 13283
tri 14993 13185 15091 13283 sw
tri 15091 13185 15189 13283 ne
rect 15189 13185 15543 13283
tri 15543 13185 15641 13283 sw
tri 15641 13185 15739 13283 ne
rect 15739 13185 16093 13283
tri 16093 13185 16191 13283 sw
tri 16191 13185 16289 13283 ne
rect 16289 13185 16643 13283
tri 16643 13185 16741 13283 sw
tri 16741 13185 16839 13283 ne
rect 16839 13185 17193 13283
tri 17193 13185 17291 13283 sw
tri 17291 13185 17389 13283 ne
rect 17389 13185 17743 13283
tri 17743 13185 17841 13283 sw
tri 17841 13185 17939 13283 ne
rect 17939 13185 18293 13283
tri 18293 13185 18391 13283 sw
tri 18391 13185 18489 13283 ne
rect 18489 13185 18843 13283
tri 18843 13185 18941 13283 sw
tri 18941 13185 19039 13283 ne
rect 19039 13185 19393 13283
tri 19393 13185 19491 13283 sw
tri 19491 13185 19589 13283 ne
rect 19589 13185 20300 13283
rect -2000 13087 241 13185
tri 241 13087 339 13185 sw
tri 339 13087 437 13185 ne
rect 437 13087 791 13185
tri 791 13087 889 13185 sw
tri 889 13087 987 13185 ne
rect 987 13087 1341 13185
tri 1341 13087 1439 13185 sw
tri 1439 13087 1537 13185 ne
rect 1537 13087 1891 13185
tri 1891 13087 1989 13185 sw
tri 1989 13087 2087 13185 ne
rect 2087 13087 2441 13185
tri 2441 13087 2539 13185 sw
tri 2539 13087 2637 13185 ne
rect 2637 13087 2991 13185
tri 2991 13087 3089 13185 sw
tri 3089 13087 3187 13185 ne
rect 3187 13087 3541 13185
tri 3541 13087 3639 13185 sw
tri 3639 13087 3737 13185 ne
rect 3737 13087 4091 13185
tri 4091 13087 4189 13185 sw
tri 4189 13087 4287 13185 ne
rect 4287 13087 4641 13185
tri 4641 13087 4739 13185 sw
tri 4739 13087 4837 13185 ne
rect 4837 13087 5191 13185
tri 5191 13087 5289 13185 sw
tri 5289 13087 5387 13185 ne
rect 5387 13087 5741 13185
tri 5741 13087 5839 13185 sw
tri 5839 13087 5937 13185 ne
rect 5937 13087 6291 13185
tri 6291 13087 6389 13185 sw
tri 6389 13087 6487 13185 ne
rect 6487 13087 6841 13185
tri 6841 13087 6939 13185 sw
tri 6939 13087 7037 13185 ne
rect 7037 13087 7391 13185
tri 7391 13087 7489 13185 sw
tri 7489 13087 7587 13185 ne
rect 7587 13087 7941 13185
tri 7941 13087 8039 13185 sw
tri 8039 13087 8137 13185 ne
rect 8137 13087 8491 13185
tri 8491 13087 8589 13185 sw
tri 8589 13087 8687 13185 ne
rect 8687 13087 9041 13185
tri 9041 13087 9139 13185 sw
tri 9139 13087 9237 13185 ne
rect 9237 13087 9591 13185
tri 9591 13087 9689 13185 sw
tri 9689 13087 9787 13185 ne
rect 9787 13087 10141 13185
tri 10141 13087 10239 13185 sw
tri 10239 13087 10337 13185 ne
rect 10337 13087 10691 13185
tri 10691 13087 10789 13185 sw
tri 10789 13087 10887 13185 ne
rect 10887 13087 11241 13185
tri 11241 13087 11339 13185 sw
tri 11339 13087 11437 13185 ne
rect 11437 13087 11791 13185
tri 11791 13087 11889 13185 sw
tri 11889 13087 11987 13185 ne
rect 11987 13087 12341 13185
tri 12341 13087 12439 13185 sw
tri 12439 13087 12537 13185 ne
rect 12537 13087 12891 13185
tri 12891 13087 12989 13185 sw
tri 12989 13087 13087 13185 ne
rect 13087 13087 13441 13185
tri 13441 13087 13539 13185 sw
tri 13539 13087 13637 13185 ne
rect 13637 13087 13991 13185
tri 13991 13087 14089 13185 sw
tri 14089 13087 14187 13185 ne
rect 14187 13087 14541 13185
tri 14541 13087 14639 13185 sw
tri 14639 13087 14737 13185 ne
rect 14737 13087 15091 13185
tri 15091 13087 15189 13185 sw
tri 15189 13087 15287 13185 ne
rect 15287 13087 15641 13185
tri 15641 13087 15739 13185 sw
tri 15739 13087 15837 13185 ne
rect 15837 13087 16191 13185
tri 16191 13087 16289 13185 sw
tri 16289 13087 16387 13185 ne
rect 16387 13087 16741 13185
tri 16741 13087 16839 13185 sw
tri 16839 13087 16937 13185 ne
rect 16937 13087 17291 13185
tri 17291 13087 17389 13185 sw
tri 17389 13087 17487 13185 ne
rect 17487 13087 17841 13185
tri 17841 13087 17939 13185 sw
tri 17939 13087 18037 13185 ne
rect 18037 13087 18391 13185
tri 18391 13087 18489 13185 sw
tri 18489 13087 18587 13185 ne
rect 18587 13087 18941 13185
tri 18941 13087 19039 13185 sw
tri 19039 13087 19137 13185 ne
rect 19137 13087 19491 13185
tri 19491 13087 19589 13185 sw
tri 19589 13087 19687 13185 ne
rect 19687 13087 20300 13185
rect -2000 12989 339 13087
tri 339 12989 437 13087 sw
tri 437 12989 535 13087 ne
rect 535 12989 889 13087
tri 889 12989 987 13087 sw
tri 987 12989 1085 13087 ne
rect 1085 12989 1439 13087
tri 1439 12989 1537 13087 sw
tri 1537 12989 1635 13087 ne
rect 1635 12989 1989 13087
tri 1989 12989 2087 13087 sw
tri 2087 12989 2185 13087 ne
rect 2185 12989 2539 13087
tri 2539 12989 2637 13087 sw
tri 2637 12989 2735 13087 ne
rect 2735 12989 3089 13087
tri 3089 12989 3187 13087 sw
tri 3187 12989 3285 13087 ne
rect 3285 12989 3639 13087
tri 3639 12989 3737 13087 sw
tri 3737 12989 3835 13087 ne
rect 3835 12989 4189 13087
tri 4189 12989 4287 13087 sw
tri 4287 12989 4385 13087 ne
rect 4385 12989 4739 13087
tri 4739 12989 4837 13087 sw
tri 4837 12989 4935 13087 ne
rect 4935 12989 5289 13087
tri 5289 12989 5387 13087 sw
tri 5387 12989 5485 13087 ne
rect 5485 12989 5839 13087
tri 5839 12989 5937 13087 sw
tri 5937 12989 6035 13087 ne
rect 6035 12989 6389 13087
tri 6389 12989 6487 13087 sw
tri 6487 12989 6585 13087 ne
rect 6585 12989 6939 13087
tri 6939 12989 7037 13087 sw
tri 7037 12989 7135 13087 ne
rect 7135 12989 7489 13087
tri 7489 12989 7587 13087 sw
tri 7587 12989 7685 13087 ne
rect 7685 12989 8039 13087
tri 8039 12989 8137 13087 sw
tri 8137 12989 8235 13087 ne
rect 8235 12989 8589 13087
tri 8589 12989 8687 13087 sw
tri 8687 12989 8785 13087 ne
rect 8785 12989 9139 13087
tri 9139 12989 9237 13087 sw
tri 9237 12989 9335 13087 ne
rect 9335 12989 9689 13087
tri 9689 12989 9787 13087 sw
tri 9787 12989 9885 13087 ne
rect 9885 12989 10239 13087
tri 10239 12989 10337 13087 sw
tri 10337 12989 10435 13087 ne
rect 10435 12989 10789 13087
tri 10789 12989 10887 13087 sw
tri 10887 12989 10985 13087 ne
rect 10985 12989 11339 13087
tri 11339 12989 11437 13087 sw
tri 11437 12989 11535 13087 ne
rect 11535 12989 11889 13087
tri 11889 12989 11987 13087 sw
tri 11987 12989 12085 13087 ne
rect 12085 12989 12439 13087
tri 12439 12989 12537 13087 sw
tri 12537 12989 12635 13087 ne
rect 12635 12989 12989 13087
tri 12989 12989 13087 13087 sw
tri 13087 12989 13185 13087 ne
rect 13185 12989 13539 13087
tri 13539 12989 13637 13087 sw
tri 13637 12989 13735 13087 ne
rect 13735 12989 14089 13087
tri 14089 12989 14187 13087 sw
tri 14187 12989 14285 13087 ne
rect 14285 12989 14639 13087
tri 14639 12989 14737 13087 sw
tri 14737 12989 14835 13087 ne
rect 14835 12989 15189 13087
tri 15189 12989 15287 13087 sw
tri 15287 12989 15385 13087 ne
rect 15385 12989 15739 13087
tri 15739 12989 15837 13087 sw
tri 15837 12989 15935 13087 ne
rect 15935 12989 16289 13087
tri 16289 12989 16387 13087 sw
tri 16387 12989 16485 13087 ne
rect 16485 12989 16839 13087
tri 16839 12989 16937 13087 sw
tri 16937 12989 17035 13087 ne
rect 17035 12989 17389 13087
tri 17389 12989 17487 13087 sw
tri 17487 12989 17585 13087 ne
rect 17585 12989 17939 13087
tri 17939 12989 18037 13087 sw
tri 18037 12989 18135 13087 ne
rect 18135 12989 18489 13087
tri 18489 12989 18587 13087 sw
tri 18587 12989 18685 13087 ne
rect 18685 12989 19039 13087
tri 19039 12989 19137 13087 sw
tri 19137 12989 19235 13087 ne
rect 19235 12989 19589 13087
tri 19589 12989 19687 13087 sw
rect 20800 12989 21800 13637
rect -2000 12985 437 12989
rect -2000 12865 215 12985
rect 335 12891 437 12985
tri 437 12891 535 12989 sw
tri 535 12891 633 12989 ne
rect 633 12985 987 12989
rect 633 12891 765 12985
rect 335 12865 535 12891
rect -2000 12861 535 12865
rect -2000 12213 -1000 12861
tri 113 12763 211 12861 ne
rect 211 12813 535 12861
tri 535 12813 613 12891 sw
tri 633 12813 711 12891 ne
rect 711 12865 765 12891
rect 885 12891 987 12985
tri 987 12891 1085 12989 sw
tri 1085 12891 1183 12989 ne
rect 1183 12985 1537 12989
rect 1183 12891 1315 12985
rect 885 12865 1085 12891
rect 711 12813 1085 12865
tri 1085 12813 1163 12891 sw
tri 1183 12813 1261 12891 ne
rect 1261 12865 1315 12891
rect 1435 12891 1537 12985
tri 1537 12891 1635 12989 sw
tri 1635 12891 1733 12989 ne
rect 1733 12985 2087 12989
rect 1733 12891 1865 12985
rect 1435 12865 1635 12891
rect 1261 12813 1635 12865
tri 1635 12813 1713 12891 sw
tri 1733 12813 1811 12891 ne
rect 1811 12865 1865 12891
rect 1985 12891 2087 12985
tri 2087 12891 2185 12989 sw
tri 2185 12891 2283 12989 ne
rect 2283 12985 2637 12989
rect 2283 12891 2415 12985
rect 1985 12865 2185 12891
rect 1811 12813 2185 12865
tri 2185 12813 2263 12891 sw
tri 2283 12813 2361 12891 ne
rect 2361 12865 2415 12891
rect 2535 12891 2637 12985
tri 2637 12891 2735 12989 sw
tri 2735 12891 2833 12989 ne
rect 2833 12985 3187 12989
rect 2833 12891 2965 12985
rect 2535 12865 2735 12891
rect 2361 12813 2735 12865
tri 2735 12813 2813 12891 sw
tri 2833 12813 2911 12891 ne
rect 2911 12865 2965 12891
rect 3085 12891 3187 12985
tri 3187 12891 3285 12989 sw
tri 3285 12891 3383 12989 ne
rect 3383 12985 3737 12989
rect 3383 12891 3515 12985
rect 3085 12865 3285 12891
rect 2911 12813 3285 12865
tri 3285 12813 3363 12891 sw
tri 3383 12813 3461 12891 ne
rect 3461 12865 3515 12891
rect 3635 12891 3737 12985
tri 3737 12891 3835 12989 sw
tri 3835 12891 3933 12989 ne
rect 3933 12985 4287 12989
rect 3933 12891 4065 12985
rect 3635 12865 3835 12891
rect 3461 12813 3835 12865
tri 3835 12813 3913 12891 sw
tri 3933 12813 4011 12891 ne
rect 4011 12865 4065 12891
rect 4185 12891 4287 12985
tri 4287 12891 4385 12989 sw
tri 4385 12891 4483 12989 ne
rect 4483 12985 4837 12989
rect 4483 12891 4615 12985
rect 4185 12865 4385 12891
rect 4011 12813 4385 12865
tri 4385 12813 4463 12891 sw
tri 4483 12813 4561 12891 ne
rect 4561 12865 4615 12891
rect 4735 12891 4837 12985
tri 4837 12891 4935 12989 sw
tri 4935 12891 5033 12989 ne
rect 5033 12985 5387 12989
rect 5033 12891 5165 12985
rect 4735 12865 4935 12891
rect 4561 12813 4935 12865
tri 4935 12813 5013 12891 sw
tri 5033 12813 5111 12891 ne
rect 5111 12865 5165 12891
rect 5285 12891 5387 12985
tri 5387 12891 5485 12989 sw
tri 5485 12891 5583 12989 ne
rect 5583 12985 5937 12989
rect 5583 12891 5715 12985
rect 5285 12865 5485 12891
rect 5111 12813 5485 12865
tri 5485 12813 5563 12891 sw
tri 5583 12813 5661 12891 ne
rect 5661 12865 5715 12891
rect 5835 12891 5937 12985
tri 5937 12891 6035 12989 sw
tri 6035 12891 6133 12989 ne
rect 6133 12985 6487 12989
rect 6133 12891 6265 12985
rect 5835 12865 6035 12891
rect 5661 12813 6035 12865
tri 6035 12813 6113 12891 sw
tri 6133 12813 6211 12891 ne
rect 6211 12865 6265 12891
rect 6385 12891 6487 12985
tri 6487 12891 6585 12989 sw
tri 6585 12891 6683 12989 ne
rect 6683 12985 7037 12989
rect 6683 12891 6815 12985
rect 6385 12865 6585 12891
rect 6211 12813 6585 12865
tri 6585 12813 6663 12891 sw
tri 6683 12813 6761 12891 ne
rect 6761 12865 6815 12891
rect 6935 12891 7037 12985
tri 7037 12891 7135 12989 sw
tri 7135 12891 7233 12989 ne
rect 7233 12985 7587 12989
rect 7233 12891 7365 12985
rect 6935 12865 7135 12891
rect 6761 12813 7135 12865
tri 7135 12813 7213 12891 sw
tri 7233 12813 7311 12891 ne
rect 7311 12865 7365 12891
rect 7485 12891 7587 12985
tri 7587 12891 7685 12989 sw
tri 7685 12891 7783 12989 ne
rect 7783 12985 8137 12989
rect 7783 12891 7915 12985
rect 7485 12865 7685 12891
rect 7311 12813 7685 12865
tri 7685 12813 7763 12891 sw
tri 7783 12813 7861 12891 ne
rect 7861 12865 7915 12891
rect 8035 12891 8137 12985
tri 8137 12891 8235 12989 sw
tri 8235 12891 8333 12989 ne
rect 8333 12985 8687 12989
rect 8333 12891 8465 12985
rect 8035 12865 8235 12891
rect 7861 12813 8235 12865
tri 8235 12813 8313 12891 sw
tri 8333 12813 8411 12891 ne
rect 8411 12865 8465 12891
rect 8585 12891 8687 12985
tri 8687 12891 8785 12989 sw
tri 8785 12891 8883 12989 ne
rect 8883 12985 9237 12989
rect 8883 12891 9015 12985
rect 8585 12865 8785 12891
rect 8411 12813 8785 12865
tri 8785 12813 8863 12891 sw
tri 8883 12813 8961 12891 ne
rect 8961 12865 9015 12891
rect 9135 12891 9237 12985
tri 9237 12891 9335 12989 sw
tri 9335 12891 9433 12989 ne
rect 9433 12985 9787 12989
rect 9433 12891 9565 12985
rect 9135 12865 9335 12891
rect 8961 12813 9335 12865
tri 9335 12813 9413 12891 sw
tri 9433 12813 9511 12891 ne
rect 9511 12865 9565 12891
rect 9685 12891 9787 12985
tri 9787 12891 9885 12989 sw
tri 9885 12891 9983 12989 ne
rect 9983 12985 10337 12989
rect 9983 12891 10115 12985
rect 9685 12865 9885 12891
rect 9511 12813 9885 12865
tri 9885 12813 9963 12891 sw
tri 9983 12813 10061 12891 ne
rect 10061 12865 10115 12891
rect 10235 12891 10337 12985
tri 10337 12891 10435 12989 sw
tri 10435 12891 10533 12989 ne
rect 10533 12985 10887 12989
rect 10533 12891 10665 12985
rect 10235 12865 10435 12891
rect 10061 12813 10435 12865
tri 10435 12813 10513 12891 sw
tri 10533 12813 10611 12891 ne
rect 10611 12865 10665 12891
rect 10785 12891 10887 12985
tri 10887 12891 10985 12989 sw
tri 10985 12891 11083 12989 ne
rect 11083 12985 11437 12989
rect 11083 12891 11215 12985
rect 10785 12865 10985 12891
rect 10611 12813 10985 12865
tri 10985 12813 11063 12891 sw
tri 11083 12813 11161 12891 ne
rect 11161 12865 11215 12891
rect 11335 12891 11437 12985
tri 11437 12891 11535 12989 sw
tri 11535 12891 11633 12989 ne
rect 11633 12985 11987 12989
rect 11633 12891 11765 12985
rect 11335 12865 11535 12891
rect 11161 12813 11535 12865
tri 11535 12813 11613 12891 sw
tri 11633 12813 11711 12891 ne
rect 11711 12865 11765 12891
rect 11885 12891 11987 12985
tri 11987 12891 12085 12989 sw
tri 12085 12891 12183 12989 ne
rect 12183 12985 12537 12989
rect 12183 12891 12315 12985
rect 11885 12865 12085 12891
rect 11711 12813 12085 12865
tri 12085 12813 12163 12891 sw
tri 12183 12813 12261 12891 ne
rect 12261 12865 12315 12891
rect 12435 12891 12537 12985
tri 12537 12891 12635 12989 sw
tri 12635 12891 12733 12989 ne
rect 12733 12985 13087 12989
rect 12733 12891 12865 12985
rect 12435 12865 12635 12891
rect 12261 12813 12635 12865
tri 12635 12813 12713 12891 sw
tri 12733 12813 12811 12891 ne
rect 12811 12865 12865 12891
rect 12985 12891 13087 12985
tri 13087 12891 13185 12989 sw
tri 13185 12891 13283 12989 ne
rect 13283 12985 13637 12989
rect 13283 12891 13415 12985
rect 12985 12865 13185 12891
rect 12811 12813 13185 12865
tri 13185 12813 13263 12891 sw
tri 13283 12813 13361 12891 ne
rect 13361 12865 13415 12891
rect 13535 12891 13637 12985
tri 13637 12891 13735 12989 sw
tri 13735 12891 13833 12989 ne
rect 13833 12985 14187 12989
rect 13833 12891 13965 12985
rect 13535 12865 13735 12891
rect 13361 12813 13735 12865
tri 13735 12813 13813 12891 sw
tri 13833 12813 13911 12891 ne
rect 13911 12865 13965 12891
rect 14085 12891 14187 12985
tri 14187 12891 14285 12989 sw
tri 14285 12891 14383 12989 ne
rect 14383 12985 14737 12989
rect 14383 12891 14515 12985
rect 14085 12865 14285 12891
rect 13911 12813 14285 12865
tri 14285 12813 14363 12891 sw
tri 14383 12813 14461 12891 ne
rect 14461 12865 14515 12891
rect 14635 12891 14737 12985
tri 14737 12891 14835 12989 sw
tri 14835 12891 14933 12989 ne
rect 14933 12985 15287 12989
rect 14933 12891 15065 12985
rect 14635 12865 14835 12891
rect 14461 12813 14835 12865
tri 14835 12813 14913 12891 sw
tri 14933 12813 15011 12891 ne
rect 15011 12865 15065 12891
rect 15185 12891 15287 12985
tri 15287 12891 15385 12989 sw
tri 15385 12891 15483 12989 ne
rect 15483 12985 15837 12989
rect 15483 12891 15615 12985
rect 15185 12865 15385 12891
rect 15011 12813 15385 12865
tri 15385 12813 15463 12891 sw
tri 15483 12813 15561 12891 ne
rect 15561 12865 15615 12891
rect 15735 12891 15837 12985
tri 15837 12891 15935 12989 sw
tri 15935 12891 16033 12989 ne
rect 16033 12985 16387 12989
rect 16033 12891 16165 12985
rect 15735 12865 15935 12891
rect 15561 12813 15935 12865
tri 15935 12813 16013 12891 sw
tri 16033 12813 16111 12891 ne
rect 16111 12865 16165 12891
rect 16285 12891 16387 12985
tri 16387 12891 16485 12989 sw
tri 16485 12891 16583 12989 ne
rect 16583 12985 16937 12989
rect 16583 12891 16715 12985
rect 16285 12865 16485 12891
rect 16111 12813 16485 12865
tri 16485 12813 16563 12891 sw
tri 16583 12813 16661 12891 ne
rect 16661 12865 16715 12891
rect 16835 12891 16937 12985
tri 16937 12891 17035 12989 sw
tri 17035 12891 17133 12989 ne
rect 17133 12985 17487 12989
rect 17133 12891 17265 12985
rect 16835 12865 17035 12891
rect 16661 12813 17035 12865
tri 17035 12813 17113 12891 sw
tri 17133 12813 17211 12891 ne
rect 17211 12865 17265 12891
rect 17385 12891 17487 12985
tri 17487 12891 17585 12989 sw
tri 17585 12891 17683 12989 ne
rect 17683 12985 18037 12989
rect 17683 12891 17815 12985
rect 17385 12865 17585 12891
rect 17211 12813 17585 12865
tri 17585 12813 17663 12891 sw
tri 17683 12813 17761 12891 ne
rect 17761 12865 17815 12891
rect 17935 12891 18037 12985
tri 18037 12891 18135 12989 sw
tri 18135 12891 18233 12989 ne
rect 18233 12985 18587 12989
rect 18233 12891 18365 12985
rect 17935 12865 18135 12891
rect 17761 12813 18135 12865
tri 18135 12813 18213 12891 sw
tri 18233 12813 18311 12891 ne
rect 18311 12865 18365 12891
rect 18485 12891 18587 12985
tri 18587 12891 18685 12989 sw
tri 18685 12891 18783 12989 ne
rect 18783 12985 19137 12989
rect 18783 12891 18915 12985
rect 18485 12865 18685 12891
rect 18311 12813 18685 12865
tri 18685 12813 18763 12891 sw
tri 18783 12813 18861 12891 ne
rect 18861 12865 18915 12891
rect 19035 12891 19137 12985
tri 19137 12891 19235 12989 sw
tri 19235 12891 19333 12989 ne
rect 19333 12985 21800 12989
rect 19333 12891 19465 12985
rect 19035 12865 19235 12891
rect 18861 12813 19235 12865
tri 19235 12813 19313 12891 sw
tri 19333 12813 19411 12891 ne
rect 19411 12865 19465 12891
rect 19585 12865 21800 12985
rect 19411 12813 21800 12865
rect 211 12763 613 12813
rect -500 12713 113 12763
tri 113 12713 163 12763 sw
tri 211 12713 261 12763 ne
rect 261 12733 613 12763
tri 613 12733 693 12813 sw
tri 711 12733 791 12813 ne
rect 791 12733 1163 12813
tri 1163 12733 1243 12813 sw
tri 1261 12733 1341 12813 ne
rect 1341 12733 1713 12813
tri 1713 12733 1793 12813 sw
tri 1811 12733 1891 12813 ne
rect 1891 12733 2263 12813
tri 2263 12733 2343 12813 sw
tri 2361 12733 2441 12813 ne
rect 2441 12733 2813 12813
tri 2813 12733 2893 12813 sw
tri 2911 12733 2991 12813 ne
rect 2991 12733 3363 12813
tri 3363 12733 3443 12813 sw
tri 3461 12733 3541 12813 ne
rect 3541 12733 3913 12813
tri 3913 12733 3993 12813 sw
tri 4011 12733 4091 12813 ne
rect 4091 12733 4463 12813
tri 4463 12733 4543 12813 sw
tri 4561 12733 4641 12813 ne
rect 4641 12733 5013 12813
tri 5013 12733 5093 12813 sw
tri 5111 12733 5191 12813 ne
rect 5191 12733 5563 12813
tri 5563 12733 5643 12813 sw
tri 5661 12733 5741 12813 ne
rect 5741 12733 6113 12813
tri 6113 12733 6193 12813 sw
tri 6211 12733 6291 12813 ne
rect 6291 12733 6663 12813
tri 6663 12733 6743 12813 sw
tri 6761 12733 6841 12813 ne
rect 6841 12733 7213 12813
tri 7213 12733 7293 12813 sw
tri 7311 12733 7391 12813 ne
rect 7391 12733 7763 12813
tri 7763 12733 7843 12813 sw
tri 7861 12733 7941 12813 ne
rect 7941 12733 8313 12813
tri 8313 12733 8393 12813 sw
tri 8411 12733 8491 12813 ne
rect 8491 12733 8863 12813
tri 8863 12733 8943 12813 sw
tri 8961 12733 9041 12813 ne
rect 9041 12733 9413 12813
tri 9413 12733 9493 12813 sw
tri 9511 12733 9591 12813 ne
rect 9591 12733 9963 12813
tri 9963 12733 10043 12813 sw
tri 10061 12733 10141 12813 ne
rect 10141 12733 10513 12813
tri 10513 12733 10593 12813 sw
tri 10611 12733 10691 12813 ne
rect 10691 12733 11063 12813
tri 11063 12733 11143 12813 sw
tri 11161 12733 11241 12813 ne
rect 11241 12733 11613 12813
tri 11613 12733 11693 12813 sw
tri 11711 12733 11791 12813 ne
rect 11791 12733 12163 12813
tri 12163 12733 12243 12813 sw
tri 12261 12733 12341 12813 ne
rect 12341 12733 12713 12813
tri 12713 12733 12793 12813 sw
tri 12811 12733 12891 12813 ne
rect 12891 12733 13263 12813
tri 13263 12733 13343 12813 sw
tri 13361 12733 13441 12813 ne
rect 13441 12733 13813 12813
tri 13813 12733 13893 12813 sw
tri 13911 12733 13991 12813 ne
rect 13991 12733 14363 12813
tri 14363 12733 14443 12813 sw
tri 14461 12733 14541 12813 ne
rect 14541 12733 14913 12813
tri 14913 12733 14993 12813 sw
tri 15011 12733 15091 12813 ne
rect 15091 12733 15463 12813
tri 15463 12733 15543 12813 sw
tri 15561 12733 15641 12813 ne
rect 15641 12733 16013 12813
tri 16013 12733 16093 12813 sw
tri 16111 12733 16191 12813 ne
rect 16191 12733 16563 12813
tri 16563 12733 16643 12813 sw
tri 16661 12733 16741 12813 ne
rect 16741 12733 17113 12813
tri 17113 12733 17193 12813 sw
tri 17211 12733 17291 12813 ne
rect 17291 12733 17663 12813
tri 17663 12733 17743 12813 sw
tri 17761 12733 17841 12813 ne
rect 17841 12733 18213 12813
tri 18213 12733 18293 12813 sw
tri 18311 12733 18391 12813 ne
rect 18391 12733 18763 12813
tri 18763 12733 18843 12813 sw
tri 18861 12733 18941 12813 ne
rect 18941 12733 19313 12813
tri 19313 12733 19393 12813 sw
tri 19411 12733 19491 12813 ne
rect 19491 12733 20100 12813
rect 261 12713 693 12733
rect -500 12635 163 12713
tri 163 12635 241 12713 sw
tri 261 12635 339 12713 ne
rect 339 12635 693 12713
tri 693 12635 791 12733 sw
tri 791 12635 889 12733 ne
rect 889 12635 1243 12733
tri 1243 12635 1341 12733 sw
tri 1341 12635 1439 12733 ne
rect 1439 12635 1793 12733
tri 1793 12635 1891 12733 sw
tri 1891 12635 1989 12733 ne
rect 1989 12635 2343 12733
tri 2343 12635 2441 12733 sw
tri 2441 12635 2539 12733 ne
rect 2539 12635 2893 12733
tri 2893 12635 2991 12733 sw
tri 2991 12635 3089 12733 ne
rect 3089 12635 3443 12733
tri 3443 12635 3541 12733 sw
tri 3541 12635 3639 12733 ne
rect 3639 12635 3993 12733
tri 3993 12635 4091 12733 sw
tri 4091 12635 4189 12733 ne
rect 4189 12635 4543 12733
tri 4543 12635 4641 12733 sw
tri 4641 12635 4739 12733 ne
rect 4739 12635 5093 12733
tri 5093 12635 5191 12733 sw
tri 5191 12635 5289 12733 ne
rect 5289 12635 5643 12733
tri 5643 12635 5741 12733 sw
tri 5741 12635 5839 12733 ne
rect 5839 12635 6193 12733
tri 6193 12635 6291 12733 sw
tri 6291 12635 6389 12733 ne
rect 6389 12635 6743 12733
tri 6743 12635 6841 12733 sw
tri 6841 12635 6939 12733 ne
rect 6939 12635 7293 12733
tri 7293 12635 7391 12733 sw
tri 7391 12635 7489 12733 ne
rect 7489 12635 7843 12733
tri 7843 12635 7941 12733 sw
tri 7941 12635 8039 12733 ne
rect 8039 12635 8393 12733
tri 8393 12635 8491 12733 sw
tri 8491 12635 8589 12733 ne
rect 8589 12635 8943 12733
tri 8943 12635 9041 12733 sw
tri 9041 12635 9139 12733 ne
rect 9139 12635 9493 12733
tri 9493 12635 9591 12733 sw
tri 9591 12635 9689 12733 ne
rect 9689 12635 10043 12733
tri 10043 12635 10141 12733 sw
tri 10141 12635 10239 12733 ne
rect 10239 12635 10593 12733
tri 10593 12635 10691 12733 sw
tri 10691 12635 10789 12733 ne
rect 10789 12635 11143 12733
tri 11143 12635 11241 12733 sw
tri 11241 12635 11339 12733 ne
rect 11339 12635 11693 12733
tri 11693 12635 11791 12733 sw
tri 11791 12635 11889 12733 ne
rect 11889 12635 12243 12733
tri 12243 12635 12341 12733 sw
tri 12341 12635 12439 12733 ne
rect 12439 12635 12793 12733
tri 12793 12635 12891 12733 sw
tri 12891 12635 12989 12733 ne
rect 12989 12635 13343 12733
tri 13343 12635 13441 12733 sw
tri 13441 12635 13539 12733 ne
rect 13539 12635 13893 12733
tri 13893 12635 13991 12733 sw
tri 13991 12635 14089 12733 ne
rect 14089 12635 14443 12733
tri 14443 12635 14541 12733 sw
tri 14541 12635 14639 12733 ne
rect 14639 12635 14993 12733
tri 14993 12635 15091 12733 sw
tri 15091 12635 15189 12733 ne
rect 15189 12635 15543 12733
tri 15543 12635 15641 12733 sw
tri 15641 12635 15739 12733 ne
rect 15739 12635 16093 12733
tri 16093 12635 16191 12733 sw
tri 16191 12635 16289 12733 ne
rect 16289 12635 16643 12733
tri 16643 12635 16741 12733 sw
tri 16741 12635 16839 12733 ne
rect 16839 12635 17193 12733
tri 17193 12635 17291 12733 sw
tri 17291 12635 17389 12733 ne
rect 17389 12635 17743 12733
tri 17743 12635 17841 12733 sw
tri 17841 12635 17939 12733 ne
rect 17939 12635 18293 12733
tri 18293 12635 18391 12733 sw
tri 18391 12635 18489 12733 ne
rect 18489 12635 18843 12733
tri 18843 12635 18941 12733 sw
tri 18941 12635 19039 12733 ne
rect 19039 12635 19393 12733
tri 19393 12635 19491 12733 sw
tri 19491 12635 19589 12733 ne
rect 19589 12713 20100 12733
rect 20200 12713 21800 12813
rect 19589 12635 21800 12713
rect -500 12587 241 12635
rect -500 12487 -400 12587
rect -300 12537 241 12587
tri 241 12537 339 12635 sw
tri 339 12537 437 12635 ne
rect 437 12537 791 12635
tri 791 12537 889 12635 sw
tri 889 12537 987 12635 ne
rect 987 12537 1341 12635
tri 1341 12537 1439 12635 sw
tri 1439 12537 1537 12635 ne
rect 1537 12537 1891 12635
tri 1891 12537 1989 12635 sw
tri 1989 12537 2087 12635 ne
rect 2087 12537 2441 12635
tri 2441 12537 2539 12635 sw
tri 2539 12537 2637 12635 ne
rect 2637 12537 2991 12635
tri 2991 12537 3089 12635 sw
tri 3089 12537 3187 12635 ne
rect 3187 12537 3541 12635
tri 3541 12537 3639 12635 sw
tri 3639 12537 3737 12635 ne
rect 3737 12537 4091 12635
tri 4091 12537 4189 12635 sw
tri 4189 12537 4287 12635 ne
rect 4287 12537 4641 12635
tri 4641 12537 4739 12635 sw
tri 4739 12537 4837 12635 ne
rect 4837 12537 5191 12635
tri 5191 12537 5289 12635 sw
tri 5289 12537 5387 12635 ne
rect 5387 12537 5741 12635
tri 5741 12537 5839 12635 sw
tri 5839 12537 5937 12635 ne
rect 5937 12537 6291 12635
tri 6291 12537 6389 12635 sw
tri 6389 12537 6487 12635 ne
rect 6487 12537 6841 12635
tri 6841 12537 6939 12635 sw
tri 6939 12537 7037 12635 ne
rect 7037 12537 7391 12635
tri 7391 12537 7489 12635 sw
tri 7489 12537 7587 12635 ne
rect 7587 12537 7941 12635
tri 7941 12537 8039 12635 sw
tri 8039 12537 8137 12635 ne
rect 8137 12537 8491 12635
tri 8491 12537 8589 12635 sw
tri 8589 12537 8687 12635 ne
rect 8687 12537 9041 12635
tri 9041 12537 9139 12635 sw
tri 9139 12537 9237 12635 ne
rect 9237 12537 9591 12635
tri 9591 12537 9689 12635 sw
tri 9689 12537 9787 12635 ne
rect 9787 12537 10141 12635
tri 10141 12537 10239 12635 sw
tri 10239 12537 10337 12635 ne
rect 10337 12537 10691 12635
tri 10691 12537 10789 12635 sw
tri 10789 12537 10887 12635 ne
rect 10887 12537 11241 12635
tri 11241 12537 11339 12635 sw
tri 11339 12537 11437 12635 ne
rect 11437 12537 11791 12635
tri 11791 12537 11889 12635 sw
tri 11889 12537 11987 12635 ne
rect 11987 12537 12341 12635
tri 12341 12537 12439 12635 sw
tri 12439 12537 12537 12635 ne
rect 12537 12537 12891 12635
tri 12891 12537 12989 12635 sw
tri 12989 12537 13087 12635 ne
rect 13087 12537 13441 12635
tri 13441 12537 13539 12635 sw
tri 13539 12537 13637 12635 ne
rect 13637 12537 13991 12635
tri 13991 12537 14089 12635 sw
tri 14089 12537 14187 12635 ne
rect 14187 12537 14541 12635
tri 14541 12537 14639 12635 sw
tri 14639 12537 14737 12635 ne
rect 14737 12537 15091 12635
tri 15091 12537 15189 12635 sw
tri 15189 12537 15287 12635 ne
rect 15287 12537 15641 12635
tri 15641 12537 15739 12635 sw
tri 15739 12537 15837 12635 ne
rect 15837 12537 16191 12635
tri 16191 12537 16289 12635 sw
tri 16289 12537 16387 12635 ne
rect 16387 12537 16741 12635
tri 16741 12537 16839 12635 sw
tri 16839 12537 16937 12635 ne
rect 16937 12537 17291 12635
tri 17291 12537 17389 12635 sw
tri 17389 12537 17487 12635 ne
rect 17487 12537 17841 12635
tri 17841 12537 17939 12635 sw
tri 17939 12537 18037 12635 ne
rect 18037 12537 18391 12635
tri 18391 12537 18489 12635 sw
tri 18489 12537 18587 12635 ne
rect 18587 12537 18941 12635
tri 18941 12537 19039 12635 sw
tri 19039 12537 19137 12635 ne
rect 19137 12537 19491 12635
tri 19491 12537 19589 12635 sw
tri 19589 12537 19687 12635 ne
rect 19687 12537 21800 12635
rect -300 12487 339 12537
rect -500 12439 339 12487
tri 339 12439 437 12537 sw
tri 437 12439 535 12537 ne
rect 535 12439 889 12537
tri 889 12439 987 12537 sw
tri 987 12439 1085 12537 ne
rect 1085 12439 1439 12537
tri 1439 12439 1537 12537 sw
tri 1537 12439 1635 12537 ne
rect 1635 12439 1989 12537
tri 1989 12439 2087 12537 sw
tri 2087 12439 2185 12537 ne
rect 2185 12439 2539 12537
tri 2539 12439 2637 12537 sw
tri 2637 12439 2735 12537 ne
rect 2735 12439 3089 12537
tri 3089 12439 3187 12537 sw
tri 3187 12439 3285 12537 ne
rect 3285 12439 3639 12537
tri 3639 12439 3737 12537 sw
tri 3737 12439 3835 12537 ne
rect 3835 12439 4189 12537
tri 4189 12439 4287 12537 sw
tri 4287 12439 4385 12537 ne
rect 4385 12439 4739 12537
tri 4739 12439 4837 12537 sw
tri 4837 12439 4935 12537 ne
rect 4935 12439 5289 12537
tri 5289 12439 5387 12537 sw
tri 5387 12439 5485 12537 ne
rect 5485 12439 5839 12537
tri 5839 12439 5937 12537 sw
tri 5937 12439 6035 12537 ne
rect 6035 12439 6389 12537
tri 6389 12439 6487 12537 sw
tri 6487 12439 6585 12537 ne
rect 6585 12439 6939 12537
tri 6939 12439 7037 12537 sw
tri 7037 12439 7135 12537 ne
rect 7135 12439 7489 12537
tri 7489 12439 7587 12537 sw
tri 7587 12439 7685 12537 ne
rect 7685 12439 8039 12537
tri 8039 12439 8137 12537 sw
tri 8137 12439 8235 12537 ne
rect 8235 12439 8589 12537
tri 8589 12439 8687 12537 sw
tri 8687 12439 8785 12537 ne
rect 8785 12439 9139 12537
tri 9139 12439 9237 12537 sw
tri 9237 12439 9335 12537 ne
rect 9335 12439 9689 12537
tri 9689 12439 9787 12537 sw
tri 9787 12439 9885 12537 ne
rect 9885 12439 10239 12537
tri 10239 12439 10337 12537 sw
tri 10337 12439 10435 12537 ne
rect 10435 12439 10789 12537
tri 10789 12439 10887 12537 sw
tri 10887 12439 10985 12537 ne
rect 10985 12439 11339 12537
tri 11339 12439 11437 12537 sw
tri 11437 12439 11535 12537 ne
rect 11535 12439 11889 12537
tri 11889 12439 11987 12537 sw
tri 11987 12439 12085 12537 ne
rect 12085 12439 12439 12537
tri 12439 12439 12537 12537 sw
tri 12537 12439 12635 12537 ne
rect 12635 12439 12989 12537
tri 12989 12439 13087 12537 sw
tri 13087 12439 13185 12537 ne
rect 13185 12439 13539 12537
tri 13539 12439 13637 12537 sw
tri 13637 12439 13735 12537 ne
rect 13735 12439 14089 12537
tri 14089 12439 14187 12537 sw
tri 14187 12439 14285 12537 ne
rect 14285 12439 14639 12537
tri 14639 12439 14737 12537 sw
tri 14737 12439 14835 12537 ne
rect 14835 12439 15189 12537
tri 15189 12439 15287 12537 sw
tri 15287 12439 15385 12537 ne
rect 15385 12439 15739 12537
tri 15739 12439 15837 12537 sw
tri 15837 12439 15935 12537 ne
rect 15935 12439 16289 12537
tri 16289 12439 16387 12537 sw
tri 16387 12439 16485 12537 ne
rect 16485 12439 16839 12537
tri 16839 12439 16937 12537 sw
tri 16937 12439 17035 12537 ne
rect 17035 12439 17389 12537
tri 17389 12439 17487 12537 sw
tri 17487 12439 17585 12537 ne
rect 17585 12439 17939 12537
tri 17939 12439 18037 12537 sw
tri 18037 12439 18135 12537 ne
rect 18135 12439 18489 12537
tri 18489 12439 18587 12537 sw
tri 18587 12439 18685 12537 ne
rect 18685 12439 19039 12537
tri 19039 12439 19137 12537 sw
tri 19137 12439 19235 12537 ne
rect 19235 12439 19589 12537
tri 19589 12439 19687 12537 sw
rect -500 12435 437 12439
rect -500 12315 215 12435
rect 335 12341 437 12435
tri 437 12341 535 12439 sw
tri 535 12341 633 12439 ne
rect 633 12435 987 12439
rect 633 12341 765 12435
rect 335 12315 535 12341
rect -500 12311 535 12315
tri 535 12311 565 12341 sw
tri 633 12311 663 12341 ne
rect 663 12315 765 12341
rect 885 12341 987 12435
tri 987 12341 1085 12439 sw
tri 1085 12341 1183 12439 ne
rect 1183 12435 1537 12439
rect 1183 12341 1315 12435
rect 885 12315 1085 12341
rect 663 12311 1085 12315
tri 1085 12311 1115 12341 sw
tri 1183 12311 1213 12341 ne
rect 1213 12315 1315 12341
rect 1435 12341 1537 12435
tri 1537 12341 1635 12439 sw
tri 1635 12341 1733 12439 ne
rect 1733 12435 2087 12439
rect 1733 12341 1865 12435
rect 1435 12315 1635 12341
rect 1213 12311 1635 12315
tri 1635 12311 1665 12341 sw
tri 1733 12311 1763 12341 ne
rect 1763 12315 1865 12341
rect 1985 12341 2087 12435
tri 2087 12341 2185 12439 sw
tri 2185 12341 2283 12439 ne
rect 2283 12435 2637 12439
rect 2283 12341 2415 12435
rect 1985 12315 2185 12341
rect 1763 12311 2185 12315
tri 2185 12311 2215 12341 sw
tri 2283 12311 2313 12341 ne
rect 2313 12315 2415 12341
rect 2535 12341 2637 12435
tri 2637 12341 2735 12439 sw
tri 2735 12341 2833 12439 ne
rect 2833 12435 3187 12439
rect 2833 12341 2965 12435
rect 2535 12315 2735 12341
rect 2313 12311 2735 12315
tri 2735 12311 2765 12341 sw
tri 2833 12311 2863 12341 ne
rect 2863 12315 2965 12341
rect 3085 12341 3187 12435
tri 3187 12341 3285 12439 sw
tri 3285 12341 3383 12439 ne
rect 3383 12435 3737 12439
rect 3383 12341 3515 12435
rect 3085 12315 3285 12341
rect 2863 12311 3285 12315
tri 3285 12311 3315 12341 sw
tri 3383 12311 3413 12341 ne
rect 3413 12315 3515 12341
rect 3635 12341 3737 12435
tri 3737 12341 3835 12439 sw
tri 3835 12341 3933 12439 ne
rect 3933 12435 4287 12439
rect 3933 12341 4065 12435
rect 3635 12315 3835 12341
rect 3413 12311 3835 12315
tri 3835 12311 3865 12341 sw
tri 3933 12311 3963 12341 ne
rect 3963 12315 4065 12341
rect 4185 12341 4287 12435
tri 4287 12341 4385 12439 sw
tri 4385 12341 4483 12439 ne
rect 4483 12435 4837 12439
rect 4483 12341 4615 12435
rect 4185 12315 4385 12341
rect 3963 12311 4385 12315
tri 4385 12311 4415 12341 sw
tri 4483 12311 4513 12341 ne
rect 4513 12315 4615 12341
rect 4735 12341 4837 12435
tri 4837 12341 4935 12439 sw
tri 4935 12341 5033 12439 ne
rect 5033 12435 5387 12439
rect 5033 12341 5165 12435
rect 4735 12315 4935 12341
rect 4513 12311 4935 12315
tri 4935 12311 4965 12341 sw
tri 5033 12311 5063 12341 ne
rect 5063 12315 5165 12341
rect 5285 12341 5387 12435
tri 5387 12341 5485 12439 sw
tri 5485 12341 5583 12439 ne
rect 5583 12435 5937 12439
rect 5583 12341 5715 12435
rect 5285 12315 5485 12341
rect 5063 12311 5485 12315
tri 5485 12311 5515 12341 sw
tri 5583 12311 5613 12341 ne
rect 5613 12315 5715 12341
rect 5835 12341 5937 12435
tri 5937 12341 6035 12439 sw
tri 6035 12341 6133 12439 ne
rect 6133 12435 6487 12439
rect 6133 12341 6265 12435
rect 5835 12315 6035 12341
rect 5613 12311 6035 12315
tri 6035 12311 6065 12341 sw
tri 6133 12311 6163 12341 ne
rect 6163 12315 6265 12341
rect 6385 12341 6487 12435
tri 6487 12341 6585 12439 sw
tri 6585 12341 6683 12439 ne
rect 6683 12435 7037 12439
rect 6683 12341 6815 12435
rect 6385 12315 6585 12341
rect 6163 12311 6585 12315
tri 6585 12311 6615 12341 sw
tri 6683 12311 6713 12341 ne
rect 6713 12315 6815 12341
rect 6935 12341 7037 12435
tri 7037 12341 7135 12439 sw
tri 7135 12341 7233 12439 ne
rect 7233 12435 7587 12439
rect 7233 12341 7365 12435
rect 6935 12315 7135 12341
rect 6713 12311 7135 12315
tri 7135 12311 7165 12341 sw
tri 7233 12311 7263 12341 ne
rect 7263 12315 7365 12341
rect 7485 12341 7587 12435
tri 7587 12341 7685 12439 sw
tri 7685 12341 7783 12439 ne
rect 7783 12435 8137 12439
rect 7783 12341 7915 12435
rect 7485 12315 7685 12341
rect 7263 12311 7685 12315
tri 7685 12311 7715 12341 sw
tri 7783 12311 7813 12341 ne
rect 7813 12315 7915 12341
rect 8035 12341 8137 12435
tri 8137 12341 8235 12439 sw
tri 8235 12341 8333 12439 ne
rect 8333 12435 8687 12439
rect 8333 12341 8465 12435
rect 8035 12315 8235 12341
rect 7813 12311 8235 12315
tri 8235 12311 8265 12341 sw
tri 8333 12311 8363 12341 ne
rect 8363 12315 8465 12341
rect 8585 12341 8687 12435
tri 8687 12341 8785 12439 sw
tri 8785 12341 8883 12439 ne
rect 8883 12435 9237 12439
rect 8883 12341 9015 12435
rect 8585 12315 8785 12341
rect 8363 12311 8785 12315
tri 8785 12311 8815 12341 sw
tri 8883 12311 8913 12341 ne
rect 8913 12315 9015 12341
rect 9135 12341 9237 12435
tri 9237 12341 9335 12439 sw
tri 9335 12341 9433 12439 ne
rect 9433 12435 9787 12439
rect 9433 12341 9565 12435
rect 9135 12315 9335 12341
rect 8913 12311 9335 12315
tri 9335 12311 9365 12341 sw
tri 9433 12311 9463 12341 ne
rect 9463 12315 9565 12341
rect 9685 12341 9787 12435
tri 9787 12341 9885 12439 sw
tri 9885 12341 9983 12439 ne
rect 9983 12435 10337 12439
rect 9983 12341 10115 12435
rect 9685 12315 9885 12341
rect 9463 12311 9885 12315
tri 9885 12311 9915 12341 sw
tri 9983 12311 10013 12341 ne
rect 10013 12315 10115 12341
rect 10235 12341 10337 12435
tri 10337 12341 10435 12439 sw
tri 10435 12341 10533 12439 ne
rect 10533 12435 10887 12439
rect 10533 12341 10665 12435
rect 10235 12315 10435 12341
rect 10013 12311 10435 12315
tri 10435 12311 10465 12341 sw
tri 10533 12311 10563 12341 ne
rect 10563 12315 10665 12341
rect 10785 12341 10887 12435
tri 10887 12341 10985 12439 sw
tri 10985 12341 11083 12439 ne
rect 11083 12435 11437 12439
rect 11083 12341 11215 12435
rect 10785 12315 10985 12341
rect 10563 12311 10985 12315
tri 10985 12311 11015 12341 sw
tri 11083 12311 11113 12341 ne
rect 11113 12315 11215 12341
rect 11335 12341 11437 12435
tri 11437 12341 11535 12439 sw
tri 11535 12341 11633 12439 ne
rect 11633 12435 11987 12439
rect 11633 12341 11765 12435
rect 11335 12315 11535 12341
rect 11113 12311 11535 12315
tri 11535 12311 11565 12341 sw
tri 11633 12311 11663 12341 ne
rect 11663 12315 11765 12341
rect 11885 12341 11987 12435
tri 11987 12341 12085 12439 sw
tri 12085 12341 12183 12439 ne
rect 12183 12435 12537 12439
rect 12183 12341 12315 12435
rect 11885 12315 12085 12341
rect 11663 12311 12085 12315
tri 12085 12311 12115 12341 sw
tri 12183 12311 12213 12341 ne
rect 12213 12315 12315 12341
rect 12435 12341 12537 12435
tri 12537 12341 12635 12439 sw
tri 12635 12341 12733 12439 ne
rect 12733 12435 13087 12439
rect 12733 12341 12865 12435
rect 12435 12315 12635 12341
rect 12213 12311 12635 12315
tri 12635 12311 12665 12341 sw
tri 12733 12311 12763 12341 ne
rect 12763 12315 12865 12341
rect 12985 12341 13087 12435
tri 13087 12341 13185 12439 sw
tri 13185 12341 13283 12439 ne
rect 13283 12435 13637 12439
rect 13283 12341 13415 12435
rect 12985 12315 13185 12341
rect 12763 12311 13185 12315
tri 13185 12311 13215 12341 sw
tri 13283 12311 13313 12341 ne
rect 13313 12315 13415 12341
rect 13535 12341 13637 12435
tri 13637 12341 13735 12439 sw
tri 13735 12341 13833 12439 ne
rect 13833 12435 14187 12439
rect 13833 12341 13965 12435
rect 13535 12315 13735 12341
rect 13313 12311 13735 12315
tri 13735 12311 13765 12341 sw
tri 13833 12311 13863 12341 ne
rect 13863 12315 13965 12341
rect 14085 12341 14187 12435
tri 14187 12341 14285 12439 sw
tri 14285 12341 14383 12439 ne
rect 14383 12435 14737 12439
rect 14383 12341 14515 12435
rect 14085 12315 14285 12341
rect 13863 12311 14285 12315
tri 14285 12311 14315 12341 sw
tri 14383 12311 14413 12341 ne
rect 14413 12315 14515 12341
rect 14635 12341 14737 12435
tri 14737 12341 14835 12439 sw
tri 14835 12341 14933 12439 ne
rect 14933 12435 15287 12439
rect 14933 12341 15065 12435
rect 14635 12315 14835 12341
rect 14413 12311 14835 12315
tri 14835 12311 14865 12341 sw
tri 14933 12311 14963 12341 ne
rect 14963 12315 15065 12341
rect 15185 12341 15287 12435
tri 15287 12341 15385 12439 sw
tri 15385 12341 15483 12439 ne
rect 15483 12435 15837 12439
rect 15483 12341 15615 12435
rect 15185 12315 15385 12341
rect 14963 12311 15385 12315
tri 15385 12311 15415 12341 sw
tri 15483 12311 15513 12341 ne
rect 15513 12315 15615 12341
rect 15735 12341 15837 12435
tri 15837 12341 15935 12439 sw
tri 15935 12341 16033 12439 ne
rect 16033 12435 16387 12439
rect 16033 12341 16165 12435
rect 15735 12315 15935 12341
rect 15513 12311 15935 12315
tri 15935 12311 15965 12341 sw
tri 16033 12311 16063 12341 ne
rect 16063 12315 16165 12341
rect 16285 12341 16387 12435
tri 16387 12341 16485 12439 sw
tri 16485 12341 16583 12439 ne
rect 16583 12435 16937 12439
rect 16583 12341 16715 12435
rect 16285 12315 16485 12341
rect 16063 12311 16485 12315
tri 16485 12311 16515 12341 sw
tri 16583 12311 16613 12341 ne
rect 16613 12315 16715 12341
rect 16835 12341 16937 12435
tri 16937 12341 17035 12439 sw
tri 17035 12341 17133 12439 ne
rect 17133 12435 17487 12439
rect 17133 12341 17265 12435
rect 16835 12315 17035 12341
rect 16613 12311 17035 12315
tri 17035 12311 17065 12341 sw
tri 17133 12311 17163 12341 ne
rect 17163 12315 17265 12341
rect 17385 12341 17487 12435
tri 17487 12341 17585 12439 sw
tri 17585 12341 17683 12439 ne
rect 17683 12435 18037 12439
rect 17683 12341 17815 12435
rect 17385 12315 17585 12341
rect 17163 12311 17585 12315
tri 17585 12311 17615 12341 sw
tri 17683 12311 17713 12341 ne
rect 17713 12315 17815 12341
rect 17935 12341 18037 12435
tri 18037 12341 18135 12439 sw
tri 18135 12341 18233 12439 ne
rect 18233 12435 18587 12439
rect 18233 12341 18365 12435
rect 17935 12315 18135 12341
rect 17713 12311 18135 12315
tri 18135 12311 18165 12341 sw
tri 18233 12311 18263 12341 ne
rect 18263 12315 18365 12341
rect 18485 12341 18587 12435
tri 18587 12341 18685 12439 sw
tri 18685 12341 18783 12439 ne
rect 18783 12435 19137 12439
rect 18783 12341 18915 12435
rect 18485 12315 18685 12341
rect 18263 12311 18685 12315
tri 18685 12311 18715 12341 sw
tri 18783 12311 18813 12341 ne
rect 18813 12315 18915 12341
rect 19035 12341 19137 12435
tri 19137 12341 19235 12439 sw
tri 19235 12341 19333 12439 ne
rect 19333 12435 20300 12439
rect 19333 12341 19465 12435
rect 19035 12315 19235 12341
rect 18813 12311 19235 12315
tri 19235 12311 19265 12341 sw
tri 19333 12311 19363 12341 ne
rect 19363 12315 19465 12341
rect 19585 12315 20300 12435
rect 19363 12311 20300 12315
tri 113 12213 211 12311 ne
rect 211 12213 565 12311
tri 565 12213 663 12311 sw
tri 663 12213 761 12311 ne
rect 761 12213 1115 12311
tri 1115 12213 1213 12311 sw
tri 1213 12213 1311 12311 ne
rect 1311 12213 1665 12311
tri 1665 12213 1763 12311 sw
tri 1763 12213 1861 12311 ne
rect 1861 12213 2215 12311
tri 2215 12213 2313 12311 sw
tri 2313 12213 2411 12311 ne
rect 2411 12213 2765 12311
tri 2765 12213 2863 12311 sw
tri 2863 12213 2961 12311 ne
rect 2961 12213 3315 12311
tri 3315 12213 3413 12311 sw
tri 3413 12213 3511 12311 ne
rect 3511 12213 3865 12311
tri 3865 12213 3963 12311 sw
tri 3963 12213 4061 12311 ne
rect 4061 12213 4415 12311
tri 4415 12213 4513 12311 sw
tri 4513 12213 4611 12311 ne
rect 4611 12213 4965 12311
tri 4965 12213 5063 12311 sw
tri 5063 12213 5161 12311 ne
rect 5161 12213 5515 12311
tri 5515 12213 5613 12311 sw
tri 5613 12213 5711 12311 ne
rect 5711 12213 6065 12311
tri 6065 12213 6163 12311 sw
tri 6163 12213 6261 12311 ne
rect 6261 12213 6615 12311
tri 6615 12213 6713 12311 sw
tri 6713 12213 6811 12311 ne
rect 6811 12213 7165 12311
tri 7165 12213 7263 12311 sw
tri 7263 12213 7361 12311 ne
rect 7361 12213 7715 12311
tri 7715 12213 7813 12311 sw
tri 7813 12213 7911 12311 ne
rect 7911 12213 8265 12311
tri 8265 12213 8363 12311 sw
tri 8363 12213 8461 12311 ne
rect 8461 12213 8815 12311
tri 8815 12213 8913 12311 sw
tri 8913 12213 9011 12311 ne
rect 9011 12213 9365 12311
tri 9365 12213 9463 12311 sw
tri 9463 12213 9561 12311 ne
rect 9561 12213 9915 12311
tri 9915 12213 10013 12311 sw
tri 10013 12213 10111 12311 ne
rect 10111 12213 10465 12311
tri 10465 12213 10563 12311 sw
tri 10563 12213 10661 12311 ne
rect 10661 12213 11015 12311
tri 11015 12213 11113 12311 sw
tri 11113 12213 11211 12311 ne
rect 11211 12213 11565 12311
tri 11565 12213 11663 12311 sw
tri 11663 12213 11761 12311 ne
rect 11761 12213 12115 12311
tri 12115 12213 12213 12311 sw
tri 12213 12213 12311 12311 ne
rect 12311 12213 12665 12311
tri 12665 12213 12763 12311 sw
tri 12763 12213 12861 12311 ne
rect 12861 12213 13215 12311
tri 13215 12213 13313 12311 sw
tri 13313 12213 13411 12311 ne
rect 13411 12213 13765 12311
tri 13765 12213 13863 12311 sw
tri 13863 12213 13961 12311 ne
rect 13961 12213 14315 12311
tri 14315 12213 14413 12311 sw
tri 14413 12213 14511 12311 ne
rect 14511 12213 14865 12311
tri 14865 12213 14963 12311 sw
tri 14963 12213 15061 12311 ne
rect 15061 12213 15415 12311
tri 15415 12213 15513 12311 sw
tri 15513 12213 15611 12311 ne
rect 15611 12213 15965 12311
tri 15965 12213 16063 12311 sw
tri 16063 12213 16161 12311 ne
rect 16161 12213 16515 12311
tri 16515 12213 16613 12311 sw
tri 16613 12213 16711 12311 ne
rect 16711 12213 17065 12311
tri 17065 12213 17163 12311 sw
tri 17163 12213 17261 12311 ne
rect 17261 12213 17615 12311
tri 17615 12213 17713 12311 sw
tri 17713 12213 17811 12311 ne
rect 17811 12213 18165 12311
tri 18165 12213 18263 12311 sw
tri 18263 12213 18361 12311 ne
rect 18361 12213 18715 12311
tri 18715 12213 18813 12311 sw
tri 18813 12213 18911 12311 ne
rect 18911 12213 19265 12311
tri 19265 12213 19363 12311 sw
tri 19363 12213 19461 12311 ne
rect 19461 12213 20300 12311
rect -2000 12183 113 12213
tri 113 12183 143 12213 sw
tri 211 12183 241 12213 ne
rect 241 12183 663 12213
tri 663 12183 693 12213 sw
tri 761 12183 791 12213 ne
rect 791 12183 1213 12213
tri 1213 12183 1243 12213 sw
tri 1311 12183 1341 12213 ne
rect 1341 12183 1763 12213
tri 1763 12183 1793 12213 sw
tri 1861 12183 1891 12213 ne
rect 1891 12183 2313 12213
tri 2313 12183 2343 12213 sw
tri 2411 12183 2441 12213 ne
rect 2441 12183 2863 12213
tri 2863 12183 2893 12213 sw
tri 2961 12183 2991 12213 ne
rect 2991 12183 3413 12213
tri 3413 12183 3443 12213 sw
tri 3511 12183 3541 12213 ne
rect 3541 12183 3963 12213
tri 3963 12183 3993 12213 sw
tri 4061 12183 4091 12213 ne
rect 4091 12183 4513 12213
tri 4513 12183 4543 12213 sw
tri 4611 12183 4641 12213 ne
rect 4641 12183 5063 12213
tri 5063 12183 5093 12213 sw
tri 5161 12183 5191 12213 ne
rect 5191 12183 5613 12213
tri 5613 12183 5643 12213 sw
tri 5711 12183 5741 12213 ne
rect 5741 12183 6163 12213
tri 6163 12183 6193 12213 sw
tri 6261 12183 6291 12213 ne
rect 6291 12183 6713 12213
tri 6713 12183 6743 12213 sw
tri 6811 12183 6841 12213 ne
rect 6841 12183 7263 12213
tri 7263 12183 7293 12213 sw
tri 7361 12183 7391 12213 ne
rect 7391 12183 7813 12213
tri 7813 12183 7843 12213 sw
tri 7911 12183 7941 12213 ne
rect 7941 12183 8363 12213
tri 8363 12183 8393 12213 sw
tri 8461 12183 8491 12213 ne
rect 8491 12183 8913 12213
tri 8913 12183 8943 12213 sw
tri 9011 12183 9041 12213 ne
rect 9041 12183 9463 12213
tri 9463 12183 9493 12213 sw
tri 9561 12183 9591 12213 ne
rect 9591 12183 10013 12213
tri 10013 12183 10043 12213 sw
tri 10111 12183 10141 12213 ne
rect 10141 12183 10563 12213
tri 10563 12183 10593 12213 sw
tri 10661 12183 10691 12213 ne
rect 10691 12183 11113 12213
tri 11113 12183 11143 12213 sw
tri 11211 12183 11241 12213 ne
rect 11241 12183 11663 12213
tri 11663 12183 11693 12213 sw
tri 11761 12183 11791 12213 ne
rect 11791 12183 12213 12213
tri 12213 12183 12243 12213 sw
tri 12311 12183 12341 12213 ne
rect 12341 12183 12763 12213
tri 12763 12183 12793 12213 sw
tri 12861 12183 12891 12213 ne
rect 12891 12183 13313 12213
tri 13313 12183 13343 12213 sw
tri 13411 12183 13441 12213 ne
rect 13441 12183 13863 12213
tri 13863 12183 13893 12213 sw
tri 13961 12183 13991 12213 ne
rect 13991 12183 14413 12213
tri 14413 12183 14443 12213 sw
tri 14511 12183 14541 12213 ne
rect 14541 12183 14963 12213
tri 14963 12183 14993 12213 sw
tri 15061 12183 15091 12213 ne
rect 15091 12183 15513 12213
tri 15513 12183 15543 12213 sw
tri 15611 12183 15641 12213 ne
rect 15641 12183 16063 12213
tri 16063 12183 16093 12213 sw
tri 16161 12183 16191 12213 ne
rect 16191 12183 16613 12213
tri 16613 12183 16643 12213 sw
tri 16711 12183 16741 12213 ne
rect 16741 12183 17163 12213
tri 17163 12183 17193 12213 sw
tri 17261 12183 17291 12213 ne
rect 17291 12183 17713 12213
tri 17713 12183 17743 12213 sw
tri 17811 12183 17841 12213 ne
rect 17841 12183 18263 12213
tri 18263 12183 18293 12213 sw
tri 18361 12183 18391 12213 ne
rect 18391 12183 18813 12213
tri 18813 12183 18843 12213 sw
tri 18911 12183 18941 12213 ne
rect 18941 12183 19363 12213
tri 19363 12183 19393 12213 sw
tri 19461 12183 19491 12213 ne
rect 19491 12183 20300 12213
rect -2000 12085 143 12183
tri 143 12085 241 12183 sw
tri 241 12085 339 12183 ne
rect 339 12085 693 12183
tri 693 12085 791 12183 sw
tri 791 12085 889 12183 ne
rect 889 12085 1243 12183
tri 1243 12085 1341 12183 sw
tri 1341 12085 1439 12183 ne
rect 1439 12085 1793 12183
tri 1793 12085 1891 12183 sw
tri 1891 12085 1989 12183 ne
rect 1989 12085 2343 12183
tri 2343 12085 2441 12183 sw
tri 2441 12085 2539 12183 ne
rect 2539 12085 2893 12183
tri 2893 12085 2991 12183 sw
tri 2991 12085 3089 12183 ne
rect 3089 12085 3443 12183
tri 3443 12085 3541 12183 sw
tri 3541 12085 3639 12183 ne
rect 3639 12085 3993 12183
tri 3993 12085 4091 12183 sw
tri 4091 12085 4189 12183 ne
rect 4189 12085 4543 12183
tri 4543 12085 4641 12183 sw
tri 4641 12085 4739 12183 ne
rect 4739 12085 5093 12183
tri 5093 12085 5191 12183 sw
tri 5191 12085 5289 12183 ne
rect 5289 12085 5643 12183
tri 5643 12085 5741 12183 sw
tri 5741 12085 5839 12183 ne
rect 5839 12085 6193 12183
tri 6193 12085 6291 12183 sw
tri 6291 12085 6389 12183 ne
rect 6389 12085 6743 12183
tri 6743 12085 6841 12183 sw
tri 6841 12085 6939 12183 ne
rect 6939 12085 7293 12183
tri 7293 12085 7391 12183 sw
tri 7391 12085 7489 12183 ne
rect 7489 12085 7843 12183
tri 7843 12085 7941 12183 sw
tri 7941 12085 8039 12183 ne
rect 8039 12085 8393 12183
tri 8393 12085 8491 12183 sw
tri 8491 12085 8589 12183 ne
rect 8589 12085 8943 12183
tri 8943 12085 9041 12183 sw
tri 9041 12085 9139 12183 ne
rect 9139 12085 9493 12183
tri 9493 12085 9591 12183 sw
tri 9591 12085 9689 12183 ne
rect 9689 12085 10043 12183
tri 10043 12085 10141 12183 sw
tri 10141 12085 10239 12183 ne
rect 10239 12085 10593 12183
tri 10593 12085 10691 12183 sw
tri 10691 12085 10789 12183 ne
rect 10789 12085 11143 12183
tri 11143 12085 11241 12183 sw
tri 11241 12085 11339 12183 ne
rect 11339 12085 11693 12183
tri 11693 12085 11791 12183 sw
tri 11791 12085 11889 12183 ne
rect 11889 12085 12243 12183
tri 12243 12085 12341 12183 sw
tri 12341 12085 12439 12183 ne
rect 12439 12085 12793 12183
tri 12793 12085 12891 12183 sw
tri 12891 12085 12989 12183 ne
rect 12989 12085 13343 12183
tri 13343 12085 13441 12183 sw
tri 13441 12085 13539 12183 ne
rect 13539 12085 13893 12183
tri 13893 12085 13991 12183 sw
tri 13991 12085 14089 12183 ne
rect 14089 12085 14443 12183
tri 14443 12085 14541 12183 sw
tri 14541 12085 14639 12183 ne
rect 14639 12085 14993 12183
tri 14993 12085 15091 12183 sw
tri 15091 12085 15189 12183 ne
rect 15189 12085 15543 12183
tri 15543 12085 15641 12183 sw
tri 15641 12085 15739 12183 ne
rect 15739 12085 16093 12183
tri 16093 12085 16191 12183 sw
tri 16191 12085 16289 12183 ne
rect 16289 12085 16643 12183
tri 16643 12085 16741 12183 sw
tri 16741 12085 16839 12183 ne
rect 16839 12085 17193 12183
tri 17193 12085 17291 12183 sw
tri 17291 12085 17389 12183 ne
rect 17389 12085 17743 12183
tri 17743 12085 17841 12183 sw
tri 17841 12085 17939 12183 ne
rect 17939 12085 18293 12183
tri 18293 12085 18391 12183 sw
tri 18391 12085 18489 12183 ne
rect 18489 12085 18843 12183
tri 18843 12085 18941 12183 sw
tri 18941 12085 19039 12183 ne
rect 19039 12085 19393 12183
tri 19393 12085 19491 12183 sw
tri 19491 12085 19589 12183 ne
rect 19589 12085 20300 12183
rect -2000 11987 241 12085
tri 241 11987 339 12085 sw
tri 339 11987 437 12085 ne
rect 437 11987 791 12085
tri 791 11987 889 12085 sw
tri 889 11987 987 12085 ne
rect 987 11987 1341 12085
tri 1341 11987 1439 12085 sw
tri 1439 11987 1537 12085 ne
rect 1537 11987 1891 12085
tri 1891 11987 1989 12085 sw
tri 1989 11987 2087 12085 ne
rect 2087 11987 2441 12085
tri 2441 11987 2539 12085 sw
tri 2539 11987 2637 12085 ne
rect 2637 11987 2991 12085
tri 2991 11987 3089 12085 sw
tri 3089 11987 3187 12085 ne
rect 3187 11987 3541 12085
tri 3541 11987 3639 12085 sw
tri 3639 11987 3737 12085 ne
rect 3737 11987 4091 12085
tri 4091 11987 4189 12085 sw
tri 4189 11987 4287 12085 ne
rect 4287 11987 4641 12085
tri 4641 11987 4739 12085 sw
tri 4739 11987 4837 12085 ne
rect 4837 11987 5191 12085
tri 5191 11987 5289 12085 sw
tri 5289 11987 5387 12085 ne
rect 5387 11987 5741 12085
tri 5741 11987 5839 12085 sw
tri 5839 11987 5937 12085 ne
rect 5937 11987 6291 12085
tri 6291 11987 6389 12085 sw
tri 6389 11987 6487 12085 ne
rect 6487 11987 6841 12085
tri 6841 11987 6939 12085 sw
tri 6939 11987 7037 12085 ne
rect 7037 11987 7391 12085
tri 7391 11987 7489 12085 sw
tri 7489 11987 7587 12085 ne
rect 7587 11987 7941 12085
tri 7941 11987 8039 12085 sw
tri 8039 11987 8137 12085 ne
rect 8137 11987 8491 12085
tri 8491 11987 8589 12085 sw
tri 8589 11987 8687 12085 ne
rect 8687 11987 9041 12085
tri 9041 11987 9139 12085 sw
tri 9139 11987 9237 12085 ne
rect 9237 11987 9591 12085
tri 9591 11987 9689 12085 sw
tri 9689 11987 9787 12085 ne
rect 9787 11987 10141 12085
tri 10141 11987 10239 12085 sw
tri 10239 11987 10337 12085 ne
rect 10337 11987 10691 12085
tri 10691 11987 10789 12085 sw
tri 10789 11987 10887 12085 ne
rect 10887 11987 11241 12085
tri 11241 11987 11339 12085 sw
tri 11339 11987 11437 12085 ne
rect 11437 11987 11791 12085
tri 11791 11987 11889 12085 sw
tri 11889 11987 11987 12085 ne
rect 11987 11987 12341 12085
tri 12341 11987 12439 12085 sw
tri 12439 11987 12537 12085 ne
rect 12537 11987 12891 12085
tri 12891 11987 12989 12085 sw
tri 12989 11987 13087 12085 ne
rect 13087 11987 13441 12085
tri 13441 11987 13539 12085 sw
tri 13539 11987 13637 12085 ne
rect 13637 11987 13991 12085
tri 13991 11987 14089 12085 sw
tri 14089 11987 14187 12085 ne
rect 14187 11987 14541 12085
tri 14541 11987 14639 12085 sw
tri 14639 11987 14737 12085 ne
rect 14737 11987 15091 12085
tri 15091 11987 15189 12085 sw
tri 15189 11987 15287 12085 ne
rect 15287 11987 15641 12085
tri 15641 11987 15739 12085 sw
tri 15739 11987 15837 12085 ne
rect 15837 11987 16191 12085
tri 16191 11987 16289 12085 sw
tri 16289 11987 16387 12085 ne
rect 16387 11987 16741 12085
tri 16741 11987 16839 12085 sw
tri 16839 11987 16937 12085 ne
rect 16937 11987 17291 12085
tri 17291 11987 17389 12085 sw
tri 17389 11987 17487 12085 ne
rect 17487 11987 17841 12085
tri 17841 11987 17939 12085 sw
tri 17939 11987 18037 12085 ne
rect 18037 11987 18391 12085
tri 18391 11987 18489 12085 sw
tri 18489 11987 18587 12085 ne
rect 18587 11987 18941 12085
tri 18941 11987 19039 12085 sw
tri 19039 11987 19137 12085 ne
rect 19137 11987 19491 12085
tri 19491 11987 19589 12085 sw
tri 19589 11987 19687 12085 ne
rect 19687 11987 20300 12085
rect -2000 11889 339 11987
tri 339 11889 437 11987 sw
tri 437 11889 535 11987 ne
rect 535 11889 889 11987
tri 889 11889 987 11987 sw
tri 987 11889 1085 11987 ne
rect 1085 11889 1439 11987
tri 1439 11889 1537 11987 sw
tri 1537 11889 1635 11987 ne
rect 1635 11889 1989 11987
tri 1989 11889 2087 11987 sw
tri 2087 11889 2185 11987 ne
rect 2185 11889 2539 11987
tri 2539 11889 2637 11987 sw
tri 2637 11889 2735 11987 ne
rect 2735 11889 3089 11987
tri 3089 11889 3187 11987 sw
tri 3187 11889 3285 11987 ne
rect 3285 11889 3639 11987
tri 3639 11889 3737 11987 sw
tri 3737 11889 3835 11987 ne
rect 3835 11889 4189 11987
tri 4189 11889 4287 11987 sw
tri 4287 11889 4385 11987 ne
rect 4385 11889 4739 11987
tri 4739 11889 4837 11987 sw
tri 4837 11889 4935 11987 ne
rect 4935 11889 5289 11987
tri 5289 11889 5387 11987 sw
tri 5387 11889 5485 11987 ne
rect 5485 11889 5839 11987
tri 5839 11889 5937 11987 sw
tri 5937 11889 6035 11987 ne
rect 6035 11889 6389 11987
tri 6389 11889 6487 11987 sw
tri 6487 11889 6585 11987 ne
rect 6585 11889 6939 11987
tri 6939 11889 7037 11987 sw
tri 7037 11889 7135 11987 ne
rect 7135 11889 7489 11987
tri 7489 11889 7587 11987 sw
tri 7587 11889 7685 11987 ne
rect 7685 11889 8039 11987
tri 8039 11889 8137 11987 sw
tri 8137 11889 8235 11987 ne
rect 8235 11889 8589 11987
tri 8589 11889 8687 11987 sw
tri 8687 11889 8785 11987 ne
rect 8785 11889 9139 11987
tri 9139 11889 9237 11987 sw
tri 9237 11889 9335 11987 ne
rect 9335 11889 9689 11987
tri 9689 11889 9787 11987 sw
tri 9787 11889 9885 11987 ne
rect 9885 11889 10239 11987
tri 10239 11889 10337 11987 sw
tri 10337 11889 10435 11987 ne
rect 10435 11889 10789 11987
tri 10789 11889 10887 11987 sw
tri 10887 11889 10985 11987 ne
rect 10985 11889 11339 11987
tri 11339 11889 11437 11987 sw
tri 11437 11889 11535 11987 ne
rect 11535 11889 11889 11987
tri 11889 11889 11987 11987 sw
tri 11987 11889 12085 11987 ne
rect 12085 11889 12439 11987
tri 12439 11889 12537 11987 sw
tri 12537 11889 12635 11987 ne
rect 12635 11889 12989 11987
tri 12989 11889 13087 11987 sw
tri 13087 11889 13185 11987 ne
rect 13185 11889 13539 11987
tri 13539 11889 13637 11987 sw
tri 13637 11889 13735 11987 ne
rect 13735 11889 14089 11987
tri 14089 11889 14187 11987 sw
tri 14187 11889 14285 11987 ne
rect 14285 11889 14639 11987
tri 14639 11889 14737 11987 sw
tri 14737 11889 14835 11987 ne
rect 14835 11889 15189 11987
tri 15189 11889 15287 11987 sw
tri 15287 11889 15385 11987 ne
rect 15385 11889 15739 11987
tri 15739 11889 15837 11987 sw
tri 15837 11889 15935 11987 ne
rect 15935 11889 16289 11987
tri 16289 11889 16387 11987 sw
tri 16387 11889 16485 11987 ne
rect 16485 11889 16839 11987
tri 16839 11889 16937 11987 sw
tri 16937 11889 17035 11987 ne
rect 17035 11889 17389 11987
tri 17389 11889 17487 11987 sw
tri 17487 11889 17585 11987 ne
rect 17585 11889 17939 11987
tri 17939 11889 18037 11987 sw
tri 18037 11889 18135 11987 ne
rect 18135 11889 18489 11987
tri 18489 11889 18587 11987 sw
tri 18587 11889 18685 11987 ne
rect 18685 11889 19039 11987
tri 19039 11889 19137 11987 sw
tri 19137 11889 19235 11987 ne
rect 19235 11889 19589 11987
tri 19589 11889 19687 11987 sw
rect 20800 11889 21800 12537
rect -2000 11885 437 11889
rect -2000 11765 215 11885
rect 335 11791 437 11885
tri 437 11791 535 11889 sw
tri 535 11791 633 11889 ne
rect 633 11885 987 11889
rect 633 11791 765 11885
rect 335 11765 535 11791
rect -2000 11761 535 11765
rect -2000 11113 -1000 11761
tri 113 11663 211 11761 ne
rect 211 11713 535 11761
tri 535 11713 613 11791 sw
tri 633 11713 711 11791 ne
rect 711 11765 765 11791
rect 885 11791 987 11885
tri 987 11791 1085 11889 sw
tri 1085 11791 1183 11889 ne
rect 1183 11885 1537 11889
rect 1183 11791 1315 11885
rect 885 11765 1085 11791
rect 711 11713 1085 11765
tri 1085 11713 1163 11791 sw
tri 1183 11713 1261 11791 ne
rect 1261 11765 1315 11791
rect 1435 11791 1537 11885
tri 1537 11791 1635 11889 sw
tri 1635 11791 1733 11889 ne
rect 1733 11885 2087 11889
rect 1733 11791 1865 11885
rect 1435 11765 1635 11791
rect 1261 11713 1635 11765
tri 1635 11713 1713 11791 sw
tri 1733 11713 1811 11791 ne
rect 1811 11765 1865 11791
rect 1985 11791 2087 11885
tri 2087 11791 2185 11889 sw
tri 2185 11791 2283 11889 ne
rect 2283 11885 2637 11889
rect 2283 11791 2415 11885
rect 1985 11765 2185 11791
rect 1811 11713 2185 11765
tri 2185 11713 2263 11791 sw
tri 2283 11713 2361 11791 ne
rect 2361 11765 2415 11791
rect 2535 11791 2637 11885
tri 2637 11791 2735 11889 sw
tri 2735 11791 2833 11889 ne
rect 2833 11885 3187 11889
rect 2833 11791 2965 11885
rect 2535 11765 2735 11791
rect 2361 11713 2735 11765
tri 2735 11713 2813 11791 sw
tri 2833 11713 2911 11791 ne
rect 2911 11765 2965 11791
rect 3085 11791 3187 11885
tri 3187 11791 3285 11889 sw
tri 3285 11791 3383 11889 ne
rect 3383 11885 3737 11889
rect 3383 11791 3515 11885
rect 3085 11765 3285 11791
rect 2911 11713 3285 11765
tri 3285 11713 3363 11791 sw
tri 3383 11713 3461 11791 ne
rect 3461 11765 3515 11791
rect 3635 11791 3737 11885
tri 3737 11791 3835 11889 sw
tri 3835 11791 3933 11889 ne
rect 3933 11885 4287 11889
rect 3933 11791 4065 11885
rect 3635 11765 3835 11791
rect 3461 11713 3835 11765
tri 3835 11713 3913 11791 sw
tri 3933 11713 4011 11791 ne
rect 4011 11765 4065 11791
rect 4185 11791 4287 11885
tri 4287 11791 4385 11889 sw
tri 4385 11791 4483 11889 ne
rect 4483 11885 4837 11889
rect 4483 11791 4615 11885
rect 4185 11765 4385 11791
rect 4011 11713 4385 11765
tri 4385 11713 4463 11791 sw
tri 4483 11713 4561 11791 ne
rect 4561 11765 4615 11791
rect 4735 11791 4837 11885
tri 4837 11791 4935 11889 sw
tri 4935 11791 5033 11889 ne
rect 5033 11885 5387 11889
rect 5033 11791 5165 11885
rect 4735 11765 4935 11791
rect 4561 11713 4935 11765
tri 4935 11713 5013 11791 sw
tri 5033 11713 5111 11791 ne
rect 5111 11765 5165 11791
rect 5285 11791 5387 11885
tri 5387 11791 5485 11889 sw
tri 5485 11791 5583 11889 ne
rect 5583 11885 5937 11889
rect 5583 11791 5715 11885
rect 5285 11765 5485 11791
rect 5111 11713 5485 11765
tri 5485 11713 5563 11791 sw
tri 5583 11713 5661 11791 ne
rect 5661 11765 5715 11791
rect 5835 11791 5937 11885
tri 5937 11791 6035 11889 sw
tri 6035 11791 6133 11889 ne
rect 6133 11885 6487 11889
rect 6133 11791 6265 11885
rect 5835 11765 6035 11791
rect 5661 11713 6035 11765
tri 6035 11713 6113 11791 sw
tri 6133 11713 6211 11791 ne
rect 6211 11765 6265 11791
rect 6385 11791 6487 11885
tri 6487 11791 6585 11889 sw
tri 6585 11791 6683 11889 ne
rect 6683 11885 7037 11889
rect 6683 11791 6815 11885
rect 6385 11765 6585 11791
rect 6211 11713 6585 11765
tri 6585 11713 6663 11791 sw
tri 6683 11713 6761 11791 ne
rect 6761 11765 6815 11791
rect 6935 11791 7037 11885
tri 7037 11791 7135 11889 sw
tri 7135 11791 7233 11889 ne
rect 7233 11885 7587 11889
rect 7233 11791 7365 11885
rect 6935 11765 7135 11791
rect 6761 11713 7135 11765
tri 7135 11713 7213 11791 sw
tri 7233 11713 7311 11791 ne
rect 7311 11765 7365 11791
rect 7485 11791 7587 11885
tri 7587 11791 7685 11889 sw
tri 7685 11791 7783 11889 ne
rect 7783 11885 8137 11889
rect 7783 11791 7915 11885
rect 7485 11765 7685 11791
rect 7311 11713 7685 11765
tri 7685 11713 7763 11791 sw
tri 7783 11713 7861 11791 ne
rect 7861 11765 7915 11791
rect 8035 11791 8137 11885
tri 8137 11791 8235 11889 sw
tri 8235 11791 8333 11889 ne
rect 8333 11885 8687 11889
rect 8333 11791 8465 11885
rect 8035 11765 8235 11791
rect 7861 11713 8235 11765
tri 8235 11713 8313 11791 sw
tri 8333 11713 8411 11791 ne
rect 8411 11765 8465 11791
rect 8585 11791 8687 11885
tri 8687 11791 8785 11889 sw
tri 8785 11791 8883 11889 ne
rect 8883 11885 9237 11889
rect 8883 11791 9015 11885
rect 8585 11765 8785 11791
rect 8411 11713 8785 11765
tri 8785 11713 8863 11791 sw
tri 8883 11713 8961 11791 ne
rect 8961 11765 9015 11791
rect 9135 11791 9237 11885
tri 9237 11791 9335 11889 sw
tri 9335 11791 9433 11889 ne
rect 9433 11885 9787 11889
rect 9433 11791 9565 11885
rect 9135 11765 9335 11791
rect 8961 11713 9335 11765
tri 9335 11713 9413 11791 sw
tri 9433 11713 9511 11791 ne
rect 9511 11765 9565 11791
rect 9685 11791 9787 11885
tri 9787 11791 9885 11889 sw
tri 9885 11791 9983 11889 ne
rect 9983 11885 10337 11889
rect 9983 11791 10115 11885
rect 9685 11765 9885 11791
rect 9511 11713 9885 11765
tri 9885 11713 9963 11791 sw
tri 9983 11713 10061 11791 ne
rect 10061 11765 10115 11791
rect 10235 11791 10337 11885
tri 10337 11791 10435 11889 sw
tri 10435 11791 10533 11889 ne
rect 10533 11885 10887 11889
rect 10533 11791 10665 11885
rect 10235 11765 10435 11791
rect 10061 11713 10435 11765
tri 10435 11713 10513 11791 sw
tri 10533 11713 10611 11791 ne
rect 10611 11765 10665 11791
rect 10785 11791 10887 11885
tri 10887 11791 10985 11889 sw
tri 10985 11791 11083 11889 ne
rect 11083 11885 11437 11889
rect 11083 11791 11215 11885
rect 10785 11765 10985 11791
rect 10611 11713 10985 11765
tri 10985 11713 11063 11791 sw
tri 11083 11713 11161 11791 ne
rect 11161 11765 11215 11791
rect 11335 11791 11437 11885
tri 11437 11791 11535 11889 sw
tri 11535 11791 11633 11889 ne
rect 11633 11885 11987 11889
rect 11633 11791 11765 11885
rect 11335 11765 11535 11791
rect 11161 11713 11535 11765
tri 11535 11713 11613 11791 sw
tri 11633 11713 11711 11791 ne
rect 11711 11765 11765 11791
rect 11885 11791 11987 11885
tri 11987 11791 12085 11889 sw
tri 12085 11791 12183 11889 ne
rect 12183 11885 12537 11889
rect 12183 11791 12315 11885
rect 11885 11765 12085 11791
rect 11711 11713 12085 11765
tri 12085 11713 12163 11791 sw
tri 12183 11713 12261 11791 ne
rect 12261 11765 12315 11791
rect 12435 11791 12537 11885
tri 12537 11791 12635 11889 sw
tri 12635 11791 12733 11889 ne
rect 12733 11885 13087 11889
rect 12733 11791 12865 11885
rect 12435 11765 12635 11791
rect 12261 11713 12635 11765
tri 12635 11713 12713 11791 sw
tri 12733 11713 12811 11791 ne
rect 12811 11765 12865 11791
rect 12985 11791 13087 11885
tri 13087 11791 13185 11889 sw
tri 13185 11791 13283 11889 ne
rect 13283 11885 13637 11889
rect 13283 11791 13415 11885
rect 12985 11765 13185 11791
rect 12811 11713 13185 11765
tri 13185 11713 13263 11791 sw
tri 13283 11713 13361 11791 ne
rect 13361 11765 13415 11791
rect 13535 11791 13637 11885
tri 13637 11791 13735 11889 sw
tri 13735 11791 13833 11889 ne
rect 13833 11885 14187 11889
rect 13833 11791 13965 11885
rect 13535 11765 13735 11791
rect 13361 11713 13735 11765
tri 13735 11713 13813 11791 sw
tri 13833 11713 13911 11791 ne
rect 13911 11765 13965 11791
rect 14085 11791 14187 11885
tri 14187 11791 14285 11889 sw
tri 14285 11791 14383 11889 ne
rect 14383 11885 14737 11889
rect 14383 11791 14515 11885
rect 14085 11765 14285 11791
rect 13911 11713 14285 11765
tri 14285 11713 14363 11791 sw
tri 14383 11713 14461 11791 ne
rect 14461 11765 14515 11791
rect 14635 11791 14737 11885
tri 14737 11791 14835 11889 sw
tri 14835 11791 14933 11889 ne
rect 14933 11885 15287 11889
rect 14933 11791 15065 11885
rect 14635 11765 14835 11791
rect 14461 11713 14835 11765
tri 14835 11713 14913 11791 sw
tri 14933 11713 15011 11791 ne
rect 15011 11765 15065 11791
rect 15185 11791 15287 11885
tri 15287 11791 15385 11889 sw
tri 15385 11791 15483 11889 ne
rect 15483 11885 15837 11889
rect 15483 11791 15615 11885
rect 15185 11765 15385 11791
rect 15011 11713 15385 11765
tri 15385 11713 15463 11791 sw
tri 15483 11713 15561 11791 ne
rect 15561 11765 15615 11791
rect 15735 11791 15837 11885
tri 15837 11791 15935 11889 sw
tri 15935 11791 16033 11889 ne
rect 16033 11885 16387 11889
rect 16033 11791 16165 11885
rect 15735 11765 15935 11791
rect 15561 11713 15935 11765
tri 15935 11713 16013 11791 sw
tri 16033 11713 16111 11791 ne
rect 16111 11765 16165 11791
rect 16285 11791 16387 11885
tri 16387 11791 16485 11889 sw
tri 16485 11791 16583 11889 ne
rect 16583 11885 16937 11889
rect 16583 11791 16715 11885
rect 16285 11765 16485 11791
rect 16111 11713 16485 11765
tri 16485 11713 16563 11791 sw
tri 16583 11713 16661 11791 ne
rect 16661 11765 16715 11791
rect 16835 11791 16937 11885
tri 16937 11791 17035 11889 sw
tri 17035 11791 17133 11889 ne
rect 17133 11885 17487 11889
rect 17133 11791 17265 11885
rect 16835 11765 17035 11791
rect 16661 11713 17035 11765
tri 17035 11713 17113 11791 sw
tri 17133 11713 17211 11791 ne
rect 17211 11765 17265 11791
rect 17385 11791 17487 11885
tri 17487 11791 17585 11889 sw
tri 17585 11791 17683 11889 ne
rect 17683 11885 18037 11889
rect 17683 11791 17815 11885
rect 17385 11765 17585 11791
rect 17211 11713 17585 11765
tri 17585 11713 17663 11791 sw
tri 17683 11713 17761 11791 ne
rect 17761 11765 17815 11791
rect 17935 11791 18037 11885
tri 18037 11791 18135 11889 sw
tri 18135 11791 18233 11889 ne
rect 18233 11885 18587 11889
rect 18233 11791 18365 11885
rect 17935 11765 18135 11791
rect 17761 11713 18135 11765
tri 18135 11713 18213 11791 sw
tri 18233 11713 18311 11791 ne
rect 18311 11765 18365 11791
rect 18485 11791 18587 11885
tri 18587 11791 18685 11889 sw
tri 18685 11791 18783 11889 ne
rect 18783 11885 19137 11889
rect 18783 11791 18915 11885
rect 18485 11765 18685 11791
rect 18311 11713 18685 11765
tri 18685 11713 18763 11791 sw
tri 18783 11713 18861 11791 ne
rect 18861 11765 18915 11791
rect 19035 11791 19137 11885
tri 19137 11791 19235 11889 sw
tri 19235 11791 19333 11889 ne
rect 19333 11885 21800 11889
rect 19333 11791 19465 11885
rect 19035 11765 19235 11791
rect 18861 11713 19235 11765
tri 19235 11713 19313 11791 sw
tri 19333 11713 19411 11791 ne
rect 19411 11765 19465 11791
rect 19585 11765 21800 11885
rect 19411 11713 21800 11765
rect 211 11663 613 11713
rect -500 11613 113 11663
tri 113 11613 163 11663 sw
tri 211 11613 261 11663 ne
rect 261 11633 613 11663
tri 613 11633 693 11713 sw
tri 711 11633 791 11713 ne
rect 791 11633 1163 11713
tri 1163 11633 1243 11713 sw
tri 1261 11633 1341 11713 ne
rect 1341 11633 1713 11713
tri 1713 11633 1793 11713 sw
tri 1811 11633 1891 11713 ne
rect 1891 11633 2263 11713
tri 2263 11633 2343 11713 sw
tri 2361 11633 2441 11713 ne
rect 2441 11633 2813 11713
tri 2813 11633 2893 11713 sw
tri 2911 11633 2991 11713 ne
rect 2991 11633 3363 11713
tri 3363 11633 3443 11713 sw
tri 3461 11633 3541 11713 ne
rect 3541 11633 3913 11713
tri 3913 11633 3993 11713 sw
tri 4011 11633 4091 11713 ne
rect 4091 11633 4463 11713
tri 4463 11633 4543 11713 sw
tri 4561 11633 4641 11713 ne
rect 4641 11633 5013 11713
tri 5013 11633 5093 11713 sw
tri 5111 11633 5191 11713 ne
rect 5191 11633 5563 11713
tri 5563 11633 5643 11713 sw
tri 5661 11633 5741 11713 ne
rect 5741 11633 6113 11713
tri 6113 11633 6193 11713 sw
tri 6211 11633 6291 11713 ne
rect 6291 11633 6663 11713
tri 6663 11633 6743 11713 sw
tri 6761 11633 6841 11713 ne
rect 6841 11633 7213 11713
tri 7213 11633 7293 11713 sw
tri 7311 11633 7391 11713 ne
rect 7391 11633 7763 11713
tri 7763 11633 7843 11713 sw
tri 7861 11633 7941 11713 ne
rect 7941 11633 8313 11713
tri 8313 11633 8393 11713 sw
tri 8411 11633 8491 11713 ne
rect 8491 11633 8863 11713
tri 8863 11633 8943 11713 sw
tri 8961 11633 9041 11713 ne
rect 9041 11633 9413 11713
tri 9413 11633 9493 11713 sw
tri 9511 11633 9591 11713 ne
rect 9591 11633 9963 11713
tri 9963 11633 10043 11713 sw
tri 10061 11633 10141 11713 ne
rect 10141 11633 10513 11713
tri 10513 11633 10593 11713 sw
tri 10611 11633 10691 11713 ne
rect 10691 11633 11063 11713
tri 11063 11633 11143 11713 sw
tri 11161 11633 11241 11713 ne
rect 11241 11633 11613 11713
tri 11613 11633 11693 11713 sw
tri 11711 11633 11791 11713 ne
rect 11791 11633 12163 11713
tri 12163 11633 12243 11713 sw
tri 12261 11633 12341 11713 ne
rect 12341 11633 12713 11713
tri 12713 11633 12793 11713 sw
tri 12811 11633 12891 11713 ne
rect 12891 11633 13263 11713
tri 13263 11633 13343 11713 sw
tri 13361 11633 13441 11713 ne
rect 13441 11633 13813 11713
tri 13813 11633 13893 11713 sw
tri 13911 11633 13991 11713 ne
rect 13991 11633 14363 11713
tri 14363 11633 14443 11713 sw
tri 14461 11633 14541 11713 ne
rect 14541 11633 14913 11713
tri 14913 11633 14993 11713 sw
tri 15011 11633 15091 11713 ne
rect 15091 11633 15463 11713
tri 15463 11633 15543 11713 sw
tri 15561 11633 15641 11713 ne
rect 15641 11633 16013 11713
tri 16013 11633 16093 11713 sw
tri 16111 11633 16191 11713 ne
rect 16191 11633 16563 11713
tri 16563 11633 16643 11713 sw
tri 16661 11633 16741 11713 ne
rect 16741 11633 17113 11713
tri 17113 11633 17193 11713 sw
tri 17211 11633 17291 11713 ne
rect 17291 11633 17663 11713
tri 17663 11633 17743 11713 sw
tri 17761 11633 17841 11713 ne
rect 17841 11633 18213 11713
tri 18213 11633 18293 11713 sw
tri 18311 11633 18391 11713 ne
rect 18391 11633 18763 11713
tri 18763 11633 18843 11713 sw
tri 18861 11633 18941 11713 ne
rect 18941 11633 19313 11713
tri 19313 11633 19393 11713 sw
tri 19411 11633 19491 11713 ne
rect 19491 11633 20100 11713
rect 261 11613 693 11633
rect -500 11535 163 11613
tri 163 11535 241 11613 sw
tri 261 11535 339 11613 ne
rect 339 11535 693 11613
tri 693 11535 791 11633 sw
tri 791 11535 889 11633 ne
rect 889 11535 1243 11633
tri 1243 11535 1341 11633 sw
tri 1341 11535 1439 11633 ne
rect 1439 11535 1793 11633
tri 1793 11535 1891 11633 sw
tri 1891 11535 1989 11633 ne
rect 1989 11535 2343 11633
tri 2343 11535 2441 11633 sw
tri 2441 11535 2539 11633 ne
rect 2539 11535 2893 11633
tri 2893 11535 2991 11633 sw
tri 2991 11535 3089 11633 ne
rect 3089 11535 3443 11633
tri 3443 11535 3541 11633 sw
tri 3541 11535 3639 11633 ne
rect 3639 11535 3993 11633
tri 3993 11535 4091 11633 sw
tri 4091 11535 4189 11633 ne
rect 4189 11535 4543 11633
tri 4543 11535 4641 11633 sw
tri 4641 11535 4739 11633 ne
rect 4739 11535 5093 11633
tri 5093 11535 5191 11633 sw
tri 5191 11535 5289 11633 ne
rect 5289 11535 5643 11633
tri 5643 11535 5741 11633 sw
tri 5741 11535 5839 11633 ne
rect 5839 11535 6193 11633
tri 6193 11535 6291 11633 sw
tri 6291 11535 6389 11633 ne
rect 6389 11535 6743 11633
tri 6743 11535 6841 11633 sw
tri 6841 11535 6939 11633 ne
rect 6939 11535 7293 11633
tri 7293 11535 7391 11633 sw
tri 7391 11535 7489 11633 ne
rect 7489 11535 7843 11633
tri 7843 11535 7941 11633 sw
tri 7941 11535 8039 11633 ne
rect 8039 11535 8393 11633
tri 8393 11535 8491 11633 sw
tri 8491 11535 8589 11633 ne
rect 8589 11535 8943 11633
tri 8943 11535 9041 11633 sw
tri 9041 11535 9139 11633 ne
rect 9139 11535 9493 11633
tri 9493 11535 9591 11633 sw
tri 9591 11535 9689 11633 ne
rect 9689 11535 10043 11633
tri 10043 11535 10141 11633 sw
tri 10141 11535 10239 11633 ne
rect 10239 11535 10593 11633
tri 10593 11535 10691 11633 sw
tri 10691 11535 10789 11633 ne
rect 10789 11535 11143 11633
tri 11143 11535 11241 11633 sw
tri 11241 11535 11339 11633 ne
rect 11339 11535 11693 11633
tri 11693 11535 11791 11633 sw
tri 11791 11535 11889 11633 ne
rect 11889 11535 12243 11633
tri 12243 11535 12341 11633 sw
tri 12341 11535 12439 11633 ne
rect 12439 11535 12793 11633
tri 12793 11535 12891 11633 sw
tri 12891 11535 12989 11633 ne
rect 12989 11535 13343 11633
tri 13343 11535 13441 11633 sw
tri 13441 11535 13539 11633 ne
rect 13539 11535 13893 11633
tri 13893 11535 13991 11633 sw
tri 13991 11535 14089 11633 ne
rect 14089 11535 14443 11633
tri 14443 11535 14541 11633 sw
tri 14541 11535 14639 11633 ne
rect 14639 11535 14993 11633
tri 14993 11535 15091 11633 sw
tri 15091 11535 15189 11633 ne
rect 15189 11535 15543 11633
tri 15543 11535 15641 11633 sw
tri 15641 11535 15739 11633 ne
rect 15739 11535 16093 11633
tri 16093 11535 16191 11633 sw
tri 16191 11535 16289 11633 ne
rect 16289 11535 16643 11633
tri 16643 11535 16741 11633 sw
tri 16741 11535 16839 11633 ne
rect 16839 11535 17193 11633
tri 17193 11535 17291 11633 sw
tri 17291 11535 17389 11633 ne
rect 17389 11535 17743 11633
tri 17743 11535 17841 11633 sw
tri 17841 11535 17939 11633 ne
rect 17939 11535 18293 11633
tri 18293 11535 18391 11633 sw
tri 18391 11535 18489 11633 ne
rect 18489 11535 18843 11633
tri 18843 11535 18941 11633 sw
tri 18941 11535 19039 11633 ne
rect 19039 11535 19393 11633
tri 19393 11535 19491 11633 sw
tri 19491 11535 19589 11633 ne
rect 19589 11613 20100 11633
rect 20200 11613 21800 11713
rect 19589 11535 21800 11613
rect -500 11487 241 11535
rect -500 11387 -400 11487
rect -300 11437 241 11487
tri 241 11437 339 11535 sw
tri 339 11437 437 11535 ne
rect 437 11437 791 11535
tri 791 11437 889 11535 sw
tri 889 11437 987 11535 ne
rect 987 11437 1341 11535
tri 1341 11437 1439 11535 sw
tri 1439 11437 1537 11535 ne
rect 1537 11437 1891 11535
tri 1891 11437 1989 11535 sw
tri 1989 11437 2087 11535 ne
rect 2087 11437 2441 11535
tri 2441 11437 2539 11535 sw
tri 2539 11437 2637 11535 ne
rect 2637 11437 2991 11535
tri 2991 11437 3089 11535 sw
tri 3089 11437 3187 11535 ne
rect 3187 11437 3541 11535
tri 3541 11437 3639 11535 sw
tri 3639 11437 3737 11535 ne
rect 3737 11437 4091 11535
tri 4091 11437 4189 11535 sw
tri 4189 11437 4287 11535 ne
rect 4287 11437 4641 11535
tri 4641 11437 4739 11535 sw
tri 4739 11437 4837 11535 ne
rect 4837 11437 5191 11535
tri 5191 11437 5289 11535 sw
tri 5289 11437 5387 11535 ne
rect 5387 11437 5741 11535
tri 5741 11437 5839 11535 sw
tri 5839 11437 5937 11535 ne
rect 5937 11437 6291 11535
tri 6291 11437 6389 11535 sw
tri 6389 11437 6487 11535 ne
rect 6487 11437 6841 11535
tri 6841 11437 6939 11535 sw
tri 6939 11437 7037 11535 ne
rect 7037 11437 7391 11535
tri 7391 11437 7489 11535 sw
tri 7489 11437 7587 11535 ne
rect 7587 11437 7941 11535
tri 7941 11437 8039 11535 sw
tri 8039 11437 8137 11535 ne
rect 8137 11437 8491 11535
tri 8491 11437 8589 11535 sw
tri 8589 11437 8687 11535 ne
rect 8687 11437 9041 11535
tri 9041 11437 9139 11535 sw
tri 9139 11437 9237 11535 ne
rect 9237 11437 9591 11535
tri 9591 11437 9689 11535 sw
tri 9689 11437 9787 11535 ne
rect 9787 11437 10141 11535
tri 10141 11437 10239 11535 sw
tri 10239 11437 10337 11535 ne
rect 10337 11437 10691 11535
tri 10691 11437 10789 11535 sw
tri 10789 11437 10887 11535 ne
rect 10887 11437 11241 11535
tri 11241 11437 11339 11535 sw
tri 11339 11437 11437 11535 ne
rect 11437 11437 11791 11535
tri 11791 11437 11889 11535 sw
tri 11889 11437 11987 11535 ne
rect 11987 11437 12341 11535
tri 12341 11437 12439 11535 sw
tri 12439 11437 12537 11535 ne
rect 12537 11437 12891 11535
tri 12891 11437 12989 11535 sw
tri 12989 11437 13087 11535 ne
rect 13087 11437 13441 11535
tri 13441 11437 13539 11535 sw
tri 13539 11437 13637 11535 ne
rect 13637 11437 13991 11535
tri 13991 11437 14089 11535 sw
tri 14089 11437 14187 11535 ne
rect 14187 11437 14541 11535
tri 14541 11437 14639 11535 sw
tri 14639 11437 14737 11535 ne
rect 14737 11437 15091 11535
tri 15091 11437 15189 11535 sw
tri 15189 11437 15287 11535 ne
rect 15287 11437 15641 11535
tri 15641 11437 15739 11535 sw
tri 15739 11437 15837 11535 ne
rect 15837 11437 16191 11535
tri 16191 11437 16289 11535 sw
tri 16289 11437 16387 11535 ne
rect 16387 11437 16741 11535
tri 16741 11437 16839 11535 sw
tri 16839 11437 16937 11535 ne
rect 16937 11437 17291 11535
tri 17291 11437 17389 11535 sw
tri 17389 11437 17487 11535 ne
rect 17487 11437 17841 11535
tri 17841 11437 17939 11535 sw
tri 17939 11437 18037 11535 ne
rect 18037 11437 18391 11535
tri 18391 11437 18489 11535 sw
tri 18489 11437 18587 11535 ne
rect 18587 11437 18941 11535
tri 18941 11437 19039 11535 sw
tri 19039 11437 19137 11535 ne
rect 19137 11437 19491 11535
tri 19491 11437 19589 11535 sw
tri 19589 11437 19687 11535 ne
rect 19687 11437 21800 11535
rect -300 11387 339 11437
rect -500 11339 339 11387
tri 339 11339 437 11437 sw
tri 437 11339 535 11437 ne
rect 535 11339 889 11437
tri 889 11339 987 11437 sw
tri 987 11339 1085 11437 ne
rect 1085 11339 1439 11437
tri 1439 11339 1537 11437 sw
tri 1537 11339 1635 11437 ne
rect 1635 11339 1989 11437
tri 1989 11339 2087 11437 sw
tri 2087 11339 2185 11437 ne
rect 2185 11339 2539 11437
tri 2539 11339 2637 11437 sw
tri 2637 11339 2735 11437 ne
rect 2735 11339 3089 11437
tri 3089 11339 3187 11437 sw
tri 3187 11339 3285 11437 ne
rect 3285 11339 3639 11437
tri 3639 11339 3737 11437 sw
tri 3737 11339 3835 11437 ne
rect 3835 11339 4189 11437
tri 4189 11339 4287 11437 sw
tri 4287 11339 4385 11437 ne
rect 4385 11339 4739 11437
tri 4739 11339 4837 11437 sw
tri 4837 11339 4935 11437 ne
rect 4935 11339 5289 11437
tri 5289 11339 5387 11437 sw
tri 5387 11339 5485 11437 ne
rect 5485 11339 5839 11437
tri 5839 11339 5937 11437 sw
tri 5937 11339 6035 11437 ne
rect 6035 11339 6389 11437
tri 6389 11339 6487 11437 sw
tri 6487 11339 6585 11437 ne
rect 6585 11339 6939 11437
tri 6939 11339 7037 11437 sw
tri 7037 11339 7135 11437 ne
rect 7135 11339 7489 11437
tri 7489 11339 7587 11437 sw
tri 7587 11339 7685 11437 ne
rect 7685 11339 8039 11437
tri 8039 11339 8137 11437 sw
tri 8137 11339 8235 11437 ne
rect 8235 11339 8589 11437
tri 8589 11339 8687 11437 sw
tri 8687 11339 8785 11437 ne
rect 8785 11339 9139 11437
tri 9139 11339 9237 11437 sw
tri 9237 11339 9335 11437 ne
rect 9335 11339 9689 11437
tri 9689 11339 9787 11437 sw
tri 9787 11339 9885 11437 ne
rect 9885 11339 10239 11437
tri 10239 11339 10337 11437 sw
tri 10337 11339 10435 11437 ne
rect 10435 11339 10789 11437
tri 10789 11339 10887 11437 sw
tri 10887 11339 10985 11437 ne
rect 10985 11339 11339 11437
tri 11339 11339 11437 11437 sw
tri 11437 11339 11535 11437 ne
rect 11535 11339 11889 11437
tri 11889 11339 11987 11437 sw
tri 11987 11339 12085 11437 ne
rect 12085 11339 12439 11437
tri 12439 11339 12537 11437 sw
tri 12537 11339 12635 11437 ne
rect 12635 11339 12989 11437
tri 12989 11339 13087 11437 sw
tri 13087 11339 13185 11437 ne
rect 13185 11339 13539 11437
tri 13539 11339 13637 11437 sw
tri 13637 11339 13735 11437 ne
rect 13735 11339 14089 11437
tri 14089 11339 14187 11437 sw
tri 14187 11339 14285 11437 ne
rect 14285 11339 14639 11437
tri 14639 11339 14737 11437 sw
tri 14737 11339 14835 11437 ne
rect 14835 11339 15189 11437
tri 15189 11339 15287 11437 sw
tri 15287 11339 15385 11437 ne
rect 15385 11339 15739 11437
tri 15739 11339 15837 11437 sw
tri 15837 11339 15935 11437 ne
rect 15935 11339 16289 11437
tri 16289 11339 16387 11437 sw
tri 16387 11339 16485 11437 ne
rect 16485 11339 16839 11437
tri 16839 11339 16937 11437 sw
tri 16937 11339 17035 11437 ne
rect 17035 11339 17389 11437
tri 17389 11339 17487 11437 sw
tri 17487 11339 17585 11437 ne
rect 17585 11339 17939 11437
tri 17939 11339 18037 11437 sw
tri 18037 11339 18135 11437 ne
rect 18135 11339 18489 11437
tri 18489 11339 18587 11437 sw
tri 18587 11339 18685 11437 ne
rect 18685 11339 19039 11437
tri 19039 11339 19137 11437 sw
tri 19137 11339 19235 11437 ne
rect 19235 11339 19589 11437
tri 19589 11339 19687 11437 sw
rect -500 11335 437 11339
rect -500 11215 215 11335
rect 335 11241 437 11335
tri 437 11241 535 11339 sw
tri 535 11241 633 11339 ne
rect 633 11335 987 11339
rect 633 11241 765 11335
rect 335 11215 535 11241
rect -500 11211 535 11215
tri 535 11211 565 11241 sw
tri 633 11211 663 11241 ne
rect 663 11215 765 11241
rect 885 11241 987 11335
tri 987 11241 1085 11339 sw
tri 1085 11241 1183 11339 ne
rect 1183 11335 1537 11339
rect 1183 11241 1315 11335
rect 885 11215 1085 11241
rect 663 11211 1085 11215
tri 1085 11211 1115 11241 sw
tri 1183 11211 1213 11241 ne
rect 1213 11215 1315 11241
rect 1435 11241 1537 11335
tri 1537 11241 1635 11339 sw
tri 1635 11241 1733 11339 ne
rect 1733 11335 2087 11339
rect 1733 11241 1865 11335
rect 1435 11215 1635 11241
rect 1213 11211 1635 11215
tri 1635 11211 1665 11241 sw
tri 1733 11211 1763 11241 ne
rect 1763 11215 1865 11241
rect 1985 11241 2087 11335
tri 2087 11241 2185 11339 sw
tri 2185 11241 2283 11339 ne
rect 2283 11335 2637 11339
rect 2283 11241 2415 11335
rect 1985 11215 2185 11241
rect 1763 11211 2185 11215
tri 2185 11211 2215 11241 sw
tri 2283 11211 2313 11241 ne
rect 2313 11215 2415 11241
rect 2535 11241 2637 11335
tri 2637 11241 2735 11339 sw
tri 2735 11241 2833 11339 ne
rect 2833 11335 3187 11339
rect 2833 11241 2965 11335
rect 2535 11215 2735 11241
rect 2313 11211 2735 11215
tri 2735 11211 2765 11241 sw
tri 2833 11211 2863 11241 ne
rect 2863 11215 2965 11241
rect 3085 11241 3187 11335
tri 3187 11241 3285 11339 sw
tri 3285 11241 3383 11339 ne
rect 3383 11335 3737 11339
rect 3383 11241 3515 11335
rect 3085 11215 3285 11241
rect 2863 11211 3285 11215
tri 3285 11211 3315 11241 sw
tri 3383 11211 3413 11241 ne
rect 3413 11215 3515 11241
rect 3635 11241 3737 11335
tri 3737 11241 3835 11339 sw
tri 3835 11241 3933 11339 ne
rect 3933 11335 4287 11339
rect 3933 11241 4065 11335
rect 3635 11215 3835 11241
rect 3413 11211 3835 11215
tri 3835 11211 3865 11241 sw
tri 3933 11211 3963 11241 ne
rect 3963 11215 4065 11241
rect 4185 11241 4287 11335
tri 4287 11241 4385 11339 sw
tri 4385 11241 4483 11339 ne
rect 4483 11335 4837 11339
rect 4483 11241 4615 11335
rect 4185 11215 4385 11241
rect 3963 11211 4385 11215
tri 4385 11211 4415 11241 sw
tri 4483 11211 4513 11241 ne
rect 4513 11215 4615 11241
rect 4735 11241 4837 11335
tri 4837 11241 4935 11339 sw
tri 4935 11241 5033 11339 ne
rect 5033 11335 5387 11339
rect 5033 11241 5165 11335
rect 4735 11215 4935 11241
rect 4513 11211 4935 11215
tri 4935 11211 4965 11241 sw
tri 5033 11211 5063 11241 ne
rect 5063 11215 5165 11241
rect 5285 11241 5387 11335
tri 5387 11241 5485 11339 sw
tri 5485 11241 5583 11339 ne
rect 5583 11335 5937 11339
rect 5583 11241 5715 11335
rect 5285 11215 5485 11241
rect 5063 11211 5485 11215
tri 5485 11211 5515 11241 sw
tri 5583 11211 5613 11241 ne
rect 5613 11215 5715 11241
rect 5835 11241 5937 11335
tri 5937 11241 6035 11339 sw
tri 6035 11241 6133 11339 ne
rect 6133 11335 6487 11339
rect 6133 11241 6265 11335
rect 5835 11215 6035 11241
rect 5613 11211 6035 11215
tri 6035 11211 6065 11241 sw
tri 6133 11211 6163 11241 ne
rect 6163 11215 6265 11241
rect 6385 11241 6487 11335
tri 6487 11241 6585 11339 sw
tri 6585 11241 6683 11339 ne
rect 6683 11335 7037 11339
rect 6683 11241 6815 11335
rect 6385 11215 6585 11241
rect 6163 11211 6585 11215
tri 6585 11211 6615 11241 sw
tri 6683 11211 6713 11241 ne
rect 6713 11215 6815 11241
rect 6935 11241 7037 11335
tri 7037 11241 7135 11339 sw
tri 7135 11241 7233 11339 ne
rect 7233 11335 7587 11339
rect 7233 11241 7365 11335
rect 6935 11215 7135 11241
rect 6713 11211 7135 11215
tri 7135 11211 7165 11241 sw
tri 7233 11211 7263 11241 ne
rect 7263 11215 7365 11241
rect 7485 11241 7587 11335
tri 7587 11241 7685 11339 sw
tri 7685 11241 7783 11339 ne
rect 7783 11335 8137 11339
rect 7783 11241 7915 11335
rect 7485 11215 7685 11241
rect 7263 11211 7685 11215
tri 7685 11211 7715 11241 sw
tri 7783 11211 7813 11241 ne
rect 7813 11215 7915 11241
rect 8035 11241 8137 11335
tri 8137 11241 8235 11339 sw
tri 8235 11241 8333 11339 ne
rect 8333 11335 8687 11339
rect 8333 11241 8465 11335
rect 8035 11215 8235 11241
rect 7813 11211 8235 11215
tri 8235 11211 8265 11241 sw
tri 8333 11211 8363 11241 ne
rect 8363 11215 8465 11241
rect 8585 11241 8687 11335
tri 8687 11241 8785 11339 sw
tri 8785 11241 8883 11339 ne
rect 8883 11335 9237 11339
rect 8883 11241 9015 11335
rect 8585 11215 8785 11241
rect 8363 11211 8785 11215
tri 8785 11211 8815 11241 sw
tri 8883 11211 8913 11241 ne
rect 8913 11215 9015 11241
rect 9135 11241 9237 11335
tri 9237 11241 9335 11339 sw
tri 9335 11241 9433 11339 ne
rect 9433 11335 9787 11339
rect 9433 11241 9565 11335
rect 9135 11215 9335 11241
rect 8913 11211 9335 11215
tri 9335 11211 9365 11241 sw
tri 9433 11211 9463 11241 ne
rect 9463 11215 9565 11241
rect 9685 11241 9787 11335
tri 9787 11241 9885 11339 sw
tri 9885 11241 9983 11339 ne
rect 9983 11335 10337 11339
rect 9983 11241 10115 11335
rect 9685 11215 9885 11241
rect 9463 11211 9885 11215
tri 9885 11211 9915 11241 sw
tri 9983 11211 10013 11241 ne
rect 10013 11215 10115 11241
rect 10235 11241 10337 11335
tri 10337 11241 10435 11339 sw
tri 10435 11241 10533 11339 ne
rect 10533 11335 10887 11339
rect 10533 11241 10665 11335
rect 10235 11215 10435 11241
rect 10013 11211 10435 11215
tri 10435 11211 10465 11241 sw
tri 10533 11211 10563 11241 ne
rect 10563 11215 10665 11241
rect 10785 11241 10887 11335
tri 10887 11241 10985 11339 sw
tri 10985 11241 11083 11339 ne
rect 11083 11335 11437 11339
rect 11083 11241 11215 11335
rect 10785 11215 10985 11241
rect 10563 11211 10985 11215
tri 10985 11211 11015 11241 sw
tri 11083 11211 11113 11241 ne
rect 11113 11215 11215 11241
rect 11335 11241 11437 11335
tri 11437 11241 11535 11339 sw
tri 11535 11241 11633 11339 ne
rect 11633 11335 11987 11339
rect 11633 11241 11765 11335
rect 11335 11215 11535 11241
rect 11113 11211 11535 11215
tri 11535 11211 11565 11241 sw
tri 11633 11211 11663 11241 ne
rect 11663 11215 11765 11241
rect 11885 11241 11987 11335
tri 11987 11241 12085 11339 sw
tri 12085 11241 12183 11339 ne
rect 12183 11335 12537 11339
rect 12183 11241 12315 11335
rect 11885 11215 12085 11241
rect 11663 11211 12085 11215
tri 12085 11211 12115 11241 sw
tri 12183 11211 12213 11241 ne
rect 12213 11215 12315 11241
rect 12435 11241 12537 11335
tri 12537 11241 12635 11339 sw
tri 12635 11241 12733 11339 ne
rect 12733 11335 13087 11339
rect 12733 11241 12865 11335
rect 12435 11215 12635 11241
rect 12213 11211 12635 11215
tri 12635 11211 12665 11241 sw
tri 12733 11211 12763 11241 ne
rect 12763 11215 12865 11241
rect 12985 11241 13087 11335
tri 13087 11241 13185 11339 sw
tri 13185 11241 13283 11339 ne
rect 13283 11335 13637 11339
rect 13283 11241 13415 11335
rect 12985 11215 13185 11241
rect 12763 11211 13185 11215
tri 13185 11211 13215 11241 sw
tri 13283 11211 13313 11241 ne
rect 13313 11215 13415 11241
rect 13535 11241 13637 11335
tri 13637 11241 13735 11339 sw
tri 13735 11241 13833 11339 ne
rect 13833 11335 14187 11339
rect 13833 11241 13965 11335
rect 13535 11215 13735 11241
rect 13313 11211 13735 11215
tri 13735 11211 13765 11241 sw
tri 13833 11211 13863 11241 ne
rect 13863 11215 13965 11241
rect 14085 11241 14187 11335
tri 14187 11241 14285 11339 sw
tri 14285 11241 14383 11339 ne
rect 14383 11335 14737 11339
rect 14383 11241 14515 11335
rect 14085 11215 14285 11241
rect 13863 11211 14285 11215
tri 14285 11211 14315 11241 sw
tri 14383 11211 14413 11241 ne
rect 14413 11215 14515 11241
rect 14635 11241 14737 11335
tri 14737 11241 14835 11339 sw
tri 14835 11241 14933 11339 ne
rect 14933 11335 15287 11339
rect 14933 11241 15065 11335
rect 14635 11215 14835 11241
rect 14413 11211 14835 11215
tri 14835 11211 14865 11241 sw
tri 14933 11211 14963 11241 ne
rect 14963 11215 15065 11241
rect 15185 11241 15287 11335
tri 15287 11241 15385 11339 sw
tri 15385 11241 15483 11339 ne
rect 15483 11335 15837 11339
rect 15483 11241 15615 11335
rect 15185 11215 15385 11241
rect 14963 11211 15385 11215
tri 15385 11211 15415 11241 sw
tri 15483 11211 15513 11241 ne
rect 15513 11215 15615 11241
rect 15735 11241 15837 11335
tri 15837 11241 15935 11339 sw
tri 15935 11241 16033 11339 ne
rect 16033 11335 16387 11339
rect 16033 11241 16165 11335
rect 15735 11215 15935 11241
rect 15513 11211 15935 11215
tri 15935 11211 15965 11241 sw
tri 16033 11211 16063 11241 ne
rect 16063 11215 16165 11241
rect 16285 11241 16387 11335
tri 16387 11241 16485 11339 sw
tri 16485 11241 16583 11339 ne
rect 16583 11335 16937 11339
rect 16583 11241 16715 11335
rect 16285 11215 16485 11241
rect 16063 11211 16485 11215
tri 16485 11211 16515 11241 sw
tri 16583 11211 16613 11241 ne
rect 16613 11215 16715 11241
rect 16835 11241 16937 11335
tri 16937 11241 17035 11339 sw
tri 17035 11241 17133 11339 ne
rect 17133 11335 17487 11339
rect 17133 11241 17265 11335
rect 16835 11215 17035 11241
rect 16613 11211 17035 11215
tri 17035 11211 17065 11241 sw
tri 17133 11211 17163 11241 ne
rect 17163 11215 17265 11241
rect 17385 11241 17487 11335
tri 17487 11241 17585 11339 sw
tri 17585 11241 17683 11339 ne
rect 17683 11335 18037 11339
rect 17683 11241 17815 11335
rect 17385 11215 17585 11241
rect 17163 11211 17585 11215
tri 17585 11211 17615 11241 sw
tri 17683 11211 17713 11241 ne
rect 17713 11215 17815 11241
rect 17935 11241 18037 11335
tri 18037 11241 18135 11339 sw
tri 18135 11241 18233 11339 ne
rect 18233 11335 18587 11339
rect 18233 11241 18365 11335
rect 17935 11215 18135 11241
rect 17713 11211 18135 11215
tri 18135 11211 18165 11241 sw
tri 18233 11211 18263 11241 ne
rect 18263 11215 18365 11241
rect 18485 11241 18587 11335
tri 18587 11241 18685 11339 sw
tri 18685 11241 18783 11339 ne
rect 18783 11335 19137 11339
rect 18783 11241 18915 11335
rect 18485 11215 18685 11241
rect 18263 11211 18685 11215
tri 18685 11211 18715 11241 sw
tri 18783 11211 18813 11241 ne
rect 18813 11215 18915 11241
rect 19035 11241 19137 11335
tri 19137 11241 19235 11339 sw
tri 19235 11241 19333 11339 ne
rect 19333 11335 20300 11339
rect 19333 11241 19465 11335
rect 19035 11215 19235 11241
rect 18813 11211 19235 11215
tri 19235 11211 19265 11241 sw
tri 19333 11211 19363 11241 ne
rect 19363 11215 19465 11241
rect 19585 11215 20300 11335
rect 19363 11211 20300 11215
tri 113 11113 211 11211 ne
rect 211 11113 565 11211
tri 565 11113 663 11211 sw
tri 663 11113 761 11211 ne
rect 761 11113 1115 11211
tri 1115 11113 1213 11211 sw
tri 1213 11113 1311 11211 ne
rect 1311 11113 1665 11211
tri 1665 11113 1763 11211 sw
tri 1763 11113 1861 11211 ne
rect 1861 11113 2215 11211
tri 2215 11113 2313 11211 sw
tri 2313 11113 2411 11211 ne
rect 2411 11113 2765 11211
tri 2765 11113 2863 11211 sw
tri 2863 11113 2961 11211 ne
rect 2961 11113 3315 11211
tri 3315 11113 3413 11211 sw
tri 3413 11113 3511 11211 ne
rect 3511 11113 3865 11211
tri 3865 11113 3963 11211 sw
tri 3963 11113 4061 11211 ne
rect 4061 11113 4415 11211
tri 4415 11113 4513 11211 sw
tri 4513 11113 4611 11211 ne
rect 4611 11113 4965 11211
tri 4965 11113 5063 11211 sw
tri 5063 11113 5161 11211 ne
rect 5161 11113 5515 11211
tri 5515 11113 5613 11211 sw
tri 5613 11113 5711 11211 ne
rect 5711 11113 6065 11211
tri 6065 11113 6163 11211 sw
tri 6163 11113 6261 11211 ne
rect 6261 11113 6615 11211
tri 6615 11113 6713 11211 sw
tri 6713 11113 6811 11211 ne
rect 6811 11113 7165 11211
tri 7165 11113 7263 11211 sw
tri 7263 11113 7361 11211 ne
rect 7361 11113 7715 11211
tri 7715 11113 7813 11211 sw
tri 7813 11113 7911 11211 ne
rect 7911 11113 8265 11211
tri 8265 11113 8363 11211 sw
tri 8363 11113 8461 11211 ne
rect 8461 11113 8815 11211
tri 8815 11113 8913 11211 sw
tri 8913 11113 9011 11211 ne
rect 9011 11113 9365 11211
tri 9365 11113 9463 11211 sw
tri 9463 11113 9561 11211 ne
rect 9561 11113 9915 11211
tri 9915 11113 10013 11211 sw
tri 10013 11113 10111 11211 ne
rect 10111 11113 10465 11211
tri 10465 11113 10563 11211 sw
tri 10563 11113 10661 11211 ne
rect 10661 11113 11015 11211
tri 11015 11113 11113 11211 sw
tri 11113 11113 11211 11211 ne
rect 11211 11113 11565 11211
tri 11565 11113 11663 11211 sw
tri 11663 11113 11761 11211 ne
rect 11761 11113 12115 11211
tri 12115 11113 12213 11211 sw
tri 12213 11113 12311 11211 ne
rect 12311 11113 12665 11211
tri 12665 11113 12763 11211 sw
tri 12763 11113 12861 11211 ne
rect 12861 11113 13215 11211
tri 13215 11113 13313 11211 sw
tri 13313 11113 13411 11211 ne
rect 13411 11113 13765 11211
tri 13765 11113 13863 11211 sw
tri 13863 11113 13961 11211 ne
rect 13961 11113 14315 11211
tri 14315 11113 14413 11211 sw
tri 14413 11113 14511 11211 ne
rect 14511 11113 14865 11211
tri 14865 11113 14963 11211 sw
tri 14963 11113 15061 11211 ne
rect 15061 11113 15415 11211
tri 15415 11113 15513 11211 sw
tri 15513 11113 15611 11211 ne
rect 15611 11113 15965 11211
tri 15965 11113 16063 11211 sw
tri 16063 11113 16161 11211 ne
rect 16161 11113 16515 11211
tri 16515 11113 16613 11211 sw
tri 16613 11113 16711 11211 ne
rect 16711 11113 17065 11211
tri 17065 11113 17163 11211 sw
tri 17163 11113 17261 11211 ne
rect 17261 11113 17615 11211
tri 17615 11113 17713 11211 sw
tri 17713 11113 17811 11211 ne
rect 17811 11113 18165 11211
tri 18165 11113 18263 11211 sw
tri 18263 11113 18361 11211 ne
rect 18361 11113 18715 11211
tri 18715 11113 18813 11211 sw
tri 18813 11113 18911 11211 ne
rect 18911 11113 19265 11211
tri 19265 11113 19363 11211 sw
tri 19363 11113 19461 11211 ne
rect 19461 11113 20300 11211
rect -2000 11083 113 11113
tri 113 11083 143 11113 sw
tri 211 11083 241 11113 ne
rect 241 11083 663 11113
tri 663 11083 693 11113 sw
tri 761 11083 791 11113 ne
rect 791 11083 1213 11113
tri 1213 11083 1243 11113 sw
tri 1311 11083 1341 11113 ne
rect 1341 11083 1763 11113
tri 1763 11083 1793 11113 sw
tri 1861 11083 1891 11113 ne
rect 1891 11083 2313 11113
tri 2313 11083 2343 11113 sw
tri 2411 11083 2441 11113 ne
rect 2441 11083 2863 11113
tri 2863 11083 2893 11113 sw
tri 2961 11083 2991 11113 ne
rect 2991 11083 3413 11113
tri 3413 11083 3443 11113 sw
tri 3511 11083 3541 11113 ne
rect 3541 11083 3963 11113
tri 3963 11083 3993 11113 sw
tri 4061 11083 4091 11113 ne
rect 4091 11083 4513 11113
tri 4513 11083 4543 11113 sw
tri 4611 11083 4641 11113 ne
rect 4641 11083 5063 11113
tri 5063 11083 5093 11113 sw
tri 5161 11083 5191 11113 ne
rect 5191 11083 5613 11113
tri 5613 11083 5643 11113 sw
tri 5711 11083 5741 11113 ne
rect 5741 11083 6163 11113
tri 6163 11083 6193 11113 sw
tri 6261 11083 6291 11113 ne
rect 6291 11083 6713 11113
tri 6713 11083 6743 11113 sw
tri 6811 11083 6841 11113 ne
rect 6841 11083 7263 11113
tri 7263 11083 7293 11113 sw
tri 7361 11083 7391 11113 ne
rect 7391 11083 7813 11113
tri 7813 11083 7843 11113 sw
tri 7911 11083 7941 11113 ne
rect 7941 11083 8363 11113
tri 8363 11083 8393 11113 sw
tri 8461 11083 8491 11113 ne
rect 8491 11083 8913 11113
tri 8913 11083 8943 11113 sw
tri 9011 11083 9041 11113 ne
rect 9041 11083 9463 11113
tri 9463 11083 9493 11113 sw
tri 9561 11083 9591 11113 ne
rect 9591 11083 10013 11113
tri 10013 11083 10043 11113 sw
tri 10111 11083 10141 11113 ne
rect 10141 11083 10563 11113
tri 10563 11083 10593 11113 sw
tri 10661 11083 10691 11113 ne
rect 10691 11083 11113 11113
tri 11113 11083 11143 11113 sw
tri 11211 11083 11241 11113 ne
rect 11241 11083 11663 11113
tri 11663 11083 11693 11113 sw
tri 11761 11083 11791 11113 ne
rect 11791 11083 12213 11113
tri 12213 11083 12243 11113 sw
tri 12311 11083 12341 11113 ne
rect 12341 11083 12763 11113
tri 12763 11083 12793 11113 sw
tri 12861 11083 12891 11113 ne
rect 12891 11083 13313 11113
tri 13313 11083 13343 11113 sw
tri 13411 11083 13441 11113 ne
rect 13441 11083 13863 11113
tri 13863 11083 13893 11113 sw
tri 13961 11083 13991 11113 ne
rect 13991 11083 14413 11113
tri 14413 11083 14443 11113 sw
tri 14511 11083 14541 11113 ne
rect 14541 11083 14963 11113
tri 14963 11083 14993 11113 sw
tri 15061 11083 15091 11113 ne
rect 15091 11083 15513 11113
tri 15513 11083 15543 11113 sw
tri 15611 11083 15641 11113 ne
rect 15641 11083 16063 11113
tri 16063 11083 16093 11113 sw
tri 16161 11083 16191 11113 ne
rect 16191 11083 16613 11113
tri 16613 11083 16643 11113 sw
tri 16711 11083 16741 11113 ne
rect 16741 11083 17163 11113
tri 17163 11083 17193 11113 sw
tri 17261 11083 17291 11113 ne
rect 17291 11083 17713 11113
tri 17713 11083 17743 11113 sw
tri 17811 11083 17841 11113 ne
rect 17841 11083 18263 11113
tri 18263 11083 18293 11113 sw
tri 18361 11083 18391 11113 ne
rect 18391 11083 18813 11113
tri 18813 11083 18843 11113 sw
tri 18911 11083 18941 11113 ne
rect 18941 11083 19363 11113
tri 19363 11083 19393 11113 sw
tri 19461 11083 19491 11113 ne
rect 19491 11083 20300 11113
rect -2000 10985 143 11083
tri 143 10985 241 11083 sw
tri 241 10985 339 11083 ne
rect 339 10985 693 11083
tri 693 10985 791 11083 sw
tri 791 10985 889 11083 ne
rect 889 10985 1243 11083
tri 1243 10985 1341 11083 sw
tri 1341 10985 1439 11083 ne
rect 1439 10985 1793 11083
tri 1793 10985 1891 11083 sw
tri 1891 10985 1989 11083 ne
rect 1989 10985 2343 11083
tri 2343 10985 2441 11083 sw
tri 2441 10985 2539 11083 ne
rect 2539 10985 2893 11083
tri 2893 10985 2991 11083 sw
tri 2991 10985 3089 11083 ne
rect 3089 10985 3443 11083
tri 3443 10985 3541 11083 sw
tri 3541 10985 3639 11083 ne
rect 3639 10985 3993 11083
tri 3993 10985 4091 11083 sw
tri 4091 10985 4189 11083 ne
rect 4189 10985 4543 11083
tri 4543 10985 4641 11083 sw
tri 4641 10985 4739 11083 ne
rect 4739 10985 5093 11083
tri 5093 10985 5191 11083 sw
tri 5191 10985 5289 11083 ne
rect 5289 10985 5643 11083
tri 5643 10985 5741 11083 sw
tri 5741 10985 5839 11083 ne
rect 5839 10985 6193 11083
tri 6193 10985 6291 11083 sw
tri 6291 10985 6389 11083 ne
rect 6389 10985 6743 11083
tri 6743 10985 6841 11083 sw
tri 6841 10985 6939 11083 ne
rect 6939 10985 7293 11083
tri 7293 10985 7391 11083 sw
tri 7391 10985 7489 11083 ne
rect 7489 10985 7843 11083
tri 7843 10985 7941 11083 sw
tri 7941 10985 8039 11083 ne
rect 8039 10985 8393 11083
tri 8393 10985 8491 11083 sw
tri 8491 10985 8589 11083 ne
rect 8589 10985 8943 11083
tri 8943 10985 9041 11083 sw
tri 9041 10985 9139 11083 ne
rect 9139 10985 9493 11083
tri 9493 10985 9591 11083 sw
tri 9591 10985 9689 11083 ne
rect 9689 10985 10043 11083
tri 10043 10985 10141 11083 sw
tri 10141 10985 10239 11083 ne
rect 10239 10985 10593 11083
tri 10593 10985 10691 11083 sw
tri 10691 10985 10789 11083 ne
rect 10789 10985 11143 11083
tri 11143 10985 11241 11083 sw
tri 11241 10985 11339 11083 ne
rect 11339 10985 11693 11083
tri 11693 10985 11791 11083 sw
tri 11791 10985 11889 11083 ne
rect 11889 10985 12243 11083
tri 12243 10985 12341 11083 sw
tri 12341 10985 12439 11083 ne
rect 12439 10985 12793 11083
tri 12793 10985 12891 11083 sw
tri 12891 10985 12989 11083 ne
rect 12989 10985 13343 11083
tri 13343 10985 13441 11083 sw
tri 13441 10985 13539 11083 ne
rect 13539 10985 13893 11083
tri 13893 10985 13991 11083 sw
tri 13991 10985 14089 11083 ne
rect 14089 10985 14443 11083
tri 14443 10985 14541 11083 sw
tri 14541 10985 14639 11083 ne
rect 14639 10985 14993 11083
tri 14993 10985 15091 11083 sw
tri 15091 10985 15189 11083 ne
rect 15189 10985 15543 11083
tri 15543 10985 15641 11083 sw
tri 15641 10985 15739 11083 ne
rect 15739 10985 16093 11083
tri 16093 10985 16191 11083 sw
tri 16191 10985 16289 11083 ne
rect 16289 10985 16643 11083
tri 16643 10985 16741 11083 sw
tri 16741 10985 16839 11083 ne
rect 16839 10985 17193 11083
tri 17193 10985 17291 11083 sw
tri 17291 10985 17389 11083 ne
rect 17389 10985 17743 11083
tri 17743 10985 17841 11083 sw
tri 17841 10985 17939 11083 ne
rect 17939 10985 18293 11083
tri 18293 10985 18391 11083 sw
tri 18391 10985 18489 11083 ne
rect 18489 10985 18843 11083
tri 18843 10985 18941 11083 sw
tri 18941 10985 19039 11083 ne
rect 19039 10985 19393 11083
tri 19393 10985 19491 11083 sw
tri 19491 10985 19589 11083 ne
rect 19589 10985 20300 11083
rect -2000 10887 241 10985
tri 241 10887 339 10985 sw
tri 339 10887 437 10985 ne
rect 437 10887 791 10985
tri 791 10887 889 10985 sw
tri 889 10887 987 10985 ne
rect 987 10887 1341 10985
tri 1341 10887 1439 10985 sw
tri 1439 10887 1537 10985 ne
rect 1537 10887 1891 10985
tri 1891 10887 1989 10985 sw
tri 1989 10887 2087 10985 ne
rect 2087 10887 2441 10985
tri 2441 10887 2539 10985 sw
tri 2539 10887 2637 10985 ne
rect 2637 10887 2991 10985
tri 2991 10887 3089 10985 sw
tri 3089 10887 3187 10985 ne
rect 3187 10887 3541 10985
tri 3541 10887 3639 10985 sw
tri 3639 10887 3737 10985 ne
rect 3737 10887 4091 10985
tri 4091 10887 4189 10985 sw
tri 4189 10887 4287 10985 ne
rect 4287 10887 4641 10985
tri 4641 10887 4739 10985 sw
tri 4739 10887 4837 10985 ne
rect 4837 10887 5191 10985
tri 5191 10887 5289 10985 sw
tri 5289 10887 5387 10985 ne
rect 5387 10887 5741 10985
tri 5741 10887 5839 10985 sw
tri 5839 10887 5937 10985 ne
rect 5937 10887 6291 10985
tri 6291 10887 6389 10985 sw
tri 6389 10887 6487 10985 ne
rect 6487 10887 6841 10985
tri 6841 10887 6939 10985 sw
tri 6939 10887 7037 10985 ne
rect 7037 10887 7391 10985
tri 7391 10887 7489 10985 sw
tri 7489 10887 7587 10985 ne
rect 7587 10887 7941 10985
tri 7941 10887 8039 10985 sw
tri 8039 10887 8137 10985 ne
rect 8137 10887 8491 10985
tri 8491 10887 8589 10985 sw
tri 8589 10887 8687 10985 ne
rect 8687 10887 9041 10985
tri 9041 10887 9139 10985 sw
tri 9139 10887 9237 10985 ne
rect 9237 10887 9591 10985
tri 9591 10887 9689 10985 sw
tri 9689 10887 9787 10985 ne
rect 9787 10887 10141 10985
tri 10141 10887 10239 10985 sw
tri 10239 10887 10337 10985 ne
rect 10337 10887 10691 10985
tri 10691 10887 10789 10985 sw
tri 10789 10887 10887 10985 ne
rect 10887 10887 11241 10985
tri 11241 10887 11339 10985 sw
tri 11339 10887 11437 10985 ne
rect 11437 10887 11791 10985
tri 11791 10887 11889 10985 sw
tri 11889 10887 11987 10985 ne
rect 11987 10887 12341 10985
tri 12341 10887 12439 10985 sw
tri 12439 10887 12537 10985 ne
rect 12537 10887 12891 10985
tri 12891 10887 12989 10985 sw
tri 12989 10887 13087 10985 ne
rect 13087 10887 13441 10985
tri 13441 10887 13539 10985 sw
tri 13539 10887 13637 10985 ne
rect 13637 10887 13991 10985
tri 13991 10887 14089 10985 sw
tri 14089 10887 14187 10985 ne
rect 14187 10887 14541 10985
tri 14541 10887 14639 10985 sw
tri 14639 10887 14737 10985 ne
rect 14737 10887 15091 10985
tri 15091 10887 15189 10985 sw
tri 15189 10887 15287 10985 ne
rect 15287 10887 15641 10985
tri 15641 10887 15739 10985 sw
tri 15739 10887 15837 10985 ne
rect 15837 10887 16191 10985
tri 16191 10887 16289 10985 sw
tri 16289 10887 16387 10985 ne
rect 16387 10887 16741 10985
tri 16741 10887 16839 10985 sw
tri 16839 10887 16937 10985 ne
rect 16937 10887 17291 10985
tri 17291 10887 17389 10985 sw
tri 17389 10887 17487 10985 ne
rect 17487 10887 17841 10985
tri 17841 10887 17939 10985 sw
tri 17939 10887 18037 10985 ne
rect 18037 10887 18391 10985
tri 18391 10887 18489 10985 sw
tri 18489 10887 18587 10985 ne
rect 18587 10887 18941 10985
tri 18941 10887 19039 10985 sw
tri 19039 10887 19137 10985 ne
rect 19137 10887 19491 10985
tri 19491 10887 19589 10985 sw
tri 19589 10887 19687 10985 ne
rect 19687 10887 20300 10985
rect -2000 10789 339 10887
tri 339 10789 437 10887 sw
tri 437 10789 535 10887 ne
rect 535 10789 889 10887
tri 889 10789 987 10887 sw
tri 987 10789 1085 10887 ne
rect 1085 10789 1439 10887
tri 1439 10789 1537 10887 sw
tri 1537 10789 1635 10887 ne
rect 1635 10789 1989 10887
tri 1989 10789 2087 10887 sw
tri 2087 10789 2185 10887 ne
rect 2185 10789 2539 10887
tri 2539 10789 2637 10887 sw
tri 2637 10789 2735 10887 ne
rect 2735 10789 3089 10887
tri 3089 10789 3187 10887 sw
tri 3187 10789 3285 10887 ne
rect 3285 10789 3639 10887
tri 3639 10789 3737 10887 sw
tri 3737 10789 3835 10887 ne
rect 3835 10789 4189 10887
tri 4189 10789 4287 10887 sw
tri 4287 10789 4385 10887 ne
rect 4385 10789 4739 10887
tri 4739 10789 4837 10887 sw
tri 4837 10789 4935 10887 ne
rect 4935 10789 5289 10887
tri 5289 10789 5387 10887 sw
tri 5387 10789 5485 10887 ne
rect 5485 10789 5839 10887
tri 5839 10789 5937 10887 sw
tri 5937 10789 6035 10887 ne
rect 6035 10789 6389 10887
tri 6389 10789 6487 10887 sw
tri 6487 10789 6585 10887 ne
rect 6585 10789 6939 10887
tri 6939 10789 7037 10887 sw
tri 7037 10789 7135 10887 ne
rect 7135 10789 7489 10887
tri 7489 10789 7587 10887 sw
tri 7587 10789 7685 10887 ne
rect 7685 10789 8039 10887
tri 8039 10789 8137 10887 sw
tri 8137 10789 8235 10887 ne
rect 8235 10789 8589 10887
tri 8589 10789 8687 10887 sw
tri 8687 10789 8785 10887 ne
rect 8785 10789 9139 10887
tri 9139 10789 9237 10887 sw
tri 9237 10789 9335 10887 ne
rect 9335 10789 9689 10887
tri 9689 10789 9787 10887 sw
tri 9787 10789 9885 10887 ne
rect 9885 10789 10239 10887
tri 10239 10789 10337 10887 sw
tri 10337 10789 10435 10887 ne
rect 10435 10789 10789 10887
tri 10789 10789 10887 10887 sw
tri 10887 10789 10985 10887 ne
rect 10985 10789 11339 10887
tri 11339 10789 11437 10887 sw
tri 11437 10789 11535 10887 ne
rect 11535 10789 11889 10887
tri 11889 10789 11987 10887 sw
tri 11987 10789 12085 10887 ne
rect 12085 10789 12439 10887
tri 12439 10789 12537 10887 sw
tri 12537 10789 12635 10887 ne
rect 12635 10789 12989 10887
tri 12989 10789 13087 10887 sw
tri 13087 10789 13185 10887 ne
rect 13185 10789 13539 10887
tri 13539 10789 13637 10887 sw
tri 13637 10789 13735 10887 ne
rect 13735 10789 14089 10887
tri 14089 10789 14187 10887 sw
tri 14187 10789 14285 10887 ne
rect 14285 10789 14639 10887
tri 14639 10789 14737 10887 sw
tri 14737 10789 14835 10887 ne
rect 14835 10789 15189 10887
tri 15189 10789 15287 10887 sw
tri 15287 10789 15385 10887 ne
rect 15385 10789 15739 10887
tri 15739 10789 15837 10887 sw
tri 15837 10789 15935 10887 ne
rect 15935 10789 16289 10887
tri 16289 10789 16387 10887 sw
tri 16387 10789 16485 10887 ne
rect 16485 10789 16839 10887
tri 16839 10789 16937 10887 sw
tri 16937 10789 17035 10887 ne
rect 17035 10789 17389 10887
tri 17389 10789 17487 10887 sw
tri 17487 10789 17585 10887 ne
rect 17585 10789 17939 10887
tri 17939 10789 18037 10887 sw
tri 18037 10789 18135 10887 ne
rect 18135 10789 18489 10887
tri 18489 10789 18587 10887 sw
tri 18587 10789 18685 10887 ne
rect 18685 10789 19039 10887
tri 19039 10789 19137 10887 sw
tri 19137 10789 19235 10887 ne
rect 19235 10789 19589 10887
tri 19589 10789 19687 10887 sw
rect 20800 10789 21800 11437
rect -2000 10785 437 10789
rect -2000 10665 215 10785
rect 335 10691 437 10785
tri 437 10691 535 10789 sw
tri 535 10691 633 10789 ne
rect 633 10785 987 10789
rect 633 10691 765 10785
rect 335 10665 535 10691
rect -2000 10661 535 10665
rect -2000 10013 -1000 10661
tri 113 10563 211 10661 ne
rect 211 10613 535 10661
tri 535 10613 613 10691 sw
tri 633 10613 711 10691 ne
rect 711 10665 765 10691
rect 885 10691 987 10785
tri 987 10691 1085 10789 sw
tri 1085 10691 1183 10789 ne
rect 1183 10785 1537 10789
rect 1183 10691 1315 10785
rect 885 10665 1085 10691
rect 711 10613 1085 10665
tri 1085 10613 1163 10691 sw
tri 1183 10613 1261 10691 ne
rect 1261 10665 1315 10691
rect 1435 10691 1537 10785
tri 1537 10691 1635 10789 sw
tri 1635 10691 1733 10789 ne
rect 1733 10785 2087 10789
rect 1733 10691 1865 10785
rect 1435 10665 1635 10691
rect 1261 10613 1635 10665
tri 1635 10613 1713 10691 sw
tri 1733 10613 1811 10691 ne
rect 1811 10665 1865 10691
rect 1985 10691 2087 10785
tri 2087 10691 2185 10789 sw
tri 2185 10691 2283 10789 ne
rect 2283 10785 2637 10789
rect 2283 10691 2415 10785
rect 1985 10665 2185 10691
rect 1811 10613 2185 10665
tri 2185 10613 2263 10691 sw
tri 2283 10613 2361 10691 ne
rect 2361 10665 2415 10691
rect 2535 10691 2637 10785
tri 2637 10691 2735 10789 sw
tri 2735 10691 2833 10789 ne
rect 2833 10785 3187 10789
rect 2833 10691 2965 10785
rect 2535 10665 2735 10691
rect 2361 10613 2735 10665
tri 2735 10613 2813 10691 sw
tri 2833 10613 2911 10691 ne
rect 2911 10665 2965 10691
rect 3085 10691 3187 10785
tri 3187 10691 3285 10789 sw
tri 3285 10691 3383 10789 ne
rect 3383 10785 3737 10789
rect 3383 10691 3515 10785
rect 3085 10665 3285 10691
rect 2911 10613 3285 10665
tri 3285 10613 3363 10691 sw
tri 3383 10613 3461 10691 ne
rect 3461 10665 3515 10691
rect 3635 10691 3737 10785
tri 3737 10691 3835 10789 sw
tri 3835 10691 3933 10789 ne
rect 3933 10785 4287 10789
rect 3933 10691 4065 10785
rect 3635 10665 3835 10691
rect 3461 10613 3835 10665
tri 3835 10613 3913 10691 sw
tri 3933 10613 4011 10691 ne
rect 4011 10665 4065 10691
rect 4185 10691 4287 10785
tri 4287 10691 4385 10789 sw
tri 4385 10691 4483 10789 ne
rect 4483 10785 4837 10789
rect 4483 10691 4615 10785
rect 4185 10665 4385 10691
rect 4011 10613 4385 10665
tri 4385 10613 4463 10691 sw
tri 4483 10613 4561 10691 ne
rect 4561 10665 4615 10691
rect 4735 10691 4837 10785
tri 4837 10691 4935 10789 sw
tri 4935 10691 5033 10789 ne
rect 5033 10785 5387 10789
rect 5033 10691 5165 10785
rect 4735 10665 4935 10691
rect 4561 10613 4935 10665
tri 4935 10613 5013 10691 sw
tri 5033 10613 5111 10691 ne
rect 5111 10665 5165 10691
rect 5285 10691 5387 10785
tri 5387 10691 5485 10789 sw
tri 5485 10691 5583 10789 ne
rect 5583 10785 5937 10789
rect 5583 10691 5715 10785
rect 5285 10665 5485 10691
rect 5111 10613 5485 10665
tri 5485 10613 5563 10691 sw
tri 5583 10613 5661 10691 ne
rect 5661 10665 5715 10691
rect 5835 10691 5937 10785
tri 5937 10691 6035 10789 sw
tri 6035 10691 6133 10789 ne
rect 6133 10785 6487 10789
rect 6133 10691 6265 10785
rect 5835 10665 6035 10691
rect 5661 10613 6035 10665
tri 6035 10613 6113 10691 sw
tri 6133 10613 6211 10691 ne
rect 6211 10665 6265 10691
rect 6385 10691 6487 10785
tri 6487 10691 6585 10789 sw
tri 6585 10691 6683 10789 ne
rect 6683 10785 7037 10789
rect 6683 10691 6815 10785
rect 6385 10665 6585 10691
rect 6211 10613 6585 10665
tri 6585 10613 6663 10691 sw
tri 6683 10613 6761 10691 ne
rect 6761 10665 6815 10691
rect 6935 10691 7037 10785
tri 7037 10691 7135 10789 sw
tri 7135 10691 7233 10789 ne
rect 7233 10785 7587 10789
rect 7233 10691 7365 10785
rect 6935 10665 7135 10691
rect 6761 10613 7135 10665
tri 7135 10613 7213 10691 sw
tri 7233 10613 7311 10691 ne
rect 7311 10665 7365 10691
rect 7485 10691 7587 10785
tri 7587 10691 7685 10789 sw
tri 7685 10691 7783 10789 ne
rect 7783 10785 8137 10789
rect 7783 10691 7915 10785
rect 7485 10665 7685 10691
rect 7311 10613 7685 10665
tri 7685 10613 7763 10691 sw
tri 7783 10613 7861 10691 ne
rect 7861 10665 7915 10691
rect 8035 10691 8137 10785
tri 8137 10691 8235 10789 sw
tri 8235 10691 8333 10789 ne
rect 8333 10785 8687 10789
rect 8333 10691 8465 10785
rect 8035 10665 8235 10691
rect 7861 10613 8235 10665
tri 8235 10613 8313 10691 sw
tri 8333 10613 8411 10691 ne
rect 8411 10665 8465 10691
rect 8585 10691 8687 10785
tri 8687 10691 8785 10789 sw
tri 8785 10691 8883 10789 ne
rect 8883 10785 9237 10789
rect 8883 10691 9015 10785
rect 8585 10665 8785 10691
rect 8411 10613 8785 10665
tri 8785 10613 8863 10691 sw
tri 8883 10613 8961 10691 ne
rect 8961 10665 9015 10691
rect 9135 10691 9237 10785
tri 9237 10691 9335 10789 sw
tri 9335 10691 9433 10789 ne
rect 9433 10785 9787 10789
rect 9433 10691 9565 10785
rect 9135 10665 9335 10691
rect 8961 10613 9335 10665
tri 9335 10613 9413 10691 sw
tri 9433 10613 9511 10691 ne
rect 9511 10665 9565 10691
rect 9685 10691 9787 10785
tri 9787 10691 9885 10789 sw
tri 9885 10691 9983 10789 ne
rect 9983 10785 10337 10789
rect 9983 10691 10115 10785
rect 9685 10665 9885 10691
rect 9511 10613 9885 10665
tri 9885 10613 9963 10691 sw
tri 9983 10613 10061 10691 ne
rect 10061 10665 10115 10691
rect 10235 10691 10337 10785
tri 10337 10691 10435 10789 sw
tri 10435 10691 10533 10789 ne
rect 10533 10785 10887 10789
rect 10533 10691 10665 10785
rect 10235 10665 10435 10691
rect 10061 10613 10435 10665
tri 10435 10613 10513 10691 sw
tri 10533 10613 10611 10691 ne
rect 10611 10665 10665 10691
rect 10785 10691 10887 10785
tri 10887 10691 10985 10789 sw
tri 10985 10691 11083 10789 ne
rect 11083 10785 11437 10789
rect 11083 10691 11215 10785
rect 10785 10665 10985 10691
rect 10611 10613 10985 10665
tri 10985 10613 11063 10691 sw
tri 11083 10613 11161 10691 ne
rect 11161 10665 11215 10691
rect 11335 10691 11437 10785
tri 11437 10691 11535 10789 sw
tri 11535 10691 11633 10789 ne
rect 11633 10785 11987 10789
rect 11633 10691 11765 10785
rect 11335 10665 11535 10691
rect 11161 10613 11535 10665
tri 11535 10613 11613 10691 sw
tri 11633 10613 11711 10691 ne
rect 11711 10665 11765 10691
rect 11885 10691 11987 10785
tri 11987 10691 12085 10789 sw
tri 12085 10691 12183 10789 ne
rect 12183 10785 12537 10789
rect 12183 10691 12315 10785
rect 11885 10665 12085 10691
rect 11711 10613 12085 10665
tri 12085 10613 12163 10691 sw
tri 12183 10613 12261 10691 ne
rect 12261 10665 12315 10691
rect 12435 10691 12537 10785
tri 12537 10691 12635 10789 sw
tri 12635 10691 12733 10789 ne
rect 12733 10785 13087 10789
rect 12733 10691 12865 10785
rect 12435 10665 12635 10691
rect 12261 10613 12635 10665
tri 12635 10613 12713 10691 sw
tri 12733 10613 12811 10691 ne
rect 12811 10665 12865 10691
rect 12985 10691 13087 10785
tri 13087 10691 13185 10789 sw
tri 13185 10691 13283 10789 ne
rect 13283 10785 13637 10789
rect 13283 10691 13415 10785
rect 12985 10665 13185 10691
rect 12811 10613 13185 10665
tri 13185 10613 13263 10691 sw
tri 13283 10613 13361 10691 ne
rect 13361 10665 13415 10691
rect 13535 10691 13637 10785
tri 13637 10691 13735 10789 sw
tri 13735 10691 13833 10789 ne
rect 13833 10785 14187 10789
rect 13833 10691 13965 10785
rect 13535 10665 13735 10691
rect 13361 10613 13735 10665
tri 13735 10613 13813 10691 sw
tri 13833 10613 13911 10691 ne
rect 13911 10665 13965 10691
rect 14085 10691 14187 10785
tri 14187 10691 14285 10789 sw
tri 14285 10691 14383 10789 ne
rect 14383 10785 14737 10789
rect 14383 10691 14515 10785
rect 14085 10665 14285 10691
rect 13911 10613 14285 10665
tri 14285 10613 14363 10691 sw
tri 14383 10613 14461 10691 ne
rect 14461 10665 14515 10691
rect 14635 10691 14737 10785
tri 14737 10691 14835 10789 sw
tri 14835 10691 14933 10789 ne
rect 14933 10785 15287 10789
rect 14933 10691 15065 10785
rect 14635 10665 14835 10691
rect 14461 10613 14835 10665
tri 14835 10613 14913 10691 sw
tri 14933 10613 15011 10691 ne
rect 15011 10665 15065 10691
rect 15185 10691 15287 10785
tri 15287 10691 15385 10789 sw
tri 15385 10691 15483 10789 ne
rect 15483 10785 15837 10789
rect 15483 10691 15615 10785
rect 15185 10665 15385 10691
rect 15011 10613 15385 10665
tri 15385 10613 15463 10691 sw
tri 15483 10613 15561 10691 ne
rect 15561 10665 15615 10691
rect 15735 10691 15837 10785
tri 15837 10691 15935 10789 sw
tri 15935 10691 16033 10789 ne
rect 16033 10785 16387 10789
rect 16033 10691 16165 10785
rect 15735 10665 15935 10691
rect 15561 10613 15935 10665
tri 15935 10613 16013 10691 sw
tri 16033 10613 16111 10691 ne
rect 16111 10665 16165 10691
rect 16285 10691 16387 10785
tri 16387 10691 16485 10789 sw
tri 16485 10691 16583 10789 ne
rect 16583 10785 16937 10789
rect 16583 10691 16715 10785
rect 16285 10665 16485 10691
rect 16111 10613 16485 10665
tri 16485 10613 16563 10691 sw
tri 16583 10613 16661 10691 ne
rect 16661 10665 16715 10691
rect 16835 10691 16937 10785
tri 16937 10691 17035 10789 sw
tri 17035 10691 17133 10789 ne
rect 17133 10785 17487 10789
rect 17133 10691 17265 10785
rect 16835 10665 17035 10691
rect 16661 10613 17035 10665
tri 17035 10613 17113 10691 sw
tri 17133 10613 17211 10691 ne
rect 17211 10665 17265 10691
rect 17385 10691 17487 10785
tri 17487 10691 17585 10789 sw
tri 17585 10691 17683 10789 ne
rect 17683 10785 18037 10789
rect 17683 10691 17815 10785
rect 17385 10665 17585 10691
rect 17211 10613 17585 10665
tri 17585 10613 17663 10691 sw
tri 17683 10613 17761 10691 ne
rect 17761 10665 17815 10691
rect 17935 10691 18037 10785
tri 18037 10691 18135 10789 sw
tri 18135 10691 18233 10789 ne
rect 18233 10785 18587 10789
rect 18233 10691 18365 10785
rect 17935 10665 18135 10691
rect 17761 10613 18135 10665
tri 18135 10613 18213 10691 sw
tri 18233 10613 18311 10691 ne
rect 18311 10665 18365 10691
rect 18485 10691 18587 10785
tri 18587 10691 18685 10789 sw
tri 18685 10691 18783 10789 ne
rect 18783 10785 19137 10789
rect 18783 10691 18915 10785
rect 18485 10665 18685 10691
rect 18311 10613 18685 10665
tri 18685 10613 18763 10691 sw
tri 18783 10613 18861 10691 ne
rect 18861 10665 18915 10691
rect 19035 10691 19137 10785
tri 19137 10691 19235 10789 sw
tri 19235 10691 19333 10789 ne
rect 19333 10785 21800 10789
rect 19333 10691 19465 10785
rect 19035 10665 19235 10691
rect 18861 10613 19235 10665
tri 19235 10613 19313 10691 sw
tri 19333 10613 19411 10691 ne
rect 19411 10665 19465 10691
rect 19585 10665 21800 10785
rect 19411 10613 21800 10665
rect 211 10563 613 10613
rect -500 10513 113 10563
tri 113 10513 163 10563 sw
tri 211 10513 261 10563 ne
rect 261 10533 613 10563
tri 613 10533 693 10613 sw
tri 711 10533 791 10613 ne
rect 791 10533 1163 10613
tri 1163 10533 1243 10613 sw
tri 1261 10533 1341 10613 ne
rect 1341 10533 1713 10613
tri 1713 10533 1793 10613 sw
tri 1811 10533 1891 10613 ne
rect 1891 10533 2263 10613
tri 2263 10533 2343 10613 sw
tri 2361 10533 2441 10613 ne
rect 2441 10533 2813 10613
tri 2813 10533 2893 10613 sw
tri 2911 10533 2991 10613 ne
rect 2991 10533 3363 10613
tri 3363 10533 3443 10613 sw
tri 3461 10533 3541 10613 ne
rect 3541 10533 3913 10613
tri 3913 10533 3993 10613 sw
tri 4011 10533 4091 10613 ne
rect 4091 10533 4463 10613
tri 4463 10533 4543 10613 sw
tri 4561 10533 4641 10613 ne
rect 4641 10533 5013 10613
tri 5013 10533 5093 10613 sw
tri 5111 10533 5191 10613 ne
rect 5191 10533 5563 10613
tri 5563 10533 5643 10613 sw
tri 5661 10533 5741 10613 ne
rect 5741 10533 6113 10613
tri 6113 10533 6193 10613 sw
tri 6211 10533 6291 10613 ne
rect 6291 10533 6663 10613
tri 6663 10533 6743 10613 sw
tri 6761 10533 6841 10613 ne
rect 6841 10533 7213 10613
tri 7213 10533 7293 10613 sw
tri 7311 10533 7391 10613 ne
rect 7391 10533 7763 10613
tri 7763 10533 7843 10613 sw
tri 7861 10533 7941 10613 ne
rect 7941 10533 8313 10613
tri 8313 10533 8393 10613 sw
tri 8411 10533 8491 10613 ne
rect 8491 10533 8863 10613
tri 8863 10533 8943 10613 sw
tri 8961 10533 9041 10613 ne
rect 9041 10533 9413 10613
tri 9413 10533 9493 10613 sw
tri 9511 10533 9591 10613 ne
rect 9591 10533 9963 10613
tri 9963 10533 10043 10613 sw
tri 10061 10533 10141 10613 ne
rect 10141 10533 10513 10613
tri 10513 10533 10593 10613 sw
tri 10611 10533 10691 10613 ne
rect 10691 10533 11063 10613
tri 11063 10533 11143 10613 sw
tri 11161 10533 11241 10613 ne
rect 11241 10533 11613 10613
tri 11613 10533 11693 10613 sw
tri 11711 10533 11791 10613 ne
rect 11791 10533 12163 10613
tri 12163 10533 12243 10613 sw
tri 12261 10533 12341 10613 ne
rect 12341 10533 12713 10613
tri 12713 10533 12793 10613 sw
tri 12811 10533 12891 10613 ne
rect 12891 10533 13263 10613
tri 13263 10533 13343 10613 sw
tri 13361 10533 13441 10613 ne
rect 13441 10533 13813 10613
tri 13813 10533 13893 10613 sw
tri 13911 10533 13991 10613 ne
rect 13991 10533 14363 10613
tri 14363 10533 14443 10613 sw
tri 14461 10533 14541 10613 ne
rect 14541 10533 14913 10613
tri 14913 10533 14993 10613 sw
tri 15011 10533 15091 10613 ne
rect 15091 10533 15463 10613
tri 15463 10533 15543 10613 sw
tri 15561 10533 15641 10613 ne
rect 15641 10533 16013 10613
tri 16013 10533 16093 10613 sw
tri 16111 10533 16191 10613 ne
rect 16191 10533 16563 10613
tri 16563 10533 16643 10613 sw
tri 16661 10533 16741 10613 ne
rect 16741 10533 17113 10613
tri 17113 10533 17193 10613 sw
tri 17211 10533 17291 10613 ne
rect 17291 10533 17663 10613
tri 17663 10533 17743 10613 sw
tri 17761 10533 17841 10613 ne
rect 17841 10533 18213 10613
tri 18213 10533 18293 10613 sw
tri 18311 10533 18391 10613 ne
rect 18391 10533 18763 10613
tri 18763 10533 18843 10613 sw
tri 18861 10533 18941 10613 ne
rect 18941 10533 19313 10613
tri 19313 10533 19393 10613 sw
tri 19411 10533 19491 10613 ne
rect 19491 10533 20100 10613
rect 261 10513 693 10533
rect -500 10435 163 10513
tri 163 10435 241 10513 sw
tri 261 10435 339 10513 ne
rect 339 10435 693 10513
tri 693 10435 791 10533 sw
tri 791 10435 889 10533 ne
rect 889 10435 1243 10533
tri 1243 10435 1341 10533 sw
tri 1341 10435 1439 10533 ne
rect 1439 10435 1793 10533
tri 1793 10435 1891 10533 sw
tri 1891 10435 1989 10533 ne
rect 1989 10435 2343 10533
tri 2343 10435 2441 10533 sw
tri 2441 10435 2539 10533 ne
rect 2539 10435 2893 10533
tri 2893 10435 2991 10533 sw
tri 2991 10435 3089 10533 ne
rect 3089 10435 3443 10533
tri 3443 10435 3541 10533 sw
tri 3541 10435 3639 10533 ne
rect 3639 10435 3993 10533
tri 3993 10435 4091 10533 sw
tri 4091 10435 4189 10533 ne
rect 4189 10435 4543 10533
tri 4543 10435 4641 10533 sw
tri 4641 10435 4739 10533 ne
rect 4739 10435 5093 10533
tri 5093 10435 5191 10533 sw
tri 5191 10435 5289 10533 ne
rect 5289 10435 5643 10533
tri 5643 10435 5741 10533 sw
tri 5741 10435 5839 10533 ne
rect 5839 10435 6193 10533
tri 6193 10435 6291 10533 sw
tri 6291 10435 6389 10533 ne
rect 6389 10435 6743 10533
tri 6743 10435 6841 10533 sw
tri 6841 10435 6939 10533 ne
rect 6939 10435 7293 10533
tri 7293 10435 7391 10533 sw
tri 7391 10435 7489 10533 ne
rect 7489 10435 7843 10533
tri 7843 10435 7941 10533 sw
tri 7941 10435 8039 10533 ne
rect 8039 10435 8393 10533
tri 8393 10435 8491 10533 sw
tri 8491 10435 8589 10533 ne
rect 8589 10435 8943 10533
tri 8943 10435 9041 10533 sw
tri 9041 10435 9139 10533 ne
rect 9139 10435 9493 10533
tri 9493 10435 9591 10533 sw
tri 9591 10435 9689 10533 ne
rect 9689 10435 10043 10533
tri 10043 10435 10141 10533 sw
tri 10141 10435 10239 10533 ne
rect 10239 10435 10593 10533
tri 10593 10435 10691 10533 sw
tri 10691 10435 10789 10533 ne
rect 10789 10435 11143 10533
tri 11143 10435 11241 10533 sw
tri 11241 10435 11339 10533 ne
rect 11339 10435 11693 10533
tri 11693 10435 11791 10533 sw
tri 11791 10435 11889 10533 ne
rect 11889 10435 12243 10533
tri 12243 10435 12341 10533 sw
tri 12341 10435 12439 10533 ne
rect 12439 10435 12793 10533
tri 12793 10435 12891 10533 sw
tri 12891 10435 12989 10533 ne
rect 12989 10435 13343 10533
tri 13343 10435 13441 10533 sw
tri 13441 10435 13539 10533 ne
rect 13539 10435 13893 10533
tri 13893 10435 13991 10533 sw
tri 13991 10435 14089 10533 ne
rect 14089 10435 14443 10533
tri 14443 10435 14541 10533 sw
tri 14541 10435 14639 10533 ne
rect 14639 10435 14993 10533
tri 14993 10435 15091 10533 sw
tri 15091 10435 15189 10533 ne
rect 15189 10435 15543 10533
tri 15543 10435 15641 10533 sw
tri 15641 10435 15739 10533 ne
rect 15739 10435 16093 10533
tri 16093 10435 16191 10533 sw
tri 16191 10435 16289 10533 ne
rect 16289 10435 16643 10533
tri 16643 10435 16741 10533 sw
tri 16741 10435 16839 10533 ne
rect 16839 10435 17193 10533
tri 17193 10435 17291 10533 sw
tri 17291 10435 17389 10533 ne
rect 17389 10435 17743 10533
tri 17743 10435 17841 10533 sw
tri 17841 10435 17939 10533 ne
rect 17939 10435 18293 10533
tri 18293 10435 18391 10533 sw
tri 18391 10435 18489 10533 ne
rect 18489 10435 18843 10533
tri 18843 10435 18941 10533 sw
tri 18941 10435 19039 10533 ne
rect 19039 10435 19393 10533
tri 19393 10435 19491 10533 sw
tri 19491 10435 19589 10533 ne
rect 19589 10513 20100 10533
rect 20200 10513 21800 10613
rect 19589 10435 21800 10513
rect -500 10387 241 10435
rect -500 10287 -400 10387
rect -300 10337 241 10387
tri 241 10337 339 10435 sw
tri 339 10337 437 10435 ne
rect 437 10337 791 10435
tri 791 10337 889 10435 sw
tri 889 10337 987 10435 ne
rect 987 10337 1341 10435
tri 1341 10337 1439 10435 sw
tri 1439 10337 1537 10435 ne
rect 1537 10337 1891 10435
tri 1891 10337 1989 10435 sw
tri 1989 10337 2087 10435 ne
rect 2087 10337 2441 10435
tri 2441 10337 2539 10435 sw
tri 2539 10337 2637 10435 ne
rect 2637 10337 2991 10435
tri 2991 10337 3089 10435 sw
tri 3089 10337 3187 10435 ne
rect 3187 10337 3541 10435
tri 3541 10337 3639 10435 sw
tri 3639 10337 3737 10435 ne
rect 3737 10337 4091 10435
tri 4091 10337 4189 10435 sw
tri 4189 10337 4287 10435 ne
rect 4287 10337 4641 10435
tri 4641 10337 4739 10435 sw
tri 4739 10337 4837 10435 ne
rect 4837 10337 5191 10435
tri 5191 10337 5289 10435 sw
tri 5289 10337 5387 10435 ne
rect 5387 10337 5741 10435
tri 5741 10337 5839 10435 sw
tri 5839 10337 5937 10435 ne
rect 5937 10337 6291 10435
tri 6291 10337 6389 10435 sw
tri 6389 10337 6487 10435 ne
rect 6487 10337 6841 10435
tri 6841 10337 6939 10435 sw
tri 6939 10337 7037 10435 ne
rect 7037 10337 7391 10435
tri 7391 10337 7489 10435 sw
tri 7489 10337 7587 10435 ne
rect 7587 10337 7941 10435
tri 7941 10337 8039 10435 sw
tri 8039 10337 8137 10435 ne
rect 8137 10337 8491 10435
tri 8491 10337 8589 10435 sw
tri 8589 10337 8687 10435 ne
rect 8687 10337 9041 10435
tri 9041 10337 9139 10435 sw
tri 9139 10337 9237 10435 ne
rect 9237 10337 9591 10435
tri 9591 10337 9689 10435 sw
tri 9689 10337 9787 10435 ne
rect 9787 10337 10141 10435
tri 10141 10337 10239 10435 sw
tri 10239 10337 10337 10435 ne
rect 10337 10337 10691 10435
tri 10691 10337 10789 10435 sw
tri 10789 10337 10887 10435 ne
rect 10887 10337 11241 10435
tri 11241 10337 11339 10435 sw
tri 11339 10337 11437 10435 ne
rect 11437 10337 11791 10435
tri 11791 10337 11889 10435 sw
tri 11889 10337 11987 10435 ne
rect 11987 10337 12341 10435
tri 12341 10337 12439 10435 sw
tri 12439 10337 12537 10435 ne
rect 12537 10337 12891 10435
tri 12891 10337 12989 10435 sw
tri 12989 10337 13087 10435 ne
rect 13087 10337 13441 10435
tri 13441 10337 13539 10435 sw
tri 13539 10337 13637 10435 ne
rect 13637 10337 13991 10435
tri 13991 10337 14089 10435 sw
tri 14089 10337 14187 10435 ne
rect 14187 10337 14541 10435
tri 14541 10337 14639 10435 sw
tri 14639 10337 14737 10435 ne
rect 14737 10337 15091 10435
tri 15091 10337 15189 10435 sw
tri 15189 10337 15287 10435 ne
rect 15287 10337 15641 10435
tri 15641 10337 15739 10435 sw
tri 15739 10337 15837 10435 ne
rect 15837 10337 16191 10435
tri 16191 10337 16289 10435 sw
tri 16289 10337 16387 10435 ne
rect 16387 10337 16741 10435
tri 16741 10337 16839 10435 sw
tri 16839 10337 16937 10435 ne
rect 16937 10337 17291 10435
tri 17291 10337 17389 10435 sw
tri 17389 10337 17487 10435 ne
rect 17487 10337 17841 10435
tri 17841 10337 17939 10435 sw
tri 17939 10337 18037 10435 ne
rect 18037 10337 18391 10435
tri 18391 10337 18489 10435 sw
tri 18489 10337 18587 10435 ne
rect 18587 10337 18941 10435
tri 18941 10337 19039 10435 sw
tri 19039 10337 19137 10435 ne
rect 19137 10337 19491 10435
tri 19491 10337 19589 10435 sw
tri 19589 10337 19687 10435 ne
rect 19687 10337 21800 10435
rect -300 10287 339 10337
rect -500 10239 339 10287
tri 339 10239 437 10337 sw
tri 437 10239 535 10337 ne
rect 535 10239 889 10337
tri 889 10239 987 10337 sw
tri 987 10239 1085 10337 ne
rect 1085 10239 1439 10337
tri 1439 10239 1537 10337 sw
tri 1537 10239 1635 10337 ne
rect 1635 10239 1989 10337
tri 1989 10239 2087 10337 sw
tri 2087 10239 2185 10337 ne
rect 2185 10239 2539 10337
tri 2539 10239 2637 10337 sw
tri 2637 10239 2735 10337 ne
rect 2735 10239 3089 10337
tri 3089 10239 3187 10337 sw
tri 3187 10239 3285 10337 ne
rect 3285 10239 3639 10337
tri 3639 10239 3737 10337 sw
tri 3737 10239 3835 10337 ne
rect 3835 10239 4189 10337
tri 4189 10239 4287 10337 sw
tri 4287 10239 4385 10337 ne
rect 4385 10239 4739 10337
tri 4739 10239 4837 10337 sw
tri 4837 10239 4935 10337 ne
rect 4935 10239 5289 10337
tri 5289 10239 5387 10337 sw
tri 5387 10239 5485 10337 ne
rect 5485 10239 5839 10337
tri 5839 10239 5937 10337 sw
tri 5937 10239 6035 10337 ne
rect 6035 10239 6389 10337
tri 6389 10239 6487 10337 sw
tri 6487 10239 6585 10337 ne
rect 6585 10239 6939 10337
tri 6939 10239 7037 10337 sw
tri 7037 10239 7135 10337 ne
rect 7135 10239 7489 10337
tri 7489 10239 7587 10337 sw
tri 7587 10239 7685 10337 ne
rect 7685 10239 8039 10337
tri 8039 10239 8137 10337 sw
tri 8137 10239 8235 10337 ne
rect 8235 10239 8589 10337
tri 8589 10239 8687 10337 sw
tri 8687 10239 8785 10337 ne
rect 8785 10239 9139 10337
tri 9139 10239 9237 10337 sw
tri 9237 10239 9335 10337 ne
rect 9335 10239 9689 10337
tri 9689 10239 9787 10337 sw
tri 9787 10239 9885 10337 ne
rect 9885 10239 10239 10337
tri 10239 10239 10337 10337 sw
tri 10337 10239 10435 10337 ne
rect 10435 10239 10789 10337
tri 10789 10239 10887 10337 sw
tri 10887 10239 10985 10337 ne
rect 10985 10239 11339 10337
tri 11339 10239 11437 10337 sw
tri 11437 10239 11535 10337 ne
rect 11535 10239 11889 10337
tri 11889 10239 11987 10337 sw
tri 11987 10239 12085 10337 ne
rect 12085 10239 12439 10337
tri 12439 10239 12537 10337 sw
tri 12537 10239 12635 10337 ne
rect 12635 10239 12989 10337
tri 12989 10239 13087 10337 sw
tri 13087 10239 13185 10337 ne
rect 13185 10239 13539 10337
tri 13539 10239 13637 10337 sw
tri 13637 10239 13735 10337 ne
rect 13735 10239 14089 10337
tri 14089 10239 14187 10337 sw
tri 14187 10239 14285 10337 ne
rect 14285 10239 14639 10337
tri 14639 10239 14737 10337 sw
tri 14737 10239 14835 10337 ne
rect 14835 10239 15189 10337
tri 15189 10239 15287 10337 sw
tri 15287 10239 15385 10337 ne
rect 15385 10239 15739 10337
tri 15739 10239 15837 10337 sw
tri 15837 10239 15935 10337 ne
rect 15935 10239 16289 10337
tri 16289 10239 16387 10337 sw
tri 16387 10239 16485 10337 ne
rect 16485 10239 16839 10337
tri 16839 10239 16937 10337 sw
tri 16937 10239 17035 10337 ne
rect 17035 10239 17389 10337
tri 17389 10239 17487 10337 sw
tri 17487 10239 17585 10337 ne
rect 17585 10239 17939 10337
tri 17939 10239 18037 10337 sw
tri 18037 10239 18135 10337 ne
rect 18135 10239 18489 10337
tri 18489 10239 18587 10337 sw
tri 18587 10239 18685 10337 ne
rect 18685 10239 19039 10337
tri 19039 10239 19137 10337 sw
tri 19137 10239 19235 10337 ne
rect 19235 10239 19589 10337
tri 19589 10239 19687 10337 sw
rect -500 10235 437 10239
rect -500 10115 215 10235
rect 335 10141 437 10235
tri 437 10141 535 10239 sw
tri 535 10141 633 10239 ne
rect 633 10235 987 10239
rect 633 10141 765 10235
rect 335 10115 535 10141
rect -500 10111 535 10115
tri 535 10111 565 10141 sw
tri 633 10111 663 10141 ne
rect 663 10115 765 10141
rect 885 10141 987 10235
tri 987 10141 1085 10239 sw
tri 1085 10141 1183 10239 ne
rect 1183 10235 1537 10239
rect 1183 10141 1315 10235
rect 885 10115 1085 10141
rect 663 10111 1085 10115
tri 1085 10111 1115 10141 sw
tri 1183 10111 1213 10141 ne
rect 1213 10115 1315 10141
rect 1435 10141 1537 10235
tri 1537 10141 1635 10239 sw
tri 1635 10141 1733 10239 ne
rect 1733 10235 2087 10239
rect 1733 10141 1865 10235
rect 1435 10115 1635 10141
rect 1213 10111 1635 10115
tri 1635 10111 1665 10141 sw
tri 1733 10111 1763 10141 ne
rect 1763 10115 1865 10141
rect 1985 10141 2087 10235
tri 2087 10141 2185 10239 sw
tri 2185 10141 2283 10239 ne
rect 2283 10235 2637 10239
rect 2283 10141 2415 10235
rect 1985 10115 2185 10141
rect 1763 10111 2185 10115
tri 2185 10111 2215 10141 sw
tri 2283 10111 2313 10141 ne
rect 2313 10115 2415 10141
rect 2535 10141 2637 10235
tri 2637 10141 2735 10239 sw
tri 2735 10141 2833 10239 ne
rect 2833 10235 3187 10239
rect 2833 10141 2965 10235
rect 2535 10115 2735 10141
rect 2313 10111 2735 10115
tri 2735 10111 2765 10141 sw
tri 2833 10111 2863 10141 ne
rect 2863 10115 2965 10141
rect 3085 10141 3187 10235
tri 3187 10141 3285 10239 sw
tri 3285 10141 3383 10239 ne
rect 3383 10235 3737 10239
rect 3383 10141 3515 10235
rect 3085 10115 3285 10141
rect 2863 10111 3285 10115
tri 3285 10111 3315 10141 sw
tri 3383 10111 3413 10141 ne
rect 3413 10115 3515 10141
rect 3635 10141 3737 10235
tri 3737 10141 3835 10239 sw
tri 3835 10141 3933 10239 ne
rect 3933 10235 4287 10239
rect 3933 10141 4065 10235
rect 3635 10115 3835 10141
rect 3413 10111 3835 10115
tri 3835 10111 3865 10141 sw
tri 3933 10111 3963 10141 ne
rect 3963 10115 4065 10141
rect 4185 10141 4287 10235
tri 4287 10141 4385 10239 sw
tri 4385 10141 4483 10239 ne
rect 4483 10235 4837 10239
rect 4483 10141 4615 10235
rect 4185 10115 4385 10141
rect 3963 10111 4385 10115
tri 4385 10111 4415 10141 sw
tri 4483 10111 4513 10141 ne
rect 4513 10115 4615 10141
rect 4735 10141 4837 10235
tri 4837 10141 4935 10239 sw
tri 4935 10141 5033 10239 ne
rect 5033 10235 5387 10239
rect 5033 10141 5165 10235
rect 4735 10115 4935 10141
rect 4513 10111 4935 10115
tri 4935 10111 4965 10141 sw
tri 5033 10111 5063 10141 ne
rect 5063 10115 5165 10141
rect 5285 10141 5387 10235
tri 5387 10141 5485 10239 sw
tri 5485 10141 5583 10239 ne
rect 5583 10235 5937 10239
rect 5583 10141 5715 10235
rect 5285 10115 5485 10141
rect 5063 10111 5485 10115
tri 5485 10111 5515 10141 sw
tri 5583 10111 5613 10141 ne
rect 5613 10115 5715 10141
rect 5835 10141 5937 10235
tri 5937 10141 6035 10239 sw
tri 6035 10141 6133 10239 ne
rect 6133 10235 6487 10239
rect 6133 10141 6265 10235
rect 5835 10115 6035 10141
rect 5613 10111 6035 10115
tri 6035 10111 6065 10141 sw
tri 6133 10111 6163 10141 ne
rect 6163 10115 6265 10141
rect 6385 10141 6487 10235
tri 6487 10141 6585 10239 sw
tri 6585 10141 6683 10239 ne
rect 6683 10235 7037 10239
rect 6683 10141 6815 10235
rect 6385 10115 6585 10141
rect 6163 10111 6585 10115
tri 6585 10111 6615 10141 sw
tri 6683 10111 6713 10141 ne
rect 6713 10115 6815 10141
rect 6935 10141 7037 10235
tri 7037 10141 7135 10239 sw
tri 7135 10141 7233 10239 ne
rect 7233 10235 7587 10239
rect 7233 10141 7365 10235
rect 6935 10115 7135 10141
rect 6713 10111 7135 10115
tri 7135 10111 7165 10141 sw
tri 7233 10111 7263 10141 ne
rect 7263 10115 7365 10141
rect 7485 10141 7587 10235
tri 7587 10141 7685 10239 sw
tri 7685 10141 7783 10239 ne
rect 7783 10235 8137 10239
rect 7783 10141 7915 10235
rect 7485 10115 7685 10141
rect 7263 10111 7685 10115
tri 7685 10111 7715 10141 sw
tri 7783 10111 7813 10141 ne
rect 7813 10115 7915 10141
rect 8035 10141 8137 10235
tri 8137 10141 8235 10239 sw
tri 8235 10141 8333 10239 ne
rect 8333 10235 8687 10239
rect 8333 10141 8465 10235
rect 8035 10115 8235 10141
rect 7813 10111 8235 10115
tri 8235 10111 8265 10141 sw
tri 8333 10111 8363 10141 ne
rect 8363 10115 8465 10141
rect 8585 10141 8687 10235
tri 8687 10141 8785 10239 sw
tri 8785 10141 8883 10239 ne
rect 8883 10235 9237 10239
rect 8883 10141 9015 10235
rect 8585 10115 8785 10141
rect 8363 10111 8785 10115
tri 8785 10111 8815 10141 sw
tri 8883 10111 8913 10141 ne
rect 8913 10115 9015 10141
rect 9135 10141 9237 10235
tri 9237 10141 9335 10239 sw
tri 9335 10141 9433 10239 ne
rect 9433 10235 9787 10239
rect 9433 10141 9565 10235
rect 9135 10115 9335 10141
rect 8913 10111 9335 10115
tri 9335 10111 9365 10141 sw
tri 9433 10111 9463 10141 ne
rect 9463 10115 9565 10141
rect 9685 10141 9787 10235
tri 9787 10141 9885 10239 sw
tri 9885 10141 9983 10239 ne
rect 9983 10235 10337 10239
rect 9983 10141 10115 10235
rect 9685 10115 9885 10141
rect 9463 10111 9885 10115
tri 9885 10111 9915 10141 sw
tri 9983 10111 10013 10141 ne
rect 10013 10115 10115 10141
rect 10235 10141 10337 10235
tri 10337 10141 10435 10239 sw
tri 10435 10141 10533 10239 ne
rect 10533 10235 10887 10239
rect 10533 10141 10665 10235
rect 10235 10115 10435 10141
rect 10013 10111 10435 10115
tri 10435 10111 10465 10141 sw
tri 10533 10111 10563 10141 ne
rect 10563 10115 10665 10141
rect 10785 10141 10887 10235
tri 10887 10141 10985 10239 sw
tri 10985 10141 11083 10239 ne
rect 11083 10235 11437 10239
rect 11083 10141 11215 10235
rect 10785 10115 10985 10141
rect 10563 10111 10985 10115
tri 10985 10111 11015 10141 sw
tri 11083 10111 11113 10141 ne
rect 11113 10115 11215 10141
rect 11335 10141 11437 10235
tri 11437 10141 11535 10239 sw
tri 11535 10141 11633 10239 ne
rect 11633 10235 11987 10239
rect 11633 10141 11765 10235
rect 11335 10115 11535 10141
rect 11113 10111 11535 10115
tri 11535 10111 11565 10141 sw
tri 11633 10111 11663 10141 ne
rect 11663 10115 11765 10141
rect 11885 10141 11987 10235
tri 11987 10141 12085 10239 sw
tri 12085 10141 12183 10239 ne
rect 12183 10235 12537 10239
rect 12183 10141 12315 10235
rect 11885 10115 12085 10141
rect 11663 10111 12085 10115
tri 12085 10111 12115 10141 sw
tri 12183 10111 12213 10141 ne
rect 12213 10115 12315 10141
rect 12435 10141 12537 10235
tri 12537 10141 12635 10239 sw
tri 12635 10141 12733 10239 ne
rect 12733 10235 13087 10239
rect 12733 10141 12865 10235
rect 12435 10115 12635 10141
rect 12213 10111 12635 10115
tri 12635 10111 12665 10141 sw
tri 12733 10111 12763 10141 ne
rect 12763 10115 12865 10141
rect 12985 10141 13087 10235
tri 13087 10141 13185 10239 sw
tri 13185 10141 13283 10239 ne
rect 13283 10235 13637 10239
rect 13283 10141 13415 10235
rect 12985 10115 13185 10141
rect 12763 10111 13185 10115
tri 13185 10111 13215 10141 sw
tri 13283 10111 13313 10141 ne
rect 13313 10115 13415 10141
rect 13535 10141 13637 10235
tri 13637 10141 13735 10239 sw
tri 13735 10141 13833 10239 ne
rect 13833 10235 14187 10239
rect 13833 10141 13965 10235
rect 13535 10115 13735 10141
rect 13313 10111 13735 10115
tri 13735 10111 13765 10141 sw
tri 13833 10111 13863 10141 ne
rect 13863 10115 13965 10141
rect 14085 10141 14187 10235
tri 14187 10141 14285 10239 sw
tri 14285 10141 14383 10239 ne
rect 14383 10235 14737 10239
rect 14383 10141 14515 10235
rect 14085 10115 14285 10141
rect 13863 10111 14285 10115
tri 14285 10111 14315 10141 sw
tri 14383 10111 14413 10141 ne
rect 14413 10115 14515 10141
rect 14635 10141 14737 10235
tri 14737 10141 14835 10239 sw
tri 14835 10141 14933 10239 ne
rect 14933 10235 15287 10239
rect 14933 10141 15065 10235
rect 14635 10115 14835 10141
rect 14413 10111 14835 10115
tri 14835 10111 14865 10141 sw
tri 14933 10111 14963 10141 ne
rect 14963 10115 15065 10141
rect 15185 10141 15287 10235
tri 15287 10141 15385 10239 sw
tri 15385 10141 15483 10239 ne
rect 15483 10235 15837 10239
rect 15483 10141 15615 10235
rect 15185 10115 15385 10141
rect 14963 10111 15385 10115
tri 15385 10111 15415 10141 sw
tri 15483 10111 15513 10141 ne
rect 15513 10115 15615 10141
rect 15735 10141 15837 10235
tri 15837 10141 15935 10239 sw
tri 15935 10141 16033 10239 ne
rect 16033 10235 16387 10239
rect 16033 10141 16165 10235
rect 15735 10115 15935 10141
rect 15513 10111 15935 10115
tri 15935 10111 15965 10141 sw
tri 16033 10111 16063 10141 ne
rect 16063 10115 16165 10141
rect 16285 10141 16387 10235
tri 16387 10141 16485 10239 sw
tri 16485 10141 16583 10239 ne
rect 16583 10235 16937 10239
rect 16583 10141 16715 10235
rect 16285 10115 16485 10141
rect 16063 10111 16485 10115
tri 16485 10111 16515 10141 sw
tri 16583 10111 16613 10141 ne
rect 16613 10115 16715 10141
rect 16835 10141 16937 10235
tri 16937 10141 17035 10239 sw
tri 17035 10141 17133 10239 ne
rect 17133 10235 17487 10239
rect 17133 10141 17265 10235
rect 16835 10115 17035 10141
rect 16613 10111 17035 10115
tri 17035 10111 17065 10141 sw
tri 17133 10111 17163 10141 ne
rect 17163 10115 17265 10141
rect 17385 10141 17487 10235
tri 17487 10141 17585 10239 sw
tri 17585 10141 17683 10239 ne
rect 17683 10235 18037 10239
rect 17683 10141 17815 10235
rect 17385 10115 17585 10141
rect 17163 10111 17585 10115
tri 17585 10111 17615 10141 sw
tri 17683 10111 17713 10141 ne
rect 17713 10115 17815 10141
rect 17935 10141 18037 10235
tri 18037 10141 18135 10239 sw
tri 18135 10141 18233 10239 ne
rect 18233 10235 18587 10239
rect 18233 10141 18365 10235
rect 17935 10115 18135 10141
rect 17713 10111 18135 10115
tri 18135 10111 18165 10141 sw
tri 18233 10111 18263 10141 ne
rect 18263 10115 18365 10141
rect 18485 10141 18587 10235
tri 18587 10141 18685 10239 sw
tri 18685 10141 18783 10239 ne
rect 18783 10235 19137 10239
rect 18783 10141 18915 10235
rect 18485 10115 18685 10141
rect 18263 10111 18685 10115
tri 18685 10111 18715 10141 sw
tri 18783 10111 18813 10141 ne
rect 18813 10115 18915 10141
rect 19035 10141 19137 10235
tri 19137 10141 19235 10239 sw
tri 19235 10141 19333 10239 ne
rect 19333 10235 20300 10239
rect 19333 10141 19465 10235
rect 19035 10115 19235 10141
rect 18813 10111 19235 10115
tri 19235 10111 19265 10141 sw
tri 19333 10111 19363 10141 ne
rect 19363 10115 19465 10141
rect 19585 10115 20300 10235
rect 19363 10111 20300 10115
tri 113 10013 211 10111 ne
rect 211 10013 565 10111
tri 565 10013 663 10111 sw
tri 663 10013 761 10111 ne
rect 761 10013 1115 10111
tri 1115 10013 1213 10111 sw
tri 1213 10013 1311 10111 ne
rect 1311 10013 1665 10111
tri 1665 10013 1763 10111 sw
tri 1763 10013 1861 10111 ne
rect 1861 10013 2215 10111
tri 2215 10013 2313 10111 sw
tri 2313 10013 2411 10111 ne
rect 2411 10013 2765 10111
tri 2765 10013 2863 10111 sw
tri 2863 10013 2961 10111 ne
rect 2961 10013 3315 10111
tri 3315 10013 3413 10111 sw
tri 3413 10013 3511 10111 ne
rect 3511 10013 3865 10111
tri 3865 10013 3963 10111 sw
tri 3963 10013 4061 10111 ne
rect 4061 10013 4415 10111
tri 4415 10013 4513 10111 sw
tri 4513 10013 4611 10111 ne
rect 4611 10013 4965 10111
tri 4965 10013 5063 10111 sw
tri 5063 10013 5161 10111 ne
rect 5161 10013 5515 10111
tri 5515 10013 5613 10111 sw
tri 5613 10013 5711 10111 ne
rect 5711 10013 6065 10111
tri 6065 10013 6163 10111 sw
tri 6163 10013 6261 10111 ne
rect 6261 10013 6615 10111
tri 6615 10013 6713 10111 sw
tri 6713 10013 6811 10111 ne
rect 6811 10013 7165 10111
tri 7165 10013 7263 10111 sw
tri 7263 10013 7361 10111 ne
rect 7361 10013 7715 10111
tri 7715 10013 7813 10111 sw
tri 7813 10013 7911 10111 ne
rect 7911 10013 8265 10111
tri 8265 10013 8363 10111 sw
tri 8363 10013 8461 10111 ne
rect 8461 10013 8815 10111
tri 8815 10013 8913 10111 sw
tri 8913 10013 9011 10111 ne
rect 9011 10013 9365 10111
tri 9365 10013 9463 10111 sw
tri 9463 10013 9561 10111 ne
rect 9561 10013 9915 10111
tri 9915 10013 10013 10111 sw
tri 10013 10013 10111 10111 ne
rect 10111 10013 10465 10111
tri 10465 10013 10563 10111 sw
tri 10563 10013 10661 10111 ne
rect 10661 10013 11015 10111
tri 11015 10013 11113 10111 sw
tri 11113 10013 11211 10111 ne
rect 11211 10013 11565 10111
tri 11565 10013 11663 10111 sw
tri 11663 10013 11761 10111 ne
rect 11761 10013 12115 10111
tri 12115 10013 12213 10111 sw
tri 12213 10013 12311 10111 ne
rect 12311 10013 12665 10111
tri 12665 10013 12763 10111 sw
tri 12763 10013 12861 10111 ne
rect 12861 10013 13215 10111
tri 13215 10013 13313 10111 sw
tri 13313 10013 13411 10111 ne
rect 13411 10013 13765 10111
tri 13765 10013 13863 10111 sw
tri 13863 10013 13961 10111 ne
rect 13961 10013 14315 10111
tri 14315 10013 14413 10111 sw
tri 14413 10013 14511 10111 ne
rect 14511 10013 14865 10111
tri 14865 10013 14963 10111 sw
tri 14963 10013 15061 10111 ne
rect 15061 10013 15415 10111
tri 15415 10013 15513 10111 sw
tri 15513 10013 15611 10111 ne
rect 15611 10013 15965 10111
tri 15965 10013 16063 10111 sw
tri 16063 10013 16161 10111 ne
rect 16161 10013 16515 10111
tri 16515 10013 16613 10111 sw
tri 16613 10013 16711 10111 ne
rect 16711 10013 17065 10111
tri 17065 10013 17163 10111 sw
tri 17163 10013 17261 10111 ne
rect 17261 10013 17615 10111
tri 17615 10013 17713 10111 sw
tri 17713 10013 17811 10111 ne
rect 17811 10013 18165 10111
tri 18165 10013 18263 10111 sw
tri 18263 10013 18361 10111 ne
rect 18361 10013 18715 10111
tri 18715 10013 18813 10111 sw
tri 18813 10013 18911 10111 ne
rect 18911 10013 19265 10111
tri 19265 10013 19363 10111 sw
tri 19363 10013 19461 10111 ne
rect 19461 10013 20300 10111
rect -2000 9983 113 10013
tri 113 9983 143 10013 sw
tri 211 9983 241 10013 ne
rect 241 9983 663 10013
tri 663 9983 693 10013 sw
tri 761 9983 791 10013 ne
rect 791 9983 1213 10013
tri 1213 9983 1243 10013 sw
tri 1311 9983 1341 10013 ne
rect 1341 9983 1763 10013
tri 1763 9983 1793 10013 sw
tri 1861 9983 1891 10013 ne
rect 1891 9983 2313 10013
tri 2313 9983 2343 10013 sw
tri 2411 9983 2441 10013 ne
rect 2441 9983 2863 10013
tri 2863 9983 2893 10013 sw
tri 2961 9983 2991 10013 ne
rect 2991 9983 3413 10013
tri 3413 9983 3443 10013 sw
tri 3511 9983 3541 10013 ne
rect 3541 9983 3963 10013
tri 3963 9983 3993 10013 sw
tri 4061 9983 4091 10013 ne
rect 4091 9983 4513 10013
tri 4513 9983 4543 10013 sw
tri 4611 9983 4641 10013 ne
rect 4641 9983 5063 10013
tri 5063 9983 5093 10013 sw
tri 5161 9983 5191 10013 ne
rect 5191 9983 5613 10013
tri 5613 9983 5643 10013 sw
tri 5711 9983 5741 10013 ne
rect 5741 9983 6163 10013
tri 6163 9983 6193 10013 sw
tri 6261 9983 6291 10013 ne
rect 6291 9983 6713 10013
tri 6713 9983 6743 10013 sw
tri 6811 9983 6841 10013 ne
rect 6841 9983 7263 10013
tri 7263 9983 7293 10013 sw
tri 7361 9983 7391 10013 ne
rect 7391 9983 7813 10013
tri 7813 9983 7843 10013 sw
tri 7911 9983 7941 10013 ne
rect 7941 9983 8363 10013
tri 8363 9983 8393 10013 sw
tri 8461 9983 8491 10013 ne
rect 8491 9983 8913 10013
tri 8913 9983 8943 10013 sw
tri 9011 9983 9041 10013 ne
rect 9041 9983 9463 10013
tri 9463 9983 9493 10013 sw
tri 9561 9983 9591 10013 ne
rect 9591 9983 10013 10013
tri 10013 9983 10043 10013 sw
tri 10111 9983 10141 10013 ne
rect 10141 9983 10563 10013
tri 10563 9983 10593 10013 sw
tri 10661 9983 10691 10013 ne
rect 10691 9983 11113 10013
tri 11113 9983 11143 10013 sw
tri 11211 9983 11241 10013 ne
rect 11241 9983 11663 10013
tri 11663 9983 11693 10013 sw
tri 11761 9983 11791 10013 ne
rect 11791 9983 12213 10013
tri 12213 9983 12243 10013 sw
tri 12311 9983 12341 10013 ne
rect 12341 9983 12763 10013
tri 12763 9983 12793 10013 sw
tri 12861 9983 12891 10013 ne
rect 12891 9983 13313 10013
tri 13313 9983 13343 10013 sw
tri 13411 9983 13441 10013 ne
rect 13441 9983 13863 10013
tri 13863 9983 13893 10013 sw
tri 13961 9983 13991 10013 ne
rect 13991 9983 14413 10013
tri 14413 9983 14443 10013 sw
tri 14511 9983 14541 10013 ne
rect 14541 9983 14963 10013
tri 14963 9983 14993 10013 sw
tri 15061 9983 15091 10013 ne
rect 15091 9983 15513 10013
tri 15513 9983 15543 10013 sw
tri 15611 9983 15641 10013 ne
rect 15641 9983 16063 10013
tri 16063 9983 16093 10013 sw
tri 16161 9983 16191 10013 ne
rect 16191 9983 16613 10013
tri 16613 9983 16643 10013 sw
tri 16711 9983 16741 10013 ne
rect 16741 9983 17163 10013
tri 17163 9983 17193 10013 sw
tri 17261 9983 17291 10013 ne
rect 17291 9983 17713 10013
tri 17713 9983 17743 10013 sw
tri 17811 9983 17841 10013 ne
rect 17841 9983 18263 10013
tri 18263 9983 18293 10013 sw
tri 18361 9983 18391 10013 ne
rect 18391 9983 18813 10013
tri 18813 9983 18843 10013 sw
tri 18911 9983 18941 10013 ne
rect 18941 9983 19363 10013
tri 19363 9983 19393 10013 sw
tri 19461 9983 19491 10013 ne
rect 19491 9983 20300 10013
rect -2000 9885 143 9983
tri 143 9885 241 9983 sw
tri 241 9885 339 9983 ne
rect 339 9885 693 9983
tri 693 9885 791 9983 sw
tri 791 9885 889 9983 ne
rect 889 9885 1243 9983
tri 1243 9885 1341 9983 sw
tri 1341 9885 1439 9983 ne
rect 1439 9885 1793 9983
tri 1793 9885 1891 9983 sw
tri 1891 9885 1989 9983 ne
rect 1989 9885 2343 9983
tri 2343 9885 2441 9983 sw
tri 2441 9885 2539 9983 ne
rect 2539 9885 2893 9983
tri 2893 9885 2991 9983 sw
tri 2991 9885 3089 9983 ne
rect 3089 9885 3443 9983
tri 3443 9885 3541 9983 sw
tri 3541 9885 3639 9983 ne
rect 3639 9885 3993 9983
tri 3993 9885 4091 9983 sw
tri 4091 9885 4189 9983 ne
rect 4189 9885 4543 9983
tri 4543 9885 4641 9983 sw
tri 4641 9885 4739 9983 ne
rect 4739 9885 5093 9983
tri 5093 9885 5191 9983 sw
tri 5191 9885 5289 9983 ne
rect 5289 9885 5643 9983
tri 5643 9885 5741 9983 sw
tri 5741 9885 5839 9983 ne
rect 5839 9885 6193 9983
tri 6193 9885 6291 9983 sw
tri 6291 9885 6389 9983 ne
rect 6389 9885 6743 9983
tri 6743 9885 6841 9983 sw
tri 6841 9885 6939 9983 ne
rect 6939 9885 7293 9983
tri 7293 9885 7391 9983 sw
tri 7391 9885 7489 9983 ne
rect 7489 9885 7843 9983
tri 7843 9885 7941 9983 sw
tri 7941 9885 8039 9983 ne
rect 8039 9885 8393 9983
tri 8393 9885 8491 9983 sw
tri 8491 9885 8589 9983 ne
rect 8589 9885 8943 9983
tri 8943 9885 9041 9983 sw
tri 9041 9885 9139 9983 ne
rect 9139 9885 9493 9983
tri 9493 9885 9591 9983 sw
tri 9591 9885 9689 9983 ne
rect 9689 9885 10043 9983
tri 10043 9885 10141 9983 sw
tri 10141 9885 10239 9983 ne
rect 10239 9885 10593 9983
tri 10593 9885 10691 9983 sw
tri 10691 9885 10789 9983 ne
rect 10789 9885 11143 9983
tri 11143 9885 11241 9983 sw
tri 11241 9885 11339 9983 ne
rect 11339 9885 11693 9983
tri 11693 9885 11791 9983 sw
tri 11791 9885 11889 9983 ne
rect 11889 9885 12243 9983
tri 12243 9885 12341 9983 sw
tri 12341 9885 12439 9983 ne
rect 12439 9885 12793 9983
tri 12793 9885 12891 9983 sw
tri 12891 9885 12989 9983 ne
rect 12989 9885 13343 9983
tri 13343 9885 13441 9983 sw
tri 13441 9885 13539 9983 ne
rect 13539 9885 13893 9983
tri 13893 9885 13991 9983 sw
tri 13991 9885 14089 9983 ne
rect 14089 9885 14443 9983
tri 14443 9885 14541 9983 sw
tri 14541 9885 14639 9983 ne
rect 14639 9885 14993 9983
tri 14993 9885 15091 9983 sw
tri 15091 9885 15189 9983 ne
rect 15189 9885 15543 9983
tri 15543 9885 15641 9983 sw
tri 15641 9885 15739 9983 ne
rect 15739 9885 16093 9983
tri 16093 9885 16191 9983 sw
tri 16191 9885 16289 9983 ne
rect 16289 9885 16643 9983
tri 16643 9885 16741 9983 sw
tri 16741 9885 16839 9983 ne
rect 16839 9885 17193 9983
tri 17193 9885 17291 9983 sw
tri 17291 9885 17389 9983 ne
rect 17389 9885 17743 9983
tri 17743 9885 17841 9983 sw
tri 17841 9885 17939 9983 ne
rect 17939 9885 18293 9983
tri 18293 9885 18391 9983 sw
tri 18391 9885 18489 9983 ne
rect 18489 9885 18843 9983
tri 18843 9885 18941 9983 sw
tri 18941 9885 19039 9983 ne
rect 19039 9885 19393 9983
tri 19393 9885 19491 9983 sw
tri 19491 9885 19589 9983 ne
rect 19589 9885 20300 9983
rect -2000 9787 241 9885
tri 241 9787 339 9885 sw
tri 339 9787 437 9885 ne
rect 437 9787 791 9885
tri 791 9787 889 9885 sw
tri 889 9787 987 9885 ne
rect 987 9787 1341 9885
tri 1341 9787 1439 9885 sw
tri 1439 9787 1537 9885 ne
rect 1537 9787 1891 9885
tri 1891 9787 1989 9885 sw
tri 1989 9787 2087 9885 ne
rect 2087 9787 2441 9885
tri 2441 9787 2539 9885 sw
tri 2539 9787 2637 9885 ne
rect 2637 9787 2991 9885
tri 2991 9787 3089 9885 sw
tri 3089 9787 3187 9885 ne
rect 3187 9787 3541 9885
tri 3541 9787 3639 9885 sw
tri 3639 9787 3737 9885 ne
rect 3737 9787 4091 9885
tri 4091 9787 4189 9885 sw
tri 4189 9787 4287 9885 ne
rect 4287 9787 4641 9885
tri 4641 9787 4739 9885 sw
tri 4739 9787 4837 9885 ne
rect 4837 9787 5191 9885
tri 5191 9787 5289 9885 sw
tri 5289 9787 5387 9885 ne
rect 5387 9787 5741 9885
tri 5741 9787 5839 9885 sw
tri 5839 9787 5937 9885 ne
rect 5937 9787 6291 9885
tri 6291 9787 6389 9885 sw
tri 6389 9787 6487 9885 ne
rect 6487 9787 6841 9885
tri 6841 9787 6939 9885 sw
tri 6939 9787 7037 9885 ne
rect 7037 9787 7391 9885
tri 7391 9787 7489 9885 sw
tri 7489 9787 7587 9885 ne
rect 7587 9787 7941 9885
tri 7941 9787 8039 9885 sw
tri 8039 9787 8137 9885 ne
rect 8137 9787 8491 9885
tri 8491 9787 8589 9885 sw
tri 8589 9787 8687 9885 ne
rect 8687 9787 9041 9885
tri 9041 9787 9139 9885 sw
tri 9139 9787 9237 9885 ne
rect 9237 9787 9591 9885
tri 9591 9787 9689 9885 sw
tri 9689 9787 9787 9885 ne
rect 9787 9787 10141 9885
tri 10141 9787 10239 9885 sw
tri 10239 9787 10337 9885 ne
rect 10337 9787 10691 9885
tri 10691 9787 10789 9885 sw
tri 10789 9787 10887 9885 ne
rect 10887 9787 11241 9885
tri 11241 9787 11339 9885 sw
tri 11339 9787 11437 9885 ne
rect 11437 9787 11791 9885
tri 11791 9787 11889 9885 sw
tri 11889 9787 11987 9885 ne
rect 11987 9787 12341 9885
tri 12341 9787 12439 9885 sw
tri 12439 9787 12537 9885 ne
rect 12537 9787 12891 9885
tri 12891 9787 12989 9885 sw
tri 12989 9787 13087 9885 ne
rect 13087 9787 13441 9885
tri 13441 9787 13539 9885 sw
tri 13539 9787 13637 9885 ne
rect 13637 9787 13991 9885
tri 13991 9787 14089 9885 sw
tri 14089 9787 14187 9885 ne
rect 14187 9787 14541 9885
tri 14541 9787 14639 9885 sw
tri 14639 9787 14737 9885 ne
rect 14737 9787 15091 9885
tri 15091 9787 15189 9885 sw
tri 15189 9787 15287 9885 ne
rect 15287 9787 15641 9885
tri 15641 9787 15739 9885 sw
tri 15739 9787 15837 9885 ne
rect 15837 9787 16191 9885
tri 16191 9787 16289 9885 sw
tri 16289 9787 16387 9885 ne
rect 16387 9787 16741 9885
tri 16741 9787 16839 9885 sw
tri 16839 9787 16937 9885 ne
rect 16937 9787 17291 9885
tri 17291 9787 17389 9885 sw
tri 17389 9787 17487 9885 ne
rect 17487 9787 17841 9885
tri 17841 9787 17939 9885 sw
tri 17939 9787 18037 9885 ne
rect 18037 9787 18391 9885
tri 18391 9787 18489 9885 sw
tri 18489 9787 18587 9885 ne
rect 18587 9787 18941 9885
tri 18941 9787 19039 9885 sw
tri 19039 9787 19137 9885 ne
rect 19137 9787 19491 9885
tri 19491 9787 19589 9885 sw
tri 19589 9787 19687 9885 ne
rect 19687 9787 20300 9885
rect -2000 9689 339 9787
tri 339 9689 437 9787 sw
tri 437 9689 535 9787 ne
rect 535 9689 889 9787
tri 889 9689 987 9787 sw
tri 987 9689 1085 9787 ne
rect 1085 9689 1439 9787
tri 1439 9689 1537 9787 sw
tri 1537 9689 1635 9787 ne
rect 1635 9689 1989 9787
tri 1989 9689 2087 9787 sw
tri 2087 9689 2185 9787 ne
rect 2185 9689 2539 9787
tri 2539 9689 2637 9787 sw
tri 2637 9689 2735 9787 ne
rect 2735 9689 3089 9787
tri 3089 9689 3187 9787 sw
tri 3187 9689 3285 9787 ne
rect 3285 9689 3639 9787
tri 3639 9689 3737 9787 sw
tri 3737 9689 3835 9787 ne
rect 3835 9689 4189 9787
tri 4189 9689 4287 9787 sw
tri 4287 9689 4385 9787 ne
rect 4385 9689 4739 9787
tri 4739 9689 4837 9787 sw
tri 4837 9689 4935 9787 ne
rect 4935 9689 5289 9787
tri 5289 9689 5387 9787 sw
tri 5387 9689 5485 9787 ne
rect 5485 9689 5839 9787
tri 5839 9689 5937 9787 sw
tri 5937 9689 6035 9787 ne
rect 6035 9689 6389 9787
tri 6389 9689 6487 9787 sw
tri 6487 9689 6585 9787 ne
rect 6585 9689 6939 9787
tri 6939 9689 7037 9787 sw
tri 7037 9689 7135 9787 ne
rect 7135 9689 7489 9787
tri 7489 9689 7587 9787 sw
tri 7587 9689 7685 9787 ne
rect 7685 9689 8039 9787
tri 8039 9689 8137 9787 sw
tri 8137 9689 8235 9787 ne
rect 8235 9689 8589 9787
tri 8589 9689 8687 9787 sw
tri 8687 9689 8785 9787 ne
rect 8785 9689 9139 9787
tri 9139 9689 9237 9787 sw
tri 9237 9689 9335 9787 ne
rect 9335 9689 9689 9787
tri 9689 9689 9787 9787 sw
tri 9787 9689 9885 9787 ne
rect 9885 9689 10239 9787
tri 10239 9689 10337 9787 sw
tri 10337 9689 10435 9787 ne
rect 10435 9689 10789 9787
tri 10789 9689 10887 9787 sw
tri 10887 9689 10985 9787 ne
rect 10985 9689 11339 9787
tri 11339 9689 11437 9787 sw
tri 11437 9689 11535 9787 ne
rect 11535 9689 11889 9787
tri 11889 9689 11987 9787 sw
tri 11987 9689 12085 9787 ne
rect 12085 9689 12439 9787
tri 12439 9689 12537 9787 sw
tri 12537 9689 12635 9787 ne
rect 12635 9689 12989 9787
tri 12989 9689 13087 9787 sw
tri 13087 9689 13185 9787 ne
rect 13185 9689 13539 9787
tri 13539 9689 13637 9787 sw
tri 13637 9689 13735 9787 ne
rect 13735 9689 14089 9787
tri 14089 9689 14187 9787 sw
tri 14187 9689 14285 9787 ne
rect 14285 9689 14639 9787
tri 14639 9689 14737 9787 sw
tri 14737 9689 14835 9787 ne
rect 14835 9689 15189 9787
tri 15189 9689 15287 9787 sw
tri 15287 9689 15385 9787 ne
rect 15385 9689 15739 9787
tri 15739 9689 15837 9787 sw
tri 15837 9689 15935 9787 ne
rect 15935 9689 16289 9787
tri 16289 9689 16387 9787 sw
tri 16387 9689 16485 9787 ne
rect 16485 9689 16839 9787
tri 16839 9689 16937 9787 sw
tri 16937 9689 17035 9787 ne
rect 17035 9689 17389 9787
tri 17389 9689 17487 9787 sw
tri 17487 9689 17585 9787 ne
rect 17585 9689 17939 9787
tri 17939 9689 18037 9787 sw
tri 18037 9689 18135 9787 ne
rect 18135 9689 18489 9787
tri 18489 9689 18587 9787 sw
tri 18587 9689 18685 9787 ne
rect 18685 9689 19039 9787
tri 19039 9689 19137 9787 sw
tri 19137 9689 19235 9787 ne
rect 19235 9689 19589 9787
tri 19589 9689 19687 9787 sw
rect 20800 9689 21800 10337
rect -2000 9685 437 9689
rect -2000 9565 215 9685
rect 335 9591 437 9685
tri 437 9591 535 9689 sw
tri 535 9591 633 9689 ne
rect 633 9685 987 9689
rect 633 9591 765 9685
rect 335 9565 535 9591
rect -2000 9561 535 9565
rect -2000 8913 -1000 9561
tri 113 9463 211 9561 ne
rect 211 9513 535 9561
tri 535 9513 613 9591 sw
tri 633 9513 711 9591 ne
rect 711 9565 765 9591
rect 885 9591 987 9685
tri 987 9591 1085 9689 sw
tri 1085 9591 1183 9689 ne
rect 1183 9685 1537 9689
rect 1183 9591 1315 9685
rect 885 9565 1085 9591
rect 711 9513 1085 9565
tri 1085 9513 1163 9591 sw
tri 1183 9513 1261 9591 ne
rect 1261 9565 1315 9591
rect 1435 9591 1537 9685
tri 1537 9591 1635 9689 sw
tri 1635 9591 1733 9689 ne
rect 1733 9685 2087 9689
rect 1733 9591 1865 9685
rect 1435 9565 1635 9591
rect 1261 9513 1635 9565
tri 1635 9513 1713 9591 sw
tri 1733 9513 1811 9591 ne
rect 1811 9565 1865 9591
rect 1985 9591 2087 9685
tri 2087 9591 2185 9689 sw
tri 2185 9591 2283 9689 ne
rect 2283 9685 2637 9689
rect 2283 9591 2415 9685
rect 1985 9565 2185 9591
rect 1811 9513 2185 9565
tri 2185 9513 2263 9591 sw
tri 2283 9513 2361 9591 ne
rect 2361 9565 2415 9591
rect 2535 9591 2637 9685
tri 2637 9591 2735 9689 sw
tri 2735 9591 2833 9689 ne
rect 2833 9685 3187 9689
rect 2833 9591 2965 9685
rect 2535 9565 2735 9591
rect 2361 9513 2735 9565
tri 2735 9513 2813 9591 sw
tri 2833 9513 2911 9591 ne
rect 2911 9565 2965 9591
rect 3085 9591 3187 9685
tri 3187 9591 3285 9689 sw
tri 3285 9591 3383 9689 ne
rect 3383 9685 3737 9689
rect 3383 9591 3515 9685
rect 3085 9565 3285 9591
rect 2911 9513 3285 9565
tri 3285 9513 3363 9591 sw
tri 3383 9513 3461 9591 ne
rect 3461 9565 3515 9591
rect 3635 9591 3737 9685
tri 3737 9591 3835 9689 sw
tri 3835 9591 3933 9689 ne
rect 3933 9685 4287 9689
rect 3933 9591 4065 9685
rect 3635 9565 3835 9591
rect 3461 9513 3835 9565
tri 3835 9513 3913 9591 sw
tri 3933 9513 4011 9591 ne
rect 4011 9565 4065 9591
rect 4185 9591 4287 9685
tri 4287 9591 4385 9689 sw
tri 4385 9591 4483 9689 ne
rect 4483 9685 4837 9689
rect 4483 9591 4615 9685
rect 4185 9565 4385 9591
rect 4011 9513 4385 9565
tri 4385 9513 4463 9591 sw
tri 4483 9513 4561 9591 ne
rect 4561 9565 4615 9591
rect 4735 9591 4837 9685
tri 4837 9591 4935 9689 sw
tri 4935 9591 5033 9689 ne
rect 5033 9685 5387 9689
rect 5033 9591 5165 9685
rect 4735 9565 4935 9591
rect 4561 9513 4935 9565
tri 4935 9513 5013 9591 sw
tri 5033 9513 5111 9591 ne
rect 5111 9565 5165 9591
rect 5285 9591 5387 9685
tri 5387 9591 5485 9689 sw
tri 5485 9591 5583 9689 ne
rect 5583 9685 5937 9689
rect 5583 9591 5715 9685
rect 5285 9565 5485 9591
rect 5111 9513 5485 9565
tri 5485 9513 5563 9591 sw
tri 5583 9513 5661 9591 ne
rect 5661 9565 5715 9591
rect 5835 9591 5937 9685
tri 5937 9591 6035 9689 sw
tri 6035 9591 6133 9689 ne
rect 6133 9685 6487 9689
rect 6133 9591 6265 9685
rect 5835 9565 6035 9591
rect 5661 9513 6035 9565
tri 6035 9513 6113 9591 sw
tri 6133 9513 6211 9591 ne
rect 6211 9565 6265 9591
rect 6385 9591 6487 9685
tri 6487 9591 6585 9689 sw
tri 6585 9591 6683 9689 ne
rect 6683 9685 7037 9689
rect 6683 9591 6815 9685
rect 6385 9565 6585 9591
rect 6211 9513 6585 9565
tri 6585 9513 6663 9591 sw
tri 6683 9513 6761 9591 ne
rect 6761 9565 6815 9591
rect 6935 9591 7037 9685
tri 7037 9591 7135 9689 sw
tri 7135 9591 7233 9689 ne
rect 7233 9685 7587 9689
rect 7233 9591 7365 9685
rect 6935 9565 7135 9591
rect 6761 9513 7135 9565
tri 7135 9513 7213 9591 sw
tri 7233 9513 7311 9591 ne
rect 7311 9565 7365 9591
rect 7485 9591 7587 9685
tri 7587 9591 7685 9689 sw
tri 7685 9591 7783 9689 ne
rect 7783 9685 8137 9689
rect 7783 9591 7915 9685
rect 7485 9565 7685 9591
rect 7311 9513 7685 9565
tri 7685 9513 7763 9591 sw
tri 7783 9513 7861 9591 ne
rect 7861 9565 7915 9591
rect 8035 9591 8137 9685
tri 8137 9591 8235 9689 sw
tri 8235 9591 8333 9689 ne
rect 8333 9685 8687 9689
rect 8333 9591 8465 9685
rect 8035 9565 8235 9591
rect 7861 9513 8235 9565
tri 8235 9513 8313 9591 sw
tri 8333 9513 8411 9591 ne
rect 8411 9565 8465 9591
rect 8585 9591 8687 9685
tri 8687 9591 8785 9689 sw
tri 8785 9591 8883 9689 ne
rect 8883 9685 9237 9689
rect 8883 9591 9015 9685
rect 8585 9565 8785 9591
rect 8411 9513 8785 9565
tri 8785 9513 8863 9591 sw
tri 8883 9513 8961 9591 ne
rect 8961 9565 9015 9591
rect 9135 9591 9237 9685
tri 9237 9591 9335 9689 sw
tri 9335 9591 9433 9689 ne
rect 9433 9685 9787 9689
rect 9433 9591 9565 9685
rect 9135 9565 9335 9591
rect 8961 9513 9335 9565
tri 9335 9513 9413 9591 sw
tri 9433 9513 9511 9591 ne
rect 9511 9565 9565 9591
rect 9685 9591 9787 9685
tri 9787 9591 9885 9689 sw
tri 9885 9591 9983 9689 ne
rect 9983 9685 10337 9689
rect 9983 9591 10115 9685
rect 9685 9565 9885 9591
rect 9511 9513 9885 9565
tri 9885 9513 9963 9591 sw
tri 9983 9513 10061 9591 ne
rect 10061 9565 10115 9591
rect 10235 9591 10337 9685
tri 10337 9591 10435 9689 sw
tri 10435 9591 10533 9689 ne
rect 10533 9685 10887 9689
rect 10533 9591 10665 9685
rect 10235 9565 10435 9591
rect 10061 9513 10435 9565
tri 10435 9513 10513 9591 sw
tri 10533 9513 10611 9591 ne
rect 10611 9565 10665 9591
rect 10785 9591 10887 9685
tri 10887 9591 10985 9689 sw
tri 10985 9591 11083 9689 ne
rect 11083 9685 11437 9689
rect 11083 9591 11215 9685
rect 10785 9565 10985 9591
rect 10611 9513 10985 9565
tri 10985 9513 11063 9591 sw
tri 11083 9513 11161 9591 ne
rect 11161 9565 11215 9591
rect 11335 9591 11437 9685
tri 11437 9591 11535 9689 sw
tri 11535 9591 11633 9689 ne
rect 11633 9685 11987 9689
rect 11633 9591 11765 9685
rect 11335 9565 11535 9591
rect 11161 9513 11535 9565
tri 11535 9513 11613 9591 sw
tri 11633 9513 11711 9591 ne
rect 11711 9565 11765 9591
rect 11885 9591 11987 9685
tri 11987 9591 12085 9689 sw
tri 12085 9591 12183 9689 ne
rect 12183 9685 12537 9689
rect 12183 9591 12315 9685
rect 11885 9565 12085 9591
rect 11711 9513 12085 9565
tri 12085 9513 12163 9591 sw
tri 12183 9513 12261 9591 ne
rect 12261 9565 12315 9591
rect 12435 9591 12537 9685
tri 12537 9591 12635 9689 sw
tri 12635 9591 12733 9689 ne
rect 12733 9685 13087 9689
rect 12733 9591 12865 9685
rect 12435 9565 12635 9591
rect 12261 9513 12635 9565
tri 12635 9513 12713 9591 sw
tri 12733 9513 12811 9591 ne
rect 12811 9565 12865 9591
rect 12985 9591 13087 9685
tri 13087 9591 13185 9689 sw
tri 13185 9591 13283 9689 ne
rect 13283 9685 13637 9689
rect 13283 9591 13415 9685
rect 12985 9565 13185 9591
rect 12811 9513 13185 9565
tri 13185 9513 13263 9591 sw
tri 13283 9513 13361 9591 ne
rect 13361 9565 13415 9591
rect 13535 9591 13637 9685
tri 13637 9591 13735 9689 sw
tri 13735 9591 13833 9689 ne
rect 13833 9685 14187 9689
rect 13833 9591 13965 9685
rect 13535 9565 13735 9591
rect 13361 9513 13735 9565
tri 13735 9513 13813 9591 sw
tri 13833 9513 13911 9591 ne
rect 13911 9565 13965 9591
rect 14085 9591 14187 9685
tri 14187 9591 14285 9689 sw
tri 14285 9591 14383 9689 ne
rect 14383 9685 14737 9689
rect 14383 9591 14515 9685
rect 14085 9565 14285 9591
rect 13911 9513 14285 9565
tri 14285 9513 14363 9591 sw
tri 14383 9513 14461 9591 ne
rect 14461 9565 14515 9591
rect 14635 9591 14737 9685
tri 14737 9591 14835 9689 sw
tri 14835 9591 14933 9689 ne
rect 14933 9685 15287 9689
rect 14933 9591 15065 9685
rect 14635 9565 14835 9591
rect 14461 9513 14835 9565
tri 14835 9513 14913 9591 sw
tri 14933 9513 15011 9591 ne
rect 15011 9565 15065 9591
rect 15185 9591 15287 9685
tri 15287 9591 15385 9689 sw
tri 15385 9591 15483 9689 ne
rect 15483 9685 15837 9689
rect 15483 9591 15615 9685
rect 15185 9565 15385 9591
rect 15011 9513 15385 9565
tri 15385 9513 15463 9591 sw
tri 15483 9513 15561 9591 ne
rect 15561 9565 15615 9591
rect 15735 9591 15837 9685
tri 15837 9591 15935 9689 sw
tri 15935 9591 16033 9689 ne
rect 16033 9685 16387 9689
rect 16033 9591 16165 9685
rect 15735 9565 15935 9591
rect 15561 9513 15935 9565
tri 15935 9513 16013 9591 sw
tri 16033 9513 16111 9591 ne
rect 16111 9565 16165 9591
rect 16285 9591 16387 9685
tri 16387 9591 16485 9689 sw
tri 16485 9591 16583 9689 ne
rect 16583 9685 16937 9689
rect 16583 9591 16715 9685
rect 16285 9565 16485 9591
rect 16111 9513 16485 9565
tri 16485 9513 16563 9591 sw
tri 16583 9513 16661 9591 ne
rect 16661 9565 16715 9591
rect 16835 9591 16937 9685
tri 16937 9591 17035 9689 sw
tri 17035 9591 17133 9689 ne
rect 17133 9685 17487 9689
rect 17133 9591 17265 9685
rect 16835 9565 17035 9591
rect 16661 9513 17035 9565
tri 17035 9513 17113 9591 sw
tri 17133 9513 17211 9591 ne
rect 17211 9565 17265 9591
rect 17385 9591 17487 9685
tri 17487 9591 17585 9689 sw
tri 17585 9591 17683 9689 ne
rect 17683 9685 18037 9689
rect 17683 9591 17815 9685
rect 17385 9565 17585 9591
rect 17211 9513 17585 9565
tri 17585 9513 17663 9591 sw
tri 17683 9513 17761 9591 ne
rect 17761 9565 17815 9591
rect 17935 9591 18037 9685
tri 18037 9591 18135 9689 sw
tri 18135 9591 18233 9689 ne
rect 18233 9685 18587 9689
rect 18233 9591 18365 9685
rect 17935 9565 18135 9591
rect 17761 9513 18135 9565
tri 18135 9513 18213 9591 sw
tri 18233 9513 18311 9591 ne
rect 18311 9565 18365 9591
rect 18485 9591 18587 9685
tri 18587 9591 18685 9689 sw
tri 18685 9591 18783 9689 ne
rect 18783 9685 19137 9689
rect 18783 9591 18915 9685
rect 18485 9565 18685 9591
rect 18311 9513 18685 9565
tri 18685 9513 18763 9591 sw
tri 18783 9513 18861 9591 ne
rect 18861 9565 18915 9591
rect 19035 9591 19137 9685
tri 19137 9591 19235 9689 sw
tri 19235 9591 19333 9689 ne
rect 19333 9685 21800 9689
rect 19333 9591 19465 9685
rect 19035 9565 19235 9591
rect 18861 9513 19235 9565
tri 19235 9513 19313 9591 sw
tri 19333 9513 19411 9591 ne
rect 19411 9565 19465 9591
rect 19585 9565 21800 9685
rect 19411 9513 21800 9565
rect 211 9463 613 9513
rect -500 9413 113 9463
tri 113 9413 163 9463 sw
tri 211 9413 261 9463 ne
rect 261 9433 613 9463
tri 613 9433 693 9513 sw
tri 711 9433 791 9513 ne
rect 791 9433 1163 9513
tri 1163 9433 1243 9513 sw
tri 1261 9433 1341 9513 ne
rect 1341 9433 1713 9513
tri 1713 9433 1793 9513 sw
tri 1811 9433 1891 9513 ne
rect 1891 9433 2263 9513
tri 2263 9433 2343 9513 sw
tri 2361 9433 2441 9513 ne
rect 2441 9433 2813 9513
tri 2813 9433 2893 9513 sw
tri 2911 9433 2991 9513 ne
rect 2991 9433 3363 9513
tri 3363 9433 3443 9513 sw
tri 3461 9433 3541 9513 ne
rect 3541 9433 3913 9513
tri 3913 9433 3993 9513 sw
tri 4011 9433 4091 9513 ne
rect 4091 9433 4463 9513
tri 4463 9433 4543 9513 sw
tri 4561 9433 4641 9513 ne
rect 4641 9433 5013 9513
tri 5013 9433 5093 9513 sw
tri 5111 9433 5191 9513 ne
rect 5191 9433 5563 9513
tri 5563 9433 5643 9513 sw
tri 5661 9433 5741 9513 ne
rect 5741 9433 6113 9513
tri 6113 9433 6193 9513 sw
tri 6211 9433 6291 9513 ne
rect 6291 9433 6663 9513
tri 6663 9433 6743 9513 sw
tri 6761 9433 6841 9513 ne
rect 6841 9433 7213 9513
tri 7213 9433 7293 9513 sw
tri 7311 9433 7391 9513 ne
rect 7391 9433 7763 9513
tri 7763 9433 7843 9513 sw
tri 7861 9433 7941 9513 ne
rect 7941 9433 8313 9513
tri 8313 9433 8393 9513 sw
tri 8411 9433 8491 9513 ne
rect 8491 9433 8863 9513
tri 8863 9433 8943 9513 sw
tri 8961 9433 9041 9513 ne
rect 9041 9433 9413 9513
tri 9413 9433 9493 9513 sw
tri 9511 9433 9591 9513 ne
rect 9591 9433 9963 9513
tri 9963 9433 10043 9513 sw
tri 10061 9433 10141 9513 ne
rect 10141 9433 10513 9513
tri 10513 9433 10593 9513 sw
tri 10611 9433 10691 9513 ne
rect 10691 9433 11063 9513
tri 11063 9433 11143 9513 sw
tri 11161 9433 11241 9513 ne
rect 11241 9433 11613 9513
tri 11613 9433 11693 9513 sw
tri 11711 9433 11791 9513 ne
rect 11791 9433 12163 9513
tri 12163 9433 12243 9513 sw
tri 12261 9433 12341 9513 ne
rect 12341 9433 12713 9513
tri 12713 9433 12793 9513 sw
tri 12811 9433 12891 9513 ne
rect 12891 9433 13263 9513
tri 13263 9433 13343 9513 sw
tri 13361 9433 13441 9513 ne
rect 13441 9433 13813 9513
tri 13813 9433 13893 9513 sw
tri 13911 9433 13991 9513 ne
rect 13991 9433 14363 9513
tri 14363 9433 14443 9513 sw
tri 14461 9433 14541 9513 ne
rect 14541 9433 14913 9513
tri 14913 9433 14993 9513 sw
tri 15011 9433 15091 9513 ne
rect 15091 9433 15463 9513
tri 15463 9433 15543 9513 sw
tri 15561 9433 15641 9513 ne
rect 15641 9433 16013 9513
tri 16013 9433 16093 9513 sw
tri 16111 9433 16191 9513 ne
rect 16191 9433 16563 9513
tri 16563 9433 16643 9513 sw
tri 16661 9433 16741 9513 ne
rect 16741 9433 17113 9513
tri 17113 9433 17193 9513 sw
tri 17211 9433 17291 9513 ne
rect 17291 9433 17663 9513
tri 17663 9433 17743 9513 sw
tri 17761 9433 17841 9513 ne
rect 17841 9433 18213 9513
tri 18213 9433 18293 9513 sw
tri 18311 9433 18391 9513 ne
rect 18391 9433 18763 9513
tri 18763 9433 18843 9513 sw
tri 18861 9433 18941 9513 ne
rect 18941 9433 19313 9513
tri 19313 9433 19393 9513 sw
tri 19411 9433 19491 9513 ne
rect 19491 9433 20100 9513
rect 261 9413 693 9433
rect -500 9335 163 9413
tri 163 9335 241 9413 sw
tri 261 9335 339 9413 ne
rect 339 9335 693 9413
tri 693 9335 791 9433 sw
tri 791 9335 889 9433 ne
rect 889 9335 1243 9433
tri 1243 9335 1341 9433 sw
tri 1341 9335 1439 9433 ne
rect 1439 9335 1793 9433
tri 1793 9335 1891 9433 sw
tri 1891 9335 1989 9433 ne
rect 1989 9335 2343 9433
tri 2343 9335 2441 9433 sw
tri 2441 9335 2539 9433 ne
rect 2539 9335 2893 9433
tri 2893 9335 2991 9433 sw
tri 2991 9335 3089 9433 ne
rect 3089 9335 3443 9433
tri 3443 9335 3541 9433 sw
tri 3541 9335 3639 9433 ne
rect 3639 9335 3993 9433
tri 3993 9335 4091 9433 sw
tri 4091 9335 4189 9433 ne
rect 4189 9335 4543 9433
tri 4543 9335 4641 9433 sw
tri 4641 9335 4739 9433 ne
rect 4739 9335 5093 9433
tri 5093 9335 5191 9433 sw
tri 5191 9335 5289 9433 ne
rect 5289 9335 5643 9433
tri 5643 9335 5741 9433 sw
tri 5741 9335 5839 9433 ne
rect 5839 9335 6193 9433
tri 6193 9335 6291 9433 sw
tri 6291 9335 6389 9433 ne
rect 6389 9335 6743 9433
tri 6743 9335 6841 9433 sw
tri 6841 9335 6939 9433 ne
rect 6939 9335 7293 9433
tri 7293 9335 7391 9433 sw
tri 7391 9335 7489 9433 ne
rect 7489 9335 7843 9433
tri 7843 9335 7941 9433 sw
tri 7941 9335 8039 9433 ne
rect 8039 9335 8393 9433
tri 8393 9335 8491 9433 sw
tri 8491 9335 8589 9433 ne
rect 8589 9335 8943 9433
tri 8943 9335 9041 9433 sw
tri 9041 9335 9139 9433 ne
rect 9139 9335 9493 9433
tri 9493 9335 9591 9433 sw
tri 9591 9335 9689 9433 ne
rect 9689 9335 10043 9433
tri 10043 9335 10141 9433 sw
tri 10141 9335 10239 9433 ne
rect 10239 9335 10593 9433
tri 10593 9335 10691 9433 sw
tri 10691 9335 10789 9433 ne
rect 10789 9335 11143 9433
tri 11143 9335 11241 9433 sw
tri 11241 9335 11339 9433 ne
rect 11339 9335 11693 9433
tri 11693 9335 11791 9433 sw
tri 11791 9335 11889 9433 ne
rect 11889 9335 12243 9433
tri 12243 9335 12341 9433 sw
tri 12341 9335 12439 9433 ne
rect 12439 9335 12793 9433
tri 12793 9335 12891 9433 sw
tri 12891 9335 12989 9433 ne
rect 12989 9335 13343 9433
tri 13343 9335 13441 9433 sw
tri 13441 9335 13539 9433 ne
rect 13539 9335 13893 9433
tri 13893 9335 13991 9433 sw
tri 13991 9335 14089 9433 ne
rect 14089 9335 14443 9433
tri 14443 9335 14541 9433 sw
tri 14541 9335 14639 9433 ne
rect 14639 9335 14993 9433
tri 14993 9335 15091 9433 sw
tri 15091 9335 15189 9433 ne
rect 15189 9335 15543 9433
tri 15543 9335 15641 9433 sw
tri 15641 9335 15739 9433 ne
rect 15739 9335 16093 9433
tri 16093 9335 16191 9433 sw
tri 16191 9335 16289 9433 ne
rect 16289 9335 16643 9433
tri 16643 9335 16741 9433 sw
tri 16741 9335 16839 9433 ne
rect 16839 9335 17193 9433
tri 17193 9335 17291 9433 sw
tri 17291 9335 17389 9433 ne
rect 17389 9335 17743 9433
tri 17743 9335 17841 9433 sw
tri 17841 9335 17939 9433 ne
rect 17939 9335 18293 9433
tri 18293 9335 18391 9433 sw
tri 18391 9335 18489 9433 ne
rect 18489 9335 18843 9433
tri 18843 9335 18941 9433 sw
tri 18941 9335 19039 9433 ne
rect 19039 9335 19393 9433
tri 19393 9335 19491 9433 sw
tri 19491 9335 19589 9433 ne
rect 19589 9413 20100 9433
rect 20200 9413 21800 9513
rect 19589 9335 21800 9413
rect -500 9287 241 9335
rect -500 9187 -400 9287
rect -300 9237 241 9287
tri 241 9237 339 9335 sw
tri 339 9237 437 9335 ne
rect 437 9237 791 9335
tri 791 9237 889 9335 sw
tri 889 9237 987 9335 ne
rect 987 9237 1341 9335
tri 1341 9237 1439 9335 sw
tri 1439 9237 1537 9335 ne
rect 1537 9237 1891 9335
tri 1891 9237 1989 9335 sw
tri 1989 9237 2087 9335 ne
rect 2087 9237 2441 9335
tri 2441 9237 2539 9335 sw
tri 2539 9237 2637 9335 ne
rect 2637 9237 2991 9335
tri 2991 9237 3089 9335 sw
tri 3089 9237 3187 9335 ne
rect 3187 9237 3541 9335
tri 3541 9237 3639 9335 sw
tri 3639 9237 3737 9335 ne
rect 3737 9237 4091 9335
tri 4091 9237 4189 9335 sw
tri 4189 9237 4287 9335 ne
rect 4287 9237 4641 9335
tri 4641 9237 4739 9335 sw
tri 4739 9237 4837 9335 ne
rect 4837 9237 5191 9335
tri 5191 9237 5289 9335 sw
tri 5289 9237 5387 9335 ne
rect 5387 9237 5741 9335
tri 5741 9237 5839 9335 sw
tri 5839 9237 5937 9335 ne
rect 5937 9237 6291 9335
tri 6291 9237 6389 9335 sw
tri 6389 9237 6487 9335 ne
rect 6487 9237 6841 9335
tri 6841 9237 6939 9335 sw
tri 6939 9237 7037 9335 ne
rect 7037 9237 7391 9335
tri 7391 9237 7489 9335 sw
tri 7489 9237 7587 9335 ne
rect 7587 9237 7941 9335
tri 7941 9237 8039 9335 sw
tri 8039 9237 8137 9335 ne
rect 8137 9237 8491 9335
tri 8491 9237 8589 9335 sw
tri 8589 9237 8687 9335 ne
rect 8687 9237 9041 9335
tri 9041 9237 9139 9335 sw
tri 9139 9237 9237 9335 ne
rect 9237 9237 9591 9335
tri 9591 9237 9689 9335 sw
tri 9689 9237 9787 9335 ne
rect 9787 9237 10141 9335
tri 10141 9237 10239 9335 sw
tri 10239 9237 10337 9335 ne
rect 10337 9237 10691 9335
tri 10691 9237 10789 9335 sw
tri 10789 9237 10887 9335 ne
rect 10887 9237 11241 9335
tri 11241 9237 11339 9335 sw
tri 11339 9237 11437 9335 ne
rect 11437 9237 11791 9335
tri 11791 9237 11889 9335 sw
tri 11889 9237 11987 9335 ne
rect 11987 9237 12341 9335
tri 12341 9237 12439 9335 sw
tri 12439 9237 12537 9335 ne
rect 12537 9237 12891 9335
tri 12891 9237 12989 9335 sw
tri 12989 9237 13087 9335 ne
rect 13087 9237 13441 9335
tri 13441 9237 13539 9335 sw
tri 13539 9237 13637 9335 ne
rect 13637 9237 13991 9335
tri 13991 9237 14089 9335 sw
tri 14089 9237 14187 9335 ne
rect 14187 9237 14541 9335
tri 14541 9237 14639 9335 sw
tri 14639 9237 14737 9335 ne
rect 14737 9237 15091 9335
tri 15091 9237 15189 9335 sw
tri 15189 9237 15287 9335 ne
rect 15287 9237 15641 9335
tri 15641 9237 15739 9335 sw
tri 15739 9237 15837 9335 ne
rect 15837 9237 16191 9335
tri 16191 9237 16289 9335 sw
tri 16289 9237 16387 9335 ne
rect 16387 9237 16741 9335
tri 16741 9237 16839 9335 sw
tri 16839 9237 16937 9335 ne
rect 16937 9237 17291 9335
tri 17291 9237 17389 9335 sw
tri 17389 9237 17487 9335 ne
rect 17487 9237 17841 9335
tri 17841 9237 17939 9335 sw
tri 17939 9237 18037 9335 ne
rect 18037 9237 18391 9335
tri 18391 9237 18489 9335 sw
tri 18489 9237 18587 9335 ne
rect 18587 9237 18941 9335
tri 18941 9237 19039 9335 sw
tri 19039 9237 19137 9335 ne
rect 19137 9237 19491 9335
tri 19491 9237 19589 9335 sw
tri 19589 9237 19687 9335 ne
rect 19687 9237 21800 9335
rect -300 9187 339 9237
rect -500 9139 339 9187
tri 339 9139 437 9237 sw
tri 437 9139 535 9237 ne
rect 535 9139 889 9237
tri 889 9139 987 9237 sw
tri 987 9139 1085 9237 ne
rect 1085 9139 1439 9237
tri 1439 9139 1537 9237 sw
tri 1537 9139 1635 9237 ne
rect 1635 9139 1989 9237
tri 1989 9139 2087 9237 sw
tri 2087 9139 2185 9237 ne
rect 2185 9139 2539 9237
tri 2539 9139 2637 9237 sw
tri 2637 9139 2735 9237 ne
rect 2735 9139 3089 9237
tri 3089 9139 3187 9237 sw
tri 3187 9139 3285 9237 ne
rect 3285 9139 3639 9237
tri 3639 9139 3737 9237 sw
tri 3737 9139 3835 9237 ne
rect 3835 9139 4189 9237
tri 4189 9139 4287 9237 sw
tri 4287 9139 4385 9237 ne
rect 4385 9139 4739 9237
tri 4739 9139 4837 9237 sw
tri 4837 9139 4935 9237 ne
rect 4935 9139 5289 9237
tri 5289 9139 5387 9237 sw
tri 5387 9139 5485 9237 ne
rect 5485 9139 5839 9237
tri 5839 9139 5937 9237 sw
tri 5937 9139 6035 9237 ne
rect 6035 9139 6389 9237
tri 6389 9139 6487 9237 sw
tri 6487 9139 6585 9237 ne
rect 6585 9139 6939 9237
tri 6939 9139 7037 9237 sw
tri 7037 9139 7135 9237 ne
rect 7135 9139 7489 9237
tri 7489 9139 7587 9237 sw
tri 7587 9139 7685 9237 ne
rect 7685 9139 8039 9237
tri 8039 9139 8137 9237 sw
tri 8137 9139 8235 9237 ne
rect 8235 9139 8589 9237
tri 8589 9139 8687 9237 sw
tri 8687 9139 8785 9237 ne
rect 8785 9139 9139 9237
tri 9139 9139 9237 9237 sw
tri 9237 9139 9335 9237 ne
rect 9335 9139 9689 9237
tri 9689 9139 9787 9237 sw
tri 9787 9139 9885 9237 ne
rect 9885 9139 10239 9237
tri 10239 9139 10337 9237 sw
tri 10337 9139 10435 9237 ne
rect 10435 9139 10789 9237
tri 10789 9139 10887 9237 sw
tri 10887 9139 10985 9237 ne
rect 10985 9139 11339 9237
tri 11339 9139 11437 9237 sw
tri 11437 9139 11535 9237 ne
rect 11535 9139 11889 9237
tri 11889 9139 11987 9237 sw
tri 11987 9139 12085 9237 ne
rect 12085 9139 12439 9237
tri 12439 9139 12537 9237 sw
tri 12537 9139 12635 9237 ne
rect 12635 9139 12989 9237
tri 12989 9139 13087 9237 sw
tri 13087 9139 13185 9237 ne
rect 13185 9139 13539 9237
tri 13539 9139 13637 9237 sw
tri 13637 9139 13735 9237 ne
rect 13735 9139 14089 9237
tri 14089 9139 14187 9237 sw
tri 14187 9139 14285 9237 ne
rect 14285 9139 14639 9237
tri 14639 9139 14737 9237 sw
tri 14737 9139 14835 9237 ne
rect 14835 9139 15189 9237
tri 15189 9139 15287 9237 sw
tri 15287 9139 15385 9237 ne
rect 15385 9139 15739 9237
tri 15739 9139 15837 9237 sw
tri 15837 9139 15935 9237 ne
rect 15935 9139 16289 9237
tri 16289 9139 16387 9237 sw
tri 16387 9139 16485 9237 ne
rect 16485 9139 16839 9237
tri 16839 9139 16937 9237 sw
tri 16937 9139 17035 9237 ne
rect 17035 9139 17389 9237
tri 17389 9139 17487 9237 sw
tri 17487 9139 17585 9237 ne
rect 17585 9139 17939 9237
tri 17939 9139 18037 9237 sw
tri 18037 9139 18135 9237 ne
rect 18135 9139 18489 9237
tri 18489 9139 18587 9237 sw
tri 18587 9139 18685 9237 ne
rect 18685 9139 19039 9237
tri 19039 9139 19137 9237 sw
tri 19137 9139 19235 9237 ne
rect 19235 9139 19589 9237
tri 19589 9139 19687 9237 sw
rect -500 9135 437 9139
rect -500 9015 215 9135
rect 335 9041 437 9135
tri 437 9041 535 9139 sw
tri 535 9041 633 9139 ne
rect 633 9135 987 9139
rect 633 9041 765 9135
rect 335 9015 535 9041
rect -500 9011 535 9015
tri 535 9011 565 9041 sw
tri 633 9011 663 9041 ne
rect 663 9015 765 9041
rect 885 9041 987 9135
tri 987 9041 1085 9139 sw
tri 1085 9041 1183 9139 ne
rect 1183 9135 1537 9139
rect 1183 9041 1315 9135
rect 885 9015 1085 9041
rect 663 9011 1085 9015
tri 1085 9011 1115 9041 sw
tri 1183 9011 1213 9041 ne
rect 1213 9015 1315 9041
rect 1435 9041 1537 9135
tri 1537 9041 1635 9139 sw
tri 1635 9041 1733 9139 ne
rect 1733 9135 2087 9139
rect 1733 9041 1865 9135
rect 1435 9015 1635 9041
rect 1213 9011 1635 9015
tri 1635 9011 1665 9041 sw
tri 1733 9011 1763 9041 ne
rect 1763 9015 1865 9041
rect 1985 9041 2087 9135
tri 2087 9041 2185 9139 sw
tri 2185 9041 2283 9139 ne
rect 2283 9135 2637 9139
rect 2283 9041 2415 9135
rect 1985 9015 2185 9041
rect 1763 9011 2185 9015
tri 2185 9011 2215 9041 sw
tri 2283 9011 2313 9041 ne
rect 2313 9015 2415 9041
rect 2535 9041 2637 9135
tri 2637 9041 2735 9139 sw
tri 2735 9041 2833 9139 ne
rect 2833 9135 3187 9139
rect 2833 9041 2965 9135
rect 2535 9015 2735 9041
rect 2313 9011 2735 9015
tri 2735 9011 2765 9041 sw
tri 2833 9011 2863 9041 ne
rect 2863 9015 2965 9041
rect 3085 9041 3187 9135
tri 3187 9041 3285 9139 sw
tri 3285 9041 3383 9139 ne
rect 3383 9135 3737 9139
rect 3383 9041 3515 9135
rect 3085 9015 3285 9041
rect 2863 9011 3285 9015
tri 3285 9011 3315 9041 sw
tri 3383 9011 3413 9041 ne
rect 3413 9015 3515 9041
rect 3635 9041 3737 9135
tri 3737 9041 3835 9139 sw
tri 3835 9041 3933 9139 ne
rect 3933 9135 4287 9139
rect 3933 9041 4065 9135
rect 3635 9015 3835 9041
rect 3413 9011 3835 9015
tri 3835 9011 3865 9041 sw
tri 3933 9011 3963 9041 ne
rect 3963 9015 4065 9041
rect 4185 9041 4287 9135
tri 4287 9041 4385 9139 sw
tri 4385 9041 4483 9139 ne
rect 4483 9135 4837 9139
rect 4483 9041 4615 9135
rect 4185 9015 4385 9041
rect 3963 9011 4385 9015
tri 4385 9011 4415 9041 sw
tri 4483 9011 4513 9041 ne
rect 4513 9015 4615 9041
rect 4735 9041 4837 9135
tri 4837 9041 4935 9139 sw
tri 4935 9041 5033 9139 ne
rect 5033 9135 5387 9139
rect 5033 9041 5165 9135
rect 4735 9015 4935 9041
rect 4513 9011 4935 9015
tri 4935 9011 4965 9041 sw
tri 5033 9011 5063 9041 ne
rect 5063 9015 5165 9041
rect 5285 9041 5387 9135
tri 5387 9041 5485 9139 sw
tri 5485 9041 5583 9139 ne
rect 5583 9135 5937 9139
rect 5583 9041 5715 9135
rect 5285 9015 5485 9041
rect 5063 9011 5485 9015
tri 5485 9011 5515 9041 sw
tri 5583 9011 5613 9041 ne
rect 5613 9015 5715 9041
rect 5835 9041 5937 9135
tri 5937 9041 6035 9139 sw
tri 6035 9041 6133 9139 ne
rect 6133 9135 6487 9139
rect 6133 9041 6265 9135
rect 5835 9015 6035 9041
rect 5613 9011 6035 9015
tri 6035 9011 6065 9041 sw
tri 6133 9011 6163 9041 ne
rect 6163 9015 6265 9041
rect 6385 9041 6487 9135
tri 6487 9041 6585 9139 sw
tri 6585 9041 6683 9139 ne
rect 6683 9135 7037 9139
rect 6683 9041 6815 9135
rect 6385 9015 6585 9041
rect 6163 9011 6585 9015
tri 6585 9011 6615 9041 sw
tri 6683 9011 6713 9041 ne
rect 6713 9015 6815 9041
rect 6935 9041 7037 9135
tri 7037 9041 7135 9139 sw
tri 7135 9041 7233 9139 ne
rect 7233 9135 7587 9139
rect 7233 9041 7365 9135
rect 6935 9015 7135 9041
rect 6713 9011 7135 9015
tri 7135 9011 7165 9041 sw
tri 7233 9011 7263 9041 ne
rect 7263 9015 7365 9041
rect 7485 9041 7587 9135
tri 7587 9041 7685 9139 sw
tri 7685 9041 7783 9139 ne
rect 7783 9135 8137 9139
rect 7783 9041 7915 9135
rect 7485 9015 7685 9041
rect 7263 9011 7685 9015
tri 7685 9011 7715 9041 sw
tri 7783 9011 7813 9041 ne
rect 7813 9015 7915 9041
rect 8035 9041 8137 9135
tri 8137 9041 8235 9139 sw
tri 8235 9041 8333 9139 ne
rect 8333 9135 8687 9139
rect 8333 9041 8465 9135
rect 8035 9015 8235 9041
rect 7813 9011 8235 9015
tri 8235 9011 8265 9041 sw
tri 8333 9011 8363 9041 ne
rect 8363 9015 8465 9041
rect 8585 9041 8687 9135
tri 8687 9041 8785 9139 sw
tri 8785 9041 8883 9139 ne
rect 8883 9135 9237 9139
rect 8883 9041 9015 9135
rect 8585 9015 8785 9041
rect 8363 9011 8785 9015
tri 8785 9011 8815 9041 sw
tri 8883 9011 8913 9041 ne
rect 8913 9015 9015 9041
rect 9135 9041 9237 9135
tri 9237 9041 9335 9139 sw
tri 9335 9041 9433 9139 ne
rect 9433 9135 9787 9139
rect 9433 9041 9565 9135
rect 9135 9015 9335 9041
rect 8913 9011 9335 9015
tri 9335 9011 9365 9041 sw
tri 9433 9011 9463 9041 ne
rect 9463 9015 9565 9041
rect 9685 9041 9787 9135
tri 9787 9041 9885 9139 sw
tri 9885 9041 9983 9139 ne
rect 9983 9135 10337 9139
rect 9983 9041 10115 9135
rect 9685 9015 9885 9041
rect 9463 9011 9885 9015
tri 9885 9011 9915 9041 sw
tri 9983 9011 10013 9041 ne
rect 10013 9015 10115 9041
rect 10235 9041 10337 9135
tri 10337 9041 10435 9139 sw
tri 10435 9041 10533 9139 ne
rect 10533 9135 10887 9139
rect 10533 9041 10665 9135
rect 10235 9015 10435 9041
rect 10013 9011 10435 9015
tri 10435 9011 10465 9041 sw
tri 10533 9011 10563 9041 ne
rect 10563 9015 10665 9041
rect 10785 9041 10887 9135
tri 10887 9041 10985 9139 sw
tri 10985 9041 11083 9139 ne
rect 11083 9135 11437 9139
rect 11083 9041 11215 9135
rect 10785 9015 10985 9041
rect 10563 9011 10985 9015
tri 10985 9011 11015 9041 sw
tri 11083 9011 11113 9041 ne
rect 11113 9015 11215 9041
rect 11335 9041 11437 9135
tri 11437 9041 11535 9139 sw
tri 11535 9041 11633 9139 ne
rect 11633 9135 11987 9139
rect 11633 9041 11765 9135
rect 11335 9015 11535 9041
rect 11113 9011 11535 9015
tri 11535 9011 11565 9041 sw
tri 11633 9011 11663 9041 ne
rect 11663 9015 11765 9041
rect 11885 9041 11987 9135
tri 11987 9041 12085 9139 sw
tri 12085 9041 12183 9139 ne
rect 12183 9135 12537 9139
rect 12183 9041 12315 9135
rect 11885 9015 12085 9041
rect 11663 9011 12085 9015
tri 12085 9011 12115 9041 sw
tri 12183 9011 12213 9041 ne
rect 12213 9015 12315 9041
rect 12435 9041 12537 9135
tri 12537 9041 12635 9139 sw
tri 12635 9041 12733 9139 ne
rect 12733 9135 13087 9139
rect 12733 9041 12865 9135
rect 12435 9015 12635 9041
rect 12213 9011 12635 9015
tri 12635 9011 12665 9041 sw
tri 12733 9011 12763 9041 ne
rect 12763 9015 12865 9041
rect 12985 9041 13087 9135
tri 13087 9041 13185 9139 sw
tri 13185 9041 13283 9139 ne
rect 13283 9135 13637 9139
rect 13283 9041 13415 9135
rect 12985 9015 13185 9041
rect 12763 9011 13185 9015
tri 13185 9011 13215 9041 sw
tri 13283 9011 13313 9041 ne
rect 13313 9015 13415 9041
rect 13535 9041 13637 9135
tri 13637 9041 13735 9139 sw
tri 13735 9041 13833 9139 ne
rect 13833 9135 14187 9139
rect 13833 9041 13965 9135
rect 13535 9015 13735 9041
rect 13313 9011 13735 9015
tri 13735 9011 13765 9041 sw
tri 13833 9011 13863 9041 ne
rect 13863 9015 13965 9041
rect 14085 9041 14187 9135
tri 14187 9041 14285 9139 sw
tri 14285 9041 14383 9139 ne
rect 14383 9135 14737 9139
rect 14383 9041 14515 9135
rect 14085 9015 14285 9041
rect 13863 9011 14285 9015
tri 14285 9011 14315 9041 sw
tri 14383 9011 14413 9041 ne
rect 14413 9015 14515 9041
rect 14635 9041 14737 9135
tri 14737 9041 14835 9139 sw
tri 14835 9041 14933 9139 ne
rect 14933 9135 15287 9139
rect 14933 9041 15065 9135
rect 14635 9015 14835 9041
rect 14413 9011 14835 9015
tri 14835 9011 14865 9041 sw
tri 14933 9011 14963 9041 ne
rect 14963 9015 15065 9041
rect 15185 9041 15287 9135
tri 15287 9041 15385 9139 sw
tri 15385 9041 15483 9139 ne
rect 15483 9135 15837 9139
rect 15483 9041 15615 9135
rect 15185 9015 15385 9041
rect 14963 9011 15385 9015
tri 15385 9011 15415 9041 sw
tri 15483 9011 15513 9041 ne
rect 15513 9015 15615 9041
rect 15735 9041 15837 9135
tri 15837 9041 15935 9139 sw
tri 15935 9041 16033 9139 ne
rect 16033 9135 16387 9139
rect 16033 9041 16165 9135
rect 15735 9015 15935 9041
rect 15513 9011 15935 9015
tri 15935 9011 15965 9041 sw
tri 16033 9011 16063 9041 ne
rect 16063 9015 16165 9041
rect 16285 9041 16387 9135
tri 16387 9041 16485 9139 sw
tri 16485 9041 16583 9139 ne
rect 16583 9135 16937 9139
rect 16583 9041 16715 9135
rect 16285 9015 16485 9041
rect 16063 9011 16485 9015
tri 16485 9011 16515 9041 sw
tri 16583 9011 16613 9041 ne
rect 16613 9015 16715 9041
rect 16835 9041 16937 9135
tri 16937 9041 17035 9139 sw
tri 17035 9041 17133 9139 ne
rect 17133 9135 17487 9139
rect 17133 9041 17265 9135
rect 16835 9015 17035 9041
rect 16613 9011 17035 9015
tri 17035 9011 17065 9041 sw
tri 17133 9011 17163 9041 ne
rect 17163 9015 17265 9041
rect 17385 9041 17487 9135
tri 17487 9041 17585 9139 sw
tri 17585 9041 17683 9139 ne
rect 17683 9135 18037 9139
rect 17683 9041 17815 9135
rect 17385 9015 17585 9041
rect 17163 9011 17585 9015
tri 17585 9011 17615 9041 sw
tri 17683 9011 17713 9041 ne
rect 17713 9015 17815 9041
rect 17935 9041 18037 9135
tri 18037 9041 18135 9139 sw
tri 18135 9041 18233 9139 ne
rect 18233 9135 18587 9139
rect 18233 9041 18365 9135
rect 17935 9015 18135 9041
rect 17713 9011 18135 9015
tri 18135 9011 18165 9041 sw
tri 18233 9011 18263 9041 ne
rect 18263 9015 18365 9041
rect 18485 9041 18587 9135
tri 18587 9041 18685 9139 sw
tri 18685 9041 18783 9139 ne
rect 18783 9135 19137 9139
rect 18783 9041 18915 9135
rect 18485 9015 18685 9041
rect 18263 9011 18685 9015
tri 18685 9011 18715 9041 sw
tri 18783 9011 18813 9041 ne
rect 18813 9015 18915 9041
rect 19035 9041 19137 9135
tri 19137 9041 19235 9139 sw
tri 19235 9041 19333 9139 ne
rect 19333 9135 20300 9139
rect 19333 9041 19465 9135
rect 19035 9015 19235 9041
rect 18813 9011 19235 9015
tri 19235 9011 19265 9041 sw
tri 19333 9011 19363 9041 ne
rect 19363 9015 19465 9041
rect 19585 9015 20300 9135
rect 19363 9011 20300 9015
tri 113 8913 211 9011 ne
rect 211 8913 565 9011
tri 565 8913 663 9011 sw
tri 663 8913 761 9011 ne
rect 761 8913 1115 9011
tri 1115 8913 1213 9011 sw
tri 1213 8913 1311 9011 ne
rect 1311 8913 1665 9011
tri 1665 8913 1763 9011 sw
tri 1763 8913 1861 9011 ne
rect 1861 8913 2215 9011
tri 2215 8913 2313 9011 sw
tri 2313 8913 2411 9011 ne
rect 2411 8913 2765 9011
tri 2765 8913 2863 9011 sw
tri 2863 8913 2961 9011 ne
rect 2961 8913 3315 9011
tri 3315 8913 3413 9011 sw
tri 3413 8913 3511 9011 ne
rect 3511 8913 3865 9011
tri 3865 8913 3963 9011 sw
tri 3963 8913 4061 9011 ne
rect 4061 8913 4415 9011
tri 4415 8913 4513 9011 sw
tri 4513 8913 4611 9011 ne
rect 4611 8913 4965 9011
tri 4965 8913 5063 9011 sw
tri 5063 8913 5161 9011 ne
rect 5161 8913 5515 9011
tri 5515 8913 5613 9011 sw
tri 5613 8913 5711 9011 ne
rect 5711 8913 6065 9011
tri 6065 8913 6163 9011 sw
tri 6163 8913 6261 9011 ne
rect 6261 8913 6615 9011
tri 6615 8913 6713 9011 sw
tri 6713 8913 6811 9011 ne
rect 6811 8913 7165 9011
tri 7165 8913 7263 9011 sw
tri 7263 8913 7361 9011 ne
rect 7361 8913 7715 9011
tri 7715 8913 7813 9011 sw
tri 7813 8913 7911 9011 ne
rect 7911 8913 8265 9011
tri 8265 8913 8363 9011 sw
tri 8363 8913 8461 9011 ne
rect 8461 8913 8815 9011
tri 8815 8913 8913 9011 sw
tri 8913 8913 9011 9011 ne
rect 9011 8913 9365 9011
tri 9365 8913 9463 9011 sw
tri 9463 8913 9561 9011 ne
rect 9561 8913 9915 9011
tri 9915 8913 10013 9011 sw
tri 10013 8913 10111 9011 ne
rect 10111 8913 10465 9011
tri 10465 8913 10563 9011 sw
tri 10563 8913 10661 9011 ne
rect 10661 8913 11015 9011
tri 11015 8913 11113 9011 sw
tri 11113 8913 11211 9011 ne
rect 11211 8913 11565 9011
tri 11565 8913 11663 9011 sw
tri 11663 8913 11761 9011 ne
rect 11761 8913 12115 9011
tri 12115 8913 12213 9011 sw
tri 12213 8913 12311 9011 ne
rect 12311 8913 12665 9011
tri 12665 8913 12763 9011 sw
tri 12763 8913 12861 9011 ne
rect 12861 8913 13215 9011
tri 13215 8913 13313 9011 sw
tri 13313 8913 13411 9011 ne
rect 13411 8913 13765 9011
tri 13765 8913 13863 9011 sw
tri 13863 8913 13961 9011 ne
rect 13961 8913 14315 9011
tri 14315 8913 14413 9011 sw
tri 14413 8913 14511 9011 ne
rect 14511 8913 14865 9011
tri 14865 8913 14963 9011 sw
tri 14963 8913 15061 9011 ne
rect 15061 8913 15415 9011
tri 15415 8913 15513 9011 sw
tri 15513 8913 15611 9011 ne
rect 15611 8913 15965 9011
tri 15965 8913 16063 9011 sw
tri 16063 8913 16161 9011 ne
rect 16161 8913 16515 9011
tri 16515 8913 16613 9011 sw
tri 16613 8913 16711 9011 ne
rect 16711 8913 17065 9011
tri 17065 8913 17163 9011 sw
tri 17163 8913 17261 9011 ne
rect 17261 8913 17615 9011
tri 17615 8913 17713 9011 sw
tri 17713 8913 17811 9011 ne
rect 17811 8913 18165 9011
tri 18165 8913 18263 9011 sw
tri 18263 8913 18361 9011 ne
rect 18361 8913 18715 9011
tri 18715 8913 18813 9011 sw
tri 18813 8913 18911 9011 ne
rect 18911 8913 19265 9011
tri 19265 8913 19363 9011 sw
tri 19363 8913 19461 9011 ne
rect 19461 8913 20300 9011
rect -2000 8883 113 8913
tri 113 8883 143 8913 sw
tri 211 8883 241 8913 ne
rect 241 8883 663 8913
tri 663 8883 693 8913 sw
tri 761 8883 791 8913 ne
rect 791 8883 1213 8913
tri 1213 8883 1243 8913 sw
tri 1311 8883 1341 8913 ne
rect 1341 8883 1763 8913
tri 1763 8883 1793 8913 sw
tri 1861 8883 1891 8913 ne
rect 1891 8883 2313 8913
tri 2313 8883 2343 8913 sw
tri 2411 8883 2441 8913 ne
rect 2441 8883 2863 8913
tri 2863 8883 2893 8913 sw
tri 2961 8883 2991 8913 ne
rect 2991 8883 3413 8913
tri 3413 8883 3443 8913 sw
tri 3511 8883 3541 8913 ne
rect 3541 8883 3963 8913
tri 3963 8883 3993 8913 sw
tri 4061 8883 4091 8913 ne
rect 4091 8883 4513 8913
tri 4513 8883 4543 8913 sw
tri 4611 8883 4641 8913 ne
rect 4641 8883 5063 8913
tri 5063 8883 5093 8913 sw
tri 5161 8883 5191 8913 ne
rect 5191 8883 5613 8913
tri 5613 8883 5643 8913 sw
tri 5711 8883 5741 8913 ne
rect 5741 8883 6163 8913
tri 6163 8883 6193 8913 sw
tri 6261 8883 6291 8913 ne
rect 6291 8883 6713 8913
tri 6713 8883 6743 8913 sw
tri 6811 8883 6841 8913 ne
rect 6841 8883 7263 8913
tri 7263 8883 7293 8913 sw
tri 7361 8883 7391 8913 ne
rect 7391 8883 7813 8913
tri 7813 8883 7843 8913 sw
tri 7911 8883 7941 8913 ne
rect 7941 8883 8363 8913
tri 8363 8883 8393 8913 sw
tri 8461 8883 8491 8913 ne
rect 8491 8883 8913 8913
tri 8913 8883 8943 8913 sw
tri 9011 8883 9041 8913 ne
rect 9041 8883 9463 8913
tri 9463 8883 9493 8913 sw
tri 9561 8883 9591 8913 ne
rect 9591 8883 10013 8913
tri 10013 8883 10043 8913 sw
tri 10111 8883 10141 8913 ne
rect 10141 8883 10563 8913
tri 10563 8883 10593 8913 sw
tri 10661 8883 10691 8913 ne
rect 10691 8883 11113 8913
tri 11113 8883 11143 8913 sw
tri 11211 8883 11241 8913 ne
rect 11241 8883 11663 8913
tri 11663 8883 11693 8913 sw
tri 11761 8883 11791 8913 ne
rect 11791 8883 12213 8913
tri 12213 8883 12243 8913 sw
tri 12311 8883 12341 8913 ne
rect 12341 8883 12763 8913
tri 12763 8883 12793 8913 sw
tri 12861 8883 12891 8913 ne
rect 12891 8883 13313 8913
tri 13313 8883 13343 8913 sw
tri 13411 8883 13441 8913 ne
rect 13441 8883 13863 8913
tri 13863 8883 13893 8913 sw
tri 13961 8883 13991 8913 ne
rect 13991 8883 14413 8913
tri 14413 8883 14443 8913 sw
tri 14511 8883 14541 8913 ne
rect 14541 8883 14963 8913
tri 14963 8883 14993 8913 sw
tri 15061 8883 15091 8913 ne
rect 15091 8883 15513 8913
tri 15513 8883 15543 8913 sw
tri 15611 8883 15641 8913 ne
rect 15641 8883 16063 8913
tri 16063 8883 16093 8913 sw
tri 16161 8883 16191 8913 ne
rect 16191 8883 16613 8913
tri 16613 8883 16643 8913 sw
tri 16711 8883 16741 8913 ne
rect 16741 8883 17163 8913
tri 17163 8883 17193 8913 sw
tri 17261 8883 17291 8913 ne
rect 17291 8883 17713 8913
tri 17713 8883 17743 8913 sw
tri 17811 8883 17841 8913 ne
rect 17841 8883 18263 8913
tri 18263 8883 18293 8913 sw
tri 18361 8883 18391 8913 ne
rect 18391 8883 18813 8913
tri 18813 8883 18843 8913 sw
tri 18911 8883 18941 8913 ne
rect 18941 8883 19363 8913
tri 19363 8883 19393 8913 sw
tri 19461 8883 19491 8913 ne
rect 19491 8883 20300 8913
rect -2000 8785 143 8883
tri 143 8785 241 8883 sw
tri 241 8785 339 8883 ne
rect 339 8785 693 8883
tri 693 8785 791 8883 sw
tri 791 8785 889 8883 ne
rect 889 8785 1243 8883
tri 1243 8785 1341 8883 sw
tri 1341 8785 1439 8883 ne
rect 1439 8785 1793 8883
tri 1793 8785 1891 8883 sw
tri 1891 8785 1989 8883 ne
rect 1989 8785 2343 8883
tri 2343 8785 2441 8883 sw
tri 2441 8785 2539 8883 ne
rect 2539 8785 2893 8883
tri 2893 8785 2991 8883 sw
tri 2991 8785 3089 8883 ne
rect 3089 8785 3443 8883
tri 3443 8785 3541 8883 sw
tri 3541 8785 3639 8883 ne
rect 3639 8785 3993 8883
tri 3993 8785 4091 8883 sw
tri 4091 8785 4189 8883 ne
rect 4189 8785 4543 8883
tri 4543 8785 4641 8883 sw
tri 4641 8785 4739 8883 ne
rect 4739 8785 5093 8883
tri 5093 8785 5191 8883 sw
tri 5191 8785 5289 8883 ne
rect 5289 8785 5643 8883
tri 5643 8785 5741 8883 sw
tri 5741 8785 5839 8883 ne
rect 5839 8785 6193 8883
tri 6193 8785 6291 8883 sw
tri 6291 8785 6389 8883 ne
rect 6389 8785 6743 8883
tri 6743 8785 6841 8883 sw
tri 6841 8785 6939 8883 ne
rect 6939 8785 7293 8883
tri 7293 8785 7391 8883 sw
tri 7391 8785 7489 8883 ne
rect 7489 8785 7843 8883
tri 7843 8785 7941 8883 sw
tri 7941 8785 8039 8883 ne
rect 8039 8785 8393 8883
tri 8393 8785 8491 8883 sw
tri 8491 8785 8589 8883 ne
rect 8589 8785 8943 8883
tri 8943 8785 9041 8883 sw
tri 9041 8785 9139 8883 ne
rect 9139 8785 9493 8883
tri 9493 8785 9591 8883 sw
tri 9591 8785 9689 8883 ne
rect 9689 8785 10043 8883
tri 10043 8785 10141 8883 sw
tri 10141 8785 10239 8883 ne
rect 10239 8785 10593 8883
tri 10593 8785 10691 8883 sw
tri 10691 8785 10789 8883 ne
rect 10789 8785 11143 8883
tri 11143 8785 11241 8883 sw
tri 11241 8785 11339 8883 ne
rect 11339 8785 11693 8883
tri 11693 8785 11791 8883 sw
tri 11791 8785 11889 8883 ne
rect 11889 8785 12243 8883
tri 12243 8785 12341 8883 sw
tri 12341 8785 12439 8883 ne
rect 12439 8785 12793 8883
tri 12793 8785 12891 8883 sw
tri 12891 8785 12989 8883 ne
rect 12989 8785 13343 8883
tri 13343 8785 13441 8883 sw
tri 13441 8785 13539 8883 ne
rect 13539 8785 13893 8883
tri 13893 8785 13991 8883 sw
tri 13991 8785 14089 8883 ne
rect 14089 8785 14443 8883
tri 14443 8785 14541 8883 sw
tri 14541 8785 14639 8883 ne
rect 14639 8785 14993 8883
tri 14993 8785 15091 8883 sw
tri 15091 8785 15189 8883 ne
rect 15189 8785 15543 8883
tri 15543 8785 15641 8883 sw
tri 15641 8785 15739 8883 ne
rect 15739 8785 16093 8883
tri 16093 8785 16191 8883 sw
tri 16191 8785 16289 8883 ne
rect 16289 8785 16643 8883
tri 16643 8785 16741 8883 sw
tri 16741 8785 16839 8883 ne
rect 16839 8785 17193 8883
tri 17193 8785 17291 8883 sw
tri 17291 8785 17389 8883 ne
rect 17389 8785 17743 8883
tri 17743 8785 17841 8883 sw
tri 17841 8785 17939 8883 ne
rect 17939 8785 18293 8883
tri 18293 8785 18391 8883 sw
tri 18391 8785 18489 8883 ne
rect 18489 8785 18843 8883
tri 18843 8785 18941 8883 sw
tri 18941 8785 19039 8883 ne
rect 19039 8785 19393 8883
tri 19393 8785 19491 8883 sw
tri 19491 8785 19589 8883 ne
rect 19589 8785 20300 8883
rect -2000 8687 241 8785
tri 241 8687 339 8785 sw
tri 339 8687 437 8785 ne
rect 437 8687 791 8785
tri 791 8687 889 8785 sw
tri 889 8687 987 8785 ne
rect 987 8687 1341 8785
tri 1341 8687 1439 8785 sw
tri 1439 8687 1537 8785 ne
rect 1537 8687 1891 8785
tri 1891 8687 1989 8785 sw
tri 1989 8687 2087 8785 ne
rect 2087 8687 2441 8785
tri 2441 8687 2539 8785 sw
tri 2539 8687 2637 8785 ne
rect 2637 8687 2991 8785
tri 2991 8687 3089 8785 sw
tri 3089 8687 3187 8785 ne
rect 3187 8687 3541 8785
tri 3541 8687 3639 8785 sw
tri 3639 8687 3737 8785 ne
rect 3737 8687 4091 8785
tri 4091 8687 4189 8785 sw
tri 4189 8687 4287 8785 ne
rect 4287 8687 4641 8785
tri 4641 8687 4739 8785 sw
tri 4739 8687 4837 8785 ne
rect 4837 8687 5191 8785
tri 5191 8687 5289 8785 sw
tri 5289 8687 5387 8785 ne
rect 5387 8687 5741 8785
tri 5741 8687 5839 8785 sw
tri 5839 8687 5937 8785 ne
rect 5937 8687 6291 8785
tri 6291 8687 6389 8785 sw
tri 6389 8687 6487 8785 ne
rect 6487 8687 6841 8785
tri 6841 8687 6939 8785 sw
tri 6939 8687 7037 8785 ne
rect 7037 8687 7391 8785
tri 7391 8687 7489 8785 sw
tri 7489 8687 7587 8785 ne
rect 7587 8687 7941 8785
tri 7941 8687 8039 8785 sw
tri 8039 8687 8137 8785 ne
rect 8137 8687 8491 8785
tri 8491 8687 8589 8785 sw
tri 8589 8687 8687 8785 ne
rect 8687 8687 9041 8785
tri 9041 8687 9139 8785 sw
tri 9139 8687 9237 8785 ne
rect 9237 8687 9591 8785
tri 9591 8687 9689 8785 sw
tri 9689 8687 9787 8785 ne
rect 9787 8687 10141 8785
tri 10141 8687 10239 8785 sw
tri 10239 8687 10337 8785 ne
rect 10337 8687 10691 8785
tri 10691 8687 10789 8785 sw
tri 10789 8687 10887 8785 ne
rect 10887 8687 11241 8785
tri 11241 8687 11339 8785 sw
tri 11339 8687 11437 8785 ne
rect 11437 8687 11791 8785
tri 11791 8687 11889 8785 sw
tri 11889 8687 11987 8785 ne
rect 11987 8687 12341 8785
tri 12341 8687 12439 8785 sw
tri 12439 8687 12537 8785 ne
rect 12537 8687 12891 8785
tri 12891 8687 12989 8785 sw
tri 12989 8687 13087 8785 ne
rect 13087 8687 13441 8785
tri 13441 8687 13539 8785 sw
tri 13539 8687 13637 8785 ne
rect 13637 8687 13991 8785
tri 13991 8687 14089 8785 sw
tri 14089 8687 14187 8785 ne
rect 14187 8687 14541 8785
tri 14541 8687 14639 8785 sw
tri 14639 8687 14737 8785 ne
rect 14737 8687 15091 8785
tri 15091 8687 15189 8785 sw
tri 15189 8687 15287 8785 ne
rect 15287 8687 15641 8785
tri 15641 8687 15739 8785 sw
tri 15739 8687 15837 8785 ne
rect 15837 8687 16191 8785
tri 16191 8687 16289 8785 sw
tri 16289 8687 16387 8785 ne
rect 16387 8687 16741 8785
tri 16741 8687 16839 8785 sw
tri 16839 8687 16937 8785 ne
rect 16937 8687 17291 8785
tri 17291 8687 17389 8785 sw
tri 17389 8687 17487 8785 ne
rect 17487 8687 17841 8785
tri 17841 8687 17939 8785 sw
tri 17939 8687 18037 8785 ne
rect 18037 8687 18391 8785
tri 18391 8687 18489 8785 sw
tri 18489 8687 18587 8785 ne
rect 18587 8687 18941 8785
tri 18941 8687 19039 8785 sw
tri 19039 8687 19137 8785 ne
rect 19137 8687 19491 8785
tri 19491 8687 19589 8785 sw
tri 19589 8687 19687 8785 ne
rect 19687 8687 20300 8785
rect -2000 8589 339 8687
tri 339 8589 437 8687 sw
tri 437 8589 535 8687 ne
rect 535 8589 889 8687
tri 889 8589 987 8687 sw
tri 987 8589 1085 8687 ne
rect 1085 8589 1439 8687
tri 1439 8589 1537 8687 sw
tri 1537 8589 1635 8687 ne
rect 1635 8589 1989 8687
tri 1989 8589 2087 8687 sw
tri 2087 8589 2185 8687 ne
rect 2185 8589 2539 8687
tri 2539 8589 2637 8687 sw
tri 2637 8589 2735 8687 ne
rect 2735 8589 3089 8687
tri 3089 8589 3187 8687 sw
tri 3187 8589 3285 8687 ne
rect 3285 8589 3639 8687
tri 3639 8589 3737 8687 sw
tri 3737 8589 3835 8687 ne
rect 3835 8589 4189 8687
tri 4189 8589 4287 8687 sw
tri 4287 8589 4385 8687 ne
rect 4385 8589 4739 8687
tri 4739 8589 4837 8687 sw
tri 4837 8589 4935 8687 ne
rect 4935 8589 5289 8687
tri 5289 8589 5387 8687 sw
tri 5387 8589 5485 8687 ne
rect 5485 8589 5839 8687
tri 5839 8589 5937 8687 sw
tri 5937 8589 6035 8687 ne
rect 6035 8589 6389 8687
tri 6389 8589 6487 8687 sw
tri 6487 8589 6585 8687 ne
rect 6585 8589 6939 8687
tri 6939 8589 7037 8687 sw
tri 7037 8589 7135 8687 ne
rect 7135 8589 7489 8687
tri 7489 8589 7587 8687 sw
tri 7587 8589 7685 8687 ne
rect 7685 8589 8039 8687
tri 8039 8589 8137 8687 sw
tri 8137 8589 8235 8687 ne
rect 8235 8589 8589 8687
tri 8589 8589 8687 8687 sw
tri 8687 8589 8785 8687 ne
rect 8785 8589 9139 8687
tri 9139 8589 9237 8687 sw
tri 9237 8589 9335 8687 ne
rect 9335 8589 9689 8687
tri 9689 8589 9787 8687 sw
tri 9787 8589 9885 8687 ne
rect 9885 8589 10239 8687
tri 10239 8589 10337 8687 sw
tri 10337 8589 10435 8687 ne
rect 10435 8589 10789 8687
tri 10789 8589 10887 8687 sw
tri 10887 8589 10985 8687 ne
rect 10985 8589 11339 8687
tri 11339 8589 11437 8687 sw
tri 11437 8589 11535 8687 ne
rect 11535 8589 11889 8687
tri 11889 8589 11987 8687 sw
tri 11987 8589 12085 8687 ne
rect 12085 8589 12439 8687
tri 12439 8589 12537 8687 sw
tri 12537 8589 12635 8687 ne
rect 12635 8589 12989 8687
tri 12989 8589 13087 8687 sw
tri 13087 8589 13185 8687 ne
rect 13185 8589 13539 8687
tri 13539 8589 13637 8687 sw
tri 13637 8589 13735 8687 ne
rect 13735 8589 14089 8687
tri 14089 8589 14187 8687 sw
tri 14187 8589 14285 8687 ne
rect 14285 8589 14639 8687
tri 14639 8589 14737 8687 sw
tri 14737 8589 14835 8687 ne
rect 14835 8589 15189 8687
tri 15189 8589 15287 8687 sw
tri 15287 8589 15385 8687 ne
rect 15385 8589 15739 8687
tri 15739 8589 15837 8687 sw
tri 15837 8589 15935 8687 ne
rect 15935 8589 16289 8687
tri 16289 8589 16387 8687 sw
tri 16387 8589 16485 8687 ne
rect 16485 8589 16839 8687
tri 16839 8589 16937 8687 sw
tri 16937 8589 17035 8687 ne
rect 17035 8589 17389 8687
tri 17389 8589 17487 8687 sw
tri 17487 8589 17585 8687 ne
rect 17585 8589 17939 8687
tri 17939 8589 18037 8687 sw
tri 18037 8589 18135 8687 ne
rect 18135 8589 18489 8687
tri 18489 8589 18587 8687 sw
tri 18587 8589 18685 8687 ne
rect 18685 8589 19039 8687
tri 19039 8589 19137 8687 sw
tri 19137 8589 19235 8687 ne
rect 19235 8589 19589 8687
tri 19589 8589 19687 8687 sw
rect 20800 8589 21800 9237
rect -2000 8585 437 8589
rect -2000 8465 215 8585
rect 335 8491 437 8585
tri 437 8491 535 8589 sw
tri 535 8491 633 8589 ne
rect 633 8585 987 8589
rect 633 8491 765 8585
rect 335 8465 535 8491
rect -2000 8461 535 8465
rect -2000 7813 -1000 8461
tri 113 8363 211 8461 ne
rect 211 8413 535 8461
tri 535 8413 613 8491 sw
tri 633 8413 711 8491 ne
rect 711 8465 765 8491
rect 885 8491 987 8585
tri 987 8491 1085 8589 sw
tri 1085 8491 1183 8589 ne
rect 1183 8585 1537 8589
rect 1183 8491 1315 8585
rect 885 8465 1085 8491
rect 711 8413 1085 8465
tri 1085 8413 1163 8491 sw
tri 1183 8413 1261 8491 ne
rect 1261 8465 1315 8491
rect 1435 8491 1537 8585
tri 1537 8491 1635 8589 sw
tri 1635 8491 1733 8589 ne
rect 1733 8585 2087 8589
rect 1733 8491 1865 8585
rect 1435 8465 1635 8491
rect 1261 8413 1635 8465
tri 1635 8413 1713 8491 sw
tri 1733 8413 1811 8491 ne
rect 1811 8465 1865 8491
rect 1985 8491 2087 8585
tri 2087 8491 2185 8589 sw
tri 2185 8491 2283 8589 ne
rect 2283 8585 2637 8589
rect 2283 8491 2415 8585
rect 1985 8465 2185 8491
rect 1811 8413 2185 8465
tri 2185 8413 2263 8491 sw
tri 2283 8413 2361 8491 ne
rect 2361 8465 2415 8491
rect 2535 8491 2637 8585
tri 2637 8491 2735 8589 sw
tri 2735 8491 2833 8589 ne
rect 2833 8585 3187 8589
rect 2833 8491 2965 8585
rect 2535 8465 2735 8491
rect 2361 8413 2735 8465
tri 2735 8413 2813 8491 sw
tri 2833 8413 2911 8491 ne
rect 2911 8465 2965 8491
rect 3085 8491 3187 8585
tri 3187 8491 3285 8589 sw
tri 3285 8491 3383 8589 ne
rect 3383 8585 3737 8589
rect 3383 8491 3515 8585
rect 3085 8465 3285 8491
rect 2911 8413 3285 8465
tri 3285 8413 3363 8491 sw
tri 3383 8413 3461 8491 ne
rect 3461 8465 3515 8491
rect 3635 8491 3737 8585
tri 3737 8491 3835 8589 sw
tri 3835 8491 3933 8589 ne
rect 3933 8585 4287 8589
rect 3933 8491 4065 8585
rect 3635 8465 3835 8491
rect 3461 8413 3835 8465
tri 3835 8413 3913 8491 sw
tri 3933 8413 4011 8491 ne
rect 4011 8465 4065 8491
rect 4185 8491 4287 8585
tri 4287 8491 4385 8589 sw
tri 4385 8491 4483 8589 ne
rect 4483 8585 4837 8589
rect 4483 8491 4615 8585
rect 4185 8465 4385 8491
rect 4011 8413 4385 8465
tri 4385 8413 4463 8491 sw
tri 4483 8413 4561 8491 ne
rect 4561 8465 4615 8491
rect 4735 8491 4837 8585
tri 4837 8491 4935 8589 sw
tri 4935 8491 5033 8589 ne
rect 5033 8585 5387 8589
rect 5033 8491 5165 8585
rect 4735 8465 4935 8491
rect 4561 8413 4935 8465
tri 4935 8413 5013 8491 sw
tri 5033 8413 5111 8491 ne
rect 5111 8465 5165 8491
rect 5285 8491 5387 8585
tri 5387 8491 5485 8589 sw
tri 5485 8491 5583 8589 ne
rect 5583 8585 5937 8589
rect 5583 8491 5715 8585
rect 5285 8465 5485 8491
rect 5111 8413 5485 8465
tri 5485 8413 5563 8491 sw
tri 5583 8413 5661 8491 ne
rect 5661 8465 5715 8491
rect 5835 8491 5937 8585
tri 5937 8491 6035 8589 sw
tri 6035 8491 6133 8589 ne
rect 6133 8585 6487 8589
rect 6133 8491 6265 8585
rect 5835 8465 6035 8491
rect 5661 8413 6035 8465
tri 6035 8413 6113 8491 sw
tri 6133 8413 6211 8491 ne
rect 6211 8465 6265 8491
rect 6385 8491 6487 8585
tri 6487 8491 6585 8589 sw
tri 6585 8491 6683 8589 ne
rect 6683 8585 7037 8589
rect 6683 8491 6815 8585
rect 6385 8465 6585 8491
rect 6211 8413 6585 8465
tri 6585 8413 6663 8491 sw
tri 6683 8413 6761 8491 ne
rect 6761 8465 6815 8491
rect 6935 8491 7037 8585
tri 7037 8491 7135 8589 sw
tri 7135 8491 7233 8589 ne
rect 7233 8585 7587 8589
rect 7233 8491 7365 8585
rect 6935 8465 7135 8491
rect 6761 8413 7135 8465
tri 7135 8413 7213 8491 sw
tri 7233 8413 7311 8491 ne
rect 7311 8465 7365 8491
rect 7485 8491 7587 8585
tri 7587 8491 7685 8589 sw
tri 7685 8491 7783 8589 ne
rect 7783 8585 8137 8589
rect 7783 8491 7915 8585
rect 7485 8465 7685 8491
rect 7311 8413 7685 8465
tri 7685 8413 7763 8491 sw
tri 7783 8413 7861 8491 ne
rect 7861 8465 7915 8491
rect 8035 8491 8137 8585
tri 8137 8491 8235 8589 sw
tri 8235 8491 8333 8589 ne
rect 8333 8585 8687 8589
rect 8333 8491 8465 8585
rect 8035 8465 8235 8491
rect 7861 8413 8235 8465
tri 8235 8413 8313 8491 sw
tri 8333 8413 8411 8491 ne
rect 8411 8465 8465 8491
rect 8585 8491 8687 8585
tri 8687 8491 8785 8589 sw
tri 8785 8491 8883 8589 ne
rect 8883 8585 9237 8589
rect 8883 8491 9015 8585
rect 8585 8465 8785 8491
rect 8411 8413 8785 8465
tri 8785 8413 8863 8491 sw
tri 8883 8413 8961 8491 ne
rect 8961 8465 9015 8491
rect 9135 8491 9237 8585
tri 9237 8491 9335 8589 sw
tri 9335 8491 9433 8589 ne
rect 9433 8585 9787 8589
rect 9433 8491 9565 8585
rect 9135 8465 9335 8491
rect 8961 8413 9335 8465
tri 9335 8413 9413 8491 sw
tri 9433 8413 9511 8491 ne
rect 9511 8465 9565 8491
rect 9685 8491 9787 8585
tri 9787 8491 9885 8589 sw
tri 9885 8491 9983 8589 ne
rect 9983 8585 10337 8589
rect 9983 8491 10115 8585
rect 9685 8465 9885 8491
rect 9511 8413 9885 8465
tri 9885 8413 9963 8491 sw
tri 9983 8413 10061 8491 ne
rect 10061 8465 10115 8491
rect 10235 8491 10337 8585
tri 10337 8491 10435 8589 sw
tri 10435 8491 10533 8589 ne
rect 10533 8585 10887 8589
rect 10533 8491 10665 8585
rect 10235 8465 10435 8491
rect 10061 8413 10435 8465
tri 10435 8413 10513 8491 sw
tri 10533 8413 10611 8491 ne
rect 10611 8465 10665 8491
rect 10785 8491 10887 8585
tri 10887 8491 10985 8589 sw
tri 10985 8491 11083 8589 ne
rect 11083 8585 11437 8589
rect 11083 8491 11215 8585
rect 10785 8465 10985 8491
rect 10611 8413 10985 8465
tri 10985 8413 11063 8491 sw
tri 11083 8413 11161 8491 ne
rect 11161 8465 11215 8491
rect 11335 8491 11437 8585
tri 11437 8491 11535 8589 sw
tri 11535 8491 11633 8589 ne
rect 11633 8585 11987 8589
rect 11633 8491 11765 8585
rect 11335 8465 11535 8491
rect 11161 8413 11535 8465
tri 11535 8413 11613 8491 sw
tri 11633 8413 11711 8491 ne
rect 11711 8465 11765 8491
rect 11885 8491 11987 8585
tri 11987 8491 12085 8589 sw
tri 12085 8491 12183 8589 ne
rect 12183 8585 12537 8589
rect 12183 8491 12315 8585
rect 11885 8465 12085 8491
rect 11711 8413 12085 8465
tri 12085 8413 12163 8491 sw
tri 12183 8413 12261 8491 ne
rect 12261 8465 12315 8491
rect 12435 8491 12537 8585
tri 12537 8491 12635 8589 sw
tri 12635 8491 12733 8589 ne
rect 12733 8585 13087 8589
rect 12733 8491 12865 8585
rect 12435 8465 12635 8491
rect 12261 8413 12635 8465
tri 12635 8413 12713 8491 sw
tri 12733 8413 12811 8491 ne
rect 12811 8465 12865 8491
rect 12985 8491 13087 8585
tri 13087 8491 13185 8589 sw
tri 13185 8491 13283 8589 ne
rect 13283 8585 13637 8589
rect 13283 8491 13415 8585
rect 12985 8465 13185 8491
rect 12811 8413 13185 8465
tri 13185 8413 13263 8491 sw
tri 13283 8413 13361 8491 ne
rect 13361 8465 13415 8491
rect 13535 8491 13637 8585
tri 13637 8491 13735 8589 sw
tri 13735 8491 13833 8589 ne
rect 13833 8585 14187 8589
rect 13833 8491 13965 8585
rect 13535 8465 13735 8491
rect 13361 8413 13735 8465
tri 13735 8413 13813 8491 sw
tri 13833 8413 13911 8491 ne
rect 13911 8465 13965 8491
rect 14085 8491 14187 8585
tri 14187 8491 14285 8589 sw
tri 14285 8491 14383 8589 ne
rect 14383 8585 14737 8589
rect 14383 8491 14515 8585
rect 14085 8465 14285 8491
rect 13911 8413 14285 8465
tri 14285 8413 14363 8491 sw
tri 14383 8413 14461 8491 ne
rect 14461 8465 14515 8491
rect 14635 8491 14737 8585
tri 14737 8491 14835 8589 sw
tri 14835 8491 14933 8589 ne
rect 14933 8585 15287 8589
rect 14933 8491 15065 8585
rect 14635 8465 14835 8491
rect 14461 8413 14835 8465
tri 14835 8413 14913 8491 sw
tri 14933 8413 15011 8491 ne
rect 15011 8465 15065 8491
rect 15185 8491 15287 8585
tri 15287 8491 15385 8589 sw
tri 15385 8491 15483 8589 ne
rect 15483 8585 15837 8589
rect 15483 8491 15615 8585
rect 15185 8465 15385 8491
rect 15011 8413 15385 8465
tri 15385 8413 15463 8491 sw
tri 15483 8413 15561 8491 ne
rect 15561 8465 15615 8491
rect 15735 8491 15837 8585
tri 15837 8491 15935 8589 sw
tri 15935 8491 16033 8589 ne
rect 16033 8585 16387 8589
rect 16033 8491 16165 8585
rect 15735 8465 15935 8491
rect 15561 8413 15935 8465
tri 15935 8413 16013 8491 sw
tri 16033 8413 16111 8491 ne
rect 16111 8465 16165 8491
rect 16285 8491 16387 8585
tri 16387 8491 16485 8589 sw
tri 16485 8491 16583 8589 ne
rect 16583 8585 16937 8589
rect 16583 8491 16715 8585
rect 16285 8465 16485 8491
rect 16111 8413 16485 8465
tri 16485 8413 16563 8491 sw
tri 16583 8413 16661 8491 ne
rect 16661 8465 16715 8491
rect 16835 8491 16937 8585
tri 16937 8491 17035 8589 sw
tri 17035 8491 17133 8589 ne
rect 17133 8585 17487 8589
rect 17133 8491 17265 8585
rect 16835 8465 17035 8491
rect 16661 8413 17035 8465
tri 17035 8413 17113 8491 sw
tri 17133 8413 17211 8491 ne
rect 17211 8465 17265 8491
rect 17385 8491 17487 8585
tri 17487 8491 17585 8589 sw
tri 17585 8491 17683 8589 ne
rect 17683 8585 18037 8589
rect 17683 8491 17815 8585
rect 17385 8465 17585 8491
rect 17211 8413 17585 8465
tri 17585 8413 17663 8491 sw
tri 17683 8413 17761 8491 ne
rect 17761 8465 17815 8491
rect 17935 8491 18037 8585
tri 18037 8491 18135 8589 sw
tri 18135 8491 18233 8589 ne
rect 18233 8585 18587 8589
rect 18233 8491 18365 8585
rect 17935 8465 18135 8491
rect 17761 8413 18135 8465
tri 18135 8413 18213 8491 sw
tri 18233 8413 18311 8491 ne
rect 18311 8465 18365 8491
rect 18485 8491 18587 8585
tri 18587 8491 18685 8589 sw
tri 18685 8491 18783 8589 ne
rect 18783 8585 19137 8589
rect 18783 8491 18915 8585
rect 18485 8465 18685 8491
rect 18311 8413 18685 8465
tri 18685 8413 18763 8491 sw
tri 18783 8413 18861 8491 ne
rect 18861 8465 18915 8491
rect 19035 8491 19137 8585
tri 19137 8491 19235 8589 sw
tri 19235 8491 19333 8589 ne
rect 19333 8585 21800 8589
rect 19333 8491 19465 8585
rect 19035 8465 19235 8491
rect 18861 8413 19235 8465
tri 19235 8413 19313 8491 sw
tri 19333 8413 19411 8491 ne
rect 19411 8465 19465 8491
rect 19585 8465 21800 8585
rect 19411 8413 21800 8465
rect 211 8363 613 8413
rect -500 8313 113 8363
tri 113 8313 163 8363 sw
tri 211 8313 261 8363 ne
rect 261 8333 613 8363
tri 613 8333 693 8413 sw
tri 711 8333 791 8413 ne
rect 791 8333 1163 8413
tri 1163 8333 1243 8413 sw
tri 1261 8333 1341 8413 ne
rect 1341 8333 1713 8413
tri 1713 8333 1793 8413 sw
tri 1811 8333 1891 8413 ne
rect 1891 8333 2263 8413
tri 2263 8333 2343 8413 sw
tri 2361 8333 2441 8413 ne
rect 2441 8333 2813 8413
tri 2813 8333 2893 8413 sw
tri 2911 8333 2991 8413 ne
rect 2991 8333 3363 8413
tri 3363 8333 3443 8413 sw
tri 3461 8333 3541 8413 ne
rect 3541 8333 3913 8413
tri 3913 8333 3993 8413 sw
tri 4011 8333 4091 8413 ne
rect 4091 8333 4463 8413
tri 4463 8333 4543 8413 sw
tri 4561 8333 4641 8413 ne
rect 4641 8333 5013 8413
tri 5013 8333 5093 8413 sw
tri 5111 8333 5191 8413 ne
rect 5191 8333 5563 8413
tri 5563 8333 5643 8413 sw
tri 5661 8333 5741 8413 ne
rect 5741 8333 6113 8413
tri 6113 8333 6193 8413 sw
tri 6211 8333 6291 8413 ne
rect 6291 8333 6663 8413
tri 6663 8333 6743 8413 sw
tri 6761 8333 6841 8413 ne
rect 6841 8333 7213 8413
tri 7213 8333 7293 8413 sw
tri 7311 8333 7391 8413 ne
rect 7391 8333 7763 8413
tri 7763 8333 7843 8413 sw
tri 7861 8333 7941 8413 ne
rect 7941 8333 8313 8413
tri 8313 8333 8393 8413 sw
tri 8411 8333 8491 8413 ne
rect 8491 8333 8863 8413
tri 8863 8333 8943 8413 sw
tri 8961 8333 9041 8413 ne
rect 9041 8333 9413 8413
tri 9413 8333 9493 8413 sw
tri 9511 8333 9591 8413 ne
rect 9591 8333 9963 8413
tri 9963 8333 10043 8413 sw
tri 10061 8333 10141 8413 ne
rect 10141 8333 10513 8413
tri 10513 8333 10593 8413 sw
tri 10611 8333 10691 8413 ne
rect 10691 8333 11063 8413
tri 11063 8333 11143 8413 sw
tri 11161 8333 11241 8413 ne
rect 11241 8333 11613 8413
tri 11613 8333 11693 8413 sw
tri 11711 8333 11791 8413 ne
rect 11791 8333 12163 8413
tri 12163 8333 12243 8413 sw
tri 12261 8333 12341 8413 ne
rect 12341 8333 12713 8413
tri 12713 8333 12793 8413 sw
tri 12811 8333 12891 8413 ne
rect 12891 8333 13263 8413
tri 13263 8333 13343 8413 sw
tri 13361 8333 13441 8413 ne
rect 13441 8333 13813 8413
tri 13813 8333 13893 8413 sw
tri 13911 8333 13991 8413 ne
rect 13991 8333 14363 8413
tri 14363 8333 14443 8413 sw
tri 14461 8333 14541 8413 ne
rect 14541 8333 14913 8413
tri 14913 8333 14993 8413 sw
tri 15011 8333 15091 8413 ne
rect 15091 8333 15463 8413
tri 15463 8333 15543 8413 sw
tri 15561 8333 15641 8413 ne
rect 15641 8333 16013 8413
tri 16013 8333 16093 8413 sw
tri 16111 8333 16191 8413 ne
rect 16191 8333 16563 8413
tri 16563 8333 16643 8413 sw
tri 16661 8333 16741 8413 ne
rect 16741 8333 17113 8413
tri 17113 8333 17193 8413 sw
tri 17211 8333 17291 8413 ne
rect 17291 8333 17663 8413
tri 17663 8333 17743 8413 sw
tri 17761 8333 17841 8413 ne
rect 17841 8333 18213 8413
tri 18213 8333 18293 8413 sw
tri 18311 8333 18391 8413 ne
rect 18391 8333 18763 8413
tri 18763 8333 18843 8413 sw
tri 18861 8333 18941 8413 ne
rect 18941 8333 19313 8413
tri 19313 8333 19393 8413 sw
tri 19411 8333 19491 8413 ne
rect 19491 8333 20100 8413
rect 261 8313 693 8333
rect -500 8235 163 8313
tri 163 8235 241 8313 sw
tri 261 8235 339 8313 ne
rect 339 8235 693 8313
tri 693 8235 791 8333 sw
tri 791 8235 889 8333 ne
rect 889 8235 1243 8333
tri 1243 8235 1341 8333 sw
tri 1341 8235 1439 8333 ne
rect 1439 8235 1793 8333
tri 1793 8235 1891 8333 sw
tri 1891 8235 1989 8333 ne
rect 1989 8235 2343 8333
tri 2343 8235 2441 8333 sw
tri 2441 8235 2539 8333 ne
rect 2539 8235 2893 8333
tri 2893 8235 2991 8333 sw
tri 2991 8235 3089 8333 ne
rect 3089 8235 3443 8333
tri 3443 8235 3541 8333 sw
tri 3541 8235 3639 8333 ne
rect 3639 8235 3993 8333
tri 3993 8235 4091 8333 sw
tri 4091 8235 4189 8333 ne
rect 4189 8235 4543 8333
tri 4543 8235 4641 8333 sw
tri 4641 8235 4739 8333 ne
rect 4739 8235 5093 8333
tri 5093 8235 5191 8333 sw
tri 5191 8235 5289 8333 ne
rect 5289 8235 5643 8333
tri 5643 8235 5741 8333 sw
tri 5741 8235 5839 8333 ne
rect 5839 8235 6193 8333
tri 6193 8235 6291 8333 sw
tri 6291 8235 6389 8333 ne
rect 6389 8235 6743 8333
tri 6743 8235 6841 8333 sw
tri 6841 8235 6939 8333 ne
rect 6939 8235 7293 8333
tri 7293 8235 7391 8333 sw
tri 7391 8235 7489 8333 ne
rect 7489 8235 7843 8333
tri 7843 8235 7941 8333 sw
tri 7941 8235 8039 8333 ne
rect 8039 8235 8393 8333
tri 8393 8235 8491 8333 sw
tri 8491 8235 8589 8333 ne
rect 8589 8235 8943 8333
tri 8943 8235 9041 8333 sw
tri 9041 8235 9139 8333 ne
rect 9139 8235 9493 8333
tri 9493 8235 9591 8333 sw
tri 9591 8235 9689 8333 ne
rect 9689 8235 10043 8333
tri 10043 8235 10141 8333 sw
tri 10141 8235 10239 8333 ne
rect 10239 8235 10593 8333
tri 10593 8235 10691 8333 sw
tri 10691 8235 10789 8333 ne
rect 10789 8235 11143 8333
tri 11143 8235 11241 8333 sw
tri 11241 8235 11339 8333 ne
rect 11339 8235 11693 8333
tri 11693 8235 11791 8333 sw
tri 11791 8235 11889 8333 ne
rect 11889 8235 12243 8333
tri 12243 8235 12341 8333 sw
tri 12341 8235 12439 8333 ne
rect 12439 8235 12793 8333
tri 12793 8235 12891 8333 sw
tri 12891 8235 12989 8333 ne
rect 12989 8235 13343 8333
tri 13343 8235 13441 8333 sw
tri 13441 8235 13539 8333 ne
rect 13539 8235 13893 8333
tri 13893 8235 13991 8333 sw
tri 13991 8235 14089 8333 ne
rect 14089 8235 14443 8333
tri 14443 8235 14541 8333 sw
tri 14541 8235 14639 8333 ne
rect 14639 8235 14993 8333
tri 14993 8235 15091 8333 sw
tri 15091 8235 15189 8333 ne
rect 15189 8235 15543 8333
tri 15543 8235 15641 8333 sw
tri 15641 8235 15739 8333 ne
rect 15739 8235 16093 8333
tri 16093 8235 16191 8333 sw
tri 16191 8235 16289 8333 ne
rect 16289 8235 16643 8333
tri 16643 8235 16741 8333 sw
tri 16741 8235 16839 8333 ne
rect 16839 8235 17193 8333
tri 17193 8235 17291 8333 sw
tri 17291 8235 17389 8333 ne
rect 17389 8235 17743 8333
tri 17743 8235 17841 8333 sw
tri 17841 8235 17939 8333 ne
rect 17939 8235 18293 8333
tri 18293 8235 18391 8333 sw
tri 18391 8235 18489 8333 ne
rect 18489 8235 18843 8333
tri 18843 8235 18941 8333 sw
tri 18941 8235 19039 8333 ne
rect 19039 8235 19393 8333
tri 19393 8235 19491 8333 sw
tri 19491 8235 19589 8333 ne
rect 19589 8313 20100 8333
rect 20200 8313 21800 8413
rect 19589 8235 21800 8313
rect -500 8187 241 8235
rect -500 8087 -400 8187
rect -300 8137 241 8187
tri 241 8137 339 8235 sw
tri 339 8137 437 8235 ne
rect 437 8137 791 8235
tri 791 8137 889 8235 sw
tri 889 8137 987 8235 ne
rect 987 8137 1341 8235
tri 1341 8137 1439 8235 sw
tri 1439 8137 1537 8235 ne
rect 1537 8137 1891 8235
tri 1891 8137 1989 8235 sw
tri 1989 8137 2087 8235 ne
rect 2087 8137 2441 8235
tri 2441 8137 2539 8235 sw
tri 2539 8137 2637 8235 ne
rect 2637 8137 2991 8235
tri 2991 8137 3089 8235 sw
tri 3089 8137 3187 8235 ne
rect 3187 8137 3541 8235
tri 3541 8137 3639 8235 sw
tri 3639 8137 3737 8235 ne
rect 3737 8137 4091 8235
tri 4091 8137 4189 8235 sw
tri 4189 8137 4287 8235 ne
rect 4287 8137 4641 8235
tri 4641 8137 4739 8235 sw
tri 4739 8137 4837 8235 ne
rect 4837 8137 5191 8235
tri 5191 8137 5289 8235 sw
tri 5289 8137 5387 8235 ne
rect 5387 8137 5741 8235
tri 5741 8137 5839 8235 sw
tri 5839 8137 5937 8235 ne
rect 5937 8137 6291 8235
tri 6291 8137 6389 8235 sw
tri 6389 8137 6487 8235 ne
rect 6487 8137 6841 8235
tri 6841 8137 6939 8235 sw
tri 6939 8137 7037 8235 ne
rect 7037 8137 7391 8235
tri 7391 8137 7489 8235 sw
tri 7489 8137 7587 8235 ne
rect 7587 8137 7941 8235
tri 7941 8137 8039 8235 sw
tri 8039 8137 8137 8235 ne
rect 8137 8137 8491 8235
tri 8491 8137 8589 8235 sw
tri 8589 8137 8687 8235 ne
rect 8687 8137 9041 8235
tri 9041 8137 9139 8235 sw
tri 9139 8137 9237 8235 ne
rect 9237 8137 9591 8235
tri 9591 8137 9689 8235 sw
tri 9689 8137 9787 8235 ne
rect 9787 8137 10141 8235
tri 10141 8137 10239 8235 sw
tri 10239 8137 10337 8235 ne
rect 10337 8137 10691 8235
tri 10691 8137 10789 8235 sw
tri 10789 8137 10887 8235 ne
rect 10887 8137 11241 8235
tri 11241 8137 11339 8235 sw
tri 11339 8137 11437 8235 ne
rect 11437 8137 11791 8235
tri 11791 8137 11889 8235 sw
tri 11889 8137 11987 8235 ne
rect 11987 8137 12341 8235
tri 12341 8137 12439 8235 sw
tri 12439 8137 12537 8235 ne
rect 12537 8137 12891 8235
tri 12891 8137 12989 8235 sw
tri 12989 8137 13087 8235 ne
rect 13087 8137 13441 8235
tri 13441 8137 13539 8235 sw
tri 13539 8137 13637 8235 ne
rect 13637 8137 13991 8235
tri 13991 8137 14089 8235 sw
tri 14089 8137 14187 8235 ne
rect 14187 8137 14541 8235
tri 14541 8137 14639 8235 sw
tri 14639 8137 14737 8235 ne
rect 14737 8137 15091 8235
tri 15091 8137 15189 8235 sw
tri 15189 8137 15287 8235 ne
rect 15287 8137 15641 8235
tri 15641 8137 15739 8235 sw
tri 15739 8137 15837 8235 ne
rect 15837 8137 16191 8235
tri 16191 8137 16289 8235 sw
tri 16289 8137 16387 8235 ne
rect 16387 8137 16741 8235
tri 16741 8137 16839 8235 sw
tri 16839 8137 16937 8235 ne
rect 16937 8137 17291 8235
tri 17291 8137 17389 8235 sw
tri 17389 8137 17487 8235 ne
rect 17487 8137 17841 8235
tri 17841 8137 17939 8235 sw
tri 17939 8137 18037 8235 ne
rect 18037 8137 18391 8235
tri 18391 8137 18489 8235 sw
tri 18489 8137 18587 8235 ne
rect 18587 8137 18941 8235
tri 18941 8137 19039 8235 sw
tri 19039 8137 19137 8235 ne
rect 19137 8137 19491 8235
tri 19491 8137 19589 8235 sw
tri 19589 8137 19687 8235 ne
rect 19687 8137 21800 8235
rect -300 8087 339 8137
rect -500 8039 339 8087
tri 339 8039 437 8137 sw
tri 437 8039 535 8137 ne
rect 535 8039 889 8137
tri 889 8039 987 8137 sw
tri 987 8039 1085 8137 ne
rect 1085 8039 1439 8137
tri 1439 8039 1537 8137 sw
tri 1537 8039 1635 8137 ne
rect 1635 8039 1989 8137
tri 1989 8039 2087 8137 sw
tri 2087 8039 2185 8137 ne
rect 2185 8039 2539 8137
tri 2539 8039 2637 8137 sw
tri 2637 8039 2735 8137 ne
rect 2735 8039 3089 8137
tri 3089 8039 3187 8137 sw
tri 3187 8039 3285 8137 ne
rect 3285 8039 3639 8137
tri 3639 8039 3737 8137 sw
tri 3737 8039 3835 8137 ne
rect 3835 8039 4189 8137
tri 4189 8039 4287 8137 sw
tri 4287 8039 4385 8137 ne
rect 4385 8039 4739 8137
tri 4739 8039 4837 8137 sw
tri 4837 8039 4935 8137 ne
rect 4935 8039 5289 8137
tri 5289 8039 5387 8137 sw
tri 5387 8039 5485 8137 ne
rect 5485 8039 5839 8137
tri 5839 8039 5937 8137 sw
tri 5937 8039 6035 8137 ne
rect 6035 8039 6389 8137
tri 6389 8039 6487 8137 sw
tri 6487 8039 6585 8137 ne
rect 6585 8039 6939 8137
tri 6939 8039 7037 8137 sw
tri 7037 8039 7135 8137 ne
rect 7135 8039 7489 8137
tri 7489 8039 7587 8137 sw
tri 7587 8039 7685 8137 ne
rect 7685 8039 8039 8137
tri 8039 8039 8137 8137 sw
tri 8137 8039 8235 8137 ne
rect 8235 8039 8589 8137
tri 8589 8039 8687 8137 sw
tri 8687 8039 8785 8137 ne
rect 8785 8039 9139 8137
tri 9139 8039 9237 8137 sw
tri 9237 8039 9335 8137 ne
rect 9335 8039 9689 8137
tri 9689 8039 9787 8137 sw
tri 9787 8039 9885 8137 ne
rect 9885 8039 10239 8137
tri 10239 8039 10337 8137 sw
tri 10337 8039 10435 8137 ne
rect 10435 8039 10789 8137
tri 10789 8039 10887 8137 sw
tri 10887 8039 10985 8137 ne
rect 10985 8039 11339 8137
tri 11339 8039 11437 8137 sw
tri 11437 8039 11535 8137 ne
rect 11535 8039 11889 8137
tri 11889 8039 11987 8137 sw
tri 11987 8039 12085 8137 ne
rect 12085 8039 12439 8137
tri 12439 8039 12537 8137 sw
tri 12537 8039 12635 8137 ne
rect 12635 8039 12989 8137
tri 12989 8039 13087 8137 sw
tri 13087 8039 13185 8137 ne
rect 13185 8039 13539 8137
tri 13539 8039 13637 8137 sw
tri 13637 8039 13735 8137 ne
rect 13735 8039 14089 8137
tri 14089 8039 14187 8137 sw
tri 14187 8039 14285 8137 ne
rect 14285 8039 14639 8137
tri 14639 8039 14737 8137 sw
tri 14737 8039 14835 8137 ne
rect 14835 8039 15189 8137
tri 15189 8039 15287 8137 sw
tri 15287 8039 15385 8137 ne
rect 15385 8039 15739 8137
tri 15739 8039 15837 8137 sw
tri 15837 8039 15935 8137 ne
rect 15935 8039 16289 8137
tri 16289 8039 16387 8137 sw
tri 16387 8039 16485 8137 ne
rect 16485 8039 16839 8137
tri 16839 8039 16937 8137 sw
tri 16937 8039 17035 8137 ne
rect 17035 8039 17389 8137
tri 17389 8039 17487 8137 sw
tri 17487 8039 17585 8137 ne
rect 17585 8039 17939 8137
tri 17939 8039 18037 8137 sw
tri 18037 8039 18135 8137 ne
rect 18135 8039 18489 8137
tri 18489 8039 18587 8137 sw
tri 18587 8039 18685 8137 ne
rect 18685 8039 19039 8137
tri 19039 8039 19137 8137 sw
tri 19137 8039 19235 8137 ne
rect 19235 8039 19589 8137
tri 19589 8039 19687 8137 sw
rect -500 8035 437 8039
rect -500 7915 215 8035
rect 335 7941 437 8035
tri 437 7941 535 8039 sw
tri 535 7941 633 8039 ne
rect 633 8035 987 8039
rect 633 7941 765 8035
rect 335 7915 535 7941
rect -500 7911 535 7915
tri 535 7911 565 7941 sw
tri 633 7911 663 7941 ne
rect 663 7915 765 7941
rect 885 7941 987 8035
tri 987 7941 1085 8039 sw
tri 1085 7941 1183 8039 ne
rect 1183 8035 1537 8039
rect 1183 7941 1315 8035
rect 885 7915 1085 7941
rect 663 7911 1085 7915
tri 1085 7911 1115 7941 sw
tri 1183 7911 1213 7941 ne
rect 1213 7915 1315 7941
rect 1435 7941 1537 8035
tri 1537 7941 1635 8039 sw
tri 1635 7941 1733 8039 ne
rect 1733 8035 2087 8039
rect 1733 7941 1865 8035
rect 1435 7915 1635 7941
rect 1213 7911 1635 7915
tri 1635 7911 1665 7941 sw
tri 1733 7911 1763 7941 ne
rect 1763 7915 1865 7941
rect 1985 7941 2087 8035
tri 2087 7941 2185 8039 sw
tri 2185 7941 2283 8039 ne
rect 2283 8035 2637 8039
rect 2283 7941 2415 8035
rect 1985 7915 2185 7941
rect 1763 7911 2185 7915
tri 2185 7911 2215 7941 sw
tri 2283 7911 2313 7941 ne
rect 2313 7915 2415 7941
rect 2535 7941 2637 8035
tri 2637 7941 2735 8039 sw
tri 2735 7941 2833 8039 ne
rect 2833 8035 3187 8039
rect 2833 7941 2965 8035
rect 2535 7915 2735 7941
rect 2313 7911 2735 7915
tri 2735 7911 2765 7941 sw
tri 2833 7911 2863 7941 ne
rect 2863 7915 2965 7941
rect 3085 7941 3187 8035
tri 3187 7941 3285 8039 sw
tri 3285 7941 3383 8039 ne
rect 3383 8035 3737 8039
rect 3383 7941 3515 8035
rect 3085 7915 3285 7941
rect 2863 7911 3285 7915
tri 3285 7911 3315 7941 sw
tri 3383 7911 3413 7941 ne
rect 3413 7915 3515 7941
rect 3635 7941 3737 8035
tri 3737 7941 3835 8039 sw
tri 3835 7941 3933 8039 ne
rect 3933 8035 4287 8039
rect 3933 7941 4065 8035
rect 3635 7915 3835 7941
rect 3413 7911 3835 7915
tri 3835 7911 3865 7941 sw
tri 3933 7911 3963 7941 ne
rect 3963 7915 4065 7941
rect 4185 7941 4287 8035
tri 4287 7941 4385 8039 sw
tri 4385 7941 4483 8039 ne
rect 4483 8035 4837 8039
rect 4483 7941 4615 8035
rect 4185 7915 4385 7941
rect 3963 7911 4385 7915
tri 4385 7911 4415 7941 sw
tri 4483 7911 4513 7941 ne
rect 4513 7915 4615 7941
rect 4735 7941 4837 8035
tri 4837 7941 4935 8039 sw
tri 4935 7941 5033 8039 ne
rect 5033 8035 5387 8039
rect 5033 7941 5165 8035
rect 4735 7915 4935 7941
rect 4513 7911 4935 7915
tri 4935 7911 4965 7941 sw
tri 5033 7911 5063 7941 ne
rect 5063 7915 5165 7941
rect 5285 7941 5387 8035
tri 5387 7941 5485 8039 sw
tri 5485 7941 5583 8039 ne
rect 5583 8035 5937 8039
rect 5583 7941 5715 8035
rect 5285 7915 5485 7941
rect 5063 7911 5485 7915
tri 5485 7911 5515 7941 sw
tri 5583 7911 5613 7941 ne
rect 5613 7915 5715 7941
rect 5835 7941 5937 8035
tri 5937 7941 6035 8039 sw
tri 6035 7941 6133 8039 ne
rect 6133 8035 6487 8039
rect 6133 7941 6265 8035
rect 5835 7915 6035 7941
rect 5613 7911 6035 7915
tri 6035 7911 6065 7941 sw
tri 6133 7911 6163 7941 ne
rect 6163 7915 6265 7941
rect 6385 7941 6487 8035
tri 6487 7941 6585 8039 sw
tri 6585 7941 6683 8039 ne
rect 6683 8035 7037 8039
rect 6683 7941 6815 8035
rect 6385 7915 6585 7941
rect 6163 7911 6585 7915
tri 6585 7911 6615 7941 sw
tri 6683 7911 6713 7941 ne
rect 6713 7915 6815 7941
rect 6935 7941 7037 8035
tri 7037 7941 7135 8039 sw
tri 7135 7941 7233 8039 ne
rect 7233 8035 7587 8039
rect 7233 7941 7365 8035
rect 6935 7915 7135 7941
rect 6713 7911 7135 7915
tri 7135 7911 7165 7941 sw
tri 7233 7911 7263 7941 ne
rect 7263 7915 7365 7941
rect 7485 7941 7587 8035
tri 7587 7941 7685 8039 sw
tri 7685 7941 7783 8039 ne
rect 7783 8035 8137 8039
rect 7783 7941 7915 8035
rect 7485 7915 7685 7941
rect 7263 7911 7685 7915
tri 7685 7911 7715 7941 sw
tri 7783 7911 7813 7941 ne
rect 7813 7915 7915 7941
rect 8035 7941 8137 8035
tri 8137 7941 8235 8039 sw
tri 8235 7941 8333 8039 ne
rect 8333 8035 8687 8039
rect 8333 7941 8465 8035
rect 8035 7915 8235 7941
rect 7813 7911 8235 7915
tri 8235 7911 8265 7941 sw
tri 8333 7911 8363 7941 ne
rect 8363 7915 8465 7941
rect 8585 7941 8687 8035
tri 8687 7941 8785 8039 sw
tri 8785 7941 8883 8039 ne
rect 8883 8035 9237 8039
rect 8883 7941 9015 8035
rect 8585 7915 8785 7941
rect 8363 7911 8785 7915
tri 8785 7911 8815 7941 sw
tri 8883 7911 8913 7941 ne
rect 8913 7915 9015 7941
rect 9135 7941 9237 8035
tri 9237 7941 9335 8039 sw
tri 9335 7941 9433 8039 ne
rect 9433 8035 9787 8039
rect 9433 7941 9565 8035
rect 9135 7915 9335 7941
rect 8913 7911 9335 7915
tri 9335 7911 9365 7941 sw
tri 9433 7911 9463 7941 ne
rect 9463 7915 9565 7941
rect 9685 7941 9787 8035
tri 9787 7941 9885 8039 sw
tri 9885 7941 9983 8039 ne
rect 9983 8035 10337 8039
rect 9983 7941 10115 8035
rect 9685 7915 9885 7941
rect 9463 7911 9885 7915
tri 9885 7911 9915 7941 sw
tri 9983 7911 10013 7941 ne
rect 10013 7915 10115 7941
rect 10235 7941 10337 8035
tri 10337 7941 10435 8039 sw
tri 10435 7941 10533 8039 ne
rect 10533 8035 10887 8039
rect 10533 7941 10665 8035
rect 10235 7915 10435 7941
rect 10013 7911 10435 7915
tri 10435 7911 10465 7941 sw
tri 10533 7911 10563 7941 ne
rect 10563 7915 10665 7941
rect 10785 7941 10887 8035
tri 10887 7941 10985 8039 sw
tri 10985 7941 11083 8039 ne
rect 11083 8035 11437 8039
rect 11083 7941 11215 8035
rect 10785 7915 10985 7941
rect 10563 7911 10985 7915
tri 10985 7911 11015 7941 sw
tri 11083 7911 11113 7941 ne
rect 11113 7915 11215 7941
rect 11335 7941 11437 8035
tri 11437 7941 11535 8039 sw
tri 11535 7941 11633 8039 ne
rect 11633 8035 11987 8039
rect 11633 7941 11765 8035
rect 11335 7915 11535 7941
rect 11113 7911 11535 7915
tri 11535 7911 11565 7941 sw
tri 11633 7911 11663 7941 ne
rect 11663 7915 11765 7941
rect 11885 7941 11987 8035
tri 11987 7941 12085 8039 sw
tri 12085 7941 12183 8039 ne
rect 12183 8035 12537 8039
rect 12183 7941 12315 8035
rect 11885 7915 12085 7941
rect 11663 7911 12085 7915
tri 12085 7911 12115 7941 sw
tri 12183 7911 12213 7941 ne
rect 12213 7915 12315 7941
rect 12435 7941 12537 8035
tri 12537 7941 12635 8039 sw
tri 12635 7941 12733 8039 ne
rect 12733 8035 13087 8039
rect 12733 7941 12865 8035
rect 12435 7915 12635 7941
rect 12213 7911 12635 7915
tri 12635 7911 12665 7941 sw
tri 12733 7911 12763 7941 ne
rect 12763 7915 12865 7941
rect 12985 7941 13087 8035
tri 13087 7941 13185 8039 sw
tri 13185 7941 13283 8039 ne
rect 13283 8035 13637 8039
rect 13283 7941 13415 8035
rect 12985 7915 13185 7941
rect 12763 7911 13185 7915
tri 13185 7911 13215 7941 sw
tri 13283 7911 13313 7941 ne
rect 13313 7915 13415 7941
rect 13535 7941 13637 8035
tri 13637 7941 13735 8039 sw
tri 13735 7941 13833 8039 ne
rect 13833 8035 14187 8039
rect 13833 7941 13965 8035
rect 13535 7915 13735 7941
rect 13313 7911 13735 7915
tri 13735 7911 13765 7941 sw
tri 13833 7911 13863 7941 ne
rect 13863 7915 13965 7941
rect 14085 7941 14187 8035
tri 14187 7941 14285 8039 sw
tri 14285 7941 14383 8039 ne
rect 14383 8035 14737 8039
rect 14383 7941 14515 8035
rect 14085 7915 14285 7941
rect 13863 7911 14285 7915
tri 14285 7911 14315 7941 sw
tri 14383 7911 14413 7941 ne
rect 14413 7915 14515 7941
rect 14635 7941 14737 8035
tri 14737 7941 14835 8039 sw
tri 14835 7941 14933 8039 ne
rect 14933 8035 15287 8039
rect 14933 7941 15065 8035
rect 14635 7915 14835 7941
rect 14413 7911 14835 7915
tri 14835 7911 14865 7941 sw
tri 14933 7911 14963 7941 ne
rect 14963 7915 15065 7941
rect 15185 7941 15287 8035
tri 15287 7941 15385 8039 sw
tri 15385 7941 15483 8039 ne
rect 15483 8035 15837 8039
rect 15483 7941 15615 8035
rect 15185 7915 15385 7941
rect 14963 7911 15385 7915
tri 15385 7911 15415 7941 sw
tri 15483 7911 15513 7941 ne
rect 15513 7915 15615 7941
rect 15735 7941 15837 8035
tri 15837 7941 15935 8039 sw
tri 15935 7941 16033 8039 ne
rect 16033 8035 16387 8039
rect 16033 7941 16165 8035
rect 15735 7915 15935 7941
rect 15513 7911 15935 7915
tri 15935 7911 15965 7941 sw
tri 16033 7911 16063 7941 ne
rect 16063 7915 16165 7941
rect 16285 7941 16387 8035
tri 16387 7941 16485 8039 sw
tri 16485 7941 16583 8039 ne
rect 16583 8035 16937 8039
rect 16583 7941 16715 8035
rect 16285 7915 16485 7941
rect 16063 7911 16485 7915
tri 16485 7911 16515 7941 sw
tri 16583 7911 16613 7941 ne
rect 16613 7915 16715 7941
rect 16835 7941 16937 8035
tri 16937 7941 17035 8039 sw
tri 17035 7941 17133 8039 ne
rect 17133 8035 17487 8039
rect 17133 7941 17265 8035
rect 16835 7915 17035 7941
rect 16613 7911 17035 7915
tri 17035 7911 17065 7941 sw
tri 17133 7911 17163 7941 ne
rect 17163 7915 17265 7941
rect 17385 7941 17487 8035
tri 17487 7941 17585 8039 sw
tri 17585 7941 17683 8039 ne
rect 17683 8035 18037 8039
rect 17683 7941 17815 8035
rect 17385 7915 17585 7941
rect 17163 7911 17585 7915
tri 17585 7911 17615 7941 sw
tri 17683 7911 17713 7941 ne
rect 17713 7915 17815 7941
rect 17935 7941 18037 8035
tri 18037 7941 18135 8039 sw
tri 18135 7941 18233 8039 ne
rect 18233 8035 18587 8039
rect 18233 7941 18365 8035
rect 17935 7915 18135 7941
rect 17713 7911 18135 7915
tri 18135 7911 18165 7941 sw
tri 18233 7911 18263 7941 ne
rect 18263 7915 18365 7941
rect 18485 7941 18587 8035
tri 18587 7941 18685 8039 sw
tri 18685 7941 18783 8039 ne
rect 18783 8035 19137 8039
rect 18783 7941 18915 8035
rect 18485 7915 18685 7941
rect 18263 7911 18685 7915
tri 18685 7911 18715 7941 sw
tri 18783 7911 18813 7941 ne
rect 18813 7915 18915 7941
rect 19035 7941 19137 8035
tri 19137 7941 19235 8039 sw
tri 19235 7941 19333 8039 ne
rect 19333 8035 20300 8039
rect 19333 7941 19465 8035
rect 19035 7915 19235 7941
rect 18813 7911 19235 7915
tri 19235 7911 19265 7941 sw
tri 19333 7911 19363 7941 ne
rect 19363 7915 19465 7941
rect 19585 7915 20300 8035
rect 19363 7911 20300 7915
tri 113 7813 211 7911 ne
rect 211 7813 565 7911
tri 565 7813 663 7911 sw
tri 663 7813 761 7911 ne
rect 761 7813 1115 7911
tri 1115 7813 1213 7911 sw
tri 1213 7813 1311 7911 ne
rect 1311 7813 1665 7911
tri 1665 7813 1763 7911 sw
tri 1763 7813 1861 7911 ne
rect 1861 7813 2215 7911
tri 2215 7813 2313 7911 sw
tri 2313 7813 2411 7911 ne
rect 2411 7813 2765 7911
tri 2765 7813 2863 7911 sw
tri 2863 7813 2961 7911 ne
rect 2961 7813 3315 7911
tri 3315 7813 3413 7911 sw
tri 3413 7813 3511 7911 ne
rect 3511 7813 3865 7911
tri 3865 7813 3963 7911 sw
tri 3963 7813 4061 7911 ne
rect 4061 7813 4415 7911
tri 4415 7813 4513 7911 sw
tri 4513 7813 4611 7911 ne
rect 4611 7813 4965 7911
tri 4965 7813 5063 7911 sw
tri 5063 7813 5161 7911 ne
rect 5161 7813 5515 7911
tri 5515 7813 5613 7911 sw
tri 5613 7813 5711 7911 ne
rect 5711 7813 6065 7911
tri 6065 7813 6163 7911 sw
tri 6163 7813 6261 7911 ne
rect 6261 7813 6615 7911
tri 6615 7813 6713 7911 sw
tri 6713 7813 6811 7911 ne
rect 6811 7813 7165 7911
tri 7165 7813 7263 7911 sw
tri 7263 7813 7361 7911 ne
rect 7361 7813 7715 7911
tri 7715 7813 7813 7911 sw
tri 7813 7813 7911 7911 ne
rect 7911 7813 8265 7911
tri 8265 7813 8363 7911 sw
tri 8363 7813 8461 7911 ne
rect 8461 7813 8815 7911
tri 8815 7813 8913 7911 sw
tri 8913 7813 9011 7911 ne
rect 9011 7813 9365 7911
tri 9365 7813 9463 7911 sw
tri 9463 7813 9561 7911 ne
rect 9561 7813 9915 7911
tri 9915 7813 10013 7911 sw
tri 10013 7813 10111 7911 ne
rect 10111 7813 10465 7911
tri 10465 7813 10563 7911 sw
tri 10563 7813 10661 7911 ne
rect 10661 7813 11015 7911
tri 11015 7813 11113 7911 sw
tri 11113 7813 11211 7911 ne
rect 11211 7813 11565 7911
tri 11565 7813 11663 7911 sw
tri 11663 7813 11761 7911 ne
rect 11761 7813 12115 7911
tri 12115 7813 12213 7911 sw
tri 12213 7813 12311 7911 ne
rect 12311 7813 12665 7911
tri 12665 7813 12763 7911 sw
tri 12763 7813 12861 7911 ne
rect 12861 7813 13215 7911
tri 13215 7813 13313 7911 sw
tri 13313 7813 13411 7911 ne
rect 13411 7813 13765 7911
tri 13765 7813 13863 7911 sw
tri 13863 7813 13961 7911 ne
rect 13961 7813 14315 7911
tri 14315 7813 14413 7911 sw
tri 14413 7813 14511 7911 ne
rect 14511 7813 14865 7911
tri 14865 7813 14963 7911 sw
tri 14963 7813 15061 7911 ne
rect 15061 7813 15415 7911
tri 15415 7813 15513 7911 sw
tri 15513 7813 15611 7911 ne
rect 15611 7813 15965 7911
tri 15965 7813 16063 7911 sw
tri 16063 7813 16161 7911 ne
rect 16161 7813 16515 7911
tri 16515 7813 16613 7911 sw
tri 16613 7813 16711 7911 ne
rect 16711 7813 17065 7911
tri 17065 7813 17163 7911 sw
tri 17163 7813 17261 7911 ne
rect 17261 7813 17615 7911
tri 17615 7813 17713 7911 sw
tri 17713 7813 17811 7911 ne
rect 17811 7813 18165 7911
tri 18165 7813 18263 7911 sw
tri 18263 7813 18361 7911 ne
rect 18361 7813 18715 7911
tri 18715 7813 18813 7911 sw
tri 18813 7813 18911 7911 ne
rect 18911 7813 19265 7911
tri 19265 7813 19363 7911 sw
tri 19363 7813 19461 7911 ne
rect 19461 7813 20300 7911
rect -2000 7783 113 7813
tri 113 7783 143 7813 sw
tri 211 7783 241 7813 ne
rect 241 7783 663 7813
tri 663 7783 693 7813 sw
tri 761 7783 791 7813 ne
rect 791 7783 1213 7813
tri 1213 7783 1243 7813 sw
tri 1311 7783 1341 7813 ne
rect 1341 7783 1763 7813
tri 1763 7783 1793 7813 sw
tri 1861 7783 1891 7813 ne
rect 1891 7783 2313 7813
tri 2313 7783 2343 7813 sw
tri 2411 7783 2441 7813 ne
rect 2441 7783 2863 7813
tri 2863 7783 2893 7813 sw
tri 2961 7783 2991 7813 ne
rect 2991 7783 3413 7813
tri 3413 7783 3443 7813 sw
tri 3511 7783 3541 7813 ne
rect 3541 7783 3963 7813
tri 3963 7783 3993 7813 sw
tri 4061 7783 4091 7813 ne
rect 4091 7783 4513 7813
tri 4513 7783 4543 7813 sw
tri 4611 7783 4641 7813 ne
rect 4641 7783 5063 7813
tri 5063 7783 5093 7813 sw
tri 5161 7783 5191 7813 ne
rect 5191 7783 5613 7813
tri 5613 7783 5643 7813 sw
tri 5711 7783 5741 7813 ne
rect 5741 7783 6163 7813
tri 6163 7783 6193 7813 sw
tri 6261 7783 6291 7813 ne
rect 6291 7783 6713 7813
tri 6713 7783 6743 7813 sw
tri 6811 7783 6841 7813 ne
rect 6841 7783 7263 7813
tri 7263 7783 7293 7813 sw
tri 7361 7783 7391 7813 ne
rect 7391 7783 7813 7813
tri 7813 7783 7843 7813 sw
tri 7911 7783 7941 7813 ne
rect 7941 7783 8363 7813
tri 8363 7783 8393 7813 sw
tri 8461 7783 8491 7813 ne
rect 8491 7783 8913 7813
tri 8913 7783 8943 7813 sw
tri 9011 7783 9041 7813 ne
rect 9041 7783 9463 7813
tri 9463 7783 9493 7813 sw
tri 9561 7783 9591 7813 ne
rect 9591 7783 10013 7813
tri 10013 7783 10043 7813 sw
tri 10111 7783 10141 7813 ne
rect 10141 7783 10563 7813
tri 10563 7783 10593 7813 sw
tri 10661 7783 10691 7813 ne
rect 10691 7783 11113 7813
tri 11113 7783 11143 7813 sw
tri 11211 7783 11241 7813 ne
rect 11241 7783 11663 7813
tri 11663 7783 11693 7813 sw
tri 11761 7783 11791 7813 ne
rect 11791 7783 12213 7813
tri 12213 7783 12243 7813 sw
tri 12311 7783 12341 7813 ne
rect 12341 7783 12763 7813
tri 12763 7783 12793 7813 sw
tri 12861 7783 12891 7813 ne
rect 12891 7783 13313 7813
tri 13313 7783 13343 7813 sw
tri 13411 7783 13441 7813 ne
rect 13441 7783 13863 7813
tri 13863 7783 13893 7813 sw
tri 13961 7783 13991 7813 ne
rect 13991 7783 14413 7813
tri 14413 7783 14443 7813 sw
tri 14511 7783 14541 7813 ne
rect 14541 7783 14963 7813
tri 14963 7783 14993 7813 sw
tri 15061 7783 15091 7813 ne
rect 15091 7783 15513 7813
tri 15513 7783 15543 7813 sw
tri 15611 7783 15641 7813 ne
rect 15641 7783 16063 7813
tri 16063 7783 16093 7813 sw
tri 16161 7783 16191 7813 ne
rect 16191 7783 16613 7813
tri 16613 7783 16643 7813 sw
tri 16711 7783 16741 7813 ne
rect 16741 7783 17163 7813
tri 17163 7783 17193 7813 sw
tri 17261 7783 17291 7813 ne
rect 17291 7783 17713 7813
tri 17713 7783 17743 7813 sw
tri 17811 7783 17841 7813 ne
rect 17841 7783 18263 7813
tri 18263 7783 18293 7813 sw
tri 18361 7783 18391 7813 ne
rect 18391 7783 18813 7813
tri 18813 7783 18843 7813 sw
tri 18911 7783 18941 7813 ne
rect 18941 7783 19363 7813
tri 19363 7783 19393 7813 sw
tri 19461 7783 19491 7813 ne
rect 19491 7783 20300 7813
rect -2000 7685 143 7783
tri 143 7685 241 7783 sw
tri 241 7685 339 7783 ne
rect 339 7685 693 7783
tri 693 7685 791 7783 sw
tri 791 7685 889 7783 ne
rect 889 7685 1243 7783
tri 1243 7685 1341 7783 sw
tri 1341 7685 1439 7783 ne
rect 1439 7685 1793 7783
tri 1793 7685 1891 7783 sw
tri 1891 7685 1989 7783 ne
rect 1989 7685 2343 7783
tri 2343 7685 2441 7783 sw
tri 2441 7685 2539 7783 ne
rect 2539 7685 2893 7783
tri 2893 7685 2991 7783 sw
tri 2991 7685 3089 7783 ne
rect 3089 7685 3443 7783
tri 3443 7685 3541 7783 sw
tri 3541 7685 3639 7783 ne
rect 3639 7685 3993 7783
tri 3993 7685 4091 7783 sw
tri 4091 7685 4189 7783 ne
rect 4189 7685 4543 7783
tri 4543 7685 4641 7783 sw
tri 4641 7685 4739 7783 ne
rect 4739 7685 5093 7783
tri 5093 7685 5191 7783 sw
tri 5191 7685 5289 7783 ne
rect 5289 7685 5643 7783
tri 5643 7685 5741 7783 sw
tri 5741 7685 5839 7783 ne
rect 5839 7685 6193 7783
tri 6193 7685 6291 7783 sw
tri 6291 7685 6389 7783 ne
rect 6389 7685 6743 7783
tri 6743 7685 6841 7783 sw
tri 6841 7685 6939 7783 ne
rect 6939 7685 7293 7783
tri 7293 7685 7391 7783 sw
tri 7391 7685 7489 7783 ne
rect 7489 7685 7843 7783
tri 7843 7685 7941 7783 sw
tri 7941 7685 8039 7783 ne
rect 8039 7685 8393 7783
tri 8393 7685 8491 7783 sw
tri 8491 7685 8589 7783 ne
rect 8589 7685 8943 7783
tri 8943 7685 9041 7783 sw
tri 9041 7685 9139 7783 ne
rect 9139 7685 9493 7783
tri 9493 7685 9591 7783 sw
tri 9591 7685 9689 7783 ne
rect 9689 7685 10043 7783
tri 10043 7685 10141 7783 sw
tri 10141 7685 10239 7783 ne
rect 10239 7685 10593 7783
tri 10593 7685 10691 7783 sw
tri 10691 7685 10789 7783 ne
rect 10789 7685 11143 7783
tri 11143 7685 11241 7783 sw
tri 11241 7685 11339 7783 ne
rect 11339 7685 11693 7783
tri 11693 7685 11791 7783 sw
tri 11791 7685 11889 7783 ne
rect 11889 7685 12243 7783
tri 12243 7685 12341 7783 sw
tri 12341 7685 12439 7783 ne
rect 12439 7685 12793 7783
tri 12793 7685 12891 7783 sw
tri 12891 7685 12989 7783 ne
rect 12989 7685 13343 7783
tri 13343 7685 13441 7783 sw
tri 13441 7685 13539 7783 ne
rect 13539 7685 13893 7783
tri 13893 7685 13991 7783 sw
tri 13991 7685 14089 7783 ne
rect 14089 7685 14443 7783
tri 14443 7685 14541 7783 sw
tri 14541 7685 14639 7783 ne
rect 14639 7685 14993 7783
tri 14993 7685 15091 7783 sw
tri 15091 7685 15189 7783 ne
rect 15189 7685 15543 7783
tri 15543 7685 15641 7783 sw
tri 15641 7685 15739 7783 ne
rect 15739 7685 16093 7783
tri 16093 7685 16191 7783 sw
tri 16191 7685 16289 7783 ne
rect 16289 7685 16643 7783
tri 16643 7685 16741 7783 sw
tri 16741 7685 16839 7783 ne
rect 16839 7685 17193 7783
tri 17193 7685 17291 7783 sw
tri 17291 7685 17389 7783 ne
rect 17389 7685 17743 7783
tri 17743 7685 17841 7783 sw
tri 17841 7685 17939 7783 ne
rect 17939 7685 18293 7783
tri 18293 7685 18391 7783 sw
tri 18391 7685 18489 7783 ne
rect 18489 7685 18843 7783
tri 18843 7685 18941 7783 sw
tri 18941 7685 19039 7783 ne
rect 19039 7685 19393 7783
tri 19393 7685 19491 7783 sw
tri 19491 7685 19589 7783 ne
rect 19589 7685 20300 7783
rect -2000 7587 241 7685
tri 241 7587 339 7685 sw
tri 339 7587 437 7685 ne
rect 437 7587 791 7685
tri 791 7587 889 7685 sw
tri 889 7587 987 7685 ne
rect 987 7587 1341 7685
tri 1341 7587 1439 7685 sw
tri 1439 7587 1537 7685 ne
rect 1537 7587 1891 7685
tri 1891 7587 1989 7685 sw
tri 1989 7587 2087 7685 ne
rect 2087 7587 2441 7685
tri 2441 7587 2539 7685 sw
tri 2539 7587 2637 7685 ne
rect 2637 7587 2991 7685
tri 2991 7587 3089 7685 sw
tri 3089 7587 3187 7685 ne
rect 3187 7587 3541 7685
tri 3541 7587 3639 7685 sw
tri 3639 7587 3737 7685 ne
rect 3737 7587 4091 7685
tri 4091 7587 4189 7685 sw
tri 4189 7587 4287 7685 ne
rect 4287 7587 4641 7685
tri 4641 7587 4739 7685 sw
tri 4739 7587 4837 7685 ne
rect 4837 7587 5191 7685
tri 5191 7587 5289 7685 sw
tri 5289 7587 5387 7685 ne
rect 5387 7587 5741 7685
tri 5741 7587 5839 7685 sw
tri 5839 7587 5937 7685 ne
rect 5937 7587 6291 7685
tri 6291 7587 6389 7685 sw
tri 6389 7587 6487 7685 ne
rect 6487 7587 6841 7685
tri 6841 7587 6939 7685 sw
tri 6939 7587 7037 7685 ne
rect 7037 7587 7391 7685
tri 7391 7587 7489 7685 sw
tri 7489 7587 7587 7685 ne
rect 7587 7587 7941 7685
tri 7941 7587 8039 7685 sw
tri 8039 7587 8137 7685 ne
rect 8137 7587 8491 7685
tri 8491 7587 8589 7685 sw
tri 8589 7587 8687 7685 ne
rect 8687 7587 9041 7685
tri 9041 7587 9139 7685 sw
tri 9139 7587 9237 7685 ne
rect 9237 7587 9591 7685
tri 9591 7587 9689 7685 sw
tri 9689 7587 9787 7685 ne
rect 9787 7587 10141 7685
tri 10141 7587 10239 7685 sw
tri 10239 7587 10337 7685 ne
rect 10337 7587 10691 7685
tri 10691 7587 10789 7685 sw
tri 10789 7587 10887 7685 ne
rect 10887 7587 11241 7685
tri 11241 7587 11339 7685 sw
tri 11339 7587 11437 7685 ne
rect 11437 7587 11791 7685
tri 11791 7587 11889 7685 sw
tri 11889 7587 11987 7685 ne
rect 11987 7587 12341 7685
tri 12341 7587 12439 7685 sw
tri 12439 7587 12537 7685 ne
rect 12537 7587 12891 7685
tri 12891 7587 12989 7685 sw
tri 12989 7587 13087 7685 ne
rect 13087 7587 13441 7685
tri 13441 7587 13539 7685 sw
tri 13539 7587 13637 7685 ne
rect 13637 7587 13991 7685
tri 13991 7587 14089 7685 sw
tri 14089 7587 14187 7685 ne
rect 14187 7587 14541 7685
tri 14541 7587 14639 7685 sw
tri 14639 7587 14737 7685 ne
rect 14737 7587 15091 7685
tri 15091 7587 15189 7685 sw
tri 15189 7587 15287 7685 ne
rect 15287 7587 15641 7685
tri 15641 7587 15739 7685 sw
tri 15739 7587 15837 7685 ne
rect 15837 7587 16191 7685
tri 16191 7587 16289 7685 sw
tri 16289 7587 16387 7685 ne
rect 16387 7587 16741 7685
tri 16741 7587 16839 7685 sw
tri 16839 7587 16937 7685 ne
rect 16937 7587 17291 7685
tri 17291 7587 17389 7685 sw
tri 17389 7587 17487 7685 ne
rect 17487 7587 17841 7685
tri 17841 7587 17939 7685 sw
tri 17939 7587 18037 7685 ne
rect 18037 7587 18391 7685
tri 18391 7587 18489 7685 sw
tri 18489 7587 18587 7685 ne
rect 18587 7587 18941 7685
tri 18941 7587 19039 7685 sw
tri 19039 7587 19137 7685 ne
rect 19137 7587 19491 7685
tri 19491 7587 19589 7685 sw
tri 19589 7587 19687 7685 ne
rect 19687 7587 20300 7685
rect -2000 7489 339 7587
tri 339 7489 437 7587 sw
tri 437 7489 535 7587 ne
rect 535 7489 889 7587
tri 889 7489 987 7587 sw
tri 987 7489 1085 7587 ne
rect 1085 7489 1439 7587
tri 1439 7489 1537 7587 sw
tri 1537 7489 1635 7587 ne
rect 1635 7489 1989 7587
tri 1989 7489 2087 7587 sw
tri 2087 7489 2185 7587 ne
rect 2185 7489 2539 7587
tri 2539 7489 2637 7587 sw
tri 2637 7489 2735 7587 ne
rect 2735 7489 3089 7587
tri 3089 7489 3187 7587 sw
tri 3187 7489 3285 7587 ne
rect 3285 7489 3639 7587
tri 3639 7489 3737 7587 sw
tri 3737 7489 3835 7587 ne
rect 3835 7489 4189 7587
tri 4189 7489 4287 7587 sw
tri 4287 7489 4385 7587 ne
rect 4385 7489 4739 7587
tri 4739 7489 4837 7587 sw
tri 4837 7489 4935 7587 ne
rect 4935 7489 5289 7587
tri 5289 7489 5387 7587 sw
tri 5387 7489 5485 7587 ne
rect 5485 7489 5839 7587
tri 5839 7489 5937 7587 sw
tri 5937 7489 6035 7587 ne
rect 6035 7489 6389 7587
tri 6389 7489 6487 7587 sw
tri 6487 7489 6585 7587 ne
rect 6585 7489 6939 7587
tri 6939 7489 7037 7587 sw
tri 7037 7489 7135 7587 ne
rect 7135 7489 7489 7587
tri 7489 7489 7587 7587 sw
tri 7587 7489 7685 7587 ne
rect 7685 7489 8039 7587
tri 8039 7489 8137 7587 sw
tri 8137 7489 8235 7587 ne
rect 8235 7489 8589 7587
tri 8589 7489 8687 7587 sw
tri 8687 7489 8785 7587 ne
rect 8785 7489 9139 7587
tri 9139 7489 9237 7587 sw
tri 9237 7489 9335 7587 ne
rect 9335 7489 9689 7587
tri 9689 7489 9787 7587 sw
tri 9787 7489 9885 7587 ne
rect 9885 7489 10239 7587
tri 10239 7489 10337 7587 sw
tri 10337 7489 10435 7587 ne
rect 10435 7489 10789 7587
tri 10789 7489 10887 7587 sw
tri 10887 7489 10985 7587 ne
rect 10985 7489 11339 7587
tri 11339 7489 11437 7587 sw
tri 11437 7489 11535 7587 ne
rect 11535 7489 11889 7587
tri 11889 7489 11987 7587 sw
tri 11987 7489 12085 7587 ne
rect 12085 7489 12439 7587
tri 12439 7489 12537 7587 sw
tri 12537 7489 12635 7587 ne
rect 12635 7489 12989 7587
tri 12989 7489 13087 7587 sw
tri 13087 7489 13185 7587 ne
rect 13185 7489 13539 7587
tri 13539 7489 13637 7587 sw
tri 13637 7489 13735 7587 ne
rect 13735 7489 14089 7587
tri 14089 7489 14187 7587 sw
tri 14187 7489 14285 7587 ne
rect 14285 7489 14639 7587
tri 14639 7489 14737 7587 sw
tri 14737 7489 14835 7587 ne
rect 14835 7489 15189 7587
tri 15189 7489 15287 7587 sw
tri 15287 7489 15385 7587 ne
rect 15385 7489 15739 7587
tri 15739 7489 15837 7587 sw
tri 15837 7489 15935 7587 ne
rect 15935 7489 16289 7587
tri 16289 7489 16387 7587 sw
tri 16387 7489 16485 7587 ne
rect 16485 7489 16839 7587
tri 16839 7489 16937 7587 sw
tri 16937 7489 17035 7587 ne
rect 17035 7489 17389 7587
tri 17389 7489 17487 7587 sw
tri 17487 7489 17585 7587 ne
rect 17585 7489 17939 7587
tri 17939 7489 18037 7587 sw
tri 18037 7489 18135 7587 ne
rect 18135 7489 18489 7587
tri 18489 7489 18587 7587 sw
tri 18587 7489 18685 7587 ne
rect 18685 7489 19039 7587
tri 19039 7489 19137 7587 sw
tri 19137 7489 19235 7587 ne
rect 19235 7489 19589 7587
tri 19589 7489 19687 7587 sw
rect 20800 7489 21800 8137
rect -2000 7485 437 7489
rect -2000 7365 215 7485
rect 335 7391 437 7485
tri 437 7391 535 7489 sw
tri 535 7391 633 7489 ne
rect 633 7485 987 7489
rect 633 7391 765 7485
rect 335 7365 535 7391
rect -2000 7361 535 7365
rect -2000 6713 -1000 7361
tri 113 7263 211 7361 ne
rect 211 7313 535 7361
tri 535 7313 613 7391 sw
tri 633 7313 711 7391 ne
rect 711 7365 765 7391
rect 885 7391 987 7485
tri 987 7391 1085 7489 sw
tri 1085 7391 1183 7489 ne
rect 1183 7485 1537 7489
rect 1183 7391 1315 7485
rect 885 7365 1085 7391
rect 711 7313 1085 7365
tri 1085 7313 1163 7391 sw
tri 1183 7313 1261 7391 ne
rect 1261 7365 1315 7391
rect 1435 7391 1537 7485
tri 1537 7391 1635 7489 sw
tri 1635 7391 1733 7489 ne
rect 1733 7485 2087 7489
rect 1733 7391 1865 7485
rect 1435 7365 1635 7391
rect 1261 7313 1635 7365
tri 1635 7313 1713 7391 sw
tri 1733 7313 1811 7391 ne
rect 1811 7365 1865 7391
rect 1985 7391 2087 7485
tri 2087 7391 2185 7489 sw
tri 2185 7391 2283 7489 ne
rect 2283 7485 2637 7489
rect 2283 7391 2415 7485
rect 1985 7365 2185 7391
rect 1811 7313 2185 7365
tri 2185 7313 2263 7391 sw
tri 2283 7313 2361 7391 ne
rect 2361 7365 2415 7391
rect 2535 7391 2637 7485
tri 2637 7391 2735 7489 sw
tri 2735 7391 2833 7489 ne
rect 2833 7485 3187 7489
rect 2833 7391 2965 7485
rect 2535 7365 2735 7391
rect 2361 7313 2735 7365
tri 2735 7313 2813 7391 sw
tri 2833 7313 2911 7391 ne
rect 2911 7365 2965 7391
rect 3085 7391 3187 7485
tri 3187 7391 3285 7489 sw
tri 3285 7391 3383 7489 ne
rect 3383 7485 3737 7489
rect 3383 7391 3515 7485
rect 3085 7365 3285 7391
rect 2911 7313 3285 7365
tri 3285 7313 3363 7391 sw
tri 3383 7313 3461 7391 ne
rect 3461 7365 3515 7391
rect 3635 7391 3737 7485
tri 3737 7391 3835 7489 sw
tri 3835 7391 3933 7489 ne
rect 3933 7485 4287 7489
rect 3933 7391 4065 7485
rect 3635 7365 3835 7391
rect 3461 7313 3835 7365
tri 3835 7313 3913 7391 sw
tri 3933 7313 4011 7391 ne
rect 4011 7365 4065 7391
rect 4185 7391 4287 7485
tri 4287 7391 4385 7489 sw
tri 4385 7391 4483 7489 ne
rect 4483 7485 4837 7489
rect 4483 7391 4615 7485
rect 4185 7365 4385 7391
rect 4011 7313 4385 7365
tri 4385 7313 4463 7391 sw
tri 4483 7313 4561 7391 ne
rect 4561 7365 4615 7391
rect 4735 7391 4837 7485
tri 4837 7391 4935 7489 sw
tri 4935 7391 5033 7489 ne
rect 5033 7485 5387 7489
rect 5033 7391 5165 7485
rect 4735 7365 4935 7391
rect 4561 7313 4935 7365
tri 4935 7313 5013 7391 sw
tri 5033 7313 5111 7391 ne
rect 5111 7365 5165 7391
rect 5285 7391 5387 7485
tri 5387 7391 5485 7489 sw
tri 5485 7391 5583 7489 ne
rect 5583 7485 5937 7489
rect 5583 7391 5715 7485
rect 5285 7365 5485 7391
rect 5111 7313 5485 7365
tri 5485 7313 5563 7391 sw
tri 5583 7313 5661 7391 ne
rect 5661 7365 5715 7391
rect 5835 7391 5937 7485
tri 5937 7391 6035 7489 sw
tri 6035 7391 6133 7489 ne
rect 6133 7485 6487 7489
rect 6133 7391 6265 7485
rect 5835 7365 6035 7391
rect 5661 7313 6035 7365
tri 6035 7313 6113 7391 sw
tri 6133 7313 6211 7391 ne
rect 6211 7365 6265 7391
rect 6385 7391 6487 7485
tri 6487 7391 6585 7489 sw
tri 6585 7391 6683 7489 ne
rect 6683 7485 7037 7489
rect 6683 7391 6815 7485
rect 6385 7365 6585 7391
rect 6211 7313 6585 7365
tri 6585 7313 6663 7391 sw
tri 6683 7313 6761 7391 ne
rect 6761 7365 6815 7391
rect 6935 7391 7037 7485
tri 7037 7391 7135 7489 sw
tri 7135 7391 7233 7489 ne
rect 7233 7485 7587 7489
rect 7233 7391 7365 7485
rect 6935 7365 7135 7391
rect 6761 7313 7135 7365
tri 7135 7313 7213 7391 sw
tri 7233 7313 7311 7391 ne
rect 7311 7365 7365 7391
rect 7485 7391 7587 7485
tri 7587 7391 7685 7489 sw
tri 7685 7391 7783 7489 ne
rect 7783 7485 8137 7489
rect 7783 7391 7915 7485
rect 7485 7365 7685 7391
rect 7311 7313 7685 7365
tri 7685 7313 7763 7391 sw
tri 7783 7313 7861 7391 ne
rect 7861 7365 7915 7391
rect 8035 7391 8137 7485
tri 8137 7391 8235 7489 sw
tri 8235 7391 8333 7489 ne
rect 8333 7485 8687 7489
rect 8333 7391 8465 7485
rect 8035 7365 8235 7391
rect 7861 7313 8235 7365
tri 8235 7313 8313 7391 sw
tri 8333 7313 8411 7391 ne
rect 8411 7365 8465 7391
rect 8585 7391 8687 7485
tri 8687 7391 8785 7489 sw
tri 8785 7391 8883 7489 ne
rect 8883 7485 9237 7489
rect 8883 7391 9015 7485
rect 8585 7365 8785 7391
rect 8411 7313 8785 7365
tri 8785 7313 8863 7391 sw
tri 8883 7313 8961 7391 ne
rect 8961 7365 9015 7391
rect 9135 7391 9237 7485
tri 9237 7391 9335 7489 sw
tri 9335 7391 9433 7489 ne
rect 9433 7485 9787 7489
rect 9433 7391 9565 7485
rect 9135 7365 9335 7391
rect 8961 7313 9335 7365
tri 9335 7313 9413 7391 sw
tri 9433 7313 9511 7391 ne
rect 9511 7365 9565 7391
rect 9685 7391 9787 7485
tri 9787 7391 9885 7489 sw
tri 9885 7391 9983 7489 ne
rect 9983 7485 10337 7489
rect 9983 7391 10115 7485
rect 9685 7365 9885 7391
rect 9511 7313 9885 7365
tri 9885 7313 9963 7391 sw
tri 9983 7313 10061 7391 ne
rect 10061 7365 10115 7391
rect 10235 7391 10337 7485
tri 10337 7391 10435 7489 sw
tri 10435 7391 10533 7489 ne
rect 10533 7485 10887 7489
rect 10533 7391 10665 7485
rect 10235 7365 10435 7391
rect 10061 7313 10435 7365
tri 10435 7313 10513 7391 sw
tri 10533 7313 10611 7391 ne
rect 10611 7365 10665 7391
rect 10785 7391 10887 7485
tri 10887 7391 10985 7489 sw
tri 10985 7391 11083 7489 ne
rect 11083 7485 11437 7489
rect 11083 7391 11215 7485
rect 10785 7365 10985 7391
rect 10611 7313 10985 7365
tri 10985 7313 11063 7391 sw
tri 11083 7313 11161 7391 ne
rect 11161 7365 11215 7391
rect 11335 7391 11437 7485
tri 11437 7391 11535 7489 sw
tri 11535 7391 11633 7489 ne
rect 11633 7485 11987 7489
rect 11633 7391 11765 7485
rect 11335 7365 11535 7391
rect 11161 7313 11535 7365
tri 11535 7313 11613 7391 sw
tri 11633 7313 11711 7391 ne
rect 11711 7365 11765 7391
rect 11885 7391 11987 7485
tri 11987 7391 12085 7489 sw
tri 12085 7391 12183 7489 ne
rect 12183 7485 12537 7489
rect 12183 7391 12315 7485
rect 11885 7365 12085 7391
rect 11711 7313 12085 7365
tri 12085 7313 12163 7391 sw
tri 12183 7313 12261 7391 ne
rect 12261 7365 12315 7391
rect 12435 7391 12537 7485
tri 12537 7391 12635 7489 sw
tri 12635 7391 12733 7489 ne
rect 12733 7485 13087 7489
rect 12733 7391 12865 7485
rect 12435 7365 12635 7391
rect 12261 7313 12635 7365
tri 12635 7313 12713 7391 sw
tri 12733 7313 12811 7391 ne
rect 12811 7365 12865 7391
rect 12985 7391 13087 7485
tri 13087 7391 13185 7489 sw
tri 13185 7391 13283 7489 ne
rect 13283 7485 13637 7489
rect 13283 7391 13415 7485
rect 12985 7365 13185 7391
rect 12811 7313 13185 7365
tri 13185 7313 13263 7391 sw
tri 13283 7313 13361 7391 ne
rect 13361 7365 13415 7391
rect 13535 7391 13637 7485
tri 13637 7391 13735 7489 sw
tri 13735 7391 13833 7489 ne
rect 13833 7485 14187 7489
rect 13833 7391 13965 7485
rect 13535 7365 13735 7391
rect 13361 7313 13735 7365
tri 13735 7313 13813 7391 sw
tri 13833 7313 13911 7391 ne
rect 13911 7365 13965 7391
rect 14085 7391 14187 7485
tri 14187 7391 14285 7489 sw
tri 14285 7391 14383 7489 ne
rect 14383 7485 14737 7489
rect 14383 7391 14515 7485
rect 14085 7365 14285 7391
rect 13911 7313 14285 7365
tri 14285 7313 14363 7391 sw
tri 14383 7313 14461 7391 ne
rect 14461 7365 14515 7391
rect 14635 7391 14737 7485
tri 14737 7391 14835 7489 sw
tri 14835 7391 14933 7489 ne
rect 14933 7485 15287 7489
rect 14933 7391 15065 7485
rect 14635 7365 14835 7391
rect 14461 7313 14835 7365
tri 14835 7313 14913 7391 sw
tri 14933 7313 15011 7391 ne
rect 15011 7365 15065 7391
rect 15185 7391 15287 7485
tri 15287 7391 15385 7489 sw
tri 15385 7391 15483 7489 ne
rect 15483 7485 15837 7489
rect 15483 7391 15615 7485
rect 15185 7365 15385 7391
rect 15011 7313 15385 7365
tri 15385 7313 15463 7391 sw
tri 15483 7313 15561 7391 ne
rect 15561 7365 15615 7391
rect 15735 7391 15837 7485
tri 15837 7391 15935 7489 sw
tri 15935 7391 16033 7489 ne
rect 16033 7485 16387 7489
rect 16033 7391 16165 7485
rect 15735 7365 15935 7391
rect 15561 7313 15935 7365
tri 15935 7313 16013 7391 sw
tri 16033 7313 16111 7391 ne
rect 16111 7365 16165 7391
rect 16285 7391 16387 7485
tri 16387 7391 16485 7489 sw
tri 16485 7391 16583 7489 ne
rect 16583 7485 16937 7489
rect 16583 7391 16715 7485
rect 16285 7365 16485 7391
rect 16111 7313 16485 7365
tri 16485 7313 16563 7391 sw
tri 16583 7313 16661 7391 ne
rect 16661 7365 16715 7391
rect 16835 7391 16937 7485
tri 16937 7391 17035 7489 sw
tri 17035 7391 17133 7489 ne
rect 17133 7485 17487 7489
rect 17133 7391 17265 7485
rect 16835 7365 17035 7391
rect 16661 7313 17035 7365
tri 17035 7313 17113 7391 sw
tri 17133 7313 17211 7391 ne
rect 17211 7365 17265 7391
rect 17385 7391 17487 7485
tri 17487 7391 17585 7489 sw
tri 17585 7391 17683 7489 ne
rect 17683 7485 18037 7489
rect 17683 7391 17815 7485
rect 17385 7365 17585 7391
rect 17211 7313 17585 7365
tri 17585 7313 17663 7391 sw
tri 17683 7313 17761 7391 ne
rect 17761 7365 17815 7391
rect 17935 7391 18037 7485
tri 18037 7391 18135 7489 sw
tri 18135 7391 18233 7489 ne
rect 18233 7485 18587 7489
rect 18233 7391 18365 7485
rect 17935 7365 18135 7391
rect 17761 7313 18135 7365
tri 18135 7313 18213 7391 sw
tri 18233 7313 18311 7391 ne
rect 18311 7365 18365 7391
rect 18485 7391 18587 7485
tri 18587 7391 18685 7489 sw
tri 18685 7391 18783 7489 ne
rect 18783 7485 19137 7489
rect 18783 7391 18915 7485
rect 18485 7365 18685 7391
rect 18311 7313 18685 7365
tri 18685 7313 18763 7391 sw
tri 18783 7313 18861 7391 ne
rect 18861 7365 18915 7391
rect 19035 7391 19137 7485
tri 19137 7391 19235 7489 sw
tri 19235 7391 19333 7489 ne
rect 19333 7485 21800 7489
rect 19333 7391 19465 7485
rect 19035 7365 19235 7391
rect 18861 7313 19235 7365
tri 19235 7313 19313 7391 sw
tri 19333 7313 19411 7391 ne
rect 19411 7365 19465 7391
rect 19585 7365 21800 7485
rect 19411 7313 21800 7365
rect 211 7263 613 7313
rect -500 7213 113 7263
tri 113 7213 163 7263 sw
tri 211 7213 261 7263 ne
rect 261 7233 613 7263
tri 613 7233 693 7313 sw
tri 711 7233 791 7313 ne
rect 791 7233 1163 7313
tri 1163 7233 1243 7313 sw
tri 1261 7233 1341 7313 ne
rect 1341 7233 1713 7313
tri 1713 7233 1793 7313 sw
tri 1811 7233 1891 7313 ne
rect 1891 7233 2263 7313
tri 2263 7233 2343 7313 sw
tri 2361 7233 2441 7313 ne
rect 2441 7233 2813 7313
tri 2813 7233 2893 7313 sw
tri 2911 7233 2991 7313 ne
rect 2991 7233 3363 7313
tri 3363 7233 3443 7313 sw
tri 3461 7233 3541 7313 ne
rect 3541 7233 3913 7313
tri 3913 7233 3993 7313 sw
tri 4011 7233 4091 7313 ne
rect 4091 7233 4463 7313
tri 4463 7233 4543 7313 sw
tri 4561 7233 4641 7313 ne
rect 4641 7233 5013 7313
tri 5013 7233 5093 7313 sw
tri 5111 7233 5191 7313 ne
rect 5191 7233 5563 7313
tri 5563 7233 5643 7313 sw
tri 5661 7233 5741 7313 ne
rect 5741 7233 6113 7313
tri 6113 7233 6193 7313 sw
tri 6211 7233 6291 7313 ne
rect 6291 7233 6663 7313
tri 6663 7233 6743 7313 sw
tri 6761 7233 6841 7313 ne
rect 6841 7233 7213 7313
tri 7213 7233 7293 7313 sw
tri 7311 7233 7391 7313 ne
rect 7391 7233 7763 7313
tri 7763 7233 7843 7313 sw
tri 7861 7233 7941 7313 ne
rect 7941 7233 8313 7313
tri 8313 7233 8393 7313 sw
tri 8411 7233 8491 7313 ne
rect 8491 7233 8863 7313
tri 8863 7233 8943 7313 sw
tri 8961 7233 9041 7313 ne
rect 9041 7233 9413 7313
tri 9413 7233 9493 7313 sw
tri 9511 7233 9591 7313 ne
rect 9591 7233 9963 7313
tri 9963 7233 10043 7313 sw
tri 10061 7233 10141 7313 ne
rect 10141 7233 10513 7313
tri 10513 7233 10593 7313 sw
tri 10611 7233 10691 7313 ne
rect 10691 7233 11063 7313
tri 11063 7233 11143 7313 sw
tri 11161 7233 11241 7313 ne
rect 11241 7233 11613 7313
tri 11613 7233 11693 7313 sw
tri 11711 7233 11791 7313 ne
rect 11791 7233 12163 7313
tri 12163 7233 12243 7313 sw
tri 12261 7233 12341 7313 ne
rect 12341 7233 12713 7313
tri 12713 7233 12793 7313 sw
tri 12811 7233 12891 7313 ne
rect 12891 7233 13263 7313
tri 13263 7233 13343 7313 sw
tri 13361 7233 13441 7313 ne
rect 13441 7233 13813 7313
tri 13813 7233 13893 7313 sw
tri 13911 7233 13991 7313 ne
rect 13991 7233 14363 7313
tri 14363 7233 14443 7313 sw
tri 14461 7233 14541 7313 ne
rect 14541 7233 14913 7313
tri 14913 7233 14993 7313 sw
tri 15011 7233 15091 7313 ne
rect 15091 7233 15463 7313
tri 15463 7233 15543 7313 sw
tri 15561 7233 15641 7313 ne
rect 15641 7233 16013 7313
tri 16013 7233 16093 7313 sw
tri 16111 7233 16191 7313 ne
rect 16191 7233 16563 7313
tri 16563 7233 16643 7313 sw
tri 16661 7233 16741 7313 ne
rect 16741 7233 17113 7313
tri 17113 7233 17193 7313 sw
tri 17211 7233 17291 7313 ne
rect 17291 7233 17663 7313
tri 17663 7233 17743 7313 sw
tri 17761 7233 17841 7313 ne
rect 17841 7233 18213 7313
tri 18213 7233 18293 7313 sw
tri 18311 7233 18391 7313 ne
rect 18391 7233 18763 7313
tri 18763 7233 18843 7313 sw
tri 18861 7233 18941 7313 ne
rect 18941 7233 19313 7313
tri 19313 7233 19393 7313 sw
tri 19411 7233 19491 7313 ne
rect 19491 7233 20100 7313
rect 261 7213 693 7233
rect -500 7135 163 7213
tri 163 7135 241 7213 sw
tri 261 7135 339 7213 ne
rect 339 7135 693 7213
tri 693 7135 791 7233 sw
tri 791 7135 889 7233 ne
rect 889 7135 1243 7233
tri 1243 7135 1341 7233 sw
tri 1341 7135 1439 7233 ne
rect 1439 7135 1793 7233
tri 1793 7135 1891 7233 sw
tri 1891 7135 1989 7233 ne
rect 1989 7135 2343 7233
tri 2343 7135 2441 7233 sw
tri 2441 7135 2539 7233 ne
rect 2539 7135 2893 7233
tri 2893 7135 2991 7233 sw
tri 2991 7135 3089 7233 ne
rect 3089 7135 3443 7233
tri 3443 7135 3541 7233 sw
tri 3541 7135 3639 7233 ne
rect 3639 7135 3993 7233
tri 3993 7135 4091 7233 sw
tri 4091 7135 4189 7233 ne
rect 4189 7135 4543 7233
tri 4543 7135 4641 7233 sw
tri 4641 7135 4739 7233 ne
rect 4739 7135 5093 7233
tri 5093 7135 5191 7233 sw
tri 5191 7135 5289 7233 ne
rect 5289 7135 5643 7233
tri 5643 7135 5741 7233 sw
tri 5741 7135 5839 7233 ne
rect 5839 7135 6193 7233
tri 6193 7135 6291 7233 sw
tri 6291 7135 6389 7233 ne
rect 6389 7135 6743 7233
tri 6743 7135 6841 7233 sw
tri 6841 7135 6939 7233 ne
rect 6939 7135 7293 7233
tri 7293 7135 7391 7233 sw
tri 7391 7135 7489 7233 ne
rect 7489 7135 7843 7233
tri 7843 7135 7941 7233 sw
tri 7941 7135 8039 7233 ne
rect 8039 7135 8393 7233
tri 8393 7135 8491 7233 sw
tri 8491 7135 8589 7233 ne
rect 8589 7135 8943 7233
tri 8943 7135 9041 7233 sw
tri 9041 7135 9139 7233 ne
rect 9139 7135 9493 7233
tri 9493 7135 9591 7233 sw
tri 9591 7135 9689 7233 ne
rect 9689 7135 10043 7233
tri 10043 7135 10141 7233 sw
tri 10141 7135 10239 7233 ne
rect 10239 7135 10593 7233
tri 10593 7135 10691 7233 sw
tri 10691 7135 10789 7233 ne
rect 10789 7135 11143 7233
tri 11143 7135 11241 7233 sw
tri 11241 7135 11339 7233 ne
rect 11339 7135 11693 7233
tri 11693 7135 11791 7233 sw
tri 11791 7135 11889 7233 ne
rect 11889 7135 12243 7233
tri 12243 7135 12341 7233 sw
tri 12341 7135 12439 7233 ne
rect 12439 7135 12793 7233
tri 12793 7135 12891 7233 sw
tri 12891 7135 12989 7233 ne
rect 12989 7135 13343 7233
tri 13343 7135 13441 7233 sw
tri 13441 7135 13539 7233 ne
rect 13539 7135 13893 7233
tri 13893 7135 13991 7233 sw
tri 13991 7135 14089 7233 ne
rect 14089 7135 14443 7233
tri 14443 7135 14541 7233 sw
tri 14541 7135 14639 7233 ne
rect 14639 7135 14993 7233
tri 14993 7135 15091 7233 sw
tri 15091 7135 15189 7233 ne
rect 15189 7135 15543 7233
tri 15543 7135 15641 7233 sw
tri 15641 7135 15739 7233 ne
rect 15739 7135 16093 7233
tri 16093 7135 16191 7233 sw
tri 16191 7135 16289 7233 ne
rect 16289 7135 16643 7233
tri 16643 7135 16741 7233 sw
tri 16741 7135 16839 7233 ne
rect 16839 7135 17193 7233
tri 17193 7135 17291 7233 sw
tri 17291 7135 17389 7233 ne
rect 17389 7135 17743 7233
tri 17743 7135 17841 7233 sw
tri 17841 7135 17939 7233 ne
rect 17939 7135 18293 7233
tri 18293 7135 18391 7233 sw
tri 18391 7135 18489 7233 ne
rect 18489 7135 18843 7233
tri 18843 7135 18941 7233 sw
tri 18941 7135 19039 7233 ne
rect 19039 7135 19393 7233
tri 19393 7135 19491 7233 sw
tri 19491 7135 19589 7233 ne
rect 19589 7213 20100 7233
rect 20200 7213 21800 7313
rect 19589 7135 21800 7213
rect -500 7087 241 7135
rect -500 6987 -400 7087
rect -300 7037 241 7087
tri 241 7037 339 7135 sw
tri 339 7037 437 7135 ne
rect 437 7037 791 7135
tri 791 7037 889 7135 sw
tri 889 7037 987 7135 ne
rect 987 7037 1341 7135
tri 1341 7037 1439 7135 sw
tri 1439 7037 1537 7135 ne
rect 1537 7037 1891 7135
tri 1891 7037 1989 7135 sw
tri 1989 7037 2087 7135 ne
rect 2087 7037 2441 7135
tri 2441 7037 2539 7135 sw
tri 2539 7037 2637 7135 ne
rect 2637 7037 2991 7135
tri 2991 7037 3089 7135 sw
tri 3089 7037 3187 7135 ne
rect 3187 7037 3541 7135
tri 3541 7037 3639 7135 sw
tri 3639 7037 3737 7135 ne
rect 3737 7037 4091 7135
tri 4091 7037 4189 7135 sw
tri 4189 7037 4287 7135 ne
rect 4287 7037 4641 7135
tri 4641 7037 4739 7135 sw
tri 4739 7037 4837 7135 ne
rect 4837 7037 5191 7135
tri 5191 7037 5289 7135 sw
tri 5289 7037 5387 7135 ne
rect 5387 7037 5741 7135
tri 5741 7037 5839 7135 sw
tri 5839 7037 5937 7135 ne
rect 5937 7037 6291 7135
tri 6291 7037 6389 7135 sw
tri 6389 7037 6487 7135 ne
rect 6487 7037 6841 7135
tri 6841 7037 6939 7135 sw
tri 6939 7037 7037 7135 ne
rect 7037 7037 7391 7135
tri 7391 7037 7489 7135 sw
tri 7489 7037 7587 7135 ne
rect 7587 7037 7941 7135
tri 7941 7037 8039 7135 sw
tri 8039 7037 8137 7135 ne
rect 8137 7037 8491 7135
tri 8491 7037 8589 7135 sw
tri 8589 7037 8687 7135 ne
rect 8687 7037 9041 7135
tri 9041 7037 9139 7135 sw
tri 9139 7037 9237 7135 ne
rect 9237 7037 9591 7135
tri 9591 7037 9689 7135 sw
tri 9689 7037 9787 7135 ne
rect 9787 7037 10141 7135
tri 10141 7037 10239 7135 sw
tri 10239 7037 10337 7135 ne
rect 10337 7037 10691 7135
tri 10691 7037 10789 7135 sw
tri 10789 7037 10887 7135 ne
rect 10887 7037 11241 7135
tri 11241 7037 11339 7135 sw
tri 11339 7037 11437 7135 ne
rect 11437 7037 11791 7135
tri 11791 7037 11889 7135 sw
tri 11889 7037 11987 7135 ne
rect 11987 7037 12341 7135
tri 12341 7037 12439 7135 sw
tri 12439 7037 12537 7135 ne
rect 12537 7037 12891 7135
tri 12891 7037 12989 7135 sw
tri 12989 7037 13087 7135 ne
rect 13087 7037 13441 7135
tri 13441 7037 13539 7135 sw
tri 13539 7037 13637 7135 ne
rect 13637 7037 13991 7135
tri 13991 7037 14089 7135 sw
tri 14089 7037 14187 7135 ne
rect 14187 7037 14541 7135
tri 14541 7037 14639 7135 sw
tri 14639 7037 14737 7135 ne
rect 14737 7037 15091 7135
tri 15091 7037 15189 7135 sw
tri 15189 7037 15287 7135 ne
rect 15287 7037 15641 7135
tri 15641 7037 15739 7135 sw
tri 15739 7037 15837 7135 ne
rect 15837 7037 16191 7135
tri 16191 7037 16289 7135 sw
tri 16289 7037 16387 7135 ne
rect 16387 7037 16741 7135
tri 16741 7037 16839 7135 sw
tri 16839 7037 16937 7135 ne
rect 16937 7037 17291 7135
tri 17291 7037 17389 7135 sw
tri 17389 7037 17487 7135 ne
rect 17487 7037 17841 7135
tri 17841 7037 17939 7135 sw
tri 17939 7037 18037 7135 ne
rect 18037 7037 18391 7135
tri 18391 7037 18489 7135 sw
tri 18489 7037 18587 7135 ne
rect 18587 7037 18941 7135
tri 18941 7037 19039 7135 sw
tri 19039 7037 19137 7135 ne
rect 19137 7037 19491 7135
tri 19491 7037 19589 7135 sw
tri 19589 7037 19687 7135 ne
rect 19687 7037 21800 7135
rect -300 6987 339 7037
rect -500 6939 339 6987
tri 339 6939 437 7037 sw
tri 437 6939 535 7037 ne
rect 535 6939 889 7037
tri 889 6939 987 7037 sw
tri 987 6939 1085 7037 ne
rect 1085 6939 1439 7037
tri 1439 6939 1537 7037 sw
tri 1537 6939 1635 7037 ne
rect 1635 6939 1989 7037
tri 1989 6939 2087 7037 sw
tri 2087 6939 2185 7037 ne
rect 2185 6939 2539 7037
tri 2539 6939 2637 7037 sw
tri 2637 6939 2735 7037 ne
rect 2735 6939 3089 7037
tri 3089 6939 3187 7037 sw
tri 3187 6939 3285 7037 ne
rect 3285 6939 3639 7037
tri 3639 6939 3737 7037 sw
tri 3737 6939 3835 7037 ne
rect 3835 6939 4189 7037
tri 4189 6939 4287 7037 sw
tri 4287 6939 4385 7037 ne
rect 4385 6939 4739 7037
tri 4739 6939 4837 7037 sw
tri 4837 6939 4935 7037 ne
rect 4935 6939 5289 7037
tri 5289 6939 5387 7037 sw
tri 5387 6939 5485 7037 ne
rect 5485 6939 5839 7037
tri 5839 6939 5937 7037 sw
tri 5937 6939 6035 7037 ne
rect 6035 6939 6389 7037
tri 6389 6939 6487 7037 sw
tri 6487 6939 6585 7037 ne
rect 6585 6939 6939 7037
tri 6939 6939 7037 7037 sw
tri 7037 6939 7135 7037 ne
rect 7135 6939 7489 7037
tri 7489 6939 7587 7037 sw
tri 7587 6939 7685 7037 ne
rect 7685 6939 8039 7037
tri 8039 6939 8137 7037 sw
tri 8137 6939 8235 7037 ne
rect 8235 6939 8589 7037
tri 8589 6939 8687 7037 sw
tri 8687 6939 8785 7037 ne
rect 8785 6939 9139 7037
tri 9139 6939 9237 7037 sw
tri 9237 6939 9335 7037 ne
rect 9335 6939 9689 7037
tri 9689 6939 9787 7037 sw
tri 9787 6939 9885 7037 ne
rect 9885 6939 10239 7037
tri 10239 6939 10337 7037 sw
tri 10337 6939 10435 7037 ne
rect 10435 6939 10789 7037
tri 10789 6939 10887 7037 sw
tri 10887 6939 10985 7037 ne
rect 10985 6939 11339 7037
tri 11339 6939 11437 7037 sw
tri 11437 6939 11535 7037 ne
rect 11535 6939 11889 7037
tri 11889 6939 11987 7037 sw
tri 11987 6939 12085 7037 ne
rect 12085 6939 12439 7037
tri 12439 6939 12537 7037 sw
tri 12537 6939 12635 7037 ne
rect 12635 6939 12989 7037
tri 12989 6939 13087 7037 sw
tri 13087 6939 13185 7037 ne
rect 13185 6939 13539 7037
tri 13539 6939 13637 7037 sw
tri 13637 6939 13735 7037 ne
rect 13735 6939 14089 7037
tri 14089 6939 14187 7037 sw
tri 14187 6939 14285 7037 ne
rect 14285 6939 14639 7037
tri 14639 6939 14737 7037 sw
tri 14737 6939 14835 7037 ne
rect 14835 6939 15189 7037
tri 15189 6939 15287 7037 sw
tri 15287 6939 15385 7037 ne
rect 15385 6939 15739 7037
tri 15739 6939 15837 7037 sw
tri 15837 6939 15935 7037 ne
rect 15935 6939 16289 7037
tri 16289 6939 16387 7037 sw
tri 16387 6939 16485 7037 ne
rect 16485 6939 16839 7037
tri 16839 6939 16937 7037 sw
tri 16937 6939 17035 7037 ne
rect 17035 6939 17389 7037
tri 17389 6939 17487 7037 sw
tri 17487 6939 17585 7037 ne
rect 17585 6939 17939 7037
tri 17939 6939 18037 7037 sw
tri 18037 6939 18135 7037 ne
rect 18135 6939 18489 7037
tri 18489 6939 18587 7037 sw
tri 18587 6939 18685 7037 ne
rect 18685 6939 19039 7037
tri 19039 6939 19137 7037 sw
tri 19137 6939 19235 7037 ne
rect 19235 6939 19589 7037
tri 19589 6939 19687 7037 sw
rect -500 6935 437 6939
rect -500 6815 215 6935
rect 335 6841 437 6935
tri 437 6841 535 6939 sw
tri 535 6841 633 6939 ne
rect 633 6935 987 6939
rect 633 6841 765 6935
rect 335 6815 535 6841
rect -500 6811 535 6815
tri 535 6811 565 6841 sw
tri 633 6811 663 6841 ne
rect 663 6815 765 6841
rect 885 6841 987 6935
tri 987 6841 1085 6939 sw
tri 1085 6841 1183 6939 ne
rect 1183 6935 1537 6939
rect 1183 6841 1315 6935
rect 885 6815 1085 6841
rect 663 6811 1085 6815
tri 1085 6811 1115 6841 sw
tri 1183 6811 1213 6841 ne
rect 1213 6815 1315 6841
rect 1435 6841 1537 6935
tri 1537 6841 1635 6939 sw
tri 1635 6841 1733 6939 ne
rect 1733 6935 2087 6939
rect 1733 6841 1865 6935
rect 1435 6815 1635 6841
rect 1213 6811 1635 6815
tri 1635 6811 1665 6841 sw
tri 1733 6811 1763 6841 ne
rect 1763 6815 1865 6841
rect 1985 6841 2087 6935
tri 2087 6841 2185 6939 sw
tri 2185 6841 2283 6939 ne
rect 2283 6935 2637 6939
rect 2283 6841 2415 6935
rect 1985 6815 2185 6841
rect 1763 6811 2185 6815
tri 2185 6811 2215 6841 sw
tri 2283 6811 2313 6841 ne
rect 2313 6815 2415 6841
rect 2535 6841 2637 6935
tri 2637 6841 2735 6939 sw
tri 2735 6841 2833 6939 ne
rect 2833 6935 3187 6939
rect 2833 6841 2965 6935
rect 2535 6815 2735 6841
rect 2313 6811 2735 6815
tri 2735 6811 2765 6841 sw
tri 2833 6811 2863 6841 ne
rect 2863 6815 2965 6841
rect 3085 6841 3187 6935
tri 3187 6841 3285 6939 sw
tri 3285 6841 3383 6939 ne
rect 3383 6935 3737 6939
rect 3383 6841 3515 6935
rect 3085 6815 3285 6841
rect 2863 6811 3285 6815
tri 3285 6811 3315 6841 sw
tri 3383 6811 3413 6841 ne
rect 3413 6815 3515 6841
rect 3635 6841 3737 6935
tri 3737 6841 3835 6939 sw
tri 3835 6841 3933 6939 ne
rect 3933 6935 4287 6939
rect 3933 6841 4065 6935
rect 3635 6815 3835 6841
rect 3413 6811 3835 6815
tri 3835 6811 3865 6841 sw
tri 3933 6811 3963 6841 ne
rect 3963 6815 4065 6841
rect 4185 6841 4287 6935
tri 4287 6841 4385 6939 sw
tri 4385 6841 4483 6939 ne
rect 4483 6935 4837 6939
rect 4483 6841 4615 6935
rect 4185 6815 4385 6841
rect 3963 6811 4385 6815
tri 4385 6811 4415 6841 sw
tri 4483 6811 4513 6841 ne
rect 4513 6815 4615 6841
rect 4735 6841 4837 6935
tri 4837 6841 4935 6939 sw
tri 4935 6841 5033 6939 ne
rect 5033 6935 5387 6939
rect 5033 6841 5165 6935
rect 4735 6815 4935 6841
rect 4513 6811 4935 6815
tri 4935 6811 4965 6841 sw
tri 5033 6811 5063 6841 ne
rect 5063 6815 5165 6841
rect 5285 6841 5387 6935
tri 5387 6841 5485 6939 sw
tri 5485 6841 5583 6939 ne
rect 5583 6935 5937 6939
rect 5583 6841 5715 6935
rect 5285 6815 5485 6841
rect 5063 6811 5485 6815
tri 5485 6811 5515 6841 sw
tri 5583 6811 5613 6841 ne
rect 5613 6815 5715 6841
rect 5835 6841 5937 6935
tri 5937 6841 6035 6939 sw
tri 6035 6841 6133 6939 ne
rect 6133 6935 6487 6939
rect 6133 6841 6265 6935
rect 5835 6815 6035 6841
rect 5613 6811 6035 6815
tri 6035 6811 6065 6841 sw
tri 6133 6811 6163 6841 ne
rect 6163 6815 6265 6841
rect 6385 6841 6487 6935
tri 6487 6841 6585 6939 sw
tri 6585 6841 6683 6939 ne
rect 6683 6935 7037 6939
rect 6683 6841 6815 6935
rect 6385 6815 6585 6841
rect 6163 6811 6585 6815
tri 6585 6811 6615 6841 sw
tri 6683 6811 6713 6841 ne
rect 6713 6815 6815 6841
rect 6935 6841 7037 6935
tri 7037 6841 7135 6939 sw
tri 7135 6841 7233 6939 ne
rect 7233 6935 7587 6939
rect 7233 6841 7365 6935
rect 6935 6815 7135 6841
rect 6713 6811 7135 6815
tri 7135 6811 7165 6841 sw
tri 7233 6811 7263 6841 ne
rect 7263 6815 7365 6841
rect 7485 6841 7587 6935
tri 7587 6841 7685 6939 sw
tri 7685 6841 7783 6939 ne
rect 7783 6935 8137 6939
rect 7783 6841 7915 6935
rect 7485 6815 7685 6841
rect 7263 6811 7685 6815
tri 7685 6811 7715 6841 sw
tri 7783 6811 7813 6841 ne
rect 7813 6815 7915 6841
rect 8035 6841 8137 6935
tri 8137 6841 8235 6939 sw
tri 8235 6841 8333 6939 ne
rect 8333 6935 8687 6939
rect 8333 6841 8465 6935
rect 8035 6815 8235 6841
rect 7813 6811 8235 6815
tri 8235 6811 8265 6841 sw
tri 8333 6811 8363 6841 ne
rect 8363 6815 8465 6841
rect 8585 6841 8687 6935
tri 8687 6841 8785 6939 sw
tri 8785 6841 8883 6939 ne
rect 8883 6935 9237 6939
rect 8883 6841 9015 6935
rect 8585 6815 8785 6841
rect 8363 6811 8785 6815
tri 8785 6811 8815 6841 sw
tri 8883 6811 8913 6841 ne
rect 8913 6815 9015 6841
rect 9135 6841 9237 6935
tri 9237 6841 9335 6939 sw
tri 9335 6841 9433 6939 ne
rect 9433 6935 9787 6939
rect 9433 6841 9565 6935
rect 9135 6815 9335 6841
rect 8913 6811 9335 6815
tri 9335 6811 9365 6841 sw
tri 9433 6811 9463 6841 ne
rect 9463 6815 9565 6841
rect 9685 6841 9787 6935
tri 9787 6841 9885 6939 sw
tri 9885 6841 9983 6939 ne
rect 9983 6935 10337 6939
rect 9983 6841 10115 6935
rect 9685 6815 9885 6841
rect 9463 6811 9885 6815
tri 9885 6811 9915 6841 sw
tri 9983 6811 10013 6841 ne
rect 10013 6815 10115 6841
rect 10235 6841 10337 6935
tri 10337 6841 10435 6939 sw
tri 10435 6841 10533 6939 ne
rect 10533 6935 10887 6939
rect 10533 6841 10665 6935
rect 10235 6815 10435 6841
rect 10013 6811 10435 6815
tri 10435 6811 10465 6841 sw
tri 10533 6811 10563 6841 ne
rect 10563 6815 10665 6841
rect 10785 6841 10887 6935
tri 10887 6841 10985 6939 sw
tri 10985 6841 11083 6939 ne
rect 11083 6935 11437 6939
rect 11083 6841 11215 6935
rect 10785 6815 10985 6841
rect 10563 6811 10985 6815
tri 10985 6811 11015 6841 sw
tri 11083 6811 11113 6841 ne
rect 11113 6815 11215 6841
rect 11335 6841 11437 6935
tri 11437 6841 11535 6939 sw
tri 11535 6841 11633 6939 ne
rect 11633 6935 11987 6939
rect 11633 6841 11765 6935
rect 11335 6815 11535 6841
rect 11113 6811 11535 6815
tri 11535 6811 11565 6841 sw
tri 11633 6811 11663 6841 ne
rect 11663 6815 11765 6841
rect 11885 6841 11987 6935
tri 11987 6841 12085 6939 sw
tri 12085 6841 12183 6939 ne
rect 12183 6935 12537 6939
rect 12183 6841 12315 6935
rect 11885 6815 12085 6841
rect 11663 6811 12085 6815
tri 12085 6811 12115 6841 sw
tri 12183 6811 12213 6841 ne
rect 12213 6815 12315 6841
rect 12435 6841 12537 6935
tri 12537 6841 12635 6939 sw
tri 12635 6841 12733 6939 ne
rect 12733 6935 13087 6939
rect 12733 6841 12865 6935
rect 12435 6815 12635 6841
rect 12213 6811 12635 6815
tri 12635 6811 12665 6841 sw
tri 12733 6811 12763 6841 ne
rect 12763 6815 12865 6841
rect 12985 6841 13087 6935
tri 13087 6841 13185 6939 sw
tri 13185 6841 13283 6939 ne
rect 13283 6935 13637 6939
rect 13283 6841 13415 6935
rect 12985 6815 13185 6841
rect 12763 6811 13185 6815
tri 13185 6811 13215 6841 sw
tri 13283 6811 13313 6841 ne
rect 13313 6815 13415 6841
rect 13535 6841 13637 6935
tri 13637 6841 13735 6939 sw
tri 13735 6841 13833 6939 ne
rect 13833 6935 14187 6939
rect 13833 6841 13965 6935
rect 13535 6815 13735 6841
rect 13313 6811 13735 6815
tri 13735 6811 13765 6841 sw
tri 13833 6811 13863 6841 ne
rect 13863 6815 13965 6841
rect 14085 6841 14187 6935
tri 14187 6841 14285 6939 sw
tri 14285 6841 14383 6939 ne
rect 14383 6935 14737 6939
rect 14383 6841 14515 6935
rect 14085 6815 14285 6841
rect 13863 6811 14285 6815
tri 14285 6811 14315 6841 sw
tri 14383 6811 14413 6841 ne
rect 14413 6815 14515 6841
rect 14635 6841 14737 6935
tri 14737 6841 14835 6939 sw
tri 14835 6841 14933 6939 ne
rect 14933 6935 15287 6939
rect 14933 6841 15065 6935
rect 14635 6815 14835 6841
rect 14413 6811 14835 6815
tri 14835 6811 14865 6841 sw
tri 14933 6811 14963 6841 ne
rect 14963 6815 15065 6841
rect 15185 6841 15287 6935
tri 15287 6841 15385 6939 sw
tri 15385 6841 15483 6939 ne
rect 15483 6935 15837 6939
rect 15483 6841 15615 6935
rect 15185 6815 15385 6841
rect 14963 6811 15385 6815
tri 15385 6811 15415 6841 sw
tri 15483 6811 15513 6841 ne
rect 15513 6815 15615 6841
rect 15735 6841 15837 6935
tri 15837 6841 15935 6939 sw
tri 15935 6841 16033 6939 ne
rect 16033 6935 16387 6939
rect 16033 6841 16165 6935
rect 15735 6815 15935 6841
rect 15513 6811 15935 6815
tri 15935 6811 15965 6841 sw
tri 16033 6811 16063 6841 ne
rect 16063 6815 16165 6841
rect 16285 6841 16387 6935
tri 16387 6841 16485 6939 sw
tri 16485 6841 16583 6939 ne
rect 16583 6935 16937 6939
rect 16583 6841 16715 6935
rect 16285 6815 16485 6841
rect 16063 6811 16485 6815
tri 16485 6811 16515 6841 sw
tri 16583 6811 16613 6841 ne
rect 16613 6815 16715 6841
rect 16835 6841 16937 6935
tri 16937 6841 17035 6939 sw
tri 17035 6841 17133 6939 ne
rect 17133 6935 17487 6939
rect 17133 6841 17265 6935
rect 16835 6815 17035 6841
rect 16613 6811 17035 6815
tri 17035 6811 17065 6841 sw
tri 17133 6811 17163 6841 ne
rect 17163 6815 17265 6841
rect 17385 6841 17487 6935
tri 17487 6841 17585 6939 sw
tri 17585 6841 17683 6939 ne
rect 17683 6935 18037 6939
rect 17683 6841 17815 6935
rect 17385 6815 17585 6841
rect 17163 6811 17585 6815
tri 17585 6811 17615 6841 sw
tri 17683 6811 17713 6841 ne
rect 17713 6815 17815 6841
rect 17935 6841 18037 6935
tri 18037 6841 18135 6939 sw
tri 18135 6841 18233 6939 ne
rect 18233 6935 18587 6939
rect 18233 6841 18365 6935
rect 17935 6815 18135 6841
rect 17713 6811 18135 6815
tri 18135 6811 18165 6841 sw
tri 18233 6811 18263 6841 ne
rect 18263 6815 18365 6841
rect 18485 6841 18587 6935
tri 18587 6841 18685 6939 sw
tri 18685 6841 18783 6939 ne
rect 18783 6935 19137 6939
rect 18783 6841 18915 6935
rect 18485 6815 18685 6841
rect 18263 6811 18685 6815
tri 18685 6811 18715 6841 sw
tri 18783 6811 18813 6841 ne
rect 18813 6815 18915 6841
rect 19035 6841 19137 6935
tri 19137 6841 19235 6939 sw
tri 19235 6841 19333 6939 ne
rect 19333 6935 20300 6939
rect 19333 6841 19465 6935
rect 19035 6815 19235 6841
rect 18813 6811 19235 6815
tri 19235 6811 19265 6841 sw
tri 19333 6811 19363 6841 ne
rect 19363 6815 19465 6841
rect 19585 6815 20300 6935
rect 19363 6811 20300 6815
tri 113 6713 211 6811 ne
rect 211 6713 565 6811
tri 565 6713 663 6811 sw
tri 663 6713 761 6811 ne
rect 761 6713 1115 6811
tri 1115 6713 1213 6811 sw
tri 1213 6713 1311 6811 ne
rect 1311 6713 1665 6811
tri 1665 6713 1763 6811 sw
tri 1763 6713 1861 6811 ne
rect 1861 6713 2215 6811
tri 2215 6713 2313 6811 sw
tri 2313 6713 2411 6811 ne
rect 2411 6713 2765 6811
tri 2765 6713 2863 6811 sw
tri 2863 6713 2961 6811 ne
rect 2961 6713 3315 6811
tri 3315 6713 3413 6811 sw
tri 3413 6713 3511 6811 ne
rect 3511 6713 3865 6811
tri 3865 6713 3963 6811 sw
tri 3963 6713 4061 6811 ne
rect 4061 6713 4415 6811
tri 4415 6713 4513 6811 sw
tri 4513 6713 4611 6811 ne
rect 4611 6713 4965 6811
tri 4965 6713 5063 6811 sw
tri 5063 6713 5161 6811 ne
rect 5161 6713 5515 6811
tri 5515 6713 5613 6811 sw
tri 5613 6713 5711 6811 ne
rect 5711 6713 6065 6811
tri 6065 6713 6163 6811 sw
tri 6163 6713 6261 6811 ne
rect 6261 6713 6615 6811
tri 6615 6713 6713 6811 sw
tri 6713 6713 6811 6811 ne
rect 6811 6713 7165 6811
tri 7165 6713 7263 6811 sw
tri 7263 6713 7361 6811 ne
rect 7361 6713 7715 6811
tri 7715 6713 7813 6811 sw
tri 7813 6713 7911 6811 ne
rect 7911 6713 8265 6811
tri 8265 6713 8363 6811 sw
tri 8363 6713 8461 6811 ne
rect 8461 6713 8815 6811
tri 8815 6713 8913 6811 sw
tri 8913 6713 9011 6811 ne
rect 9011 6713 9365 6811
tri 9365 6713 9463 6811 sw
tri 9463 6713 9561 6811 ne
rect 9561 6713 9915 6811
tri 9915 6713 10013 6811 sw
tri 10013 6713 10111 6811 ne
rect 10111 6713 10465 6811
tri 10465 6713 10563 6811 sw
tri 10563 6713 10661 6811 ne
rect 10661 6713 11015 6811
tri 11015 6713 11113 6811 sw
tri 11113 6713 11211 6811 ne
rect 11211 6713 11565 6811
tri 11565 6713 11663 6811 sw
tri 11663 6713 11761 6811 ne
rect 11761 6713 12115 6811
tri 12115 6713 12213 6811 sw
tri 12213 6713 12311 6811 ne
rect 12311 6713 12665 6811
tri 12665 6713 12763 6811 sw
tri 12763 6713 12861 6811 ne
rect 12861 6713 13215 6811
tri 13215 6713 13313 6811 sw
tri 13313 6713 13411 6811 ne
rect 13411 6713 13765 6811
tri 13765 6713 13863 6811 sw
tri 13863 6713 13961 6811 ne
rect 13961 6713 14315 6811
tri 14315 6713 14413 6811 sw
tri 14413 6713 14511 6811 ne
rect 14511 6713 14865 6811
tri 14865 6713 14963 6811 sw
tri 14963 6713 15061 6811 ne
rect 15061 6713 15415 6811
tri 15415 6713 15513 6811 sw
tri 15513 6713 15611 6811 ne
rect 15611 6713 15965 6811
tri 15965 6713 16063 6811 sw
tri 16063 6713 16161 6811 ne
rect 16161 6713 16515 6811
tri 16515 6713 16613 6811 sw
tri 16613 6713 16711 6811 ne
rect 16711 6713 17065 6811
tri 17065 6713 17163 6811 sw
tri 17163 6713 17261 6811 ne
rect 17261 6713 17615 6811
tri 17615 6713 17713 6811 sw
tri 17713 6713 17811 6811 ne
rect 17811 6713 18165 6811
tri 18165 6713 18263 6811 sw
tri 18263 6713 18361 6811 ne
rect 18361 6713 18715 6811
tri 18715 6713 18813 6811 sw
tri 18813 6713 18911 6811 ne
rect 18911 6713 19265 6811
tri 19265 6713 19363 6811 sw
tri 19363 6713 19461 6811 ne
rect 19461 6713 20300 6811
rect -2000 6683 113 6713
tri 113 6683 143 6713 sw
tri 211 6683 241 6713 ne
rect 241 6683 663 6713
tri 663 6683 693 6713 sw
tri 761 6683 791 6713 ne
rect 791 6683 1213 6713
tri 1213 6683 1243 6713 sw
tri 1311 6683 1341 6713 ne
rect 1341 6683 1763 6713
tri 1763 6683 1793 6713 sw
tri 1861 6683 1891 6713 ne
rect 1891 6683 2313 6713
tri 2313 6683 2343 6713 sw
tri 2411 6683 2441 6713 ne
rect 2441 6683 2863 6713
tri 2863 6683 2893 6713 sw
tri 2961 6683 2991 6713 ne
rect 2991 6683 3413 6713
tri 3413 6683 3443 6713 sw
tri 3511 6683 3541 6713 ne
rect 3541 6683 3963 6713
tri 3963 6683 3993 6713 sw
tri 4061 6683 4091 6713 ne
rect 4091 6683 4513 6713
tri 4513 6683 4543 6713 sw
tri 4611 6683 4641 6713 ne
rect 4641 6683 5063 6713
tri 5063 6683 5093 6713 sw
tri 5161 6683 5191 6713 ne
rect 5191 6683 5613 6713
tri 5613 6683 5643 6713 sw
tri 5711 6683 5741 6713 ne
rect 5741 6683 6163 6713
tri 6163 6683 6193 6713 sw
tri 6261 6683 6291 6713 ne
rect 6291 6683 6713 6713
tri 6713 6683 6743 6713 sw
tri 6811 6683 6841 6713 ne
rect 6841 6683 7263 6713
tri 7263 6683 7293 6713 sw
tri 7361 6683 7391 6713 ne
rect 7391 6683 7813 6713
tri 7813 6683 7843 6713 sw
tri 7911 6683 7941 6713 ne
rect 7941 6683 8363 6713
tri 8363 6683 8393 6713 sw
tri 8461 6683 8491 6713 ne
rect 8491 6683 8913 6713
tri 8913 6683 8943 6713 sw
tri 9011 6683 9041 6713 ne
rect 9041 6683 9463 6713
tri 9463 6683 9493 6713 sw
tri 9561 6683 9591 6713 ne
rect 9591 6683 10013 6713
tri 10013 6683 10043 6713 sw
tri 10111 6683 10141 6713 ne
rect 10141 6683 10563 6713
tri 10563 6683 10593 6713 sw
tri 10661 6683 10691 6713 ne
rect 10691 6683 11113 6713
tri 11113 6683 11143 6713 sw
tri 11211 6683 11241 6713 ne
rect 11241 6683 11663 6713
tri 11663 6683 11693 6713 sw
tri 11761 6683 11791 6713 ne
rect 11791 6683 12213 6713
tri 12213 6683 12243 6713 sw
tri 12311 6683 12341 6713 ne
rect 12341 6683 12763 6713
tri 12763 6683 12793 6713 sw
tri 12861 6683 12891 6713 ne
rect 12891 6683 13313 6713
tri 13313 6683 13343 6713 sw
tri 13411 6683 13441 6713 ne
rect 13441 6683 13863 6713
tri 13863 6683 13893 6713 sw
tri 13961 6683 13991 6713 ne
rect 13991 6683 14413 6713
tri 14413 6683 14443 6713 sw
tri 14511 6683 14541 6713 ne
rect 14541 6683 14963 6713
tri 14963 6683 14993 6713 sw
tri 15061 6683 15091 6713 ne
rect 15091 6683 15513 6713
tri 15513 6683 15543 6713 sw
tri 15611 6683 15641 6713 ne
rect 15641 6683 16063 6713
tri 16063 6683 16093 6713 sw
tri 16161 6683 16191 6713 ne
rect 16191 6683 16613 6713
tri 16613 6683 16643 6713 sw
tri 16711 6683 16741 6713 ne
rect 16741 6683 17163 6713
tri 17163 6683 17193 6713 sw
tri 17261 6683 17291 6713 ne
rect 17291 6683 17713 6713
tri 17713 6683 17743 6713 sw
tri 17811 6683 17841 6713 ne
rect 17841 6683 18263 6713
tri 18263 6683 18293 6713 sw
tri 18361 6683 18391 6713 ne
rect 18391 6683 18813 6713
tri 18813 6683 18843 6713 sw
tri 18911 6683 18941 6713 ne
rect 18941 6683 19363 6713
tri 19363 6683 19393 6713 sw
tri 19461 6683 19491 6713 ne
rect 19491 6683 20300 6713
rect -2000 6585 143 6683
tri 143 6585 241 6683 sw
tri 241 6585 339 6683 ne
rect 339 6585 693 6683
tri 693 6585 791 6683 sw
tri 791 6585 889 6683 ne
rect 889 6585 1243 6683
tri 1243 6585 1341 6683 sw
tri 1341 6585 1439 6683 ne
rect 1439 6585 1793 6683
tri 1793 6585 1891 6683 sw
tri 1891 6585 1989 6683 ne
rect 1989 6585 2343 6683
tri 2343 6585 2441 6683 sw
tri 2441 6585 2539 6683 ne
rect 2539 6585 2893 6683
tri 2893 6585 2991 6683 sw
tri 2991 6585 3089 6683 ne
rect 3089 6585 3443 6683
tri 3443 6585 3541 6683 sw
tri 3541 6585 3639 6683 ne
rect 3639 6585 3993 6683
tri 3993 6585 4091 6683 sw
tri 4091 6585 4189 6683 ne
rect 4189 6585 4543 6683
tri 4543 6585 4641 6683 sw
tri 4641 6585 4739 6683 ne
rect 4739 6585 5093 6683
tri 5093 6585 5191 6683 sw
tri 5191 6585 5289 6683 ne
rect 5289 6585 5643 6683
tri 5643 6585 5741 6683 sw
tri 5741 6585 5839 6683 ne
rect 5839 6585 6193 6683
tri 6193 6585 6291 6683 sw
tri 6291 6585 6389 6683 ne
rect 6389 6585 6743 6683
tri 6743 6585 6841 6683 sw
tri 6841 6585 6939 6683 ne
rect 6939 6585 7293 6683
tri 7293 6585 7391 6683 sw
tri 7391 6585 7489 6683 ne
rect 7489 6585 7843 6683
tri 7843 6585 7941 6683 sw
tri 7941 6585 8039 6683 ne
rect 8039 6585 8393 6683
tri 8393 6585 8491 6683 sw
tri 8491 6585 8589 6683 ne
rect 8589 6585 8943 6683
tri 8943 6585 9041 6683 sw
tri 9041 6585 9139 6683 ne
rect 9139 6585 9493 6683
tri 9493 6585 9591 6683 sw
tri 9591 6585 9689 6683 ne
rect 9689 6585 10043 6683
tri 10043 6585 10141 6683 sw
tri 10141 6585 10239 6683 ne
rect 10239 6585 10593 6683
tri 10593 6585 10691 6683 sw
tri 10691 6585 10789 6683 ne
rect 10789 6585 11143 6683
tri 11143 6585 11241 6683 sw
tri 11241 6585 11339 6683 ne
rect 11339 6585 11693 6683
tri 11693 6585 11791 6683 sw
tri 11791 6585 11889 6683 ne
rect 11889 6585 12243 6683
tri 12243 6585 12341 6683 sw
tri 12341 6585 12439 6683 ne
rect 12439 6585 12793 6683
tri 12793 6585 12891 6683 sw
tri 12891 6585 12989 6683 ne
rect 12989 6585 13343 6683
tri 13343 6585 13441 6683 sw
tri 13441 6585 13539 6683 ne
rect 13539 6585 13893 6683
tri 13893 6585 13991 6683 sw
tri 13991 6585 14089 6683 ne
rect 14089 6585 14443 6683
tri 14443 6585 14541 6683 sw
tri 14541 6585 14639 6683 ne
rect 14639 6585 14993 6683
tri 14993 6585 15091 6683 sw
tri 15091 6585 15189 6683 ne
rect 15189 6585 15543 6683
tri 15543 6585 15641 6683 sw
tri 15641 6585 15739 6683 ne
rect 15739 6585 16093 6683
tri 16093 6585 16191 6683 sw
tri 16191 6585 16289 6683 ne
rect 16289 6585 16643 6683
tri 16643 6585 16741 6683 sw
tri 16741 6585 16839 6683 ne
rect 16839 6585 17193 6683
tri 17193 6585 17291 6683 sw
tri 17291 6585 17389 6683 ne
rect 17389 6585 17743 6683
tri 17743 6585 17841 6683 sw
tri 17841 6585 17939 6683 ne
rect 17939 6585 18293 6683
tri 18293 6585 18391 6683 sw
tri 18391 6585 18489 6683 ne
rect 18489 6585 18843 6683
tri 18843 6585 18941 6683 sw
tri 18941 6585 19039 6683 ne
rect 19039 6585 19393 6683
tri 19393 6585 19491 6683 sw
tri 19491 6585 19589 6683 ne
rect 19589 6585 20300 6683
rect -2000 6487 241 6585
tri 241 6487 339 6585 sw
tri 339 6487 437 6585 ne
rect 437 6487 791 6585
tri 791 6487 889 6585 sw
tri 889 6487 987 6585 ne
rect 987 6487 1341 6585
tri 1341 6487 1439 6585 sw
tri 1439 6487 1537 6585 ne
rect 1537 6487 1891 6585
tri 1891 6487 1989 6585 sw
tri 1989 6487 2087 6585 ne
rect 2087 6487 2441 6585
tri 2441 6487 2539 6585 sw
tri 2539 6487 2637 6585 ne
rect 2637 6487 2991 6585
tri 2991 6487 3089 6585 sw
tri 3089 6487 3187 6585 ne
rect 3187 6487 3541 6585
tri 3541 6487 3639 6585 sw
tri 3639 6487 3737 6585 ne
rect 3737 6487 4091 6585
tri 4091 6487 4189 6585 sw
tri 4189 6487 4287 6585 ne
rect 4287 6487 4641 6585
tri 4641 6487 4739 6585 sw
tri 4739 6487 4837 6585 ne
rect 4837 6487 5191 6585
tri 5191 6487 5289 6585 sw
tri 5289 6487 5387 6585 ne
rect 5387 6487 5741 6585
tri 5741 6487 5839 6585 sw
tri 5839 6487 5937 6585 ne
rect 5937 6487 6291 6585
tri 6291 6487 6389 6585 sw
tri 6389 6487 6487 6585 ne
rect 6487 6487 6841 6585
tri 6841 6487 6939 6585 sw
tri 6939 6487 7037 6585 ne
rect 7037 6487 7391 6585
tri 7391 6487 7489 6585 sw
tri 7489 6487 7587 6585 ne
rect 7587 6487 7941 6585
tri 7941 6487 8039 6585 sw
tri 8039 6487 8137 6585 ne
rect 8137 6487 8491 6585
tri 8491 6487 8589 6585 sw
tri 8589 6487 8687 6585 ne
rect 8687 6487 9041 6585
tri 9041 6487 9139 6585 sw
tri 9139 6487 9237 6585 ne
rect 9237 6487 9591 6585
tri 9591 6487 9689 6585 sw
tri 9689 6487 9787 6585 ne
rect 9787 6487 10141 6585
tri 10141 6487 10239 6585 sw
tri 10239 6487 10337 6585 ne
rect 10337 6487 10691 6585
tri 10691 6487 10789 6585 sw
tri 10789 6487 10887 6585 ne
rect 10887 6487 11241 6585
tri 11241 6487 11339 6585 sw
tri 11339 6487 11437 6585 ne
rect 11437 6487 11791 6585
tri 11791 6487 11889 6585 sw
tri 11889 6487 11987 6585 ne
rect 11987 6487 12341 6585
tri 12341 6487 12439 6585 sw
tri 12439 6487 12537 6585 ne
rect 12537 6487 12891 6585
tri 12891 6487 12989 6585 sw
tri 12989 6487 13087 6585 ne
rect 13087 6487 13441 6585
tri 13441 6487 13539 6585 sw
tri 13539 6487 13637 6585 ne
rect 13637 6487 13991 6585
tri 13991 6487 14089 6585 sw
tri 14089 6487 14187 6585 ne
rect 14187 6487 14541 6585
tri 14541 6487 14639 6585 sw
tri 14639 6487 14737 6585 ne
rect 14737 6487 15091 6585
tri 15091 6487 15189 6585 sw
tri 15189 6487 15287 6585 ne
rect 15287 6487 15641 6585
tri 15641 6487 15739 6585 sw
tri 15739 6487 15837 6585 ne
rect 15837 6487 16191 6585
tri 16191 6487 16289 6585 sw
tri 16289 6487 16387 6585 ne
rect 16387 6487 16741 6585
tri 16741 6487 16839 6585 sw
tri 16839 6487 16937 6585 ne
rect 16937 6487 17291 6585
tri 17291 6487 17389 6585 sw
tri 17389 6487 17487 6585 ne
rect 17487 6487 17841 6585
tri 17841 6487 17939 6585 sw
tri 17939 6487 18037 6585 ne
rect 18037 6487 18391 6585
tri 18391 6487 18489 6585 sw
tri 18489 6487 18587 6585 ne
rect 18587 6487 18941 6585
tri 18941 6487 19039 6585 sw
tri 19039 6487 19137 6585 ne
rect 19137 6487 19491 6585
tri 19491 6487 19589 6585 sw
tri 19589 6487 19687 6585 ne
rect 19687 6487 20300 6585
rect -2000 6389 339 6487
tri 339 6389 437 6487 sw
tri 437 6389 535 6487 ne
rect 535 6389 889 6487
tri 889 6389 987 6487 sw
tri 987 6389 1085 6487 ne
rect 1085 6389 1439 6487
tri 1439 6389 1537 6487 sw
tri 1537 6389 1635 6487 ne
rect 1635 6389 1989 6487
tri 1989 6389 2087 6487 sw
tri 2087 6389 2185 6487 ne
rect 2185 6389 2539 6487
tri 2539 6389 2637 6487 sw
tri 2637 6389 2735 6487 ne
rect 2735 6389 3089 6487
tri 3089 6389 3187 6487 sw
tri 3187 6389 3285 6487 ne
rect 3285 6389 3639 6487
tri 3639 6389 3737 6487 sw
tri 3737 6389 3835 6487 ne
rect 3835 6389 4189 6487
tri 4189 6389 4287 6487 sw
tri 4287 6389 4385 6487 ne
rect 4385 6389 4739 6487
tri 4739 6389 4837 6487 sw
tri 4837 6389 4935 6487 ne
rect 4935 6389 5289 6487
tri 5289 6389 5387 6487 sw
tri 5387 6389 5485 6487 ne
rect 5485 6389 5839 6487
tri 5839 6389 5937 6487 sw
tri 5937 6389 6035 6487 ne
rect 6035 6389 6389 6487
tri 6389 6389 6487 6487 sw
tri 6487 6389 6585 6487 ne
rect 6585 6389 6939 6487
tri 6939 6389 7037 6487 sw
tri 7037 6389 7135 6487 ne
rect 7135 6389 7489 6487
tri 7489 6389 7587 6487 sw
tri 7587 6389 7685 6487 ne
rect 7685 6389 8039 6487
tri 8039 6389 8137 6487 sw
tri 8137 6389 8235 6487 ne
rect 8235 6389 8589 6487
tri 8589 6389 8687 6487 sw
tri 8687 6389 8785 6487 ne
rect 8785 6389 9139 6487
tri 9139 6389 9237 6487 sw
tri 9237 6389 9335 6487 ne
rect 9335 6389 9689 6487
tri 9689 6389 9787 6487 sw
tri 9787 6389 9885 6487 ne
rect 9885 6389 10239 6487
tri 10239 6389 10337 6487 sw
tri 10337 6389 10435 6487 ne
rect 10435 6389 10789 6487
tri 10789 6389 10887 6487 sw
tri 10887 6389 10985 6487 ne
rect 10985 6389 11339 6487
tri 11339 6389 11437 6487 sw
tri 11437 6389 11535 6487 ne
rect 11535 6389 11889 6487
tri 11889 6389 11987 6487 sw
tri 11987 6389 12085 6487 ne
rect 12085 6389 12439 6487
tri 12439 6389 12537 6487 sw
tri 12537 6389 12635 6487 ne
rect 12635 6389 12989 6487
tri 12989 6389 13087 6487 sw
tri 13087 6389 13185 6487 ne
rect 13185 6389 13539 6487
tri 13539 6389 13637 6487 sw
tri 13637 6389 13735 6487 ne
rect 13735 6389 14089 6487
tri 14089 6389 14187 6487 sw
tri 14187 6389 14285 6487 ne
rect 14285 6389 14639 6487
tri 14639 6389 14737 6487 sw
tri 14737 6389 14835 6487 ne
rect 14835 6389 15189 6487
tri 15189 6389 15287 6487 sw
tri 15287 6389 15385 6487 ne
rect 15385 6389 15739 6487
tri 15739 6389 15837 6487 sw
tri 15837 6389 15935 6487 ne
rect 15935 6389 16289 6487
tri 16289 6389 16387 6487 sw
tri 16387 6389 16485 6487 ne
rect 16485 6389 16839 6487
tri 16839 6389 16937 6487 sw
tri 16937 6389 17035 6487 ne
rect 17035 6389 17389 6487
tri 17389 6389 17487 6487 sw
tri 17487 6389 17585 6487 ne
rect 17585 6389 17939 6487
tri 17939 6389 18037 6487 sw
tri 18037 6389 18135 6487 ne
rect 18135 6389 18489 6487
tri 18489 6389 18587 6487 sw
tri 18587 6389 18685 6487 ne
rect 18685 6389 19039 6487
tri 19039 6389 19137 6487 sw
tri 19137 6389 19235 6487 ne
rect 19235 6389 19589 6487
tri 19589 6389 19687 6487 sw
rect 20800 6389 21800 7037
rect -2000 6385 437 6389
rect -2000 6265 215 6385
rect 335 6291 437 6385
tri 437 6291 535 6389 sw
tri 535 6291 633 6389 ne
rect 633 6385 987 6389
rect 633 6291 765 6385
rect 335 6265 535 6291
rect -2000 6261 535 6265
rect -2000 5613 -1000 6261
tri 113 6163 211 6261 ne
rect 211 6213 535 6261
tri 535 6213 613 6291 sw
tri 633 6213 711 6291 ne
rect 711 6265 765 6291
rect 885 6291 987 6385
tri 987 6291 1085 6389 sw
tri 1085 6291 1183 6389 ne
rect 1183 6385 1537 6389
rect 1183 6291 1315 6385
rect 885 6265 1085 6291
rect 711 6213 1085 6265
tri 1085 6213 1163 6291 sw
tri 1183 6213 1261 6291 ne
rect 1261 6265 1315 6291
rect 1435 6291 1537 6385
tri 1537 6291 1635 6389 sw
tri 1635 6291 1733 6389 ne
rect 1733 6385 2087 6389
rect 1733 6291 1865 6385
rect 1435 6265 1635 6291
rect 1261 6213 1635 6265
tri 1635 6213 1713 6291 sw
tri 1733 6213 1811 6291 ne
rect 1811 6265 1865 6291
rect 1985 6291 2087 6385
tri 2087 6291 2185 6389 sw
tri 2185 6291 2283 6389 ne
rect 2283 6385 2637 6389
rect 2283 6291 2415 6385
rect 1985 6265 2185 6291
rect 1811 6213 2185 6265
tri 2185 6213 2263 6291 sw
tri 2283 6213 2361 6291 ne
rect 2361 6265 2415 6291
rect 2535 6291 2637 6385
tri 2637 6291 2735 6389 sw
tri 2735 6291 2833 6389 ne
rect 2833 6385 3187 6389
rect 2833 6291 2965 6385
rect 2535 6265 2735 6291
rect 2361 6213 2735 6265
tri 2735 6213 2813 6291 sw
tri 2833 6213 2911 6291 ne
rect 2911 6265 2965 6291
rect 3085 6291 3187 6385
tri 3187 6291 3285 6389 sw
tri 3285 6291 3383 6389 ne
rect 3383 6385 3737 6389
rect 3383 6291 3515 6385
rect 3085 6265 3285 6291
rect 2911 6213 3285 6265
tri 3285 6213 3363 6291 sw
tri 3383 6213 3461 6291 ne
rect 3461 6265 3515 6291
rect 3635 6291 3737 6385
tri 3737 6291 3835 6389 sw
tri 3835 6291 3933 6389 ne
rect 3933 6385 4287 6389
rect 3933 6291 4065 6385
rect 3635 6265 3835 6291
rect 3461 6213 3835 6265
tri 3835 6213 3913 6291 sw
tri 3933 6213 4011 6291 ne
rect 4011 6265 4065 6291
rect 4185 6291 4287 6385
tri 4287 6291 4385 6389 sw
tri 4385 6291 4483 6389 ne
rect 4483 6385 4837 6389
rect 4483 6291 4615 6385
rect 4185 6265 4385 6291
rect 4011 6213 4385 6265
tri 4385 6213 4463 6291 sw
tri 4483 6213 4561 6291 ne
rect 4561 6265 4615 6291
rect 4735 6291 4837 6385
tri 4837 6291 4935 6389 sw
tri 4935 6291 5033 6389 ne
rect 5033 6385 5387 6389
rect 5033 6291 5165 6385
rect 4735 6265 4935 6291
rect 4561 6213 4935 6265
tri 4935 6213 5013 6291 sw
tri 5033 6213 5111 6291 ne
rect 5111 6265 5165 6291
rect 5285 6291 5387 6385
tri 5387 6291 5485 6389 sw
tri 5485 6291 5583 6389 ne
rect 5583 6385 5937 6389
rect 5583 6291 5715 6385
rect 5285 6265 5485 6291
rect 5111 6213 5485 6265
tri 5485 6213 5563 6291 sw
tri 5583 6213 5661 6291 ne
rect 5661 6265 5715 6291
rect 5835 6291 5937 6385
tri 5937 6291 6035 6389 sw
tri 6035 6291 6133 6389 ne
rect 6133 6385 6487 6389
rect 6133 6291 6265 6385
rect 5835 6265 6035 6291
rect 5661 6213 6035 6265
tri 6035 6213 6113 6291 sw
tri 6133 6213 6211 6291 ne
rect 6211 6265 6265 6291
rect 6385 6291 6487 6385
tri 6487 6291 6585 6389 sw
tri 6585 6291 6683 6389 ne
rect 6683 6385 7037 6389
rect 6683 6291 6815 6385
rect 6385 6265 6585 6291
rect 6211 6213 6585 6265
tri 6585 6213 6663 6291 sw
tri 6683 6213 6761 6291 ne
rect 6761 6265 6815 6291
rect 6935 6291 7037 6385
tri 7037 6291 7135 6389 sw
tri 7135 6291 7233 6389 ne
rect 7233 6385 7587 6389
rect 7233 6291 7365 6385
rect 6935 6265 7135 6291
rect 6761 6213 7135 6265
tri 7135 6213 7213 6291 sw
tri 7233 6213 7311 6291 ne
rect 7311 6265 7365 6291
rect 7485 6291 7587 6385
tri 7587 6291 7685 6389 sw
tri 7685 6291 7783 6389 ne
rect 7783 6385 8137 6389
rect 7783 6291 7915 6385
rect 7485 6265 7685 6291
rect 7311 6213 7685 6265
tri 7685 6213 7763 6291 sw
tri 7783 6213 7861 6291 ne
rect 7861 6265 7915 6291
rect 8035 6291 8137 6385
tri 8137 6291 8235 6389 sw
tri 8235 6291 8333 6389 ne
rect 8333 6385 8687 6389
rect 8333 6291 8465 6385
rect 8035 6265 8235 6291
rect 7861 6213 8235 6265
tri 8235 6213 8313 6291 sw
tri 8333 6213 8411 6291 ne
rect 8411 6265 8465 6291
rect 8585 6291 8687 6385
tri 8687 6291 8785 6389 sw
tri 8785 6291 8883 6389 ne
rect 8883 6385 9237 6389
rect 8883 6291 9015 6385
rect 8585 6265 8785 6291
rect 8411 6213 8785 6265
tri 8785 6213 8863 6291 sw
tri 8883 6213 8961 6291 ne
rect 8961 6265 9015 6291
rect 9135 6291 9237 6385
tri 9237 6291 9335 6389 sw
tri 9335 6291 9433 6389 ne
rect 9433 6385 9787 6389
rect 9433 6291 9565 6385
rect 9135 6265 9335 6291
rect 8961 6213 9335 6265
tri 9335 6213 9413 6291 sw
tri 9433 6213 9511 6291 ne
rect 9511 6265 9565 6291
rect 9685 6291 9787 6385
tri 9787 6291 9885 6389 sw
tri 9885 6291 9983 6389 ne
rect 9983 6385 10337 6389
rect 9983 6291 10115 6385
rect 9685 6265 9885 6291
rect 9511 6213 9885 6265
tri 9885 6213 9963 6291 sw
tri 9983 6213 10061 6291 ne
rect 10061 6265 10115 6291
rect 10235 6291 10337 6385
tri 10337 6291 10435 6389 sw
tri 10435 6291 10533 6389 ne
rect 10533 6385 10887 6389
rect 10533 6291 10665 6385
rect 10235 6265 10435 6291
rect 10061 6213 10435 6265
tri 10435 6213 10513 6291 sw
tri 10533 6213 10611 6291 ne
rect 10611 6265 10665 6291
rect 10785 6291 10887 6385
tri 10887 6291 10985 6389 sw
tri 10985 6291 11083 6389 ne
rect 11083 6385 11437 6389
rect 11083 6291 11215 6385
rect 10785 6265 10985 6291
rect 10611 6213 10985 6265
tri 10985 6213 11063 6291 sw
tri 11083 6213 11161 6291 ne
rect 11161 6265 11215 6291
rect 11335 6291 11437 6385
tri 11437 6291 11535 6389 sw
tri 11535 6291 11633 6389 ne
rect 11633 6385 11987 6389
rect 11633 6291 11765 6385
rect 11335 6265 11535 6291
rect 11161 6213 11535 6265
tri 11535 6213 11613 6291 sw
tri 11633 6213 11711 6291 ne
rect 11711 6265 11765 6291
rect 11885 6291 11987 6385
tri 11987 6291 12085 6389 sw
tri 12085 6291 12183 6389 ne
rect 12183 6385 12537 6389
rect 12183 6291 12315 6385
rect 11885 6265 12085 6291
rect 11711 6213 12085 6265
tri 12085 6213 12163 6291 sw
tri 12183 6213 12261 6291 ne
rect 12261 6265 12315 6291
rect 12435 6291 12537 6385
tri 12537 6291 12635 6389 sw
tri 12635 6291 12733 6389 ne
rect 12733 6385 13087 6389
rect 12733 6291 12865 6385
rect 12435 6265 12635 6291
rect 12261 6213 12635 6265
tri 12635 6213 12713 6291 sw
tri 12733 6213 12811 6291 ne
rect 12811 6265 12865 6291
rect 12985 6291 13087 6385
tri 13087 6291 13185 6389 sw
tri 13185 6291 13283 6389 ne
rect 13283 6385 13637 6389
rect 13283 6291 13415 6385
rect 12985 6265 13185 6291
rect 12811 6213 13185 6265
tri 13185 6213 13263 6291 sw
tri 13283 6213 13361 6291 ne
rect 13361 6265 13415 6291
rect 13535 6291 13637 6385
tri 13637 6291 13735 6389 sw
tri 13735 6291 13833 6389 ne
rect 13833 6385 14187 6389
rect 13833 6291 13965 6385
rect 13535 6265 13735 6291
rect 13361 6213 13735 6265
tri 13735 6213 13813 6291 sw
tri 13833 6213 13911 6291 ne
rect 13911 6265 13965 6291
rect 14085 6291 14187 6385
tri 14187 6291 14285 6389 sw
tri 14285 6291 14383 6389 ne
rect 14383 6385 14737 6389
rect 14383 6291 14515 6385
rect 14085 6265 14285 6291
rect 13911 6213 14285 6265
tri 14285 6213 14363 6291 sw
tri 14383 6213 14461 6291 ne
rect 14461 6265 14515 6291
rect 14635 6291 14737 6385
tri 14737 6291 14835 6389 sw
tri 14835 6291 14933 6389 ne
rect 14933 6385 15287 6389
rect 14933 6291 15065 6385
rect 14635 6265 14835 6291
rect 14461 6213 14835 6265
tri 14835 6213 14913 6291 sw
tri 14933 6213 15011 6291 ne
rect 15011 6265 15065 6291
rect 15185 6291 15287 6385
tri 15287 6291 15385 6389 sw
tri 15385 6291 15483 6389 ne
rect 15483 6385 15837 6389
rect 15483 6291 15615 6385
rect 15185 6265 15385 6291
rect 15011 6213 15385 6265
tri 15385 6213 15463 6291 sw
tri 15483 6213 15561 6291 ne
rect 15561 6265 15615 6291
rect 15735 6291 15837 6385
tri 15837 6291 15935 6389 sw
tri 15935 6291 16033 6389 ne
rect 16033 6385 16387 6389
rect 16033 6291 16165 6385
rect 15735 6265 15935 6291
rect 15561 6213 15935 6265
tri 15935 6213 16013 6291 sw
tri 16033 6213 16111 6291 ne
rect 16111 6265 16165 6291
rect 16285 6291 16387 6385
tri 16387 6291 16485 6389 sw
tri 16485 6291 16583 6389 ne
rect 16583 6385 16937 6389
rect 16583 6291 16715 6385
rect 16285 6265 16485 6291
rect 16111 6213 16485 6265
tri 16485 6213 16563 6291 sw
tri 16583 6213 16661 6291 ne
rect 16661 6265 16715 6291
rect 16835 6291 16937 6385
tri 16937 6291 17035 6389 sw
tri 17035 6291 17133 6389 ne
rect 17133 6385 17487 6389
rect 17133 6291 17265 6385
rect 16835 6265 17035 6291
rect 16661 6213 17035 6265
tri 17035 6213 17113 6291 sw
tri 17133 6213 17211 6291 ne
rect 17211 6265 17265 6291
rect 17385 6291 17487 6385
tri 17487 6291 17585 6389 sw
tri 17585 6291 17683 6389 ne
rect 17683 6385 18037 6389
rect 17683 6291 17815 6385
rect 17385 6265 17585 6291
rect 17211 6213 17585 6265
tri 17585 6213 17663 6291 sw
tri 17683 6213 17761 6291 ne
rect 17761 6265 17815 6291
rect 17935 6291 18037 6385
tri 18037 6291 18135 6389 sw
tri 18135 6291 18233 6389 ne
rect 18233 6385 18587 6389
rect 18233 6291 18365 6385
rect 17935 6265 18135 6291
rect 17761 6213 18135 6265
tri 18135 6213 18213 6291 sw
tri 18233 6213 18311 6291 ne
rect 18311 6265 18365 6291
rect 18485 6291 18587 6385
tri 18587 6291 18685 6389 sw
tri 18685 6291 18783 6389 ne
rect 18783 6385 19137 6389
rect 18783 6291 18915 6385
rect 18485 6265 18685 6291
rect 18311 6213 18685 6265
tri 18685 6213 18763 6291 sw
tri 18783 6213 18861 6291 ne
rect 18861 6265 18915 6291
rect 19035 6291 19137 6385
tri 19137 6291 19235 6389 sw
tri 19235 6291 19333 6389 ne
rect 19333 6385 21800 6389
rect 19333 6291 19465 6385
rect 19035 6265 19235 6291
rect 18861 6213 19235 6265
tri 19235 6213 19313 6291 sw
tri 19333 6213 19411 6291 ne
rect 19411 6265 19465 6291
rect 19585 6265 21800 6385
rect 19411 6213 21800 6265
rect 211 6163 613 6213
rect -500 6113 113 6163
tri 113 6113 163 6163 sw
tri 211 6113 261 6163 ne
rect 261 6133 613 6163
tri 613 6133 693 6213 sw
tri 711 6133 791 6213 ne
rect 791 6133 1163 6213
tri 1163 6133 1243 6213 sw
tri 1261 6133 1341 6213 ne
rect 1341 6133 1713 6213
tri 1713 6133 1793 6213 sw
tri 1811 6133 1891 6213 ne
rect 1891 6133 2263 6213
tri 2263 6133 2343 6213 sw
tri 2361 6133 2441 6213 ne
rect 2441 6133 2813 6213
tri 2813 6133 2893 6213 sw
tri 2911 6133 2991 6213 ne
rect 2991 6133 3363 6213
tri 3363 6133 3443 6213 sw
tri 3461 6133 3541 6213 ne
rect 3541 6133 3913 6213
tri 3913 6133 3993 6213 sw
tri 4011 6133 4091 6213 ne
rect 4091 6133 4463 6213
tri 4463 6133 4543 6213 sw
tri 4561 6133 4641 6213 ne
rect 4641 6133 5013 6213
tri 5013 6133 5093 6213 sw
tri 5111 6133 5191 6213 ne
rect 5191 6133 5563 6213
tri 5563 6133 5643 6213 sw
tri 5661 6133 5741 6213 ne
rect 5741 6133 6113 6213
tri 6113 6133 6193 6213 sw
tri 6211 6133 6291 6213 ne
rect 6291 6133 6663 6213
tri 6663 6133 6743 6213 sw
tri 6761 6133 6841 6213 ne
rect 6841 6133 7213 6213
tri 7213 6133 7293 6213 sw
tri 7311 6133 7391 6213 ne
rect 7391 6133 7763 6213
tri 7763 6133 7843 6213 sw
tri 7861 6133 7941 6213 ne
rect 7941 6133 8313 6213
tri 8313 6133 8393 6213 sw
tri 8411 6133 8491 6213 ne
rect 8491 6133 8863 6213
tri 8863 6133 8943 6213 sw
tri 8961 6133 9041 6213 ne
rect 9041 6133 9413 6213
tri 9413 6133 9493 6213 sw
tri 9511 6133 9591 6213 ne
rect 9591 6133 9963 6213
tri 9963 6133 10043 6213 sw
tri 10061 6133 10141 6213 ne
rect 10141 6133 10513 6213
tri 10513 6133 10593 6213 sw
tri 10611 6133 10691 6213 ne
rect 10691 6133 11063 6213
tri 11063 6133 11143 6213 sw
tri 11161 6133 11241 6213 ne
rect 11241 6133 11613 6213
tri 11613 6133 11693 6213 sw
tri 11711 6133 11791 6213 ne
rect 11791 6133 12163 6213
tri 12163 6133 12243 6213 sw
tri 12261 6133 12341 6213 ne
rect 12341 6133 12713 6213
tri 12713 6133 12793 6213 sw
tri 12811 6133 12891 6213 ne
rect 12891 6133 13263 6213
tri 13263 6133 13343 6213 sw
tri 13361 6133 13441 6213 ne
rect 13441 6133 13813 6213
tri 13813 6133 13893 6213 sw
tri 13911 6133 13991 6213 ne
rect 13991 6133 14363 6213
tri 14363 6133 14443 6213 sw
tri 14461 6133 14541 6213 ne
rect 14541 6133 14913 6213
tri 14913 6133 14993 6213 sw
tri 15011 6133 15091 6213 ne
rect 15091 6133 15463 6213
tri 15463 6133 15543 6213 sw
tri 15561 6133 15641 6213 ne
rect 15641 6133 16013 6213
tri 16013 6133 16093 6213 sw
tri 16111 6133 16191 6213 ne
rect 16191 6133 16563 6213
tri 16563 6133 16643 6213 sw
tri 16661 6133 16741 6213 ne
rect 16741 6133 17113 6213
tri 17113 6133 17193 6213 sw
tri 17211 6133 17291 6213 ne
rect 17291 6133 17663 6213
tri 17663 6133 17743 6213 sw
tri 17761 6133 17841 6213 ne
rect 17841 6133 18213 6213
tri 18213 6133 18293 6213 sw
tri 18311 6133 18391 6213 ne
rect 18391 6133 18763 6213
tri 18763 6133 18843 6213 sw
tri 18861 6133 18941 6213 ne
rect 18941 6133 19313 6213
tri 19313 6133 19393 6213 sw
tri 19411 6133 19491 6213 ne
rect 19491 6133 20100 6213
rect 261 6113 693 6133
rect -500 6035 163 6113
tri 163 6035 241 6113 sw
tri 261 6035 339 6113 ne
rect 339 6035 693 6113
tri 693 6035 791 6133 sw
tri 791 6035 889 6133 ne
rect 889 6035 1243 6133
tri 1243 6035 1341 6133 sw
tri 1341 6035 1439 6133 ne
rect 1439 6035 1793 6133
tri 1793 6035 1891 6133 sw
tri 1891 6035 1989 6133 ne
rect 1989 6035 2343 6133
tri 2343 6035 2441 6133 sw
tri 2441 6035 2539 6133 ne
rect 2539 6035 2893 6133
tri 2893 6035 2991 6133 sw
tri 2991 6035 3089 6133 ne
rect 3089 6035 3443 6133
tri 3443 6035 3541 6133 sw
tri 3541 6035 3639 6133 ne
rect 3639 6035 3993 6133
tri 3993 6035 4091 6133 sw
tri 4091 6035 4189 6133 ne
rect 4189 6035 4543 6133
tri 4543 6035 4641 6133 sw
tri 4641 6035 4739 6133 ne
rect 4739 6035 5093 6133
tri 5093 6035 5191 6133 sw
tri 5191 6035 5289 6133 ne
rect 5289 6035 5643 6133
tri 5643 6035 5741 6133 sw
tri 5741 6035 5839 6133 ne
rect 5839 6035 6193 6133
tri 6193 6035 6291 6133 sw
tri 6291 6035 6389 6133 ne
rect 6389 6035 6743 6133
tri 6743 6035 6841 6133 sw
tri 6841 6035 6939 6133 ne
rect 6939 6035 7293 6133
tri 7293 6035 7391 6133 sw
tri 7391 6035 7489 6133 ne
rect 7489 6035 7843 6133
tri 7843 6035 7941 6133 sw
tri 7941 6035 8039 6133 ne
rect 8039 6035 8393 6133
tri 8393 6035 8491 6133 sw
tri 8491 6035 8589 6133 ne
rect 8589 6035 8943 6133
tri 8943 6035 9041 6133 sw
tri 9041 6035 9139 6133 ne
rect 9139 6035 9493 6133
tri 9493 6035 9591 6133 sw
tri 9591 6035 9689 6133 ne
rect 9689 6035 10043 6133
tri 10043 6035 10141 6133 sw
tri 10141 6035 10239 6133 ne
rect 10239 6035 10593 6133
tri 10593 6035 10691 6133 sw
tri 10691 6035 10789 6133 ne
rect 10789 6035 11143 6133
tri 11143 6035 11241 6133 sw
tri 11241 6035 11339 6133 ne
rect 11339 6035 11693 6133
tri 11693 6035 11791 6133 sw
tri 11791 6035 11889 6133 ne
rect 11889 6035 12243 6133
tri 12243 6035 12341 6133 sw
tri 12341 6035 12439 6133 ne
rect 12439 6035 12793 6133
tri 12793 6035 12891 6133 sw
tri 12891 6035 12989 6133 ne
rect 12989 6035 13343 6133
tri 13343 6035 13441 6133 sw
tri 13441 6035 13539 6133 ne
rect 13539 6035 13893 6133
tri 13893 6035 13991 6133 sw
tri 13991 6035 14089 6133 ne
rect 14089 6035 14443 6133
tri 14443 6035 14541 6133 sw
tri 14541 6035 14639 6133 ne
rect 14639 6035 14993 6133
tri 14993 6035 15091 6133 sw
tri 15091 6035 15189 6133 ne
rect 15189 6035 15543 6133
tri 15543 6035 15641 6133 sw
tri 15641 6035 15739 6133 ne
rect 15739 6035 16093 6133
tri 16093 6035 16191 6133 sw
tri 16191 6035 16289 6133 ne
rect 16289 6035 16643 6133
tri 16643 6035 16741 6133 sw
tri 16741 6035 16839 6133 ne
rect 16839 6035 17193 6133
tri 17193 6035 17291 6133 sw
tri 17291 6035 17389 6133 ne
rect 17389 6035 17743 6133
tri 17743 6035 17841 6133 sw
tri 17841 6035 17939 6133 ne
rect 17939 6035 18293 6133
tri 18293 6035 18391 6133 sw
tri 18391 6035 18489 6133 ne
rect 18489 6035 18843 6133
tri 18843 6035 18941 6133 sw
tri 18941 6035 19039 6133 ne
rect 19039 6035 19393 6133
tri 19393 6035 19491 6133 sw
tri 19491 6035 19589 6133 ne
rect 19589 6113 20100 6133
rect 20200 6113 21800 6213
rect 19589 6035 21800 6113
rect -500 5987 241 6035
rect -500 5887 -400 5987
rect -300 5937 241 5987
tri 241 5937 339 6035 sw
tri 339 5937 437 6035 ne
rect 437 5937 791 6035
tri 791 5937 889 6035 sw
tri 889 5937 987 6035 ne
rect 987 5937 1341 6035
tri 1341 5937 1439 6035 sw
tri 1439 5937 1537 6035 ne
rect 1537 5937 1891 6035
tri 1891 5937 1989 6035 sw
tri 1989 5937 2087 6035 ne
rect 2087 5937 2441 6035
tri 2441 5937 2539 6035 sw
tri 2539 5937 2637 6035 ne
rect 2637 5937 2991 6035
tri 2991 5937 3089 6035 sw
tri 3089 5937 3187 6035 ne
rect 3187 5937 3541 6035
tri 3541 5937 3639 6035 sw
tri 3639 5937 3737 6035 ne
rect 3737 5937 4091 6035
tri 4091 5937 4189 6035 sw
tri 4189 5937 4287 6035 ne
rect 4287 5937 4641 6035
tri 4641 5937 4739 6035 sw
tri 4739 5937 4837 6035 ne
rect 4837 5937 5191 6035
tri 5191 5937 5289 6035 sw
tri 5289 5937 5387 6035 ne
rect 5387 5937 5741 6035
tri 5741 5937 5839 6035 sw
tri 5839 5937 5937 6035 ne
rect 5937 5937 6291 6035
tri 6291 5937 6389 6035 sw
tri 6389 5937 6487 6035 ne
rect 6487 5937 6841 6035
tri 6841 5937 6939 6035 sw
tri 6939 5937 7037 6035 ne
rect 7037 5937 7391 6035
tri 7391 5937 7489 6035 sw
tri 7489 5937 7587 6035 ne
rect 7587 5937 7941 6035
tri 7941 5937 8039 6035 sw
tri 8039 5937 8137 6035 ne
rect 8137 5937 8491 6035
tri 8491 5937 8589 6035 sw
tri 8589 5937 8687 6035 ne
rect 8687 5937 9041 6035
tri 9041 5937 9139 6035 sw
tri 9139 5937 9237 6035 ne
rect 9237 5937 9591 6035
tri 9591 5937 9689 6035 sw
tri 9689 5937 9787 6035 ne
rect 9787 5937 10141 6035
tri 10141 5937 10239 6035 sw
tri 10239 5937 10337 6035 ne
rect 10337 5937 10691 6035
tri 10691 5937 10789 6035 sw
tri 10789 5937 10887 6035 ne
rect 10887 5937 11241 6035
tri 11241 5937 11339 6035 sw
tri 11339 5937 11437 6035 ne
rect 11437 5937 11791 6035
tri 11791 5937 11889 6035 sw
tri 11889 5937 11987 6035 ne
rect 11987 5937 12341 6035
tri 12341 5937 12439 6035 sw
tri 12439 5937 12537 6035 ne
rect 12537 5937 12891 6035
tri 12891 5937 12989 6035 sw
tri 12989 5937 13087 6035 ne
rect 13087 5937 13441 6035
tri 13441 5937 13539 6035 sw
tri 13539 5937 13637 6035 ne
rect 13637 5937 13991 6035
tri 13991 5937 14089 6035 sw
tri 14089 5937 14187 6035 ne
rect 14187 5937 14541 6035
tri 14541 5937 14639 6035 sw
tri 14639 5937 14737 6035 ne
rect 14737 5937 15091 6035
tri 15091 5937 15189 6035 sw
tri 15189 5937 15287 6035 ne
rect 15287 5937 15641 6035
tri 15641 5937 15739 6035 sw
tri 15739 5937 15837 6035 ne
rect 15837 5937 16191 6035
tri 16191 5937 16289 6035 sw
tri 16289 5937 16387 6035 ne
rect 16387 5937 16741 6035
tri 16741 5937 16839 6035 sw
tri 16839 5937 16937 6035 ne
rect 16937 5937 17291 6035
tri 17291 5937 17389 6035 sw
tri 17389 5937 17487 6035 ne
rect 17487 5937 17841 6035
tri 17841 5937 17939 6035 sw
tri 17939 5937 18037 6035 ne
rect 18037 5937 18391 6035
tri 18391 5937 18489 6035 sw
tri 18489 5937 18587 6035 ne
rect 18587 5937 18941 6035
tri 18941 5937 19039 6035 sw
tri 19039 5937 19137 6035 ne
rect 19137 5937 19491 6035
tri 19491 5937 19589 6035 sw
tri 19589 5937 19687 6035 ne
rect 19687 5937 21800 6035
rect -300 5887 339 5937
rect -500 5839 339 5887
tri 339 5839 437 5937 sw
tri 437 5839 535 5937 ne
rect 535 5839 889 5937
tri 889 5839 987 5937 sw
tri 987 5839 1085 5937 ne
rect 1085 5839 1439 5937
tri 1439 5839 1537 5937 sw
tri 1537 5839 1635 5937 ne
rect 1635 5839 1989 5937
tri 1989 5839 2087 5937 sw
tri 2087 5839 2185 5937 ne
rect 2185 5839 2539 5937
tri 2539 5839 2637 5937 sw
tri 2637 5839 2735 5937 ne
rect 2735 5839 3089 5937
tri 3089 5839 3187 5937 sw
tri 3187 5839 3285 5937 ne
rect 3285 5839 3639 5937
tri 3639 5839 3737 5937 sw
tri 3737 5839 3835 5937 ne
rect 3835 5839 4189 5937
tri 4189 5839 4287 5937 sw
tri 4287 5839 4385 5937 ne
rect 4385 5839 4739 5937
tri 4739 5839 4837 5937 sw
tri 4837 5839 4935 5937 ne
rect 4935 5839 5289 5937
tri 5289 5839 5387 5937 sw
tri 5387 5839 5485 5937 ne
rect 5485 5839 5839 5937
tri 5839 5839 5937 5937 sw
tri 5937 5839 6035 5937 ne
rect 6035 5839 6389 5937
tri 6389 5839 6487 5937 sw
tri 6487 5839 6585 5937 ne
rect 6585 5839 6939 5937
tri 6939 5839 7037 5937 sw
tri 7037 5839 7135 5937 ne
rect 7135 5839 7489 5937
tri 7489 5839 7587 5937 sw
tri 7587 5839 7685 5937 ne
rect 7685 5839 8039 5937
tri 8039 5839 8137 5937 sw
tri 8137 5839 8235 5937 ne
rect 8235 5839 8589 5937
tri 8589 5839 8687 5937 sw
tri 8687 5839 8785 5937 ne
rect 8785 5839 9139 5937
tri 9139 5839 9237 5937 sw
tri 9237 5839 9335 5937 ne
rect 9335 5839 9689 5937
tri 9689 5839 9787 5937 sw
tri 9787 5839 9885 5937 ne
rect 9885 5839 10239 5937
tri 10239 5839 10337 5937 sw
tri 10337 5839 10435 5937 ne
rect 10435 5839 10789 5937
tri 10789 5839 10887 5937 sw
tri 10887 5839 10985 5937 ne
rect 10985 5839 11339 5937
tri 11339 5839 11437 5937 sw
tri 11437 5839 11535 5937 ne
rect 11535 5839 11889 5937
tri 11889 5839 11987 5937 sw
tri 11987 5839 12085 5937 ne
rect 12085 5839 12439 5937
tri 12439 5839 12537 5937 sw
tri 12537 5839 12635 5937 ne
rect 12635 5839 12989 5937
tri 12989 5839 13087 5937 sw
tri 13087 5839 13185 5937 ne
rect 13185 5839 13539 5937
tri 13539 5839 13637 5937 sw
tri 13637 5839 13735 5937 ne
rect 13735 5839 14089 5937
tri 14089 5839 14187 5937 sw
tri 14187 5839 14285 5937 ne
rect 14285 5839 14639 5937
tri 14639 5839 14737 5937 sw
tri 14737 5839 14835 5937 ne
rect 14835 5839 15189 5937
tri 15189 5839 15287 5937 sw
tri 15287 5839 15385 5937 ne
rect 15385 5839 15739 5937
tri 15739 5839 15837 5937 sw
tri 15837 5839 15935 5937 ne
rect 15935 5839 16289 5937
tri 16289 5839 16387 5937 sw
tri 16387 5839 16485 5937 ne
rect 16485 5839 16839 5937
tri 16839 5839 16937 5937 sw
tri 16937 5839 17035 5937 ne
rect 17035 5839 17389 5937
tri 17389 5839 17487 5937 sw
tri 17487 5839 17585 5937 ne
rect 17585 5839 17939 5937
tri 17939 5839 18037 5937 sw
tri 18037 5839 18135 5937 ne
rect 18135 5839 18489 5937
tri 18489 5839 18587 5937 sw
tri 18587 5839 18685 5937 ne
rect 18685 5839 19039 5937
tri 19039 5839 19137 5937 sw
tri 19137 5839 19235 5937 ne
rect 19235 5839 19589 5937
tri 19589 5839 19687 5937 sw
rect -500 5835 437 5839
rect -500 5715 215 5835
rect 335 5741 437 5835
tri 437 5741 535 5839 sw
tri 535 5741 633 5839 ne
rect 633 5835 987 5839
rect 633 5741 765 5835
rect 335 5715 535 5741
rect -500 5711 535 5715
tri 535 5711 565 5741 sw
tri 633 5711 663 5741 ne
rect 663 5715 765 5741
rect 885 5741 987 5835
tri 987 5741 1085 5839 sw
tri 1085 5741 1183 5839 ne
rect 1183 5835 1537 5839
rect 1183 5741 1315 5835
rect 885 5715 1085 5741
rect 663 5711 1085 5715
tri 1085 5711 1115 5741 sw
tri 1183 5711 1213 5741 ne
rect 1213 5715 1315 5741
rect 1435 5741 1537 5835
tri 1537 5741 1635 5839 sw
tri 1635 5741 1733 5839 ne
rect 1733 5835 2087 5839
rect 1733 5741 1865 5835
rect 1435 5715 1635 5741
rect 1213 5711 1635 5715
tri 1635 5711 1665 5741 sw
tri 1733 5711 1763 5741 ne
rect 1763 5715 1865 5741
rect 1985 5741 2087 5835
tri 2087 5741 2185 5839 sw
tri 2185 5741 2283 5839 ne
rect 2283 5835 2637 5839
rect 2283 5741 2415 5835
rect 1985 5715 2185 5741
rect 1763 5711 2185 5715
tri 2185 5711 2215 5741 sw
tri 2283 5711 2313 5741 ne
rect 2313 5715 2415 5741
rect 2535 5741 2637 5835
tri 2637 5741 2735 5839 sw
tri 2735 5741 2833 5839 ne
rect 2833 5835 3187 5839
rect 2833 5741 2965 5835
rect 2535 5715 2735 5741
rect 2313 5711 2735 5715
tri 2735 5711 2765 5741 sw
tri 2833 5711 2863 5741 ne
rect 2863 5715 2965 5741
rect 3085 5741 3187 5835
tri 3187 5741 3285 5839 sw
tri 3285 5741 3383 5839 ne
rect 3383 5835 3737 5839
rect 3383 5741 3515 5835
rect 3085 5715 3285 5741
rect 2863 5711 3285 5715
tri 3285 5711 3315 5741 sw
tri 3383 5711 3413 5741 ne
rect 3413 5715 3515 5741
rect 3635 5741 3737 5835
tri 3737 5741 3835 5839 sw
tri 3835 5741 3933 5839 ne
rect 3933 5835 4287 5839
rect 3933 5741 4065 5835
rect 3635 5715 3835 5741
rect 3413 5711 3835 5715
tri 3835 5711 3865 5741 sw
tri 3933 5711 3963 5741 ne
rect 3963 5715 4065 5741
rect 4185 5741 4287 5835
tri 4287 5741 4385 5839 sw
tri 4385 5741 4483 5839 ne
rect 4483 5835 4837 5839
rect 4483 5741 4615 5835
rect 4185 5715 4385 5741
rect 3963 5711 4385 5715
tri 4385 5711 4415 5741 sw
tri 4483 5711 4513 5741 ne
rect 4513 5715 4615 5741
rect 4735 5741 4837 5835
tri 4837 5741 4935 5839 sw
tri 4935 5741 5033 5839 ne
rect 5033 5835 5387 5839
rect 5033 5741 5165 5835
rect 4735 5715 4935 5741
rect 4513 5711 4935 5715
tri 4935 5711 4965 5741 sw
tri 5033 5711 5063 5741 ne
rect 5063 5715 5165 5741
rect 5285 5741 5387 5835
tri 5387 5741 5485 5839 sw
tri 5485 5741 5583 5839 ne
rect 5583 5835 5937 5839
rect 5583 5741 5715 5835
rect 5285 5715 5485 5741
rect 5063 5711 5485 5715
tri 5485 5711 5515 5741 sw
tri 5583 5711 5613 5741 ne
rect 5613 5715 5715 5741
rect 5835 5741 5937 5835
tri 5937 5741 6035 5839 sw
tri 6035 5741 6133 5839 ne
rect 6133 5835 6487 5839
rect 6133 5741 6265 5835
rect 5835 5715 6035 5741
rect 5613 5711 6035 5715
tri 6035 5711 6065 5741 sw
tri 6133 5711 6163 5741 ne
rect 6163 5715 6265 5741
rect 6385 5741 6487 5835
tri 6487 5741 6585 5839 sw
tri 6585 5741 6683 5839 ne
rect 6683 5835 7037 5839
rect 6683 5741 6815 5835
rect 6385 5715 6585 5741
rect 6163 5711 6585 5715
tri 6585 5711 6615 5741 sw
tri 6683 5711 6713 5741 ne
rect 6713 5715 6815 5741
rect 6935 5741 7037 5835
tri 7037 5741 7135 5839 sw
tri 7135 5741 7233 5839 ne
rect 7233 5835 7587 5839
rect 7233 5741 7365 5835
rect 6935 5715 7135 5741
rect 6713 5711 7135 5715
tri 7135 5711 7165 5741 sw
tri 7233 5711 7263 5741 ne
rect 7263 5715 7365 5741
rect 7485 5741 7587 5835
tri 7587 5741 7685 5839 sw
tri 7685 5741 7783 5839 ne
rect 7783 5835 8137 5839
rect 7783 5741 7915 5835
rect 7485 5715 7685 5741
rect 7263 5711 7685 5715
tri 7685 5711 7715 5741 sw
tri 7783 5711 7813 5741 ne
rect 7813 5715 7915 5741
rect 8035 5741 8137 5835
tri 8137 5741 8235 5839 sw
tri 8235 5741 8333 5839 ne
rect 8333 5835 8687 5839
rect 8333 5741 8465 5835
rect 8035 5715 8235 5741
rect 7813 5711 8235 5715
tri 8235 5711 8265 5741 sw
tri 8333 5711 8363 5741 ne
rect 8363 5715 8465 5741
rect 8585 5741 8687 5835
tri 8687 5741 8785 5839 sw
tri 8785 5741 8883 5839 ne
rect 8883 5835 9237 5839
rect 8883 5741 9015 5835
rect 8585 5715 8785 5741
rect 8363 5711 8785 5715
tri 8785 5711 8815 5741 sw
tri 8883 5711 8913 5741 ne
rect 8913 5715 9015 5741
rect 9135 5741 9237 5835
tri 9237 5741 9335 5839 sw
tri 9335 5741 9433 5839 ne
rect 9433 5835 9787 5839
rect 9433 5741 9565 5835
rect 9135 5715 9335 5741
rect 8913 5711 9335 5715
tri 9335 5711 9365 5741 sw
tri 9433 5711 9463 5741 ne
rect 9463 5715 9565 5741
rect 9685 5741 9787 5835
tri 9787 5741 9885 5839 sw
tri 9885 5741 9983 5839 ne
rect 9983 5835 10337 5839
rect 9983 5741 10115 5835
rect 9685 5715 9885 5741
rect 9463 5711 9885 5715
tri 9885 5711 9915 5741 sw
tri 9983 5711 10013 5741 ne
rect 10013 5715 10115 5741
rect 10235 5741 10337 5835
tri 10337 5741 10435 5839 sw
tri 10435 5741 10533 5839 ne
rect 10533 5835 10887 5839
rect 10533 5741 10665 5835
rect 10235 5715 10435 5741
rect 10013 5711 10435 5715
tri 10435 5711 10465 5741 sw
tri 10533 5711 10563 5741 ne
rect 10563 5715 10665 5741
rect 10785 5741 10887 5835
tri 10887 5741 10985 5839 sw
tri 10985 5741 11083 5839 ne
rect 11083 5835 11437 5839
rect 11083 5741 11215 5835
rect 10785 5715 10985 5741
rect 10563 5711 10985 5715
tri 10985 5711 11015 5741 sw
tri 11083 5711 11113 5741 ne
rect 11113 5715 11215 5741
rect 11335 5741 11437 5835
tri 11437 5741 11535 5839 sw
tri 11535 5741 11633 5839 ne
rect 11633 5835 11987 5839
rect 11633 5741 11765 5835
rect 11335 5715 11535 5741
rect 11113 5711 11535 5715
tri 11535 5711 11565 5741 sw
tri 11633 5711 11663 5741 ne
rect 11663 5715 11765 5741
rect 11885 5741 11987 5835
tri 11987 5741 12085 5839 sw
tri 12085 5741 12183 5839 ne
rect 12183 5835 12537 5839
rect 12183 5741 12315 5835
rect 11885 5715 12085 5741
rect 11663 5711 12085 5715
tri 12085 5711 12115 5741 sw
tri 12183 5711 12213 5741 ne
rect 12213 5715 12315 5741
rect 12435 5741 12537 5835
tri 12537 5741 12635 5839 sw
tri 12635 5741 12733 5839 ne
rect 12733 5835 13087 5839
rect 12733 5741 12865 5835
rect 12435 5715 12635 5741
rect 12213 5711 12635 5715
tri 12635 5711 12665 5741 sw
tri 12733 5711 12763 5741 ne
rect 12763 5715 12865 5741
rect 12985 5741 13087 5835
tri 13087 5741 13185 5839 sw
tri 13185 5741 13283 5839 ne
rect 13283 5835 13637 5839
rect 13283 5741 13415 5835
rect 12985 5715 13185 5741
rect 12763 5711 13185 5715
tri 13185 5711 13215 5741 sw
tri 13283 5711 13313 5741 ne
rect 13313 5715 13415 5741
rect 13535 5741 13637 5835
tri 13637 5741 13735 5839 sw
tri 13735 5741 13833 5839 ne
rect 13833 5835 14187 5839
rect 13833 5741 13965 5835
rect 13535 5715 13735 5741
rect 13313 5711 13735 5715
tri 13735 5711 13765 5741 sw
tri 13833 5711 13863 5741 ne
rect 13863 5715 13965 5741
rect 14085 5741 14187 5835
tri 14187 5741 14285 5839 sw
tri 14285 5741 14383 5839 ne
rect 14383 5835 14737 5839
rect 14383 5741 14515 5835
rect 14085 5715 14285 5741
rect 13863 5711 14285 5715
tri 14285 5711 14315 5741 sw
tri 14383 5711 14413 5741 ne
rect 14413 5715 14515 5741
rect 14635 5741 14737 5835
tri 14737 5741 14835 5839 sw
tri 14835 5741 14933 5839 ne
rect 14933 5835 15287 5839
rect 14933 5741 15065 5835
rect 14635 5715 14835 5741
rect 14413 5711 14835 5715
tri 14835 5711 14865 5741 sw
tri 14933 5711 14963 5741 ne
rect 14963 5715 15065 5741
rect 15185 5741 15287 5835
tri 15287 5741 15385 5839 sw
tri 15385 5741 15483 5839 ne
rect 15483 5835 15837 5839
rect 15483 5741 15615 5835
rect 15185 5715 15385 5741
rect 14963 5711 15385 5715
tri 15385 5711 15415 5741 sw
tri 15483 5711 15513 5741 ne
rect 15513 5715 15615 5741
rect 15735 5741 15837 5835
tri 15837 5741 15935 5839 sw
tri 15935 5741 16033 5839 ne
rect 16033 5835 16387 5839
rect 16033 5741 16165 5835
rect 15735 5715 15935 5741
rect 15513 5711 15935 5715
tri 15935 5711 15965 5741 sw
tri 16033 5711 16063 5741 ne
rect 16063 5715 16165 5741
rect 16285 5741 16387 5835
tri 16387 5741 16485 5839 sw
tri 16485 5741 16583 5839 ne
rect 16583 5835 16937 5839
rect 16583 5741 16715 5835
rect 16285 5715 16485 5741
rect 16063 5711 16485 5715
tri 16485 5711 16515 5741 sw
tri 16583 5711 16613 5741 ne
rect 16613 5715 16715 5741
rect 16835 5741 16937 5835
tri 16937 5741 17035 5839 sw
tri 17035 5741 17133 5839 ne
rect 17133 5835 17487 5839
rect 17133 5741 17265 5835
rect 16835 5715 17035 5741
rect 16613 5711 17035 5715
tri 17035 5711 17065 5741 sw
tri 17133 5711 17163 5741 ne
rect 17163 5715 17265 5741
rect 17385 5741 17487 5835
tri 17487 5741 17585 5839 sw
tri 17585 5741 17683 5839 ne
rect 17683 5835 18037 5839
rect 17683 5741 17815 5835
rect 17385 5715 17585 5741
rect 17163 5711 17585 5715
tri 17585 5711 17615 5741 sw
tri 17683 5711 17713 5741 ne
rect 17713 5715 17815 5741
rect 17935 5741 18037 5835
tri 18037 5741 18135 5839 sw
tri 18135 5741 18233 5839 ne
rect 18233 5835 18587 5839
rect 18233 5741 18365 5835
rect 17935 5715 18135 5741
rect 17713 5711 18135 5715
tri 18135 5711 18165 5741 sw
tri 18233 5711 18263 5741 ne
rect 18263 5715 18365 5741
rect 18485 5741 18587 5835
tri 18587 5741 18685 5839 sw
tri 18685 5741 18783 5839 ne
rect 18783 5835 19137 5839
rect 18783 5741 18915 5835
rect 18485 5715 18685 5741
rect 18263 5711 18685 5715
tri 18685 5711 18715 5741 sw
tri 18783 5711 18813 5741 ne
rect 18813 5715 18915 5741
rect 19035 5741 19137 5835
tri 19137 5741 19235 5839 sw
tri 19235 5741 19333 5839 ne
rect 19333 5835 20300 5839
rect 19333 5741 19465 5835
rect 19035 5715 19235 5741
rect 18813 5711 19235 5715
tri 19235 5711 19265 5741 sw
tri 19333 5711 19363 5741 ne
rect 19363 5715 19465 5741
rect 19585 5715 20300 5835
rect 19363 5711 20300 5715
tri 113 5613 211 5711 ne
rect 211 5613 565 5711
tri 565 5613 663 5711 sw
tri 663 5613 761 5711 ne
rect 761 5613 1115 5711
tri 1115 5613 1213 5711 sw
tri 1213 5613 1311 5711 ne
rect 1311 5613 1665 5711
tri 1665 5613 1763 5711 sw
tri 1763 5613 1861 5711 ne
rect 1861 5613 2215 5711
tri 2215 5613 2313 5711 sw
tri 2313 5613 2411 5711 ne
rect 2411 5613 2765 5711
tri 2765 5613 2863 5711 sw
tri 2863 5613 2961 5711 ne
rect 2961 5613 3315 5711
tri 3315 5613 3413 5711 sw
tri 3413 5613 3511 5711 ne
rect 3511 5613 3865 5711
tri 3865 5613 3963 5711 sw
tri 3963 5613 4061 5711 ne
rect 4061 5613 4415 5711
tri 4415 5613 4513 5711 sw
tri 4513 5613 4611 5711 ne
rect 4611 5613 4965 5711
tri 4965 5613 5063 5711 sw
tri 5063 5613 5161 5711 ne
rect 5161 5613 5515 5711
tri 5515 5613 5613 5711 sw
tri 5613 5613 5711 5711 ne
rect 5711 5613 6065 5711
tri 6065 5613 6163 5711 sw
tri 6163 5613 6261 5711 ne
rect 6261 5613 6615 5711
tri 6615 5613 6713 5711 sw
tri 6713 5613 6811 5711 ne
rect 6811 5613 7165 5711
tri 7165 5613 7263 5711 sw
tri 7263 5613 7361 5711 ne
rect 7361 5613 7715 5711
tri 7715 5613 7813 5711 sw
tri 7813 5613 7911 5711 ne
rect 7911 5613 8265 5711
tri 8265 5613 8363 5711 sw
tri 8363 5613 8461 5711 ne
rect 8461 5613 8815 5711
tri 8815 5613 8913 5711 sw
tri 8913 5613 9011 5711 ne
rect 9011 5613 9365 5711
tri 9365 5613 9463 5711 sw
tri 9463 5613 9561 5711 ne
rect 9561 5613 9915 5711
tri 9915 5613 10013 5711 sw
tri 10013 5613 10111 5711 ne
rect 10111 5613 10465 5711
tri 10465 5613 10563 5711 sw
tri 10563 5613 10661 5711 ne
rect 10661 5613 11015 5711
tri 11015 5613 11113 5711 sw
tri 11113 5613 11211 5711 ne
rect 11211 5613 11565 5711
tri 11565 5613 11663 5711 sw
tri 11663 5613 11761 5711 ne
rect 11761 5613 12115 5711
tri 12115 5613 12213 5711 sw
tri 12213 5613 12311 5711 ne
rect 12311 5613 12665 5711
tri 12665 5613 12763 5711 sw
tri 12763 5613 12861 5711 ne
rect 12861 5613 13215 5711
tri 13215 5613 13313 5711 sw
tri 13313 5613 13411 5711 ne
rect 13411 5613 13765 5711
tri 13765 5613 13863 5711 sw
tri 13863 5613 13961 5711 ne
rect 13961 5613 14315 5711
tri 14315 5613 14413 5711 sw
tri 14413 5613 14511 5711 ne
rect 14511 5613 14865 5711
tri 14865 5613 14963 5711 sw
tri 14963 5613 15061 5711 ne
rect 15061 5613 15415 5711
tri 15415 5613 15513 5711 sw
tri 15513 5613 15611 5711 ne
rect 15611 5613 15965 5711
tri 15965 5613 16063 5711 sw
tri 16063 5613 16161 5711 ne
rect 16161 5613 16515 5711
tri 16515 5613 16613 5711 sw
tri 16613 5613 16711 5711 ne
rect 16711 5613 17065 5711
tri 17065 5613 17163 5711 sw
tri 17163 5613 17261 5711 ne
rect 17261 5613 17615 5711
tri 17615 5613 17713 5711 sw
tri 17713 5613 17811 5711 ne
rect 17811 5613 18165 5711
tri 18165 5613 18263 5711 sw
tri 18263 5613 18361 5711 ne
rect 18361 5613 18715 5711
tri 18715 5613 18813 5711 sw
tri 18813 5613 18911 5711 ne
rect 18911 5613 19265 5711
tri 19265 5613 19363 5711 sw
tri 19363 5613 19461 5711 ne
rect 19461 5613 20300 5711
rect -2000 5583 113 5613
tri 113 5583 143 5613 sw
tri 211 5583 241 5613 ne
rect 241 5583 663 5613
tri 663 5583 693 5613 sw
tri 761 5583 791 5613 ne
rect 791 5583 1213 5613
tri 1213 5583 1243 5613 sw
tri 1311 5583 1341 5613 ne
rect 1341 5583 1763 5613
tri 1763 5583 1793 5613 sw
tri 1861 5583 1891 5613 ne
rect 1891 5583 2313 5613
tri 2313 5583 2343 5613 sw
tri 2411 5583 2441 5613 ne
rect 2441 5583 2863 5613
tri 2863 5583 2893 5613 sw
tri 2961 5583 2991 5613 ne
rect 2991 5583 3413 5613
tri 3413 5583 3443 5613 sw
tri 3511 5583 3541 5613 ne
rect 3541 5583 3963 5613
tri 3963 5583 3993 5613 sw
tri 4061 5583 4091 5613 ne
rect 4091 5583 4513 5613
tri 4513 5583 4543 5613 sw
tri 4611 5583 4641 5613 ne
rect 4641 5583 5063 5613
tri 5063 5583 5093 5613 sw
tri 5161 5583 5191 5613 ne
rect 5191 5583 5613 5613
tri 5613 5583 5643 5613 sw
tri 5711 5583 5741 5613 ne
rect 5741 5583 6163 5613
tri 6163 5583 6193 5613 sw
tri 6261 5583 6291 5613 ne
rect 6291 5583 6713 5613
tri 6713 5583 6743 5613 sw
tri 6811 5583 6841 5613 ne
rect 6841 5583 7263 5613
tri 7263 5583 7293 5613 sw
tri 7361 5583 7391 5613 ne
rect 7391 5583 7813 5613
tri 7813 5583 7843 5613 sw
tri 7911 5583 7941 5613 ne
rect 7941 5583 8363 5613
tri 8363 5583 8393 5613 sw
tri 8461 5583 8491 5613 ne
rect 8491 5583 8913 5613
tri 8913 5583 8943 5613 sw
tri 9011 5583 9041 5613 ne
rect 9041 5583 9463 5613
tri 9463 5583 9493 5613 sw
tri 9561 5583 9591 5613 ne
rect 9591 5583 10013 5613
tri 10013 5583 10043 5613 sw
tri 10111 5583 10141 5613 ne
rect 10141 5583 10563 5613
tri 10563 5583 10593 5613 sw
tri 10661 5583 10691 5613 ne
rect 10691 5583 11113 5613
tri 11113 5583 11143 5613 sw
tri 11211 5583 11241 5613 ne
rect 11241 5583 11663 5613
tri 11663 5583 11693 5613 sw
tri 11761 5583 11791 5613 ne
rect 11791 5583 12213 5613
tri 12213 5583 12243 5613 sw
tri 12311 5583 12341 5613 ne
rect 12341 5583 12763 5613
tri 12763 5583 12793 5613 sw
tri 12861 5583 12891 5613 ne
rect 12891 5583 13313 5613
tri 13313 5583 13343 5613 sw
tri 13411 5583 13441 5613 ne
rect 13441 5583 13863 5613
tri 13863 5583 13893 5613 sw
tri 13961 5583 13991 5613 ne
rect 13991 5583 14413 5613
tri 14413 5583 14443 5613 sw
tri 14511 5583 14541 5613 ne
rect 14541 5583 14963 5613
tri 14963 5583 14993 5613 sw
tri 15061 5583 15091 5613 ne
rect 15091 5583 15513 5613
tri 15513 5583 15543 5613 sw
tri 15611 5583 15641 5613 ne
rect 15641 5583 16063 5613
tri 16063 5583 16093 5613 sw
tri 16161 5583 16191 5613 ne
rect 16191 5583 16613 5613
tri 16613 5583 16643 5613 sw
tri 16711 5583 16741 5613 ne
rect 16741 5583 17163 5613
tri 17163 5583 17193 5613 sw
tri 17261 5583 17291 5613 ne
rect 17291 5583 17713 5613
tri 17713 5583 17743 5613 sw
tri 17811 5583 17841 5613 ne
rect 17841 5583 18263 5613
tri 18263 5583 18293 5613 sw
tri 18361 5583 18391 5613 ne
rect 18391 5583 18813 5613
tri 18813 5583 18843 5613 sw
tri 18911 5583 18941 5613 ne
rect 18941 5583 19363 5613
tri 19363 5583 19393 5613 sw
tri 19461 5583 19491 5613 ne
rect 19491 5583 20300 5613
rect -2000 5485 143 5583
tri 143 5485 241 5583 sw
tri 241 5485 339 5583 ne
rect 339 5485 693 5583
tri 693 5485 791 5583 sw
tri 791 5485 889 5583 ne
rect 889 5485 1243 5583
tri 1243 5485 1341 5583 sw
tri 1341 5485 1439 5583 ne
rect 1439 5485 1793 5583
tri 1793 5485 1891 5583 sw
tri 1891 5485 1989 5583 ne
rect 1989 5485 2343 5583
tri 2343 5485 2441 5583 sw
tri 2441 5485 2539 5583 ne
rect 2539 5485 2893 5583
tri 2893 5485 2991 5583 sw
tri 2991 5485 3089 5583 ne
rect 3089 5485 3443 5583
tri 3443 5485 3541 5583 sw
tri 3541 5485 3639 5583 ne
rect 3639 5485 3993 5583
tri 3993 5485 4091 5583 sw
tri 4091 5485 4189 5583 ne
rect 4189 5485 4543 5583
tri 4543 5485 4641 5583 sw
tri 4641 5485 4739 5583 ne
rect 4739 5485 5093 5583
tri 5093 5485 5191 5583 sw
tri 5191 5485 5289 5583 ne
rect 5289 5485 5643 5583
tri 5643 5485 5741 5583 sw
tri 5741 5485 5839 5583 ne
rect 5839 5485 6193 5583
tri 6193 5485 6291 5583 sw
tri 6291 5485 6389 5583 ne
rect 6389 5485 6743 5583
tri 6743 5485 6841 5583 sw
tri 6841 5485 6939 5583 ne
rect 6939 5485 7293 5583
tri 7293 5485 7391 5583 sw
tri 7391 5485 7489 5583 ne
rect 7489 5485 7843 5583
tri 7843 5485 7941 5583 sw
tri 7941 5485 8039 5583 ne
rect 8039 5485 8393 5583
tri 8393 5485 8491 5583 sw
tri 8491 5485 8589 5583 ne
rect 8589 5485 8943 5583
tri 8943 5485 9041 5583 sw
tri 9041 5485 9139 5583 ne
rect 9139 5485 9493 5583
tri 9493 5485 9591 5583 sw
tri 9591 5485 9689 5583 ne
rect 9689 5485 10043 5583
tri 10043 5485 10141 5583 sw
tri 10141 5485 10239 5583 ne
rect 10239 5485 10593 5583
tri 10593 5485 10691 5583 sw
tri 10691 5485 10789 5583 ne
rect 10789 5485 11143 5583
tri 11143 5485 11241 5583 sw
tri 11241 5485 11339 5583 ne
rect 11339 5485 11693 5583
tri 11693 5485 11791 5583 sw
tri 11791 5485 11889 5583 ne
rect 11889 5485 12243 5583
tri 12243 5485 12341 5583 sw
tri 12341 5485 12439 5583 ne
rect 12439 5485 12793 5583
tri 12793 5485 12891 5583 sw
tri 12891 5485 12989 5583 ne
rect 12989 5485 13343 5583
tri 13343 5485 13441 5583 sw
tri 13441 5485 13539 5583 ne
rect 13539 5485 13893 5583
tri 13893 5485 13991 5583 sw
tri 13991 5485 14089 5583 ne
rect 14089 5485 14443 5583
tri 14443 5485 14541 5583 sw
tri 14541 5485 14639 5583 ne
rect 14639 5485 14993 5583
tri 14993 5485 15091 5583 sw
tri 15091 5485 15189 5583 ne
rect 15189 5485 15543 5583
tri 15543 5485 15641 5583 sw
tri 15641 5485 15739 5583 ne
rect 15739 5485 16093 5583
tri 16093 5485 16191 5583 sw
tri 16191 5485 16289 5583 ne
rect 16289 5485 16643 5583
tri 16643 5485 16741 5583 sw
tri 16741 5485 16839 5583 ne
rect 16839 5485 17193 5583
tri 17193 5485 17291 5583 sw
tri 17291 5485 17389 5583 ne
rect 17389 5485 17743 5583
tri 17743 5485 17841 5583 sw
tri 17841 5485 17939 5583 ne
rect 17939 5485 18293 5583
tri 18293 5485 18391 5583 sw
tri 18391 5485 18489 5583 ne
rect 18489 5485 18843 5583
tri 18843 5485 18941 5583 sw
tri 18941 5485 19039 5583 ne
rect 19039 5485 19393 5583
tri 19393 5485 19491 5583 sw
tri 19491 5485 19589 5583 ne
rect 19589 5485 20300 5583
rect -2000 5387 241 5485
tri 241 5387 339 5485 sw
tri 339 5387 437 5485 ne
rect 437 5387 791 5485
tri 791 5387 889 5485 sw
tri 889 5387 987 5485 ne
rect 987 5387 1341 5485
tri 1341 5387 1439 5485 sw
tri 1439 5387 1537 5485 ne
rect 1537 5387 1891 5485
tri 1891 5387 1989 5485 sw
tri 1989 5387 2087 5485 ne
rect 2087 5387 2441 5485
tri 2441 5387 2539 5485 sw
tri 2539 5387 2637 5485 ne
rect 2637 5387 2991 5485
tri 2991 5387 3089 5485 sw
tri 3089 5387 3187 5485 ne
rect 3187 5387 3541 5485
tri 3541 5387 3639 5485 sw
tri 3639 5387 3737 5485 ne
rect 3737 5387 4091 5485
tri 4091 5387 4189 5485 sw
tri 4189 5387 4287 5485 ne
rect 4287 5387 4641 5485
tri 4641 5387 4739 5485 sw
tri 4739 5387 4837 5485 ne
rect 4837 5387 5191 5485
tri 5191 5387 5289 5485 sw
tri 5289 5387 5387 5485 ne
rect 5387 5387 5741 5485
tri 5741 5387 5839 5485 sw
tri 5839 5387 5937 5485 ne
rect 5937 5387 6291 5485
tri 6291 5387 6389 5485 sw
tri 6389 5387 6487 5485 ne
rect 6487 5387 6841 5485
tri 6841 5387 6939 5485 sw
tri 6939 5387 7037 5485 ne
rect 7037 5387 7391 5485
tri 7391 5387 7489 5485 sw
tri 7489 5387 7587 5485 ne
rect 7587 5387 7941 5485
tri 7941 5387 8039 5485 sw
tri 8039 5387 8137 5485 ne
rect 8137 5387 8491 5485
tri 8491 5387 8589 5485 sw
tri 8589 5387 8687 5485 ne
rect 8687 5387 9041 5485
tri 9041 5387 9139 5485 sw
tri 9139 5387 9237 5485 ne
rect 9237 5387 9591 5485
tri 9591 5387 9689 5485 sw
tri 9689 5387 9787 5485 ne
rect 9787 5387 10141 5485
tri 10141 5387 10239 5485 sw
tri 10239 5387 10337 5485 ne
rect 10337 5387 10691 5485
tri 10691 5387 10789 5485 sw
tri 10789 5387 10887 5485 ne
rect 10887 5387 11241 5485
tri 11241 5387 11339 5485 sw
tri 11339 5387 11437 5485 ne
rect 11437 5387 11791 5485
tri 11791 5387 11889 5485 sw
tri 11889 5387 11987 5485 ne
rect 11987 5387 12341 5485
tri 12341 5387 12439 5485 sw
tri 12439 5387 12537 5485 ne
rect 12537 5387 12891 5485
tri 12891 5387 12989 5485 sw
tri 12989 5387 13087 5485 ne
rect 13087 5387 13441 5485
tri 13441 5387 13539 5485 sw
tri 13539 5387 13637 5485 ne
rect 13637 5387 13991 5485
tri 13991 5387 14089 5485 sw
tri 14089 5387 14187 5485 ne
rect 14187 5387 14541 5485
tri 14541 5387 14639 5485 sw
tri 14639 5387 14737 5485 ne
rect 14737 5387 15091 5485
tri 15091 5387 15189 5485 sw
tri 15189 5387 15287 5485 ne
rect 15287 5387 15641 5485
tri 15641 5387 15739 5485 sw
tri 15739 5387 15837 5485 ne
rect 15837 5387 16191 5485
tri 16191 5387 16289 5485 sw
tri 16289 5387 16387 5485 ne
rect 16387 5387 16741 5485
tri 16741 5387 16839 5485 sw
tri 16839 5387 16937 5485 ne
rect 16937 5387 17291 5485
tri 17291 5387 17389 5485 sw
tri 17389 5387 17487 5485 ne
rect 17487 5387 17841 5485
tri 17841 5387 17939 5485 sw
tri 17939 5387 18037 5485 ne
rect 18037 5387 18391 5485
tri 18391 5387 18489 5485 sw
tri 18489 5387 18587 5485 ne
rect 18587 5387 18941 5485
tri 18941 5387 19039 5485 sw
tri 19039 5387 19137 5485 ne
rect 19137 5387 19491 5485
tri 19491 5387 19589 5485 sw
tri 19589 5387 19687 5485 ne
rect 19687 5387 20300 5485
rect -2000 5289 339 5387
tri 339 5289 437 5387 sw
tri 437 5289 535 5387 ne
rect 535 5289 889 5387
tri 889 5289 987 5387 sw
tri 987 5289 1085 5387 ne
rect 1085 5289 1439 5387
tri 1439 5289 1537 5387 sw
tri 1537 5289 1635 5387 ne
rect 1635 5289 1989 5387
tri 1989 5289 2087 5387 sw
tri 2087 5289 2185 5387 ne
rect 2185 5289 2539 5387
tri 2539 5289 2637 5387 sw
tri 2637 5289 2735 5387 ne
rect 2735 5289 3089 5387
tri 3089 5289 3187 5387 sw
tri 3187 5289 3285 5387 ne
rect 3285 5289 3639 5387
tri 3639 5289 3737 5387 sw
tri 3737 5289 3835 5387 ne
rect 3835 5289 4189 5387
tri 4189 5289 4287 5387 sw
tri 4287 5289 4385 5387 ne
rect 4385 5289 4739 5387
tri 4739 5289 4837 5387 sw
tri 4837 5289 4935 5387 ne
rect 4935 5289 5289 5387
tri 5289 5289 5387 5387 sw
tri 5387 5289 5485 5387 ne
rect 5485 5289 5839 5387
tri 5839 5289 5937 5387 sw
tri 5937 5289 6035 5387 ne
rect 6035 5289 6389 5387
tri 6389 5289 6487 5387 sw
tri 6487 5289 6585 5387 ne
rect 6585 5289 6939 5387
tri 6939 5289 7037 5387 sw
tri 7037 5289 7135 5387 ne
rect 7135 5289 7489 5387
tri 7489 5289 7587 5387 sw
tri 7587 5289 7685 5387 ne
rect 7685 5289 8039 5387
tri 8039 5289 8137 5387 sw
tri 8137 5289 8235 5387 ne
rect 8235 5289 8589 5387
tri 8589 5289 8687 5387 sw
tri 8687 5289 8785 5387 ne
rect 8785 5289 9139 5387
tri 9139 5289 9237 5387 sw
tri 9237 5289 9335 5387 ne
rect 9335 5289 9689 5387
tri 9689 5289 9787 5387 sw
tri 9787 5289 9885 5387 ne
rect 9885 5289 10239 5387
tri 10239 5289 10337 5387 sw
tri 10337 5289 10435 5387 ne
rect 10435 5289 10789 5387
tri 10789 5289 10887 5387 sw
tri 10887 5289 10985 5387 ne
rect 10985 5289 11339 5387
tri 11339 5289 11437 5387 sw
tri 11437 5289 11535 5387 ne
rect 11535 5289 11889 5387
tri 11889 5289 11987 5387 sw
tri 11987 5289 12085 5387 ne
rect 12085 5289 12439 5387
tri 12439 5289 12537 5387 sw
tri 12537 5289 12635 5387 ne
rect 12635 5289 12989 5387
tri 12989 5289 13087 5387 sw
tri 13087 5289 13185 5387 ne
rect 13185 5289 13539 5387
tri 13539 5289 13637 5387 sw
tri 13637 5289 13735 5387 ne
rect 13735 5289 14089 5387
tri 14089 5289 14187 5387 sw
tri 14187 5289 14285 5387 ne
rect 14285 5289 14639 5387
tri 14639 5289 14737 5387 sw
tri 14737 5289 14835 5387 ne
rect 14835 5289 15189 5387
tri 15189 5289 15287 5387 sw
tri 15287 5289 15385 5387 ne
rect 15385 5289 15739 5387
tri 15739 5289 15837 5387 sw
tri 15837 5289 15935 5387 ne
rect 15935 5289 16289 5387
tri 16289 5289 16387 5387 sw
tri 16387 5289 16485 5387 ne
rect 16485 5289 16839 5387
tri 16839 5289 16937 5387 sw
tri 16937 5289 17035 5387 ne
rect 17035 5289 17389 5387
tri 17389 5289 17487 5387 sw
tri 17487 5289 17585 5387 ne
rect 17585 5289 17939 5387
tri 17939 5289 18037 5387 sw
tri 18037 5289 18135 5387 ne
rect 18135 5289 18489 5387
tri 18489 5289 18587 5387 sw
tri 18587 5289 18685 5387 ne
rect 18685 5289 19039 5387
tri 19039 5289 19137 5387 sw
tri 19137 5289 19235 5387 ne
rect 19235 5289 19589 5387
tri 19589 5289 19687 5387 sw
rect 20800 5289 21800 5937
rect -2000 5285 437 5289
rect -2000 5165 215 5285
rect 335 5191 437 5285
tri 437 5191 535 5289 sw
tri 535 5191 633 5289 ne
rect 633 5285 987 5289
rect 633 5191 765 5285
rect 335 5165 535 5191
rect -2000 5161 535 5165
rect -2000 4513 -1000 5161
tri 113 5063 211 5161 ne
rect 211 5113 535 5161
tri 535 5113 613 5191 sw
tri 633 5113 711 5191 ne
rect 711 5165 765 5191
rect 885 5191 987 5285
tri 987 5191 1085 5289 sw
tri 1085 5191 1183 5289 ne
rect 1183 5285 1537 5289
rect 1183 5191 1315 5285
rect 885 5165 1085 5191
rect 711 5113 1085 5165
tri 1085 5113 1163 5191 sw
tri 1183 5113 1261 5191 ne
rect 1261 5165 1315 5191
rect 1435 5191 1537 5285
tri 1537 5191 1635 5289 sw
tri 1635 5191 1733 5289 ne
rect 1733 5285 2087 5289
rect 1733 5191 1865 5285
rect 1435 5165 1635 5191
rect 1261 5113 1635 5165
tri 1635 5113 1713 5191 sw
tri 1733 5113 1811 5191 ne
rect 1811 5165 1865 5191
rect 1985 5191 2087 5285
tri 2087 5191 2185 5289 sw
tri 2185 5191 2283 5289 ne
rect 2283 5285 2637 5289
rect 2283 5191 2415 5285
rect 1985 5165 2185 5191
rect 1811 5113 2185 5165
tri 2185 5113 2263 5191 sw
tri 2283 5113 2361 5191 ne
rect 2361 5165 2415 5191
rect 2535 5191 2637 5285
tri 2637 5191 2735 5289 sw
tri 2735 5191 2833 5289 ne
rect 2833 5285 3187 5289
rect 2833 5191 2965 5285
rect 2535 5165 2735 5191
rect 2361 5113 2735 5165
tri 2735 5113 2813 5191 sw
tri 2833 5113 2911 5191 ne
rect 2911 5165 2965 5191
rect 3085 5191 3187 5285
tri 3187 5191 3285 5289 sw
tri 3285 5191 3383 5289 ne
rect 3383 5285 3737 5289
rect 3383 5191 3515 5285
rect 3085 5165 3285 5191
rect 2911 5113 3285 5165
tri 3285 5113 3363 5191 sw
tri 3383 5113 3461 5191 ne
rect 3461 5165 3515 5191
rect 3635 5191 3737 5285
tri 3737 5191 3835 5289 sw
tri 3835 5191 3933 5289 ne
rect 3933 5285 4287 5289
rect 3933 5191 4065 5285
rect 3635 5165 3835 5191
rect 3461 5113 3835 5165
tri 3835 5113 3913 5191 sw
tri 3933 5113 4011 5191 ne
rect 4011 5165 4065 5191
rect 4185 5191 4287 5285
tri 4287 5191 4385 5289 sw
tri 4385 5191 4483 5289 ne
rect 4483 5285 4837 5289
rect 4483 5191 4615 5285
rect 4185 5165 4385 5191
rect 4011 5113 4385 5165
tri 4385 5113 4463 5191 sw
tri 4483 5113 4561 5191 ne
rect 4561 5165 4615 5191
rect 4735 5191 4837 5285
tri 4837 5191 4935 5289 sw
tri 4935 5191 5033 5289 ne
rect 5033 5285 5387 5289
rect 5033 5191 5165 5285
rect 4735 5165 4935 5191
rect 4561 5113 4935 5165
tri 4935 5113 5013 5191 sw
tri 5033 5113 5111 5191 ne
rect 5111 5165 5165 5191
rect 5285 5191 5387 5285
tri 5387 5191 5485 5289 sw
tri 5485 5191 5583 5289 ne
rect 5583 5285 5937 5289
rect 5583 5191 5715 5285
rect 5285 5165 5485 5191
rect 5111 5113 5485 5165
tri 5485 5113 5563 5191 sw
tri 5583 5113 5661 5191 ne
rect 5661 5165 5715 5191
rect 5835 5191 5937 5285
tri 5937 5191 6035 5289 sw
tri 6035 5191 6133 5289 ne
rect 6133 5285 6487 5289
rect 6133 5191 6265 5285
rect 5835 5165 6035 5191
rect 5661 5113 6035 5165
tri 6035 5113 6113 5191 sw
tri 6133 5113 6211 5191 ne
rect 6211 5165 6265 5191
rect 6385 5191 6487 5285
tri 6487 5191 6585 5289 sw
tri 6585 5191 6683 5289 ne
rect 6683 5285 7037 5289
rect 6683 5191 6815 5285
rect 6385 5165 6585 5191
rect 6211 5113 6585 5165
tri 6585 5113 6663 5191 sw
tri 6683 5113 6761 5191 ne
rect 6761 5165 6815 5191
rect 6935 5191 7037 5285
tri 7037 5191 7135 5289 sw
tri 7135 5191 7233 5289 ne
rect 7233 5285 7587 5289
rect 7233 5191 7365 5285
rect 6935 5165 7135 5191
rect 6761 5113 7135 5165
tri 7135 5113 7213 5191 sw
tri 7233 5113 7311 5191 ne
rect 7311 5165 7365 5191
rect 7485 5191 7587 5285
tri 7587 5191 7685 5289 sw
tri 7685 5191 7783 5289 ne
rect 7783 5285 8137 5289
rect 7783 5191 7915 5285
rect 7485 5165 7685 5191
rect 7311 5113 7685 5165
tri 7685 5113 7763 5191 sw
tri 7783 5113 7861 5191 ne
rect 7861 5165 7915 5191
rect 8035 5191 8137 5285
tri 8137 5191 8235 5289 sw
tri 8235 5191 8333 5289 ne
rect 8333 5285 8687 5289
rect 8333 5191 8465 5285
rect 8035 5165 8235 5191
rect 7861 5113 8235 5165
tri 8235 5113 8313 5191 sw
tri 8333 5113 8411 5191 ne
rect 8411 5165 8465 5191
rect 8585 5191 8687 5285
tri 8687 5191 8785 5289 sw
tri 8785 5191 8883 5289 ne
rect 8883 5285 9237 5289
rect 8883 5191 9015 5285
rect 8585 5165 8785 5191
rect 8411 5113 8785 5165
tri 8785 5113 8863 5191 sw
tri 8883 5113 8961 5191 ne
rect 8961 5165 9015 5191
rect 9135 5191 9237 5285
tri 9237 5191 9335 5289 sw
tri 9335 5191 9433 5289 ne
rect 9433 5285 9787 5289
rect 9433 5191 9565 5285
rect 9135 5165 9335 5191
rect 8961 5113 9335 5165
tri 9335 5113 9413 5191 sw
tri 9433 5113 9511 5191 ne
rect 9511 5165 9565 5191
rect 9685 5191 9787 5285
tri 9787 5191 9885 5289 sw
tri 9885 5191 9983 5289 ne
rect 9983 5285 10337 5289
rect 9983 5191 10115 5285
rect 9685 5165 9885 5191
rect 9511 5113 9885 5165
tri 9885 5113 9963 5191 sw
tri 9983 5113 10061 5191 ne
rect 10061 5165 10115 5191
rect 10235 5191 10337 5285
tri 10337 5191 10435 5289 sw
tri 10435 5191 10533 5289 ne
rect 10533 5285 10887 5289
rect 10533 5191 10665 5285
rect 10235 5165 10435 5191
rect 10061 5113 10435 5165
tri 10435 5113 10513 5191 sw
tri 10533 5113 10611 5191 ne
rect 10611 5165 10665 5191
rect 10785 5191 10887 5285
tri 10887 5191 10985 5289 sw
tri 10985 5191 11083 5289 ne
rect 11083 5285 11437 5289
rect 11083 5191 11215 5285
rect 10785 5165 10985 5191
rect 10611 5113 10985 5165
tri 10985 5113 11063 5191 sw
tri 11083 5113 11161 5191 ne
rect 11161 5165 11215 5191
rect 11335 5191 11437 5285
tri 11437 5191 11535 5289 sw
tri 11535 5191 11633 5289 ne
rect 11633 5285 11987 5289
rect 11633 5191 11765 5285
rect 11335 5165 11535 5191
rect 11161 5113 11535 5165
tri 11535 5113 11613 5191 sw
tri 11633 5113 11711 5191 ne
rect 11711 5165 11765 5191
rect 11885 5191 11987 5285
tri 11987 5191 12085 5289 sw
tri 12085 5191 12183 5289 ne
rect 12183 5285 12537 5289
rect 12183 5191 12315 5285
rect 11885 5165 12085 5191
rect 11711 5113 12085 5165
tri 12085 5113 12163 5191 sw
tri 12183 5113 12261 5191 ne
rect 12261 5165 12315 5191
rect 12435 5191 12537 5285
tri 12537 5191 12635 5289 sw
tri 12635 5191 12733 5289 ne
rect 12733 5285 13087 5289
rect 12733 5191 12865 5285
rect 12435 5165 12635 5191
rect 12261 5113 12635 5165
tri 12635 5113 12713 5191 sw
tri 12733 5113 12811 5191 ne
rect 12811 5165 12865 5191
rect 12985 5191 13087 5285
tri 13087 5191 13185 5289 sw
tri 13185 5191 13283 5289 ne
rect 13283 5285 13637 5289
rect 13283 5191 13415 5285
rect 12985 5165 13185 5191
rect 12811 5113 13185 5165
tri 13185 5113 13263 5191 sw
tri 13283 5113 13361 5191 ne
rect 13361 5165 13415 5191
rect 13535 5191 13637 5285
tri 13637 5191 13735 5289 sw
tri 13735 5191 13833 5289 ne
rect 13833 5285 14187 5289
rect 13833 5191 13965 5285
rect 13535 5165 13735 5191
rect 13361 5113 13735 5165
tri 13735 5113 13813 5191 sw
tri 13833 5113 13911 5191 ne
rect 13911 5165 13965 5191
rect 14085 5191 14187 5285
tri 14187 5191 14285 5289 sw
tri 14285 5191 14383 5289 ne
rect 14383 5285 14737 5289
rect 14383 5191 14515 5285
rect 14085 5165 14285 5191
rect 13911 5113 14285 5165
tri 14285 5113 14363 5191 sw
tri 14383 5113 14461 5191 ne
rect 14461 5165 14515 5191
rect 14635 5191 14737 5285
tri 14737 5191 14835 5289 sw
tri 14835 5191 14933 5289 ne
rect 14933 5285 15287 5289
rect 14933 5191 15065 5285
rect 14635 5165 14835 5191
rect 14461 5113 14835 5165
tri 14835 5113 14913 5191 sw
tri 14933 5113 15011 5191 ne
rect 15011 5165 15065 5191
rect 15185 5191 15287 5285
tri 15287 5191 15385 5289 sw
tri 15385 5191 15483 5289 ne
rect 15483 5285 15837 5289
rect 15483 5191 15615 5285
rect 15185 5165 15385 5191
rect 15011 5113 15385 5165
tri 15385 5113 15463 5191 sw
tri 15483 5113 15561 5191 ne
rect 15561 5165 15615 5191
rect 15735 5191 15837 5285
tri 15837 5191 15935 5289 sw
tri 15935 5191 16033 5289 ne
rect 16033 5285 16387 5289
rect 16033 5191 16165 5285
rect 15735 5165 15935 5191
rect 15561 5113 15935 5165
tri 15935 5113 16013 5191 sw
tri 16033 5113 16111 5191 ne
rect 16111 5165 16165 5191
rect 16285 5191 16387 5285
tri 16387 5191 16485 5289 sw
tri 16485 5191 16583 5289 ne
rect 16583 5285 16937 5289
rect 16583 5191 16715 5285
rect 16285 5165 16485 5191
rect 16111 5113 16485 5165
tri 16485 5113 16563 5191 sw
tri 16583 5113 16661 5191 ne
rect 16661 5165 16715 5191
rect 16835 5191 16937 5285
tri 16937 5191 17035 5289 sw
tri 17035 5191 17133 5289 ne
rect 17133 5285 17487 5289
rect 17133 5191 17265 5285
rect 16835 5165 17035 5191
rect 16661 5113 17035 5165
tri 17035 5113 17113 5191 sw
tri 17133 5113 17211 5191 ne
rect 17211 5165 17265 5191
rect 17385 5191 17487 5285
tri 17487 5191 17585 5289 sw
tri 17585 5191 17683 5289 ne
rect 17683 5285 18037 5289
rect 17683 5191 17815 5285
rect 17385 5165 17585 5191
rect 17211 5113 17585 5165
tri 17585 5113 17663 5191 sw
tri 17683 5113 17761 5191 ne
rect 17761 5165 17815 5191
rect 17935 5191 18037 5285
tri 18037 5191 18135 5289 sw
tri 18135 5191 18233 5289 ne
rect 18233 5285 18587 5289
rect 18233 5191 18365 5285
rect 17935 5165 18135 5191
rect 17761 5113 18135 5165
tri 18135 5113 18213 5191 sw
tri 18233 5113 18311 5191 ne
rect 18311 5165 18365 5191
rect 18485 5191 18587 5285
tri 18587 5191 18685 5289 sw
tri 18685 5191 18783 5289 ne
rect 18783 5285 19137 5289
rect 18783 5191 18915 5285
rect 18485 5165 18685 5191
rect 18311 5113 18685 5165
tri 18685 5113 18763 5191 sw
tri 18783 5113 18861 5191 ne
rect 18861 5165 18915 5191
rect 19035 5191 19137 5285
tri 19137 5191 19235 5289 sw
tri 19235 5191 19333 5289 ne
rect 19333 5285 21800 5289
rect 19333 5191 19465 5285
rect 19035 5165 19235 5191
rect 18861 5113 19235 5165
tri 19235 5113 19313 5191 sw
tri 19333 5113 19411 5191 ne
rect 19411 5165 19465 5191
rect 19585 5165 21800 5285
rect 19411 5113 21800 5165
rect 211 5063 613 5113
rect -500 5013 113 5063
tri 113 5013 163 5063 sw
tri 211 5013 261 5063 ne
rect 261 5033 613 5063
tri 613 5033 693 5113 sw
tri 711 5033 791 5113 ne
rect 791 5033 1163 5113
tri 1163 5033 1243 5113 sw
tri 1261 5033 1341 5113 ne
rect 1341 5033 1713 5113
tri 1713 5033 1793 5113 sw
tri 1811 5033 1891 5113 ne
rect 1891 5033 2263 5113
tri 2263 5033 2343 5113 sw
tri 2361 5033 2441 5113 ne
rect 2441 5033 2813 5113
tri 2813 5033 2893 5113 sw
tri 2911 5033 2991 5113 ne
rect 2991 5033 3363 5113
tri 3363 5033 3443 5113 sw
tri 3461 5033 3541 5113 ne
rect 3541 5033 3913 5113
tri 3913 5033 3993 5113 sw
tri 4011 5033 4091 5113 ne
rect 4091 5033 4463 5113
tri 4463 5033 4543 5113 sw
tri 4561 5033 4641 5113 ne
rect 4641 5033 5013 5113
tri 5013 5033 5093 5113 sw
tri 5111 5033 5191 5113 ne
rect 5191 5033 5563 5113
tri 5563 5033 5643 5113 sw
tri 5661 5033 5741 5113 ne
rect 5741 5033 6113 5113
tri 6113 5033 6193 5113 sw
tri 6211 5033 6291 5113 ne
rect 6291 5033 6663 5113
tri 6663 5033 6743 5113 sw
tri 6761 5033 6841 5113 ne
rect 6841 5033 7213 5113
tri 7213 5033 7293 5113 sw
tri 7311 5033 7391 5113 ne
rect 7391 5033 7763 5113
tri 7763 5033 7843 5113 sw
tri 7861 5033 7941 5113 ne
rect 7941 5033 8313 5113
tri 8313 5033 8393 5113 sw
tri 8411 5033 8491 5113 ne
rect 8491 5033 8863 5113
tri 8863 5033 8943 5113 sw
tri 8961 5033 9041 5113 ne
rect 9041 5033 9413 5113
tri 9413 5033 9493 5113 sw
tri 9511 5033 9591 5113 ne
rect 9591 5033 9963 5113
tri 9963 5033 10043 5113 sw
tri 10061 5033 10141 5113 ne
rect 10141 5033 10513 5113
tri 10513 5033 10593 5113 sw
tri 10611 5033 10691 5113 ne
rect 10691 5033 11063 5113
tri 11063 5033 11143 5113 sw
tri 11161 5033 11241 5113 ne
rect 11241 5033 11613 5113
tri 11613 5033 11693 5113 sw
tri 11711 5033 11791 5113 ne
rect 11791 5033 12163 5113
tri 12163 5033 12243 5113 sw
tri 12261 5033 12341 5113 ne
rect 12341 5033 12713 5113
tri 12713 5033 12793 5113 sw
tri 12811 5033 12891 5113 ne
rect 12891 5033 13263 5113
tri 13263 5033 13343 5113 sw
tri 13361 5033 13441 5113 ne
rect 13441 5033 13813 5113
tri 13813 5033 13893 5113 sw
tri 13911 5033 13991 5113 ne
rect 13991 5033 14363 5113
tri 14363 5033 14443 5113 sw
tri 14461 5033 14541 5113 ne
rect 14541 5033 14913 5113
tri 14913 5033 14993 5113 sw
tri 15011 5033 15091 5113 ne
rect 15091 5033 15463 5113
tri 15463 5033 15543 5113 sw
tri 15561 5033 15641 5113 ne
rect 15641 5033 16013 5113
tri 16013 5033 16093 5113 sw
tri 16111 5033 16191 5113 ne
rect 16191 5033 16563 5113
tri 16563 5033 16643 5113 sw
tri 16661 5033 16741 5113 ne
rect 16741 5033 17113 5113
tri 17113 5033 17193 5113 sw
tri 17211 5033 17291 5113 ne
rect 17291 5033 17663 5113
tri 17663 5033 17743 5113 sw
tri 17761 5033 17841 5113 ne
rect 17841 5033 18213 5113
tri 18213 5033 18293 5113 sw
tri 18311 5033 18391 5113 ne
rect 18391 5033 18763 5113
tri 18763 5033 18843 5113 sw
tri 18861 5033 18941 5113 ne
rect 18941 5033 19313 5113
tri 19313 5033 19393 5113 sw
tri 19411 5033 19491 5113 ne
rect 19491 5033 20100 5113
rect 261 5013 693 5033
rect -500 4935 163 5013
tri 163 4935 241 5013 sw
tri 261 4935 339 5013 ne
rect 339 4935 693 5013
tri 693 4935 791 5033 sw
tri 791 4935 889 5033 ne
rect 889 4935 1243 5033
tri 1243 4935 1341 5033 sw
tri 1341 4935 1439 5033 ne
rect 1439 4935 1793 5033
tri 1793 4935 1891 5033 sw
tri 1891 4935 1989 5033 ne
rect 1989 4935 2343 5033
tri 2343 4935 2441 5033 sw
tri 2441 4935 2539 5033 ne
rect 2539 4935 2893 5033
tri 2893 4935 2991 5033 sw
tri 2991 4935 3089 5033 ne
rect 3089 4935 3443 5033
tri 3443 4935 3541 5033 sw
tri 3541 4935 3639 5033 ne
rect 3639 4935 3993 5033
tri 3993 4935 4091 5033 sw
tri 4091 4935 4189 5033 ne
rect 4189 4935 4543 5033
tri 4543 4935 4641 5033 sw
tri 4641 4935 4739 5033 ne
rect 4739 4935 5093 5033
tri 5093 4935 5191 5033 sw
tri 5191 4935 5289 5033 ne
rect 5289 4935 5643 5033
tri 5643 4935 5741 5033 sw
tri 5741 4935 5839 5033 ne
rect 5839 4935 6193 5033
tri 6193 4935 6291 5033 sw
tri 6291 4935 6389 5033 ne
rect 6389 4935 6743 5033
tri 6743 4935 6841 5033 sw
tri 6841 4935 6939 5033 ne
rect 6939 4935 7293 5033
tri 7293 4935 7391 5033 sw
tri 7391 4935 7489 5033 ne
rect 7489 4935 7843 5033
tri 7843 4935 7941 5033 sw
tri 7941 4935 8039 5033 ne
rect 8039 4935 8393 5033
tri 8393 4935 8491 5033 sw
tri 8491 4935 8589 5033 ne
rect 8589 4935 8943 5033
tri 8943 4935 9041 5033 sw
tri 9041 4935 9139 5033 ne
rect 9139 4935 9493 5033
tri 9493 4935 9591 5033 sw
tri 9591 4935 9689 5033 ne
rect 9689 4935 10043 5033
tri 10043 4935 10141 5033 sw
tri 10141 4935 10239 5033 ne
rect 10239 4935 10593 5033
tri 10593 4935 10691 5033 sw
tri 10691 4935 10789 5033 ne
rect 10789 4935 11143 5033
tri 11143 4935 11241 5033 sw
tri 11241 4935 11339 5033 ne
rect 11339 4935 11693 5033
tri 11693 4935 11791 5033 sw
tri 11791 4935 11889 5033 ne
rect 11889 4935 12243 5033
tri 12243 4935 12341 5033 sw
tri 12341 4935 12439 5033 ne
rect 12439 4935 12793 5033
tri 12793 4935 12891 5033 sw
tri 12891 4935 12989 5033 ne
rect 12989 4935 13343 5033
tri 13343 4935 13441 5033 sw
tri 13441 4935 13539 5033 ne
rect 13539 4935 13893 5033
tri 13893 4935 13991 5033 sw
tri 13991 4935 14089 5033 ne
rect 14089 4935 14443 5033
tri 14443 4935 14541 5033 sw
tri 14541 4935 14639 5033 ne
rect 14639 4935 14993 5033
tri 14993 4935 15091 5033 sw
tri 15091 4935 15189 5033 ne
rect 15189 4935 15543 5033
tri 15543 4935 15641 5033 sw
tri 15641 4935 15739 5033 ne
rect 15739 4935 16093 5033
tri 16093 4935 16191 5033 sw
tri 16191 4935 16289 5033 ne
rect 16289 4935 16643 5033
tri 16643 4935 16741 5033 sw
tri 16741 4935 16839 5033 ne
rect 16839 4935 17193 5033
tri 17193 4935 17291 5033 sw
tri 17291 4935 17389 5033 ne
rect 17389 4935 17743 5033
tri 17743 4935 17841 5033 sw
tri 17841 4935 17939 5033 ne
rect 17939 4935 18293 5033
tri 18293 4935 18391 5033 sw
tri 18391 4935 18489 5033 ne
rect 18489 4935 18843 5033
tri 18843 4935 18941 5033 sw
tri 18941 4935 19039 5033 ne
rect 19039 4935 19393 5033
tri 19393 4935 19491 5033 sw
tri 19491 4935 19589 5033 ne
rect 19589 5013 20100 5033
rect 20200 5013 21800 5113
rect 19589 4935 21800 5013
rect -500 4887 241 4935
rect -500 4787 -400 4887
rect -300 4837 241 4887
tri 241 4837 339 4935 sw
tri 339 4837 437 4935 ne
rect 437 4837 791 4935
tri 791 4837 889 4935 sw
tri 889 4837 987 4935 ne
rect 987 4837 1341 4935
tri 1341 4837 1439 4935 sw
tri 1439 4837 1537 4935 ne
rect 1537 4837 1891 4935
tri 1891 4837 1989 4935 sw
tri 1989 4837 2087 4935 ne
rect 2087 4837 2441 4935
tri 2441 4837 2539 4935 sw
tri 2539 4837 2637 4935 ne
rect 2637 4837 2991 4935
tri 2991 4837 3089 4935 sw
tri 3089 4837 3187 4935 ne
rect 3187 4837 3541 4935
tri 3541 4837 3639 4935 sw
tri 3639 4837 3737 4935 ne
rect 3737 4837 4091 4935
tri 4091 4837 4189 4935 sw
tri 4189 4837 4287 4935 ne
rect 4287 4837 4641 4935
tri 4641 4837 4739 4935 sw
tri 4739 4837 4837 4935 ne
rect 4837 4837 5191 4935
tri 5191 4837 5289 4935 sw
tri 5289 4837 5387 4935 ne
rect 5387 4837 5741 4935
tri 5741 4837 5839 4935 sw
tri 5839 4837 5937 4935 ne
rect 5937 4837 6291 4935
tri 6291 4837 6389 4935 sw
tri 6389 4837 6487 4935 ne
rect 6487 4837 6841 4935
tri 6841 4837 6939 4935 sw
tri 6939 4837 7037 4935 ne
rect 7037 4837 7391 4935
tri 7391 4837 7489 4935 sw
tri 7489 4837 7587 4935 ne
rect 7587 4837 7941 4935
tri 7941 4837 8039 4935 sw
tri 8039 4837 8137 4935 ne
rect 8137 4837 8491 4935
tri 8491 4837 8589 4935 sw
tri 8589 4837 8687 4935 ne
rect 8687 4837 9041 4935
tri 9041 4837 9139 4935 sw
tri 9139 4837 9237 4935 ne
rect 9237 4837 9591 4935
tri 9591 4837 9689 4935 sw
tri 9689 4837 9787 4935 ne
rect 9787 4837 10141 4935
tri 10141 4837 10239 4935 sw
tri 10239 4837 10337 4935 ne
rect 10337 4837 10691 4935
tri 10691 4837 10789 4935 sw
tri 10789 4837 10887 4935 ne
rect 10887 4837 11241 4935
tri 11241 4837 11339 4935 sw
tri 11339 4837 11437 4935 ne
rect 11437 4837 11791 4935
tri 11791 4837 11889 4935 sw
tri 11889 4837 11987 4935 ne
rect 11987 4837 12341 4935
tri 12341 4837 12439 4935 sw
tri 12439 4837 12537 4935 ne
rect 12537 4837 12891 4935
tri 12891 4837 12989 4935 sw
tri 12989 4837 13087 4935 ne
rect 13087 4837 13441 4935
tri 13441 4837 13539 4935 sw
tri 13539 4837 13637 4935 ne
rect 13637 4837 13991 4935
tri 13991 4837 14089 4935 sw
tri 14089 4837 14187 4935 ne
rect 14187 4837 14541 4935
tri 14541 4837 14639 4935 sw
tri 14639 4837 14737 4935 ne
rect 14737 4837 15091 4935
tri 15091 4837 15189 4935 sw
tri 15189 4837 15287 4935 ne
rect 15287 4837 15641 4935
tri 15641 4837 15739 4935 sw
tri 15739 4837 15837 4935 ne
rect 15837 4837 16191 4935
tri 16191 4837 16289 4935 sw
tri 16289 4837 16387 4935 ne
rect 16387 4837 16741 4935
tri 16741 4837 16839 4935 sw
tri 16839 4837 16937 4935 ne
rect 16937 4837 17291 4935
tri 17291 4837 17389 4935 sw
tri 17389 4837 17487 4935 ne
rect 17487 4837 17841 4935
tri 17841 4837 17939 4935 sw
tri 17939 4837 18037 4935 ne
rect 18037 4837 18391 4935
tri 18391 4837 18489 4935 sw
tri 18489 4837 18587 4935 ne
rect 18587 4837 18941 4935
tri 18941 4837 19039 4935 sw
tri 19039 4837 19137 4935 ne
rect 19137 4837 19491 4935
tri 19491 4837 19589 4935 sw
tri 19589 4837 19687 4935 ne
rect 19687 4837 21800 4935
rect -300 4787 339 4837
rect -500 4739 339 4787
tri 339 4739 437 4837 sw
tri 437 4739 535 4837 ne
rect 535 4739 889 4837
tri 889 4739 987 4837 sw
tri 987 4739 1085 4837 ne
rect 1085 4739 1439 4837
tri 1439 4739 1537 4837 sw
tri 1537 4739 1635 4837 ne
rect 1635 4739 1989 4837
tri 1989 4739 2087 4837 sw
tri 2087 4739 2185 4837 ne
rect 2185 4739 2539 4837
tri 2539 4739 2637 4837 sw
tri 2637 4739 2735 4837 ne
rect 2735 4739 3089 4837
tri 3089 4739 3187 4837 sw
tri 3187 4739 3285 4837 ne
rect 3285 4739 3639 4837
tri 3639 4739 3737 4837 sw
tri 3737 4739 3835 4837 ne
rect 3835 4739 4189 4837
tri 4189 4739 4287 4837 sw
tri 4287 4739 4385 4837 ne
rect 4385 4739 4739 4837
tri 4739 4739 4837 4837 sw
tri 4837 4739 4935 4837 ne
rect 4935 4739 5289 4837
tri 5289 4739 5387 4837 sw
tri 5387 4739 5485 4837 ne
rect 5485 4739 5839 4837
tri 5839 4739 5937 4837 sw
tri 5937 4739 6035 4837 ne
rect 6035 4739 6389 4837
tri 6389 4739 6487 4837 sw
tri 6487 4739 6585 4837 ne
rect 6585 4739 6939 4837
tri 6939 4739 7037 4837 sw
tri 7037 4739 7135 4837 ne
rect 7135 4739 7489 4837
tri 7489 4739 7587 4837 sw
tri 7587 4739 7685 4837 ne
rect 7685 4739 8039 4837
tri 8039 4739 8137 4837 sw
tri 8137 4739 8235 4837 ne
rect 8235 4739 8589 4837
tri 8589 4739 8687 4837 sw
tri 8687 4739 8785 4837 ne
rect 8785 4739 9139 4837
tri 9139 4739 9237 4837 sw
tri 9237 4739 9335 4837 ne
rect 9335 4739 9689 4837
tri 9689 4739 9787 4837 sw
tri 9787 4739 9885 4837 ne
rect 9885 4739 10239 4837
tri 10239 4739 10337 4837 sw
tri 10337 4739 10435 4837 ne
rect 10435 4739 10789 4837
tri 10789 4739 10887 4837 sw
tri 10887 4739 10985 4837 ne
rect 10985 4739 11339 4837
tri 11339 4739 11437 4837 sw
tri 11437 4739 11535 4837 ne
rect 11535 4739 11889 4837
tri 11889 4739 11987 4837 sw
tri 11987 4739 12085 4837 ne
rect 12085 4739 12439 4837
tri 12439 4739 12537 4837 sw
tri 12537 4739 12635 4837 ne
rect 12635 4739 12989 4837
tri 12989 4739 13087 4837 sw
tri 13087 4739 13185 4837 ne
rect 13185 4739 13539 4837
tri 13539 4739 13637 4837 sw
tri 13637 4739 13735 4837 ne
rect 13735 4739 14089 4837
tri 14089 4739 14187 4837 sw
tri 14187 4739 14285 4837 ne
rect 14285 4739 14639 4837
tri 14639 4739 14737 4837 sw
tri 14737 4739 14835 4837 ne
rect 14835 4739 15189 4837
tri 15189 4739 15287 4837 sw
tri 15287 4739 15385 4837 ne
rect 15385 4739 15739 4837
tri 15739 4739 15837 4837 sw
tri 15837 4739 15935 4837 ne
rect 15935 4739 16289 4837
tri 16289 4739 16387 4837 sw
tri 16387 4739 16485 4837 ne
rect 16485 4739 16839 4837
tri 16839 4739 16937 4837 sw
tri 16937 4739 17035 4837 ne
rect 17035 4739 17389 4837
tri 17389 4739 17487 4837 sw
tri 17487 4739 17585 4837 ne
rect 17585 4739 17939 4837
tri 17939 4739 18037 4837 sw
tri 18037 4739 18135 4837 ne
rect 18135 4739 18489 4837
tri 18489 4739 18587 4837 sw
tri 18587 4739 18685 4837 ne
rect 18685 4739 19039 4837
tri 19039 4739 19137 4837 sw
tri 19137 4739 19235 4837 ne
rect 19235 4739 19589 4837
tri 19589 4739 19687 4837 sw
rect -500 4735 437 4739
rect -500 4615 215 4735
rect 335 4641 437 4735
tri 437 4641 535 4739 sw
tri 535 4641 633 4739 ne
rect 633 4735 987 4739
rect 633 4641 765 4735
rect 335 4615 535 4641
rect -500 4611 535 4615
tri 535 4611 565 4641 sw
tri 633 4611 663 4641 ne
rect 663 4615 765 4641
rect 885 4641 987 4735
tri 987 4641 1085 4739 sw
tri 1085 4641 1183 4739 ne
rect 1183 4735 1537 4739
rect 1183 4641 1315 4735
rect 885 4615 1085 4641
rect 663 4611 1085 4615
tri 1085 4611 1115 4641 sw
tri 1183 4611 1213 4641 ne
rect 1213 4615 1315 4641
rect 1435 4641 1537 4735
tri 1537 4641 1635 4739 sw
tri 1635 4641 1733 4739 ne
rect 1733 4735 2087 4739
rect 1733 4641 1865 4735
rect 1435 4615 1635 4641
rect 1213 4611 1635 4615
tri 1635 4611 1665 4641 sw
tri 1733 4611 1763 4641 ne
rect 1763 4615 1865 4641
rect 1985 4641 2087 4735
tri 2087 4641 2185 4739 sw
tri 2185 4641 2283 4739 ne
rect 2283 4735 2637 4739
rect 2283 4641 2415 4735
rect 1985 4615 2185 4641
rect 1763 4611 2185 4615
tri 2185 4611 2215 4641 sw
tri 2283 4611 2313 4641 ne
rect 2313 4615 2415 4641
rect 2535 4641 2637 4735
tri 2637 4641 2735 4739 sw
tri 2735 4641 2833 4739 ne
rect 2833 4735 3187 4739
rect 2833 4641 2965 4735
rect 2535 4615 2735 4641
rect 2313 4611 2735 4615
tri 2735 4611 2765 4641 sw
tri 2833 4611 2863 4641 ne
rect 2863 4615 2965 4641
rect 3085 4641 3187 4735
tri 3187 4641 3285 4739 sw
tri 3285 4641 3383 4739 ne
rect 3383 4735 3737 4739
rect 3383 4641 3515 4735
rect 3085 4615 3285 4641
rect 2863 4611 3285 4615
tri 3285 4611 3315 4641 sw
tri 3383 4611 3413 4641 ne
rect 3413 4615 3515 4641
rect 3635 4641 3737 4735
tri 3737 4641 3835 4739 sw
tri 3835 4641 3933 4739 ne
rect 3933 4735 4287 4739
rect 3933 4641 4065 4735
rect 3635 4615 3835 4641
rect 3413 4611 3835 4615
tri 3835 4611 3865 4641 sw
tri 3933 4611 3963 4641 ne
rect 3963 4615 4065 4641
rect 4185 4641 4287 4735
tri 4287 4641 4385 4739 sw
tri 4385 4641 4483 4739 ne
rect 4483 4735 4837 4739
rect 4483 4641 4615 4735
rect 4185 4615 4385 4641
rect 3963 4611 4385 4615
tri 4385 4611 4415 4641 sw
tri 4483 4611 4513 4641 ne
rect 4513 4615 4615 4641
rect 4735 4641 4837 4735
tri 4837 4641 4935 4739 sw
tri 4935 4641 5033 4739 ne
rect 5033 4735 5387 4739
rect 5033 4641 5165 4735
rect 4735 4615 4935 4641
rect 4513 4611 4935 4615
tri 4935 4611 4965 4641 sw
tri 5033 4611 5063 4641 ne
rect 5063 4615 5165 4641
rect 5285 4641 5387 4735
tri 5387 4641 5485 4739 sw
tri 5485 4641 5583 4739 ne
rect 5583 4735 5937 4739
rect 5583 4641 5715 4735
rect 5285 4615 5485 4641
rect 5063 4611 5485 4615
tri 5485 4611 5515 4641 sw
tri 5583 4611 5613 4641 ne
rect 5613 4615 5715 4641
rect 5835 4641 5937 4735
tri 5937 4641 6035 4739 sw
tri 6035 4641 6133 4739 ne
rect 6133 4735 6487 4739
rect 6133 4641 6265 4735
rect 5835 4615 6035 4641
rect 5613 4611 6035 4615
tri 6035 4611 6065 4641 sw
tri 6133 4611 6163 4641 ne
rect 6163 4615 6265 4641
rect 6385 4641 6487 4735
tri 6487 4641 6585 4739 sw
tri 6585 4641 6683 4739 ne
rect 6683 4735 7037 4739
rect 6683 4641 6815 4735
rect 6385 4615 6585 4641
rect 6163 4611 6585 4615
tri 6585 4611 6615 4641 sw
tri 6683 4611 6713 4641 ne
rect 6713 4615 6815 4641
rect 6935 4641 7037 4735
tri 7037 4641 7135 4739 sw
tri 7135 4641 7233 4739 ne
rect 7233 4735 7587 4739
rect 7233 4641 7365 4735
rect 6935 4615 7135 4641
rect 6713 4611 7135 4615
tri 7135 4611 7165 4641 sw
tri 7233 4611 7263 4641 ne
rect 7263 4615 7365 4641
rect 7485 4641 7587 4735
tri 7587 4641 7685 4739 sw
tri 7685 4641 7783 4739 ne
rect 7783 4735 8137 4739
rect 7783 4641 7915 4735
rect 7485 4615 7685 4641
rect 7263 4611 7685 4615
tri 7685 4611 7715 4641 sw
tri 7783 4611 7813 4641 ne
rect 7813 4615 7915 4641
rect 8035 4641 8137 4735
tri 8137 4641 8235 4739 sw
tri 8235 4641 8333 4739 ne
rect 8333 4735 8687 4739
rect 8333 4641 8465 4735
rect 8035 4615 8235 4641
rect 7813 4611 8235 4615
tri 8235 4611 8265 4641 sw
tri 8333 4611 8363 4641 ne
rect 8363 4615 8465 4641
rect 8585 4641 8687 4735
tri 8687 4641 8785 4739 sw
tri 8785 4641 8883 4739 ne
rect 8883 4735 9237 4739
rect 8883 4641 9015 4735
rect 8585 4615 8785 4641
rect 8363 4611 8785 4615
tri 8785 4611 8815 4641 sw
tri 8883 4611 8913 4641 ne
rect 8913 4615 9015 4641
rect 9135 4641 9237 4735
tri 9237 4641 9335 4739 sw
tri 9335 4641 9433 4739 ne
rect 9433 4735 9787 4739
rect 9433 4641 9565 4735
rect 9135 4615 9335 4641
rect 8913 4611 9335 4615
tri 9335 4611 9365 4641 sw
tri 9433 4611 9463 4641 ne
rect 9463 4615 9565 4641
rect 9685 4641 9787 4735
tri 9787 4641 9885 4739 sw
tri 9885 4641 9983 4739 ne
rect 9983 4735 10337 4739
rect 9983 4641 10115 4735
rect 9685 4615 9885 4641
rect 9463 4611 9885 4615
tri 9885 4611 9915 4641 sw
tri 9983 4611 10013 4641 ne
rect 10013 4615 10115 4641
rect 10235 4641 10337 4735
tri 10337 4641 10435 4739 sw
tri 10435 4641 10533 4739 ne
rect 10533 4735 10887 4739
rect 10533 4641 10665 4735
rect 10235 4615 10435 4641
rect 10013 4611 10435 4615
tri 10435 4611 10465 4641 sw
tri 10533 4611 10563 4641 ne
rect 10563 4615 10665 4641
rect 10785 4641 10887 4735
tri 10887 4641 10985 4739 sw
tri 10985 4641 11083 4739 ne
rect 11083 4735 11437 4739
rect 11083 4641 11215 4735
rect 10785 4615 10985 4641
rect 10563 4611 10985 4615
tri 10985 4611 11015 4641 sw
tri 11083 4611 11113 4641 ne
rect 11113 4615 11215 4641
rect 11335 4641 11437 4735
tri 11437 4641 11535 4739 sw
tri 11535 4641 11633 4739 ne
rect 11633 4735 11987 4739
rect 11633 4641 11765 4735
rect 11335 4615 11535 4641
rect 11113 4611 11535 4615
tri 11535 4611 11565 4641 sw
tri 11633 4611 11663 4641 ne
rect 11663 4615 11765 4641
rect 11885 4641 11987 4735
tri 11987 4641 12085 4739 sw
tri 12085 4641 12183 4739 ne
rect 12183 4735 12537 4739
rect 12183 4641 12315 4735
rect 11885 4615 12085 4641
rect 11663 4611 12085 4615
tri 12085 4611 12115 4641 sw
tri 12183 4611 12213 4641 ne
rect 12213 4615 12315 4641
rect 12435 4641 12537 4735
tri 12537 4641 12635 4739 sw
tri 12635 4641 12733 4739 ne
rect 12733 4735 13087 4739
rect 12733 4641 12865 4735
rect 12435 4615 12635 4641
rect 12213 4611 12635 4615
tri 12635 4611 12665 4641 sw
tri 12733 4611 12763 4641 ne
rect 12763 4615 12865 4641
rect 12985 4641 13087 4735
tri 13087 4641 13185 4739 sw
tri 13185 4641 13283 4739 ne
rect 13283 4735 13637 4739
rect 13283 4641 13415 4735
rect 12985 4615 13185 4641
rect 12763 4611 13185 4615
tri 13185 4611 13215 4641 sw
tri 13283 4611 13313 4641 ne
rect 13313 4615 13415 4641
rect 13535 4641 13637 4735
tri 13637 4641 13735 4739 sw
tri 13735 4641 13833 4739 ne
rect 13833 4735 14187 4739
rect 13833 4641 13965 4735
rect 13535 4615 13735 4641
rect 13313 4611 13735 4615
tri 13735 4611 13765 4641 sw
tri 13833 4611 13863 4641 ne
rect 13863 4615 13965 4641
rect 14085 4641 14187 4735
tri 14187 4641 14285 4739 sw
tri 14285 4641 14383 4739 ne
rect 14383 4735 14737 4739
rect 14383 4641 14515 4735
rect 14085 4615 14285 4641
rect 13863 4611 14285 4615
tri 14285 4611 14315 4641 sw
tri 14383 4611 14413 4641 ne
rect 14413 4615 14515 4641
rect 14635 4641 14737 4735
tri 14737 4641 14835 4739 sw
tri 14835 4641 14933 4739 ne
rect 14933 4735 15287 4739
rect 14933 4641 15065 4735
rect 14635 4615 14835 4641
rect 14413 4611 14835 4615
tri 14835 4611 14865 4641 sw
tri 14933 4611 14963 4641 ne
rect 14963 4615 15065 4641
rect 15185 4641 15287 4735
tri 15287 4641 15385 4739 sw
tri 15385 4641 15483 4739 ne
rect 15483 4735 15837 4739
rect 15483 4641 15615 4735
rect 15185 4615 15385 4641
rect 14963 4611 15385 4615
tri 15385 4611 15415 4641 sw
tri 15483 4611 15513 4641 ne
rect 15513 4615 15615 4641
rect 15735 4641 15837 4735
tri 15837 4641 15935 4739 sw
tri 15935 4641 16033 4739 ne
rect 16033 4735 16387 4739
rect 16033 4641 16165 4735
rect 15735 4615 15935 4641
rect 15513 4611 15935 4615
tri 15935 4611 15965 4641 sw
tri 16033 4611 16063 4641 ne
rect 16063 4615 16165 4641
rect 16285 4641 16387 4735
tri 16387 4641 16485 4739 sw
tri 16485 4641 16583 4739 ne
rect 16583 4735 16937 4739
rect 16583 4641 16715 4735
rect 16285 4615 16485 4641
rect 16063 4611 16485 4615
tri 16485 4611 16515 4641 sw
tri 16583 4611 16613 4641 ne
rect 16613 4615 16715 4641
rect 16835 4641 16937 4735
tri 16937 4641 17035 4739 sw
tri 17035 4641 17133 4739 ne
rect 17133 4735 17487 4739
rect 17133 4641 17265 4735
rect 16835 4615 17035 4641
rect 16613 4611 17035 4615
tri 17035 4611 17065 4641 sw
tri 17133 4611 17163 4641 ne
rect 17163 4615 17265 4641
rect 17385 4641 17487 4735
tri 17487 4641 17585 4739 sw
tri 17585 4641 17683 4739 ne
rect 17683 4735 18037 4739
rect 17683 4641 17815 4735
rect 17385 4615 17585 4641
rect 17163 4611 17585 4615
tri 17585 4611 17615 4641 sw
tri 17683 4611 17713 4641 ne
rect 17713 4615 17815 4641
rect 17935 4641 18037 4735
tri 18037 4641 18135 4739 sw
tri 18135 4641 18233 4739 ne
rect 18233 4735 18587 4739
rect 18233 4641 18365 4735
rect 17935 4615 18135 4641
rect 17713 4611 18135 4615
tri 18135 4611 18165 4641 sw
tri 18233 4611 18263 4641 ne
rect 18263 4615 18365 4641
rect 18485 4641 18587 4735
tri 18587 4641 18685 4739 sw
tri 18685 4641 18783 4739 ne
rect 18783 4735 19137 4739
rect 18783 4641 18915 4735
rect 18485 4615 18685 4641
rect 18263 4611 18685 4615
tri 18685 4611 18715 4641 sw
tri 18783 4611 18813 4641 ne
rect 18813 4615 18915 4641
rect 19035 4641 19137 4735
tri 19137 4641 19235 4739 sw
tri 19235 4641 19333 4739 ne
rect 19333 4735 20300 4739
rect 19333 4641 19465 4735
rect 19035 4615 19235 4641
rect 18813 4611 19235 4615
tri 19235 4611 19265 4641 sw
tri 19333 4611 19363 4641 ne
rect 19363 4615 19465 4641
rect 19585 4615 20300 4735
rect 19363 4611 20300 4615
tri 113 4513 211 4611 ne
rect 211 4513 565 4611
tri 565 4513 663 4611 sw
tri 663 4513 761 4611 ne
rect 761 4513 1115 4611
tri 1115 4513 1213 4611 sw
tri 1213 4513 1311 4611 ne
rect 1311 4513 1665 4611
tri 1665 4513 1763 4611 sw
tri 1763 4513 1861 4611 ne
rect 1861 4513 2215 4611
tri 2215 4513 2313 4611 sw
tri 2313 4513 2411 4611 ne
rect 2411 4513 2765 4611
tri 2765 4513 2863 4611 sw
tri 2863 4513 2961 4611 ne
rect 2961 4513 3315 4611
tri 3315 4513 3413 4611 sw
tri 3413 4513 3511 4611 ne
rect 3511 4513 3865 4611
tri 3865 4513 3963 4611 sw
tri 3963 4513 4061 4611 ne
rect 4061 4513 4415 4611
tri 4415 4513 4513 4611 sw
tri 4513 4513 4611 4611 ne
rect 4611 4513 4965 4611
tri 4965 4513 5063 4611 sw
tri 5063 4513 5161 4611 ne
rect 5161 4513 5515 4611
tri 5515 4513 5613 4611 sw
tri 5613 4513 5711 4611 ne
rect 5711 4513 6065 4611
tri 6065 4513 6163 4611 sw
tri 6163 4513 6261 4611 ne
rect 6261 4513 6615 4611
tri 6615 4513 6713 4611 sw
tri 6713 4513 6811 4611 ne
rect 6811 4513 7165 4611
tri 7165 4513 7263 4611 sw
tri 7263 4513 7361 4611 ne
rect 7361 4513 7715 4611
tri 7715 4513 7813 4611 sw
tri 7813 4513 7911 4611 ne
rect 7911 4513 8265 4611
tri 8265 4513 8363 4611 sw
tri 8363 4513 8461 4611 ne
rect 8461 4513 8815 4611
tri 8815 4513 8913 4611 sw
tri 8913 4513 9011 4611 ne
rect 9011 4513 9365 4611
tri 9365 4513 9463 4611 sw
tri 9463 4513 9561 4611 ne
rect 9561 4513 9915 4611
tri 9915 4513 10013 4611 sw
tri 10013 4513 10111 4611 ne
rect 10111 4513 10465 4611
tri 10465 4513 10563 4611 sw
tri 10563 4513 10661 4611 ne
rect 10661 4513 11015 4611
tri 11015 4513 11113 4611 sw
tri 11113 4513 11211 4611 ne
rect 11211 4513 11565 4611
tri 11565 4513 11663 4611 sw
tri 11663 4513 11761 4611 ne
rect 11761 4513 12115 4611
tri 12115 4513 12213 4611 sw
tri 12213 4513 12311 4611 ne
rect 12311 4513 12665 4611
tri 12665 4513 12763 4611 sw
tri 12763 4513 12861 4611 ne
rect 12861 4513 13215 4611
tri 13215 4513 13313 4611 sw
tri 13313 4513 13411 4611 ne
rect 13411 4513 13765 4611
tri 13765 4513 13863 4611 sw
tri 13863 4513 13961 4611 ne
rect 13961 4513 14315 4611
tri 14315 4513 14413 4611 sw
tri 14413 4513 14511 4611 ne
rect 14511 4513 14865 4611
tri 14865 4513 14963 4611 sw
tri 14963 4513 15061 4611 ne
rect 15061 4513 15415 4611
tri 15415 4513 15513 4611 sw
tri 15513 4513 15611 4611 ne
rect 15611 4513 15965 4611
tri 15965 4513 16063 4611 sw
tri 16063 4513 16161 4611 ne
rect 16161 4513 16515 4611
tri 16515 4513 16613 4611 sw
tri 16613 4513 16711 4611 ne
rect 16711 4513 17065 4611
tri 17065 4513 17163 4611 sw
tri 17163 4513 17261 4611 ne
rect 17261 4513 17615 4611
tri 17615 4513 17713 4611 sw
tri 17713 4513 17811 4611 ne
rect 17811 4513 18165 4611
tri 18165 4513 18263 4611 sw
tri 18263 4513 18361 4611 ne
rect 18361 4513 18715 4611
tri 18715 4513 18813 4611 sw
tri 18813 4513 18911 4611 ne
rect 18911 4513 19265 4611
tri 19265 4513 19363 4611 sw
tri 19363 4513 19461 4611 ne
rect 19461 4513 20300 4611
rect -2000 4483 113 4513
tri 113 4483 143 4513 sw
tri 211 4483 241 4513 ne
rect 241 4483 663 4513
tri 663 4483 693 4513 sw
tri 761 4483 791 4513 ne
rect 791 4483 1213 4513
tri 1213 4483 1243 4513 sw
tri 1311 4483 1341 4513 ne
rect 1341 4483 1763 4513
tri 1763 4483 1793 4513 sw
tri 1861 4483 1891 4513 ne
rect 1891 4483 2313 4513
tri 2313 4483 2343 4513 sw
tri 2411 4483 2441 4513 ne
rect 2441 4483 2863 4513
tri 2863 4483 2893 4513 sw
tri 2961 4483 2991 4513 ne
rect 2991 4483 3413 4513
tri 3413 4483 3443 4513 sw
tri 3511 4483 3541 4513 ne
rect 3541 4483 3963 4513
tri 3963 4483 3993 4513 sw
tri 4061 4483 4091 4513 ne
rect 4091 4483 4513 4513
tri 4513 4483 4543 4513 sw
tri 4611 4483 4641 4513 ne
rect 4641 4483 5063 4513
tri 5063 4483 5093 4513 sw
tri 5161 4483 5191 4513 ne
rect 5191 4483 5613 4513
tri 5613 4483 5643 4513 sw
tri 5711 4483 5741 4513 ne
rect 5741 4483 6163 4513
tri 6163 4483 6193 4513 sw
tri 6261 4483 6291 4513 ne
rect 6291 4483 6713 4513
tri 6713 4483 6743 4513 sw
tri 6811 4483 6841 4513 ne
rect 6841 4483 7263 4513
tri 7263 4483 7293 4513 sw
tri 7361 4483 7391 4513 ne
rect 7391 4483 7813 4513
tri 7813 4483 7843 4513 sw
tri 7911 4483 7941 4513 ne
rect 7941 4483 8363 4513
tri 8363 4483 8393 4513 sw
tri 8461 4483 8491 4513 ne
rect 8491 4483 8913 4513
tri 8913 4483 8943 4513 sw
tri 9011 4483 9041 4513 ne
rect 9041 4483 9463 4513
tri 9463 4483 9493 4513 sw
tri 9561 4483 9591 4513 ne
rect 9591 4483 10013 4513
tri 10013 4483 10043 4513 sw
tri 10111 4483 10141 4513 ne
rect 10141 4483 10563 4513
tri 10563 4483 10593 4513 sw
tri 10661 4483 10691 4513 ne
rect 10691 4483 11113 4513
tri 11113 4483 11143 4513 sw
tri 11211 4483 11241 4513 ne
rect 11241 4483 11663 4513
tri 11663 4483 11693 4513 sw
tri 11761 4483 11791 4513 ne
rect 11791 4483 12213 4513
tri 12213 4483 12243 4513 sw
tri 12311 4483 12341 4513 ne
rect 12341 4483 12763 4513
tri 12763 4483 12793 4513 sw
tri 12861 4483 12891 4513 ne
rect 12891 4483 13313 4513
tri 13313 4483 13343 4513 sw
tri 13411 4483 13441 4513 ne
rect 13441 4483 13863 4513
tri 13863 4483 13893 4513 sw
tri 13961 4483 13991 4513 ne
rect 13991 4483 14413 4513
tri 14413 4483 14443 4513 sw
tri 14511 4483 14541 4513 ne
rect 14541 4483 14963 4513
tri 14963 4483 14993 4513 sw
tri 15061 4483 15091 4513 ne
rect 15091 4483 15513 4513
tri 15513 4483 15543 4513 sw
tri 15611 4483 15641 4513 ne
rect 15641 4483 16063 4513
tri 16063 4483 16093 4513 sw
tri 16161 4483 16191 4513 ne
rect 16191 4483 16613 4513
tri 16613 4483 16643 4513 sw
tri 16711 4483 16741 4513 ne
rect 16741 4483 17163 4513
tri 17163 4483 17193 4513 sw
tri 17261 4483 17291 4513 ne
rect 17291 4483 17713 4513
tri 17713 4483 17743 4513 sw
tri 17811 4483 17841 4513 ne
rect 17841 4483 18263 4513
tri 18263 4483 18293 4513 sw
tri 18361 4483 18391 4513 ne
rect 18391 4483 18813 4513
tri 18813 4483 18843 4513 sw
tri 18911 4483 18941 4513 ne
rect 18941 4483 19363 4513
tri 19363 4483 19393 4513 sw
tri 19461 4483 19491 4513 ne
rect 19491 4483 20300 4513
rect -2000 4385 143 4483
tri 143 4385 241 4483 sw
tri 241 4385 339 4483 ne
rect 339 4385 693 4483
tri 693 4385 791 4483 sw
tri 791 4385 889 4483 ne
rect 889 4385 1243 4483
tri 1243 4385 1341 4483 sw
tri 1341 4385 1439 4483 ne
rect 1439 4385 1793 4483
tri 1793 4385 1891 4483 sw
tri 1891 4385 1989 4483 ne
rect 1989 4385 2343 4483
tri 2343 4385 2441 4483 sw
tri 2441 4385 2539 4483 ne
rect 2539 4385 2893 4483
tri 2893 4385 2991 4483 sw
tri 2991 4385 3089 4483 ne
rect 3089 4385 3443 4483
tri 3443 4385 3541 4483 sw
tri 3541 4385 3639 4483 ne
rect 3639 4385 3993 4483
tri 3993 4385 4091 4483 sw
tri 4091 4385 4189 4483 ne
rect 4189 4385 4543 4483
tri 4543 4385 4641 4483 sw
tri 4641 4385 4739 4483 ne
rect 4739 4385 5093 4483
tri 5093 4385 5191 4483 sw
tri 5191 4385 5289 4483 ne
rect 5289 4385 5643 4483
tri 5643 4385 5741 4483 sw
tri 5741 4385 5839 4483 ne
rect 5839 4385 6193 4483
tri 6193 4385 6291 4483 sw
tri 6291 4385 6389 4483 ne
rect 6389 4385 6743 4483
tri 6743 4385 6841 4483 sw
tri 6841 4385 6939 4483 ne
rect 6939 4385 7293 4483
tri 7293 4385 7391 4483 sw
tri 7391 4385 7489 4483 ne
rect 7489 4385 7843 4483
tri 7843 4385 7941 4483 sw
tri 7941 4385 8039 4483 ne
rect 8039 4385 8393 4483
tri 8393 4385 8491 4483 sw
tri 8491 4385 8589 4483 ne
rect 8589 4385 8943 4483
tri 8943 4385 9041 4483 sw
tri 9041 4385 9139 4483 ne
rect 9139 4385 9493 4483
tri 9493 4385 9591 4483 sw
tri 9591 4385 9689 4483 ne
rect 9689 4385 10043 4483
tri 10043 4385 10141 4483 sw
tri 10141 4385 10239 4483 ne
rect 10239 4385 10593 4483
tri 10593 4385 10691 4483 sw
tri 10691 4385 10789 4483 ne
rect 10789 4385 11143 4483
tri 11143 4385 11241 4483 sw
tri 11241 4385 11339 4483 ne
rect 11339 4385 11693 4483
tri 11693 4385 11791 4483 sw
tri 11791 4385 11889 4483 ne
rect 11889 4385 12243 4483
tri 12243 4385 12341 4483 sw
tri 12341 4385 12439 4483 ne
rect 12439 4385 12793 4483
tri 12793 4385 12891 4483 sw
tri 12891 4385 12989 4483 ne
rect 12989 4385 13343 4483
tri 13343 4385 13441 4483 sw
tri 13441 4385 13539 4483 ne
rect 13539 4385 13893 4483
tri 13893 4385 13991 4483 sw
tri 13991 4385 14089 4483 ne
rect 14089 4385 14443 4483
tri 14443 4385 14541 4483 sw
tri 14541 4385 14639 4483 ne
rect 14639 4385 14993 4483
tri 14993 4385 15091 4483 sw
tri 15091 4385 15189 4483 ne
rect 15189 4385 15543 4483
tri 15543 4385 15641 4483 sw
tri 15641 4385 15739 4483 ne
rect 15739 4385 16093 4483
tri 16093 4385 16191 4483 sw
tri 16191 4385 16289 4483 ne
rect 16289 4385 16643 4483
tri 16643 4385 16741 4483 sw
tri 16741 4385 16839 4483 ne
rect 16839 4385 17193 4483
tri 17193 4385 17291 4483 sw
tri 17291 4385 17389 4483 ne
rect 17389 4385 17743 4483
tri 17743 4385 17841 4483 sw
tri 17841 4385 17939 4483 ne
rect 17939 4385 18293 4483
tri 18293 4385 18391 4483 sw
tri 18391 4385 18489 4483 ne
rect 18489 4385 18843 4483
tri 18843 4385 18941 4483 sw
tri 18941 4385 19039 4483 ne
rect 19039 4385 19393 4483
tri 19393 4385 19491 4483 sw
tri 19491 4385 19589 4483 ne
rect 19589 4385 20300 4483
rect -2000 4287 241 4385
tri 241 4287 339 4385 sw
tri 339 4287 437 4385 ne
rect 437 4287 791 4385
tri 791 4287 889 4385 sw
tri 889 4287 987 4385 ne
rect 987 4287 1341 4385
tri 1341 4287 1439 4385 sw
tri 1439 4287 1537 4385 ne
rect 1537 4287 1891 4385
tri 1891 4287 1989 4385 sw
tri 1989 4287 2087 4385 ne
rect 2087 4287 2441 4385
tri 2441 4287 2539 4385 sw
tri 2539 4287 2637 4385 ne
rect 2637 4287 2991 4385
tri 2991 4287 3089 4385 sw
tri 3089 4287 3187 4385 ne
rect 3187 4287 3541 4385
tri 3541 4287 3639 4385 sw
tri 3639 4287 3737 4385 ne
rect 3737 4287 4091 4385
tri 4091 4287 4189 4385 sw
tri 4189 4287 4287 4385 ne
rect 4287 4287 4641 4385
tri 4641 4287 4739 4385 sw
tri 4739 4287 4837 4385 ne
rect 4837 4287 5191 4385
tri 5191 4287 5289 4385 sw
tri 5289 4287 5387 4385 ne
rect 5387 4287 5741 4385
tri 5741 4287 5839 4385 sw
tri 5839 4287 5937 4385 ne
rect 5937 4287 6291 4385
tri 6291 4287 6389 4385 sw
tri 6389 4287 6487 4385 ne
rect 6487 4287 6841 4385
tri 6841 4287 6939 4385 sw
tri 6939 4287 7037 4385 ne
rect 7037 4287 7391 4385
tri 7391 4287 7489 4385 sw
tri 7489 4287 7587 4385 ne
rect 7587 4287 7941 4385
tri 7941 4287 8039 4385 sw
tri 8039 4287 8137 4385 ne
rect 8137 4287 8491 4385
tri 8491 4287 8589 4385 sw
tri 8589 4287 8687 4385 ne
rect 8687 4287 9041 4385
tri 9041 4287 9139 4385 sw
tri 9139 4287 9237 4385 ne
rect 9237 4287 9591 4385
tri 9591 4287 9689 4385 sw
tri 9689 4287 9787 4385 ne
rect 9787 4287 10141 4385
tri 10141 4287 10239 4385 sw
tri 10239 4287 10337 4385 ne
rect 10337 4287 10691 4385
tri 10691 4287 10789 4385 sw
tri 10789 4287 10887 4385 ne
rect 10887 4287 11241 4385
tri 11241 4287 11339 4385 sw
tri 11339 4287 11437 4385 ne
rect 11437 4287 11791 4385
tri 11791 4287 11889 4385 sw
tri 11889 4287 11987 4385 ne
rect 11987 4287 12341 4385
tri 12341 4287 12439 4385 sw
tri 12439 4287 12537 4385 ne
rect 12537 4287 12891 4385
tri 12891 4287 12989 4385 sw
tri 12989 4287 13087 4385 ne
rect 13087 4287 13441 4385
tri 13441 4287 13539 4385 sw
tri 13539 4287 13637 4385 ne
rect 13637 4287 13991 4385
tri 13991 4287 14089 4385 sw
tri 14089 4287 14187 4385 ne
rect 14187 4287 14541 4385
tri 14541 4287 14639 4385 sw
tri 14639 4287 14737 4385 ne
rect 14737 4287 15091 4385
tri 15091 4287 15189 4385 sw
tri 15189 4287 15287 4385 ne
rect 15287 4287 15641 4385
tri 15641 4287 15739 4385 sw
tri 15739 4287 15837 4385 ne
rect 15837 4287 16191 4385
tri 16191 4287 16289 4385 sw
tri 16289 4287 16387 4385 ne
rect 16387 4287 16741 4385
tri 16741 4287 16839 4385 sw
tri 16839 4287 16937 4385 ne
rect 16937 4287 17291 4385
tri 17291 4287 17389 4385 sw
tri 17389 4287 17487 4385 ne
rect 17487 4287 17841 4385
tri 17841 4287 17939 4385 sw
tri 17939 4287 18037 4385 ne
rect 18037 4287 18391 4385
tri 18391 4287 18489 4385 sw
tri 18489 4287 18587 4385 ne
rect 18587 4287 18941 4385
tri 18941 4287 19039 4385 sw
tri 19039 4287 19137 4385 ne
rect 19137 4287 19491 4385
tri 19491 4287 19589 4385 sw
tri 19589 4287 19687 4385 ne
rect 19687 4287 20300 4385
rect -2000 4189 339 4287
tri 339 4189 437 4287 sw
tri 437 4189 535 4287 ne
rect 535 4189 889 4287
tri 889 4189 987 4287 sw
tri 987 4189 1085 4287 ne
rect 1085 4189 1439 4287
tri 1439 4189 1537 4287 sw
tri 1537 4189 1635 4287 ne
rect 1635 4189 1989 4287
tri 1989 4189 2087 4287 sw
tri 2087 4189 2185 4287 ne
rect 2185 4189 2539 4287
tri 2539 4189 2637 4287 sw
tri 2637 4189 2735 4287 ne
rect 2735 4189 3089 4287
tri 3089 4189 3187 4287 sw
tri 3187 4189 3285 4287 ne
rect 3285 4189 3639 4287
tri 3639 4189 3737 4287 sw
tri 3737 4189 3835 4287 ne
rect 3835 4189 4189 4287
tri 4189 4189 4287 4287 sw
tri 4287 4189 4385 4287 ne
rect 4385 4189 4739 4287
tri 4739 4189 4837 4287 sw
tri 4837 4189 4935 4287 ne
rect 4935 4189 5289 4287
tri 5289 4189 5387 4287 sw
tri 5387 4189 5485 4287 ne
rect 5485 4189 5839 4287
tri 5839 4189 5937 4287 sw
tri 5937 4189 6035 4287 ne
rect 6035 4189 6389 4287
tri 6389 4189 6487 4287 sw
tri 6487 4189 6585 4287 ne
rect 6585 4189 6939 4287
tri 6939 4189 7037 4287 sw
tri 7037 4189 7135 4287 ne
rect 7135 4189 7489 4287
tri 7489 4189 7587 4287 sw
tri 7587 4189 7685 4287 ne
rect 7685 4189 8039 4287
tri 8039 4189 8137 4287 sw
tri 8137 4189 8235 4287 ne
rect 8235 4189 8589 4287
tri 8589 4189 8687 4287 sw
tri 8687 4189 8785 4287 ne
rect 8785 4189 9139 4287
tri 9139 4189 9237 4287 sw
tri 9237 4189 9335 4287 ne
rect 9335 4189 9689 4287
tri 9689 4189 9787 4287 sw
tri 9787 4189 9885 4287 ne
rect 9885 4189 10239 4287
tri 10239 4189 10337 4287 sw
tri 10337 4189 10435 4287 ne
rect 10435 4189 10789 4287
tri 10789 4189 10887 4287 sw
tri 10887 4189 10985 4287 ne
rect 10985 4189 11339 4287
tri 11339 4189 11437 4287 sw
tri 11437 4189 11535 4287 ne
rect 11535 4189 11889 4287
tri 11889 4189 11987 4287 sw
tri 11987 4189 12085 4287 ne
rect 12085 4189 12439 4287
tri 12439 4189 12537 4287 sw
tri 12537 4189 12635 4287 ne
rect 12635 4189 12989 4287
tri 12989 4189 13087 4287 sw
tri 13087 4189 13185 4287 ne
rect 13185 4189 13539 4287
tri 13539 4189 13637 4287 sw
tri 13637 4189 13735 4287 ne
rect 13735 4189 14089 4287
tri 14089 4189 14187 4287 sw
tri 14187 4189 14285 4287 ne
rect 14285 4189 14639 4287
tri 14639 4189 14737 4287 sw
tri 14737 4189 14835 4287 ne
rect 14835 4189 15189 4287
tri 15189 4189 15287 4287 sw
tri 15287 4189 15385 4287 ne
rect 15385 4189 15739 4287
tri 15739 4189 15837 4287 sw
tri 15837 4189 15935 4287 ne
rect 15935 4189 16289 4287
tri 16289 4189 16387 4287 sw
tri 16387 4189 16485 4287 ne
rect 16485 4189 16839 4287
tri 16839 4189 16937 4287 sw
tri 16937 4189 17035 4287 ne
rect 17035 4189 17389 4287
tri 17389 4189 17487 4287 sw
tri 17487 4189 17585 4287 ne
rect 17585 4189 17939 4287
tri 17939 4189 18037 4287 sw
tri 18037 4189 18135 4287 ne
rect 18135 4189 18489 4287
tri 18489 4189 18587 4287 sw
tri 18587 4189 18685 4287 ne
rect 18685 4189 19039 4287
tri 19039 4189 19137 4287 sw
tri 19137 4189 19235 4287 ne
rect 19235 4189 19589 4287
tri 19589 4189 19687 4287 sw
rect 20800 4189 21800 4837
rect -2000 4185 437 4189
rect -2000 4065 215 4185
rect 335 4091 437 4185
tri 437 4091 535 4189 sw
tri 535 4091 633 4189 ne
rect 633 4185 987 4189
rect 633 4091 765 4185
rect 335 4065 535 4091
rect -2000 4061 535 4065
rect -2000 3413 -1000 4061
tri 113 3963 211 4061 ne
rect 211 4013 535 4061
tri 535 4013 613 4091 sw
tri 633 4013 711 4091 ne
rect 711 4065 765 4091
rect 885 4091 987 4185
tri 987 4091 1085 4189 sw
tri 1085 4091 1183 4189 ne
rect 1183 4185 1537 4189
rect 1183 4091 1315 4185
rect 885 4065 1085 4091
rect 711 4013 1085 4065
tri 1085 4013 1163 4091 sw
tri 1183 4013 1261 4091 ne
rect 1261 4065 1315 4091
rect 1435 4091 1537 4185
tri 1537 4091 1635 4189 sw
tri 1635 4091 1733 4189 ne
rect 1733 4185 2087 4189
rect 1733 4091 1865 4185
rect 1435 4065 1635 4091
rect 1261 4013 1635 4065
tri 1635 4013 1713 4091 sw
tri 1733 4013 1811 4091 ne
rect 1811 4065 1865 4091
rect 1985 4091 2087 4185
tri 2087 4091 2185 4189 sw
tri 2185 4091 2283 4189 ne
rect 2283 4185 2637 4189
rect 2283 4091 2415 4185
rect 1985 4065 2185 4091
rect 1811 4013 2185 4065
tri 2185 4013 2263 4091 sw
tri 2283 4013 2361 4091 ne
rect 2361 4065 2415 4091
rect 2535 4091 2637 4185
tri 2637 4091 2735 4189 sw
tri 2735 4091 2833 4189 ne
rect 2833 4185 3187 4189
rect 2833 4091 2965 4185
rect 2535 4065 2735 4091
rect 2361 4013 2735 4065
tri 2735 4013 2813 4091 sw
tri 2833 4013 2911 4091 ne
rect 2911 4065 2965 4091
rect 3085 4091 3187 4185
tri 3187 4091 3285 4189 sw
tri 3285 4091 3383 4189 ne
rect 3383 4185 3737 4189
rect 3383 4091 3515 4185
rect 3085 4065 3285 4091
rect 2911 4013 3285 4065
tri 3285 4013 3363 4091 sw
tri 3383 4013 3461 4091 ne
rect 3461 4065 3515 4091
rect 3635 4091 3737 4185
tri 3737 4091 3835 4189 sw
tri 3835 4091 3933 4189 ne
rect 3933 4185 4287 4189
rect 3933 4091 4065 4185
rect 3635 4065 3835 4091
rect 3461 4013 3835 4065
tri 3835 4013 3913 4091 sw
tri 3933 4013 4011 4091 ne
rect 4011 4065 4065 4091
rect 4185 4091 4287 4185
tri 4287 4091 4385 4189 sw
tri 4385 4091 4483 4189 ne
rect 4483 4185 4837 4189
rect 4483 4091 4615 4185
rect 4185 4065 4385 4091
rect 4011 4013 4385 4065
tri 4385 4013 4463 4091 sw
tri 4483 4013 4561 4091 ne
rect 4561 4065 4615 4091
rect 4735 4091 4837 4185
tri 4837 4091 4935 4189 sw
tri 4935 4091 5033 4189 ne
rect 5033 4185 5387 4189
rect 5033 4091 5165 4185
rect 4735 4065 4935 4091
rect 4561 4013 4935 4065
tri 4935 4013 5013 4091 sw
tri 5033 4013 5111 4091 ne
rect 5111 4065 5165 4091
rect 5285 4091 5387 4185
tri 5387 4091 5485 4189 sw
tri 5485 4091 5583 4189 ne
rect 5583 4185 5937 4189
rect 5583 4091 5715 4185
rect 5285 4065 5485 4091
rect 5111 4013 5485 4065
tri 5485 4013 5563 4091 sw
tri 5583 4013 5661 4091 ne
rect 5661 4065 5715 4091
rect 5835 4091 5937 4185
tri 5937 4091 6035 4189 sw
tri 6035 4091 6133 4189 ne
rect 6133 4185 6487 4189
rect 6133 4091 6265 4185
rect 5835 4065 6035 4091
rect 5661 4013 6035 4065
tri 6035 4013 6113 4091 sw
tri 6133 4013 6211 4091 ne
rect 6211 4065 6265 4091
rect 6385 4091 6487 4185
tri 6487 4091 6585 4189 sw
tri 6585 4091 6683 4189 ne
rect 6683 4185 7037 4189
rect 6683 4091 6815 4185
rect 6385 4065 6585 4091
rect 6211 4013 6585 4065
tri 6585 4013 6663 4091 sw
tri 6683 4013 6761 4091 ne
rect 6761 4065 6815 4091
rect 6935 4091 7037 4185
tri 7037 4091 7135 4189 sw
tri 7135 4091 7233 4189 ne
rect 7233 4185 7587 4189
rect 7233 4091 7365 4185
rect 6935 4065 7135 4091
rect 6761 4013 7135 4065
tri 7135 4013 7213 4091 sw
tri 7233 4013 7311 4091 ne
rect 7311 4065 7365 4091
rect 7485 4091 7587 4185
tri 7587 4091 7685 4189 sw
tri 7685 4091 7783 4189 ne
rect 7783 4185 8137 4189
rect 7783 4091 7915 4185
rect 7485 4065 7685 4091
rect 7311 4013 7685 4065
tri 7685 4013 7763 4091 sw
tri 7783 4013 7861 4091 ne
rect 7861 4065 7915 4091
rect 8035 4091 8137 4185
tri 8137 4091 8235 4189 sw
tri 8235 4091 8333 4189 ne
rect 8333 4185 8687 4189
rect 8333 4091 8465 4185
rect 8035 4065 8235 4091
rect 7861 4013 8235 4065
tri 8235 4013 8313 4091 sw
tri 8333 4013 8411 4091 ne
rect 8411 4065 8465 4091
rect 8585 4091 8687 4185
tri 8687 4091 8785 4189 sw
tri 8785 4091 8883 4189 ne
rect 8883 4185 9237 4189
rect 8883 4091 9015 4185
rect 8585 4065 8785 4091
rect 8411 4013 8785 4065
tri 8785 4013 8863 4091 sw
tri 8883 4013 8961 4091 ne
rect 8961 4065 9015 4091
rect 9135 4091 9237 4185
tri 9237 4091 9335 4189 sw
tri 9335 4091 9433 4189 ne
rect 9433 4185 9787 4189
rect 9433 4091 9565 4185
rect 9135 4065 9335 4091
rect 8961 4013 9335 4065
tri 9335 4013 9413 4091 sw
tri 9433 4013 9511 4091 ne
rect 9511 4065 9565 4091
rect 9685 4091 9787 4185
tri 9787 4091 9885 4189 sw
tri 9885 4091 9983 4189 ne
rect 9983 4185 10337 4189
rect 9983 4091 10115 4185
rect 9685 4065 9885 4091
rect 9511 4013 9885 4065
tri 9885 4013 9963 4091 sw
tri 9983 4013 10061 4091 ne
rect 10061 4065 10115 4091
rect 10235 4091 10337 4185
tri 10337 4091 10435 4189 sw
tri 10435 4091 10533 4189 ne
rect 10533 4185 10887 4189
rect 10533 4091 10665 4185
rect 10235 4065 10435 4091
rect 10061 4013 10435 4065
tri 10435 4013 10513 4091 sw
tri 10533 4013 10611 4091 ne
rect 10611 4065 10665 4091
rect 10785 4091 10887 4185
tri 10887 4091 10985 4189 sw
tri 10985 4091 11083 4189 ne
rect 11083 4185 11437 4189
rect 11083 4091 11215 4185
rect 10785 4065 10985 4091
rect 10611 4013 10985 4065
tri 10985 4013 11063 4091 sw
tri 11083 4013 11161 4091 ne
rect 11161 4065 11215 4091
rect 11335 4091 11437 4185
tri 11437 4091 11535 4189 sw
tri 11535 4091 11633 4189 ne
rect 11633 4185 11987 4189
rect 11633 4091 11765 4185
rect 11335 4065 11535 4091
rect 11161 4013 11535 4065
tri 11535 4013 11613 4091 sw
tri 11633 4013 11711 4091 ne
rect 11711 4065 11765 4091
rect 11885 4091 11987 4185
tri 11987 4091 12085 4189 sw
tri 12085 4091 12183 4189 ne
rect 12183 4185 12537 4189
rect 12183 4091 12315 4185
rect 11885 4065 12085 4091
rect 11711 4013 12085 4065
tri 12085 4013 12163 4091 sw
tri 12183 4013 12261 4091 ne
rect 12261 4065 12315 4091
rect 12435 4091 12537 4185
tri 12537 4091 12635 4189 sw
tri 12635 4091 12733 4189 ne
rect 12733 4185 13087 4189
rect 12733 4091 12865 4185
rect 12435 4065 12635 4091
rect 12261 4013 12635 4065
tri 12635 4013 12713 4091 sw
tri 12733 4013 12811 4091 ne
rect 12811 4065 12865 4091
rect 12985 4091 13087 4185
tri 13087 4091 13185 4189 sw
tri 13185 4091 13283 4189 ne
rect 13283 4185 13637 4189
rect 13283 4091 13415 4185
rect 12985 4065 13185 4091
rect 12811 4013 13185 4065
tri 13185 4013 13263 4091 sw
tri 13283 4013 13361 4091 ne
rect 13361 4065 13415 4091
rect 13535 4091 13637 4185
tri 13637 4091 13735 4189 sw
tri 13735 4091 13833 4189 ne
rect 13833 4185 14187 4189
rect 13833 4091 13965 4185
rect 13535 4065 13735 4091
rect 13361 4013 13735 4065
tri 13735 4013 13813 4091 sw
tri 13833 4013 13911 4091 ne
rect 13911 4065 13965 4091
rect 14085 4091 14187 4185
tri 14187 4091 14285 4189 sw
tri 14285 4091 14383 4189 ne
rect 14383 4185 14737 4189
rect 14383 4091 14515 4185
rect 14085 4065 14285 4091
rect 13911 4013 14285 4065
tri 14285 4013 14363 4091 sw
tri 14383 4013 14461 4091 ne
rect 14461 4065 14515 4091
rect 14635 4091 14737 4185
tri 14737 4091 14835 4189 sw
tri 14835 4091 14933 4189 ne
rect 14933 4185 15287 4189
rect 14933 4091 15065 4185
rect 14635 4065 14835 4091
rect 14461 4013 14835 4065
tri 14835 4013 14913 4091 sw
tri 14933 4013 15011 4091 ne
rect 15011 4065 15065 4091
rect 15185 4091 15287 4185
tri 15287 4091 15385 4189 sw
tri 15385 4091 15483 4189 ne
rect 15483 4185 15837 4189
rect 15483 4091 15615 4185
rect 15185 4065 15385 4091
rect 15011 4013 15385 4065
tri 15385 4013 15463 4091 sw
tri 15483 4013 15561 4091 ne
rect 15561 4065 15615 4091
rect 15735 4091 15837 4185
tri 15837 4091 15935 4189 sw
tri 15935 4091 16033 4189 ne
rect 16033 4185 16387 4189
rect 16033 4091 16165 4185
rect 15735 4065 15935 4091
rect 15561 4013 15935 4065
tri 15935 4013 16013 4091 sw
tri 16033 4013 16111 4091 ne
rect 16111 4065 16165 4091
rect 16285 4091 16387 4185
tri 16387 4091 16485 4189 sw
tri 16485 4091 16583 4189 ne
rect 16583 4185 16937 4189
rect 16583 4091 16715 4185
rect 16285 4065 16485 4091
rect 16111 4013 16485 4065
tri 16485 4013 16563 4091 sw
tri 16583 4013 16661 4091 ne
rect 16661 4065 16715 4091
rect 16835 4091 16937 4185
tri 16937 4091 17035 4189 sw
tri 17035 4091 17133 4189 ne
rect 17133 4185 17487 4189
rect 17133 4091 17265 4185
rect 16835 4065 17035 4091
rect 16661 4013 17035 4065
tri 17035 4013 17113 4091 sw
tri 17133 4013 17211 4091 ne
rect 17211 4065 17265 4091
rect 17385 4091 17487 4185
tri 17487 4091 17585 4189 sw
tri 17585 4091 17683 4189 ne
rect 17683 4185 18037 4189
rect 17683 4091 17815 4185
rect 17385 4065 17585 4091
rect 17211 4013 17585 4065
tri 17585 4013 17663 4091 sw
tri 17683 4013 17761 4091 ne
rect 17761 4065 17815 4091
rect 17935 4091 18037 4185
tri 18037 4091 18135 4189 sw
tri 18135 4091 18233 4189 ne
rect 18233 4185 18587 4189
rect 18233 4091 18365 4185
rect 17935 4065 18135 4091
rect 17761 4013 18135 4065
tri 18135 4013 18213 4091 sw
tri 18233 4013 18311 4091 ne
rect 18311 4065 18365 4091
rect 18485 4091 18587 4185
tri 18587 4091 18685 4189 sw
tri 18685 4091 18783 4189 ne
rect 18783 4185 19137 4189
rect 18783 4091 18915 4185
rect 18485 4065 18685 4091
rect 18311 4013 18685 4065
tri 18685 4013 18763 4091 sw
tri 18783 4013 18861 4091 ne
rect 18861 4065 18915 4091
rect 19035 4091 19137 4185
tri 19137 4091 19235 4189 sw
tri 19235 4091 19333 4189 ne
rect 19333 4185 21800 4189
rect 19333 4091 19465 4185
rect 19035 4065 19235 4091
rect 18861 4013 19235 4065
tri 19235 4013 19313 4091 sw
tri 19333 4013 19411 4091 ne
rect 19411 4065 19465 4091
rect 19585 4065 21800 4185
rect 19411 4013 21800 4065
rect 211 3963 613 4013
rect -500 3913 113 3963
tri 113 3913 163 3963 sw
tri 211 3913 261 3963 ne
rect 261 3933 613 3963
tri 613 3933 693 4013 sw
tri 711 3933 791 4013 ne
rect 791 3933 1163 4013
tri 1163 3933 1243 4013 sw
tri 1261 3933 1341 4013 ne
rect 1341 3933 1713 4013
tri 1713 3933 1793 4013 sw
tri 1811 3933 1891 4013 ne
rect 1891 3933 2263 4013
tri 2263 3933 2343 4013 sw
tri 2361 3933 2441 4013 ne
rect 2441 3933 2813 4013
tri 2813 3933 2893 4013 sw
tri 2911 3933 2991 4013 ne
rect 2991 3933 3363 4013
tri 3363 3933 3443 4013 sw
tri 3461 3933 3541 4013 ne
rect 3541 3933 3913 4013
tri 3913 3933 3993 4013 sw
tri 4011 3933 4091 4013 ne
rect 4091 3933 4463 4013
tri 4463 3933 4543 4013 sw
tri 4561 3933 4641 4013 ne
rect 4641 3933 5013 4013
tri 5013 3933 5093 4013 sw
tri 5111 3933 5191 4013 ne
rect 5191 3933 5563 4013
tri 5563 3933 5643 4013 sw
tri 5661 3933 5741 4013 ne
rect 5741 3933 6113 4013
tri 6113 3933 6193 4013 sw
tri 6211 3933 6291 4013 ne
rect 6291 3933 6663 4013
tri 6663 3933 6743 4013 sw
tri 6761 3933 6841 4013 ne
rect 6841 3933 7213 4013
tri 7213 3933 7293 4013 sw
tri 7311 3933 7391 4013 ne
rect 7391 3933 7763 4013
tri 7763 3933 7843 4013 sw
tri 7861 3933 7941 4013 ne
rect 7941 3933 8313 4013
tri 8313 3933 8393 4013 sw
tri 8411 3933 8491 4013 ne
rect 8491 3933 8863 4013
tri 8863 3933 8943 4013 sw
tri 8961 3933 9041 4013 ne
rect 9041 3933 9413 4013
tri 9413 3933 9493 4013 sw
tri 9511 3933 9591 4013 ne
rect 9591 3933 9963 4013
tri 9963 3933 10043 4013 sw
tri 10061 3933 10141 4013 ne
rect 10141 3933 10513 4013
tri 10513 3933 10593 4013 sw
tri 10611 3933 10691 4013 ne
rect 10691 3933 11063 4013
tri 11063 3933 11143 4013 sw
tri 11161 3933 11241 4013 ne
rect 11241 3933 11613 4013
tri 11613 3933 11693 4013 sw
tri 11711 3933 11791 4013 ne
rect 11791 3933 12163 4013
tri 12163 3933 12243 4013 sw
tri 12261 3933 12341 4013 ne
rect 12341 3933 12713 4013
tri 12713 3933 12793 4013 sw
tri 12811 3933 12891 4013 ne
rect 12891 3933 13263 4013
tri 13263 3933 13343 4013 sw
tri 13361 3933 13441 4013 ne
rect 13441 3933 13813 4013
tri 13813 3933 13893 4013 sw
tri 13911 3933 13991 4013 ne
rect 13991 3933 14363 4013
tri 14363 3933 14443 4013 sw
tri 14461 3933 14541 4013 ne
rect 14541 3933 14913 4013
tri 14913 3933 14993 4013 sw
tri 15011 3933 15091 4013 ne
rect 15091 3933 15463 4013
tri 15463 3933 15543 4013 sw
tri 15561 3933 15641 4013 ne
rect 15641 3933 16013 4013
tri 16013 3933 16093 4013 sw
tri 16111 3933 16191 4013 ne
rect 16191 3933 16563 4013
tri 16563 3933 16643 4013 sw
tri 16661 3933 16741 4013 ne
rect 16741 3933 17113 4013
tri 17113 3933 17193 4013 sw
tri 17211 3933 17291 4013 ne
rect 17291 3933 17663 4013
tri 17663 3933 17743 4013 sw
tri 17761 3933 17841 4013 ne
rect 17841 3933 18213 4013
tri 18213 3933 18293 4013 sw
tri 18311 3933 18391 4013 ne
rect 18391 3933 18763 4013
tri 18763 3933 18843 4013 sw
tri 18861 3933 18941 4013 ne
rect 18941 3933 19313 4013
tri 19313 3933 19393 4013 sw
tri 19411 3933 19491 4013 ne
rect 19491 3933 20100 4013
rect 261 3913 693 3933
rect -500 3835 163 3913
tri 163 3835 241 3913 sw
tri 261 3835 339 3913 ne
rect 339 3835 693 3913
tri 693 3835 791 3933 sw
tri 791 3835 889 3933 ne
rect 889 3835 1243 3933
tri 1243 3835 1341 3933 sw
tri 1341 3835 1439 3933 ne
rect 1439 3835 1793 3933
tri 1793 3835 1891 3933 sw
tri 1891 3835 1989 3933 ne
rect 1989 3835 2343 3933
tri 2343 3835 2441 3933 sw
tri 2441 3835 2539 3933 ne
rect 2539 3835 2893 3933
tri 2893 3835 2991 3933 sw
tri 2991 3835 3089 3933 ne
rect 3089 3835 3443 3933
tri 3443 3835 3541 3933 sw
tri 3541 3835 3639 3933 ne
rect 3639 3835 3993 3933
tri 3993 3835 4091 3933 sw
tri 4091 3835 4189 3933 ne
rect 4189 3835 4543 3933
tri 4543 3835 4641 3933 sw
tri 4641 3835 4739 3933 ne
rect 4739 3835 5093 3933
tri 5093 3835 5191 3933 sw
tri 5191 3835 5289 3933 ne
rect 5289 3835 5643 3933
tri 5643 3835 5741 3933 sw
tri 5741 3835 5839 3933 ne
rect 5839 3835 6193 3933
tri 6193 3835 6291 3933 sw
tri 6291 3835 6389 3933 ne
rect 6389 3835 6743 3933
tri 6743 3835 6841 3933 sw
tri 6841 3835 6939 3933 ne
rect 6939 3835 7293 3933
tri 7293 3835 7391 3933 sw
tri 7391 3835 7489 3933 ne
rect 7489 3835 7843 3933
tri 7843 3835 7941 3933 sw
tri 7941 3835 8039 3933 ne
rect 8039 3835 8393 3933
tri 8393 3835 8491 3933 sw
tri 8491 3835 8589 3933 ne
rect 8589 3835 8943 3933
tri 8943 3835 9041 3933 sw
tri 9041 3835 9139 3933 ne
rect 9139 3835 9493 3933
tri 9493 3835 9591 3933 sw
tri 9591 3835 9689 3933 ne
rect 9689 3835 10043 3933
tri 10043 3835 10141 3933 sw
tri 10141 3835 10239 3933 ne
rect 10239 3835 10593 3933
tri 10593 3835 10691 3933 sw
tri 10691 3835 10789 3933 ne
rect 10789 3835 11143 3933
tri 11143 3835 11241 3933 sw
tri 11241 3835 11339 3933 ne
rect 11339 3835 11693 3933
tri 11693 3835 11791 3933 sw
tri 11791 3835 11889 3933 ne
rect 11889 3835 12243 3933
tri 12243 3835 12341 3933 sw
tri 12341 3835 12439 3933 ne
rect 12439 3835 12793 3933
tri 12793 3835 12891 3933 sw
tri 12891 3835 12989 3933 ne
rect 12989 3835 13343 3933
tri 13343 3835 13441 3933 sw
tri 13441 3835 13539 3933 ne
rect 13539 3835 13893 3933
tri 13893 3835 13991 3933 sw
tri 13991 3835 14089 3933 ne
rect 14089 3835 14443 3933
tri 14443 3835 14541 3933 sw
tri 14541 3835 14639 3933 ne
rect 14639 3835 14993 3933
tri 14993 3835 15091 3933 sw
tri 15091 3835 15189 3933 ne
rect 15189 3835 15543 3933
tri 15543 3835 15641 3933 sw
tri 15641 3835 15739 3933 ne
rect 15739 3835 16093 3933
tri 16093 3835 16191 3933 sw
tri 16191 3835 16289 3933 ne
rect 16289 3835 16643 3933
tri 16643 3835 16741 3933 sw
tri 16741 3835 16839 3933 ne
rect 16839 3835 17193 3933
tri 17193 3835 17291 3933 sw
tri 17291 3835 17389 3933 ne
rect 17389 3835 17743 3933
tri 17743 3835 17841 3933 sw
tri 17841 3835 17939 3933 ne
rect 17939 3835 18293 3933
tri 18293 3835 18391 3933 sw
tri 18391 3835 18489 3933 ne
rect 18489 3835 18843 3933
tri 18843 3835 18941 3933 sw
tri 18941 3835 19039 3933 ne
rect 19039 3835 19393 3933
tri 19393 3835 19491 3933 sw
tri 19491 3835 19589 3933 ne
rect 19589 3913 20100 3933
rect 20200 3913 21800 4013
rect 19589 3835 21800 3913
rect -500 3787 241 3835
rect -500 3687 -400 3787
rect -300 3737 241 3787
tri 241 3737 339 3835 sw
tri 339 3737 437 3835 ne
rect 437 3737 791 3835
tri 791 3737 889 3835 sw
tri 889 3737 987 3835 ne
rect 987 3737 1341 3835
tri 1341 3737 1439 3835 sw
tri 1439 3737 1537 3835 ne
rect 1537 3737 1891 3835
tri 1891 3737 1989 3835 sw
tri 1989 3737 2087 3835 ne
rect 2087 3737 2441 3835
tri 2441 3737 2539 3835 sw
tri 2539 3737 2637 3835 ne
rect 2637 3737 2991 3835
tri 2991 3737 3089 3835 sw
tri 3089 3737 3187 3835 ne
rect 3187 3737 3541 3835
tri 3541 3737 3639 3835 sw
tri 3639 3737 3737 3835 ne
rect 3737 3737 4091 3835
tri 4091 3737 4189 3835 sw
tri 4189 3737 4287 3835 ne
rect 4287 3737 4641 3835
tri 4641 3737 4739 3835 sw
tri 4739 3737 4837 3835 ne
rect 4837 3737 5191 3835
tri 5191 3737 5289 3835 sw
tri 5289 3737 5387 3835 ne
rect 5387 3737 5741 3835
tri 5741 3737 5839 3835 sw
tri 5839 3737 5937 3835 ne
rect 5937 3737 6291 3835
tri 6291 3737 6389 3835 sw
tri 6389 3737 6487 3835 ne
rect 6487 3737 6841 3835
tri 6841 3737 6939 3835 sw
tri 6939 3737 7037 3835 ne
rect 7037 3737 7391 3835
tri 7391 3737 7489 3835 sw
tri 7489 3737 7587 3835 ne
rect 7587 3737 7941 3835
tri 7941 3737 8039 3835 sw
tri 8039 3737 8137 3835 ne
rect 8137 3737 8491 3835
tri 8491 3737 8589 3835 sw
tri 8589 3737 8687 3835 ne
rect 8687 3737 9041 3835
tri 9041 3737 9139 3835 sw
tri 9139 3737 9237 3835 ne
rect 9237 3737 9591 3835
tri 9591 3737 9689 3835 sw
tri 9689 3737 9787 3835 ne
rect 9787 3737 10141 3835
tri 10141 3737 10239 3835 sw
tri 10239 3737 10337 3835 ne
rect 10337 3737 10691 3835
tri 10691 3737 10789 3835 sw
tri 10789 3737 10887 3835 ne
rect 10887 3737 11241 3835
tri 11241 3737 11339 3835 sw
tri 11339 3737 11437 3835 ne
rect 11437 3737 11791 3835
tri 11791 3737 11889 3835 sw
tri 11889 3737 11987 3835 ne
rect 11987 3737 12341 3835
tri 12341 3737 12439 3835 sw
tri 12439 3737 12537 3835 ne
rect 12537 3737 12891 3835
tri 12891 3737 12989 3835 sw
tri 12989 3737 13087 3835 ne
rect 13087 3737 13441 3835
tri 13441 3737 13539 3835 sw
tri 13539 3737 13637 3835 ne
rect 13637 3737 13991 3835
tri 13991 3737 14089 3835 sw
tri 14089 3737 14187 3835 ne
rect 14187 3737 14541 3835
tri 14541 3737 14639 3835 sw
tri 14639 3737 14737 3835 ne
rect 14737 3737 15091 3835
tri 15091 3737 15189 3835 sw
tri 15189 3737 15287 3835 ne
rect 15287 3737 15641 3835
tri 15641 3737 15739 3835 sw
tri 15739 3737 15837 3835 ne
rect 15837 3737 16191 3835
tri 16191 3737 16289 3835 sw
tri 16289 3737 16387 3835 ne
rect 16387 3737 16741 3835
tri 16741 3737 16839 3835 sw
tri 16839 3737 16937 3835 ne
rect 16937 3737 17291 3835
tri 17291 3737 17389 3835 sw
tri 17389 3737 17487 3835 ne
rect 17487 3737 17841 3835
tri 17841 3737 17939 3835 sw
tri 17939 3737 18037 3835 ne
rect 18037 3737 18391 3835
tri 18391 3737 18489 3835 sw
tri 18489 3737 18587 3835 ne
rect 18587 3737 18941 3835
tri 18941 3737 19039 3835 sw
tri 19039 3737 19137 3835 ne
rect 19137 3737 19491 3835
tri 19491 3737 19589 3835 sw
tri 19589 3737 19687 3835 ne
rect 19687 3737 21800 3835
rect -300 3687 339 3737
rect -500 3639 339 3687
tri 339 3639 437 3737 sw
tri 437 3639 535 3737 ne
rect 535 3639 889 3737
tri 889 3639 987 3737 sw
tri 987 3639 1085 3737 ne
rect 1085 3639 1439 3737
tri 1439 3639 1537 3737 sw
tri 1537 3639 1635 3737 ne
rect 1635 3639 1989 3737
tri 1989 3639 2087 3737 sw
tri 2087 3639 2185 3737 ne
rect 2185 3639 2539 3737
tri 2539 3639 2637 3737 sw
tri 2637 3639 2735 3737 ne
rect 2735 3639 3089 3737
tri 3089 3639 3187 3737 sw
tri 3187 3639 3285 3737 ne
rect 3285 3639 3639 3737
tri 3639 3639 3737 3737 sw
tri 3737 3639 3835 3737 ne
rect 3835 3639 4189 3737
tri 4189 3639 4287 3737 sw
tri 4287 3639 4385 3737 ne
rect 4385 3639 4739 3737
tri 4739 3639 4837 3737 sw
tri 4837 3639 4935 3737 ne
rect 4935 3639 5289 3737
tri 5289 3639 5387 3737 sw
tri 5387 3639 5485 3737 ne
rect 5485 3639 5839 3737
tri 5839 3639 5937 3737 sw
tri 5937 3639 6035 3737 ne
rect 6035 3639 6389 3737
tri 6389 3639 6487 3737 sw
tri 6487 3639 6585 3737 ne
rect 6585 3639 6939 3737
tri 6939 3639 7037 3737 sw
tri 7037 3639 7135 3737 ne
rect 7135 3639 7489 3737
tri 7489 3639 7587 3737 sw
tri 7587 3639 7685 3737 ne
rect 7685 3639 8039 3737
tri 8039 3639 8137 3737 sw
tri 8137 3639 8235 3737 ne
rect 8235 3639 8589 3737
tri 8589 3639 8687 3737 sw
tri 8687 3639 8785 3737 ne
rect 8785 3639 9139 3737
tri 9139 3639 9237 3737 sw
tri 9237 3639 9335 3737 ne
rect 9335 3639 9689 3737
tri 9689 3639 9787 3737 sw
tri 9787 3639 9885 3737 ne
rect 9885 3639 10239 3737
tri 10239 3639 10337 3737 sw
tri 10337 3639 10435 3737 ne
rect 10435 3639 10789 3737
tri 10789 3639 10887 3737 sw
tri 10887 3639 10985 3737 ne
rect 10985 3639 11339 3737
tri 11339 3639 11437 3737 sw
tri 11437 3639 11535 3737 ne
rect 11535 3639 11889 3737
tri 11889 3639 11987 3737 sw
tri 11987 3639 12085 3737 ne
rect 12085 3639 12439 3737
tri 12439 3639 12537 3737 sw
tri 12537 3639 12635 3737 ne
rect 12635 3639 12989 3737
tri 12989 3639 13087 3737 sw
tri 13087 3639 13185 3737 ne
rect 13185 3639 13539 3737
tri 13539 3639 13637 3737 sw
tri 13637 3639 13735 3737 ne
rect 13735 3639 14089 3737
tri 14089 3639 14187 3737 sw
tri 14187 3639 14285 3737 ne
rect 14285 3639 14639 3737
tri 14639 3639 14737 3737 sw
tri 14737 3639 14835 3737 ne
rect 14835 3639 15189 3737
tri 15189 3639 15287 3737 sw
tri 15287 3639 15385 3737 ne
rect 15385 3639 15739 3737
tri 15739 3639 15837 3737 sw
tri 15837 3639 15935 3737 ne
rect 15935 3639 16289 3737
tri 16289 3639 16387 3737 sw
tri 16387 3639 16485 3737 ne
rect 16485 3639 16839 3737
tri 16839 3639 16937 3737 sw
tri 16937 3639 17035 3737 ne
rect 17035 3639 17389 3737
tri 17389 3639 17487 3737 sw
tri 17487 3639 17585 3737 ne
rect 17585 3639 17939 3737
tri 17939 3639 18037 3737 sw
tri 18037 3639 18135 3737 ne
rect 18135 3639 18489 3737
tri 18489 3639 18587 3737 sw
tri 18587 3639 18685 3737 ne
rect 18685 3639 19039 3737
tri 19039 3639 19137 3737 sw
tri 19137 3639 19235 3737 ne
rect 19235 3639 19589 3737
tri 19589 3639 19687 3737 sw
rect -500 3635 437 3639
rect -500 3515 215 3635
rect 335 3541 437 3635
tri 437 3541 535 3639 sw
tri 535 3541 633 3639 ne
rect 633 3635 987 3639
rect 633 3541 765 3635
rect 335 3515 535 3541
rect -500 3511 535 3515
tri 535 3511 565 3541 sw
tri 633 3511 663 3541 ne
rect 663 3515 765 3541
rect 885 3541 987 3635
tri 987 3541 1085 3639 sw
tri 1085 3541 1183 3639 ne
rect 1183 3635 1537 3639
rect 1183 3541 1315 3635
rect 885 3515 1085 3541
rect 663 3511 1085 3515
tri 1085 3511 1115 3541 sw
tri 1183 3511 1213 3541 ne
rect 1213 3515 1315 3541
rect 1435 3541 1537 3635
tri 1537 3541 1635 3639 sw
tri 1635 3541 1733 3639 ne
rect 1733 3635 2087 3639
rect 1733 3541 1865 3635
rect 1435 3515 1635 3541
rect 1213 3511 1635 3515
tri 1635 3511 1665 3541 sw
tri 1733 3511 1763 3541 ne
rect 1763 3515 1865 3541
rect 1985 3541 2087 3635
tri 2087 3541 2185 3639 sw
tri 2185 3541 2283 3639 ne
rect 2283 3635 2637 3639
rect 2283 3541 2415 3635
rect 1985 3515 2185 3541
rect 1763 3511 2185 3515
tri 2185 3511 2215 3541 sw
tri 2283 3511 2313 3541 ne
rect 2313 3515 2415 3541
rect 2535 3541 2637 3635
tri 2637 3541 2735 3639 sw
tri 2735 3541 2833 3639 ne
rect 2833 3635 3187 3639
rect 2833 3541 2965 3635
rect 2535 3515 2735 3541
rect 2313 3511 2735 3515
tri 2735 3511 2765 3541 sw
tri 2833 3511 2863 3541 ne
rect 2863 3515 2965 3541
rect 3085 3541 3187 3635
tri 3187 3541 3285 3639 sw
tri 3285 3541 3383 3639 ne
rect 3383 3635 3737 3639
rect 3383 3541 3515 3635
rect 3085 3515 3285 3541
rect 2863 3511 3285 3515
tri 3285 3511 3315 3541 sw
tri 3383 3511 3413 3541 ne
rect 3413 3515 3515 3541
rect 3635 3541 3737 3635
tri 3737 3541 3835 3639 sw
tri 3835 3541 3933 3639 ne
rect 3933 3635 4287 3639
rect 3933 3541 4065 3635
rect 3635 3515 3835 3541
rect 3413 3511 3835 3515
tri 3835 3511 3865 3541 sw
tri 3933 3511 3963 3541 ne
rect 3963 3515 4065 3541
rect 4185 3541 4287 3635
tri 4287 3541 4385 3639 sw
tri 4385 3541 4483 3639 ne
rect 4483 3635 4837 3639
rect 4483 3541 4615 3635
rect 4185 3515 4385 3541
rect 3963 3511 4385 3515
tri 4385 3511 4415 3541 sw
tri 4483 3511 4513 3541 ne
rect 4513 3515 4615 3541
rect 4735 3541 4837 3635
tri 4837 3541 4935 3639 sw
tri 4935 3541 5033 3639 ne
rect 5033 3635 5387 3639
rect 5033 3541 5165 3635
rect 4735 3515 4935 3541
rect 4513 3511 4935 3515
tri 4935 3511 4965 3541 sw
tri 5033 3511 5063 3541 ne
rect 5063 3515 5165 3541
rect 5285 3541 5387 3635
tri 5387 3541 5485 3639 sw
tri 5485 3541 5583 3639 ne
rect 5583 3635 5937 3639
rect 5583 3541 5715 3635
rect 5285 3515 5485 3541
rect 5063 3511 5485 3515
tri 5485 3511 5515 3541 sw
tri 5583 3511 5613 3541 ne
rect 5613 3515 5715 3541
rect 5835 3541 5937 3635
tri 5937 3541 6035 3639 sw
tri 6035 3541 6133 3639 ne
rect 6133 3635 6487 3639
rect 6133 3541 6265 3635
rect 5835 3515 6035 3541
rect 5613 3511 6035 3515
tri 6035 3511 6065 3541 sw
tri 6133 3511 6163 3541 ne
rect 6163 3515 6265 3541
rect 6385 3541 6487 3635
tri 6487 3541 6585 3639 sw
tri 6585 3541 6683 3639 ne
rect 6683 3635 7037 3639
rect 6683 3541 6815 3635
rect 6385 3515 6585 3541
rect 6163 3511 6585 3515
tri 6585 3511 6615 3541 sw
tri 6683 3511 6713 3541 ne
rect 6713 3515 6815 3541
rect 6935 3541 7037 3635
tri 7037 3541 7135 3639 sw
tri 7135 3541 7233 3639 ne
rect 7233 3635 7587 3639
rect 7233 3541 7365 3635
rect 6935 3515 7135 3541
rect 6713 3511 7135 3515
tri 7135 3511 7165 3541 sw
tri 7233 3511 7263 3541 ne
rect 7263 3515 7365 3541
rect 7485 3541 7587 3635
tri 7587 3541 7685 3639 sw
tri 7685 3541 7783 3639 ne
rect 7783 3635 8137 3639
rect 7783 3541 7915 3635
rect 7485 3515 7685 3541
rect 7263 3511 7685 3515
tri 7685 3511 7715 3541 sw
tri 7783 3511 7813 3541 ne
rect 7813 3515 7915 3541
rect 8035 3541 8137 3635
tri 8137 3541 8235 3639 sw
tri 8235 3541 8333 3639 ne
rect 8333 3635 8687 3639
rect 8333 3541 8465 3635
rect 8035 3515 8235 3541
rect 7813 3511 8235 3515
tri 8235 3511 8265 3541 sw
tri 8333 3511 8363 3541 ne
rect 8363 3515 8465 3541
rect 8585 3541 8687 3635
tri 8687 3541 8785 3639 sw
tri 8785 3541 8883 3639 ne
rect 8883 3635 9237 3639
rect 8883 3541 9015 3635
rect 8585 3515 8785 3541
rect 8363 3511 8785 3515
tri 8785 3511 8815 3541 sw
tri 8883 3511 8913 3541 ne
rect 8913 3515 9015 3541
rect 9135 3541 9237 3635
tri 9237 3541 9335 3639 sw
tri 9335 3541 9433 3639 ne
rect 9433 3635 9787 3639
rect 9433 3541 9565 3635
rect 9135 3515 9335 3541
rect 8913 3511 9335 3515
tri 9335 3511 9365 3541 sw
tri 9433 3511 9463 3541 ne
rect 9463 3515 9565 3541
rect 9685 3541 9787 3635
tri 9787 3541 9885 3639 sw
tri 9885 3541 9983 3639 ne
rect 9983 3635 10337 3639
rect 9983 3541 10115 3635
rect 9685 3515 9885 3541
rect 9463 3511 9885 3515
tri 9885 3511 9915 3541 sw
tri 9983 3511 10013 3541 ne
rect 10013 3515 10115 3541
rect 10235 3541 10337 3635
tri 10337 3541 10435 3639 sw
tri 10435 3541 10533 3639 ne
rect 10533 3635 10887 3639
rect 10533 3541 10665 3635
rect 10235 3515 10435 3541
rect 10013 3511 10435 3515
tri 10435 3511 10465 3541 sw
tri 10533 3511 10563 3541 ne
rect 10563 3515 10665 3541
rect 10785 3541 10887 3635
tri 10887 3541 10985 3639 sw
tri 10985 3541 11083 3639 ne
rect 11083 3635 11437 3639
rect 11083 3541 11215 3635
rect 10785 3515 10985 3541
rect 10563 3511 10985 3515
tri 10985 3511 11015 3541 sw
tri 11083 3511 11113 3541 ne
rect 11113 3515 11215 3541
rect 11335 3541 11437 3635
tri 11437 3541 11535 3639 sw
tri 11535 3541 11633 3639 ne
rect 11633 3635 11987 3639
rect 11633 3541 11765 3635
rect 11335 3515 11535 3541
rect 11113 3511 11535 3515
tri 11535 3511 11565 3541 sw
tri 11633 3511 11663 3541 ne
rect 11663 3515 11765 3541
rect 11885 3541 11987 3635
tri 11987 3541 12085 3639 sw
tri 12085 3541 12183 3639 ne
rect 12183 3635 12537 3639
rect 12183 3541 12315 3635
rect 11885 3515 12085 3541
rect 11663 3511 12085 3515
tri 12085 3511 12115 3541 sw
tri 12183 3511 12213 3541 ne
rect 12213 3515 12315 3541
rect 12435 3541 12537 3635
tri 12537 3541 12635 3639 sw
tri 12635 3541 12733 3639 ne
rect 12733 3635 13087 3639
rect 12733 3541 12865 3635
rect 12435 3515 12635 3541
rect 12213 3511 12635 3515
tri 12635 3511 12665 3541 sw
tri 12733 3511 12763 3541 ne
rect 12763 3515 12865 3541
rect 12985 3541 13087 3635
tri 13087 3541 13185 3639 sw
tri 13185 3541 13283 3639 ne
rect 13283 3635 13637 3639
rect 13283 3541 13415 3635
rect 12985 3515 13185 3541
rect 12763 3511 13185 3515
tri 13185 3511 13215 3541 sw
tri 13283 3511 13313 3541 ne
rect 13313 3515 13415 3541
rect 13535 3541 13637 3635
tri 13637 3541 13735 3639 sw
tri 13735 3541 13833 3639 ne
rect 13833 3635 14187 3639
rect 13833 3541 13965 3635
rect 13535 3515 13735 3541
rect 13313 3511 13735 3515
tri 13735 3511 13765 3541 sw
tri 13833 3511 13863 3541 ne
rect 13863 3515 13965 3541
rect 14085 3541 14187 3635
tri 14187 3541 14285 3639 sw
tri 14285 3541 14383 3639 ne
rect 14383 3635 14737 3639
rect 14383 3541 14515 3635
rect 14085 3515 14285 3541
rect 13863 3511 14285 3515
tri 14285 3511 14315 3541 sw
tri 14383 3511 14413 3541 ne
rect 14413 3515 14515 3541
rect 14635 3541 14737 3635
tri 14737 3541 14835 3639 sw
tri 14835 3541 14933 3639 ne
rect 14933 3635 15287 3639
rect 14933 3541 15065 3635
rect 14635 3515 14835 3541
rect 14413 3511 14835 3515
tri 14835 3511 14865 3541 sw
tri 14933 3511 14963 3541 ne
rect 14963 3515 15065 3541
rect 15185 3541 15287 3635
tri 15287 3541 15385 3639 sw
tri 15385 3541 15483 3639 ne
rect 15483 3635 15837 3639
rect 15483 3541 15615 3635
rect 15185 3515 15385 3541
rect 14963 3511 15385 3515
tri 15385 3511 15415 3541 sw
tri 15483 3511 15513 3541 ne
rect 15513 3515 15615 3541
rect 15735 3541 15837 3635
tri 15837 3541 15935 3639 sw
tri 15935 3541 16033 3639 ne
rect 16033 3635 16387 3639
rect 16033 3541 16165 3635
rect 15735 3515 15935 3541
rect 15513 3511 15935 3515
tri 15935 3511 15965 3541 sw
tri 16033 3511 16063 3541 ne
rect 16063 3515 16165 3541
rect 16285 3541 16387 3635
tri 16387 3541 16485 3639 sw
tri 16485 3541 16583 3639 ne
rect 16583 3635 16937 3639
rect 16583 3541 16715 3635
rect 16285 3515 16485 3541
rect 16063 3511 16485 3515
tri 16485 3511 16515 3541 sw
tri 16583 3511 16613 3541 ne
rect 16613 3515 16715 3541
rect 16835 3541 16937 3635
tri 16937 3541 17035 3639 sw
tri 17035 3541 17133 3639 ne
rect 17133 3635 17487 3639
rect 17133 3541 17265 3635
rect 16835 3515 17035 3541
rect 16613 3511 17035 3515
tri 17035 3511 17065 3541 sw
tri 17133 3511 17163 3541 ne
rect 17163 3515 17265 3541
rect 17385 3541 17487 3635
tri 17487 3541 17585 3639 sw
tri 17585 3541 17683 3639 ne
rect 17683 3635 18037 3639
rect 17683 3541 17815 3635
rect 17385 3515 17585 3541
rect 17163 3511 17585 3515
tri 17585 3511 17615 3541 sw
tri 17683 3511 17713 3541 ne
rect 17713 3515 17815 3541
rect 17935 3541 18037 3635
tri 18037 3541 18135 3639 sw
tri 18135 3541 18233 3639 ne
rect 18233 3635 18587 3639
rect 18233 3541 18365 3635
rect 17935 3515 18135 3541
rect 17713 3511 18135 3515
tri 18135 3511 18165 3541 sw
tri 18233 3511 18263 3541 ne
rect 18263 3515 18365 3541
rect 18485 3541 18587 3635
tri 18587 3541 18685 3639 sw
tri 18685 3541 18783 3639 ne
rect 18783 3635 19137 3639
rect 18783 3541 18915 3635
rect 18485 3515 18685 3541
rect 18263 3511 18685 3515
tri 18685 3511 18715 3541 sw
tri 18783 3511 18813 3541 ne
rect 18813 3515 18915 3541
rect 19035 3541 19137 3635
tri 19137 3541 19235 3639 sw
tri 19235 3541 19333 3639 ne
rect 19333 3635 20300 3639
rect 19333 3541 19465 3635
rect 19035 3515 19235 3541
rect 18813 3511 19235 3515
tri 19235 3511 19265 3541 sw
tri 19333 3511 19363 3541 ne
rect 19363 3515 19465 3541
rect 19585 3515 20300 3635
rect 19363 3511 20300 3515
tri 113 3413 211 3511 ne
rect 211 3413 565 3511
tri 565 3413 663 3511 sw
tri 663 3413 761 3511 ne
rect 761 3413 1115 3511
tri 1115 3413 1213 3511 sw
tri 1213 3413 1311 3511 ne
rect 1311 3413 1665 3511
tri 1665 3413 1763 3511 sw
tri 1763 3413 1861 3511 ne
rect 1861 3413 2215 3511
tri 2215 3413 2313 3511 sw
tri 2313 3413 2411 3511 ne
rect 2411 3413 2765 3511
tri 2765 3413 2863 3511 sw
tri 2863 3413 2961 3511 ne
rect 2961 3413 3315 3511
tri 3315 3413 3413 3511 sw
tri 3413 3413 3511 3511 ne
rect 3511 3413 3865 3511
tri 3865 3413 3963 3511 sw
tri 3963 3413 4061 3511 ne
rect 4061 3413 4415 3511
tri 4415 3413 4513 3511 sw
tri 4513 3413 4611 3511 ne
rect 4611 3413 4965 3511
tri 4965 3413 5063 3511 sw
tri 5063 3413 5161 3511 ne
rect 5161 3413 5515 3511
tri 5515 3413 5613 3511 sw
tri 5613 3413 5711 3511 ne
rect 5711 3413 6065 3511
tri 6065 3413 6163 3511 sw
tri 6163 3413 6261 3511 ne
rect 6261 3413 6615 3511
tri 6615 3413 6713 3511 sw
tri 6713 3413 6811 3511 ne
rect 6811 3413 7165 3511
tri 7165 3413 7263 3511 sw
tri 7263 3413 7361 3511 ne
rect 7361 3413 7715 3511
tri 7715 3413 7813 3511 sw
tri 7813 3413 7911 3511 ne
rect 7911 3413 8265 3511
tri 8265 3413 8363 3511 sw
tri 8363 3413 8461 3511 ne
rect 8461 3413 8815 3511
tri 8815 3413 8913 3511 sw
tri 8913 3413 9011 3511 ne
rect 9011 3413 9365 3511
tri 9365 3413 9463 3511 sw
tri 9463 3413 9561 3511 ne
rect 9561 3413 9915 3511
tri 9915 3413 10013 3511 sw
tri 10013 3413 10111 3511 ne
rect 10111 3413 10465 3511
tri 10465 3413 10563 3511 sw
tri 10563 3413 10661 3511 ne
rect 10661 3413 11015 3511
tri 11015 3413 11113 3511 sw
tri 11113 3413 11211 3511 ne
rect 11211 3413 11565 3511
tri 11565 3413 11663 3511 sw
tri 11663 3413 11761 3511 ne
rect 11761 3413 12115 3511
tri 12115 3413 12213 3511 sw
tri 12213 3413 12311 3511 ne
rect 12311 3413 12665 3511
tri 12665 3413 12763 3511 sw
tri 12763 3413 12861 3511 ne
rect 12861 3413 13215 3511
tri 13215 3413 13313 3511 sw
tri 13313 3413 13411 3511 ne
rect 13411 3413 13765 3511
tri 13765 3413 13863 3511 sw
tri 13863 3413 13961 3511 ne
rect 13961 3413 14315 3511
tri 14315 3413 14413 3511 sw
tri 14413 3413 14511 3511 ne
rect 14511 3413 14865 3511
tri 14865 3413 14963 3511 sw
tri 14963 3413 15061 3511 ne
rect 15061 3413 15415 3511
tri 15415 3413 15513 3511 sw
tri 15513 3413 15611 3511 ne
rect 15611 3413 15965 3511
tri 15965 3413 16063 3511 sw
tri 16063 3413 16161 3511 ne
rect 16161 3413 16515 3511
tri 16515 3413 16613 3511 sw
tri 16613 3413 16711 3511 ne
rect 16711 3413 17065 3511
tri 17065 3413 17163 3511 sw
tri 17163 3413 17261 3511 ne
rect 17261 3413 17615 3511
tri 17615 3413 17713 3511 sw
tri 17713 3413 17811 3511 ne
rect 17811 3413 18165 3511
tri 18165 3413 18263 3511 sw
tri 18263 3413 18361 3511 ne
rect 18361 3413 18715 3511
tri 18715 3413 18813 3511 sw
tri 18813 3413 18911 3511 ne
rect 18911 3413 19265 3511
tri 19265 3413 19363 3511 sw
tri 19363 3413 19461 3511 ne
rect 19461 3413 20300 3511
rect -2000 3383 113 3413
tri 113 3383 143 3413 sw
tri 211 3383 241 3413 ne
rect 241 3383 663 3413
tri 663 3383 693 3413 sw
tri 761 3383 791 3413 ne
rect 791 3383 1213 3413
tri 1213 3383 1243 3413 sw
tri 1311 3383 1341 3413 ne
rect 1341 3383 1763 3413
tri 1763 3383 1793 3413 sw
tri 1861 3383 1891 3413 ne
rect 1891 3383 2313 3413
tri 2313 3383 2343 3413 sw
tri 2411 3383 2441 3413 ne
rect 2441 3383 2863 3413
tri 2863 3383 2893 3413 sw
tri 2961 3383 2991 3413 ne
rect 2991 3383 3413 3413
tri 3413 3383 3443 3413 sw
tri 3511 3383 3541 3413 ne
rect 3541 3383 3963 3413
tri 3963 3383 3993 3413 sw
tri 4061 3383 4091 3413 ne
rect 4091 3383 4513 3413
tri 4513 3383 4543 3413 sw
tri 4611 3383 4641 3413 ne
rect 4641 3383 5063 3413
tri 5063 3383 5093 3413 sw
tri 5161 3383 5191 3413 ne
rect 5191 3383 5613 3413
tri 5613 3383 5643 3413 sw
tri 5711 3383 5741 3413 ne
rect 5741 3383 6163 3413
tri 6163 3383 6193 3413 sw
tri 6261 3383 6291 3413 ne
rect 6291 3383 6713 3413
tri 6713 3383 6743 3413 sw
tri 6811 3383 6841 3413 ne
rect 6841 3383 7263 3413
tri 7263 3383 7293 3413 sw
tri 7361 3383 7391 3413 ne
rect 7391 3383 7813 3413
tri 7813 3383 7843 3413 sw
tri 7911 3383 7941 3413 ne
rect 7941 3383 8363 3413
tri 8363 3383 8393 3413 sw
tri 8461 3383 8491 3413 ne
rect 8491 3383 8913 3413
tri 8913 3383 8943 3413 sw
tri 9011 3383 9041 3413 ne
rect 9041 3383 9463 3413
tri 9463 3383 9493 3413 sw
tri 9561 3383 9591 3413 ne
rect 9591 3383 10013 3413
tri 10013 3383 10043 3413 sw
tri 10111 3383 10141 3413 ne
rect 10141 3383 10563 3413
tri 10563 3383 10593 3413 sw
tri 10661 3383 10691 3413 ne
rect 10691 3383 11113 3413
tri 11113 3383 11143 3413 sw
tri 11211 3383 11241 3413 ne
rect 11241 3383 11663 3413
tri 11663 3383 11693 3413 sw
tri 11761 3383 11791 3413 ne
rect 11791 3383 12213 3413
tri 12213 3383 12243 3413 sw
tri 12311 3383 12341 3413 ne
rect 12341 3383 12763 3413
tri 12763 3383 12793 3413 sw
tri 12861 3383 12891 3413 ne
rect 12891 3383 13313 3413
tri 13313 3383 13343 3413 sw
tri 13411 3383 13441 3413 ne
rect 13441 3383 13863 3413
tri 13863 3383 13893 3413 sw
tri 13961 3383 13991 3413 ne
rect 13991 3383 14413 3413
tri 14413 3383 14443 3413 sw
tri 14511 3383 14541 3413 ne
rect 14541 3383 14963 3413
tri 14963 3383 14993 3413 sw
tri 15061 3383 15091 3413 ne
rect 15091 3383 15513 3413
tri 15513 3383 15543 3413 sw
tri 15611 3383 15641 3413 ne
rect 15641 3383 16063 3413
tri 16063 3383 16093 3413 sw
tri 16161 3383 16191 3413 ne
rect 16191 3383 16613 3413
tri 16613 3383 16643 3413 sw
tri 16711 3383 16741 3413 ne
rect 16741 3383 17163 3413
tri 17163 3383 17193 3413 sw
tri 17261 3383 17291 3413 ne
rect 17291 3383 17713 3413
tri 17713 3383 17743 3413 sw
tri 17811 3383 17841 3413 ne
rect 17841 3383 18263 3413
tri 18263 3383 18293 3413 sw
tri 18361 3383 18391 3413 ne
rect 18391 3383 18813 3413
tri 18813 3383 18843 3413 sw
tri 18911 3383 18941 3413 ne
rect 18941 3383 19363 3413
tri 19363 3383 19393 3413 sw
tri 19461 3383 19491 3413 ne
rect 19491 3383 20300 3413
rect -2000 3285 143 3383
tri 143 3285 241 3383 sw
tri 241 3285 339 3383 ne
rect 339 3285 693 3383
tri 693 3285 791 3383 sw
tri 791 3285 889 3383 ne
rect 889 3285 1243 3383
tri 1243 3285 1341 3383 sw
tri 1341 3285 1439 3383 ne
rect 1439 3285 1793 3383
tri 1793 3285 1891 3383 sw
tri 1891 3285 1989 3383 ne
rect 1989 3285 2343 3383
tri 2343 3285 2441 3383 sw
tri 2441 3285 2539 3383 ne
rect 2539 3285 2893 3383
tri 2893 3285 2991 3383 sw
tri 2991 3285 3089 3383 ne
rect 3089 3285 3443 3383
tri 3443 3285 3541 3383 sw
tri 3541 3285 3639 3383 ne
rect 3639 3285 3993 3383
tri 3993 3285 4091 3383 sw
tri 4091 3285 4189 3383 ne
rect 4189 3285 4543 3383
tri 4543 3285 4641 3383 sw
tri 4641 3285 4739 3383 ne
rect 4739 3285 5093 3383
tri 5093 3285 5191 3383 sw
tri 5191 3285 5289 3383 ne
rect 5289 3285 5643 3383
tri 5643 3285 5741 3383 sw
tri 5741 3285 5839 3383 ne
rect 5839 3285 6193 3383
tri 6193 3285 6291 3383 sw
tri 6291 3285 6389 3383 ne
rect 6389 3285 6743 3383
tri 6743 3285 6841 3383 sw
tri 6841 3285 6939 3383 ne
rect 6939 3285 7293 3383
tri 7293 3285 7391 3383 sw
tri 7391 3285 7489 3383 ne
rect 7489 3285 7843 3383
tri 7843 3285 7941 3383 sw
tri 7941 3285 8039 3383 ne
rect 8039 3285 8393 3383
tri 8393 3285 8491 3383 sw
tri 8491 3285 8589 3383 ne
rect 8589 3285 8943 3383
tri 8943 3285 9041 3383 sw
tri 9041 3285 9139 3383 ne
rect 9139 3285 9493 3383
tri 9493 3285 9591 3383 sw
tri 9591 3285 9689 3383 ne
rect 9689 3285 10043 3383
tri 10043 3285 10141 3383 sw
tri 10141 3285 10239 3383 ne
rect 10239 3285 10593 3383
tri 10593 3285 10691 3383 sw
tri 10691 3285 10789 3383 ne
rect 10789 3285 11143 3383
tri 11143 3285 11241 3383 sw
tri 11241 3285 11339 3383 ne
rect 11339 3285 11693 3383
tri 11693 3285 11791 3383 sw
tri 11791 3285 11889 3383 ne
rect 11889 3285 12243 3383
tri 12243 3285 12341 3383 sw
tri 12341 3285 12439 3383 ne
rect 12439 3285 12793 3383
tri 12793 3285 12891 3383 sw
tri 12891 3285 12989 3383 ne
rect 12989 3285 13343 3383
tri 13343 3285 13441 3383 sw
tri 13441 3285 13539 3383 ne
rect 13539 3285 13893 3383
tri 13893 3285 13991 3383 sw
tri 13991 3285 14089 3383 ne
rect 14089 3285 14443 3383
tri 14443 3285 14541 3383 sw
tri 14541 3285 14639 3383 ne
rect 14639 3285 14993 3383
tri 14993 3285 15091 3383 sw
tri 15091 3285 15189 3383 ne
rect 15189 3285 15543 3383
tri 15543 3285 15641 3383 sw
tri 15641 3285 15739 3383 ne
rect 15739 3285 16093 3383
tri 16093 3285 16191 3383 sw
tri 16191 3285 16289 3383 ne
rect 16289 3285 16643 3383
tri 16643 3285 16741 3383 sw
tri 16741 3285 16839 3383 ne
rect 16839 3285 17193 3383
tri 17193 3285 17291 3383 sw
tri 17291 3285 17389 3383 ne
rect 17389 3285 17743 3383
tri 17743 3285 17841 3383 sw
tri 17841 3285 17939 3383 ne
rect 17939 3285 18293 3383
tri 18293 3285 18391 3383 sw
tri 18391 3285 18489 3383 ne
rect 18489 3285 18843 3383
tri 18843 3285 18941 3383 sw
tri 18941 3285 19039 3383 ne
rect 19039 3285 19393 3383
tri 19393 3285 19491 3383 sw
tri 19491 3285 19589 3383 ne
rect 19589 3285 20300 3383
rect -2000 3187 241 3285
tri 241 3187 339 3285 sw
tri 339 3187 437 3285 ne
rect 437 3187 791 3285
tri 791 3187 889 3285 sw
tri 889 3187 987 3285 ne
rect 987 3187 1341 3285
tri 1341 3187 1439 3285 sw
tri 1439 3187 1537 3285 ne
rect 1537 3187 1891 3285
tri 1891 3187 1989 3285 sw
tri 1989 3187 2087 3285 ne
rect 2087 3187 2441 3285
tri 2441 3187 2539 3285 sw
tri 2539 3187 2637 3285 ne
rect 2637 3187 2991 3285
tri 2991 3187 3089 3285 sw
tri 3089 3187 3187 3285 ne
rect 3187 3187 3541 3285
tri 3541 3187 3639 3285 sw
tri 3639 3187 3737 3285 ne
rect 3737 3187 4091 3285
tri 4091 3187 4189 3285 sw
tri 4189 3187 4287 3285 ne
rect 4287 3187 4641 3285
tri 4641 3187 4739 3285 sw
tri 4739 3187 4837 3285 ne
rect 4837 3187 5191 3285
tri 5191 3187 5289 3285 sw
tri 5289 3187 5387 3285 ne
rect 5387 3187 5741 3285
tri 5741 3187 5839 3285 sw
tri 5839 3187 5937 3285 ne
rect 5937 3187 6291 3285
tri 6291 3187 6389 3285 sw
tri 6389 3187 6487 3285 ne
rect 6487 3187 6841 3285
tri 6841 3187 6939 3285 sw
tri 6939 3187 7037 3285 ne
rect 7037 3187 7391 3285
tri 7391 3187 7489 3285 sw
tri 7489 3187 7587 3285 ne
rect 7587 3187 7941 3285
tri 7941 3187 8039 3285 sw
tri 8039 3187 8137 3285 ne
rect 8137 3187 8491 3285
tri 8491 3187 8589 3285 sw
tri 8589 3187 8687 3285 ne
rect 8687 3187 9041 3285
tri 9041 3187 9139 3285 sw
tri 9139 3187 9237 3285 ne
rect 9237 3187 9591 3285
tri 9591 3187 9689 3285 sw
tri 9689 3187 9787 3285 ne
rect 9787 3187 10141 3285
tri 10141 3187 10239 3285 sw
tri 10239 3187 10337 3285 ne
rect 10337 3187 10691 3285
tri 10691 3187 10789 3285 sw
tri 10789 3187 10887 3285 ne
rect 10887 3187 11241 3285
tri 11241 3187 11339 3285 sw
tri 11339 3187 11437 3285 ne
rect 11437 3187 11791 3285
tri 11791 3187 11889 3285 sw
tri 11889 3187 11987 3285 ne
rect 11987 3187 12341 3285
tri 12341 3187 12439 3285 sw
tri 12439 3187 12537 3285 ne
rect 12537 3187 12891 3285
tri 12891 3187 12989 3285 sw
tri 12989 3187 13087 3285 ne
rect 13087 3187 13441 3285
tri 13441 3187 13539 3285 sw
tri 13539 3187 13637 3285 ne
rect 13637 3187 13991 3285
tri 13991 3187 14089 3285 sw
tri 14089 3187 14187 3285 ne
rect 14187 3187 14541 3285
tri 14541 3187 14639 3285 sw
tri 14639 3187 14737 3285 ne
rect 14737 3187 15091 3285
tri 15091 3187 15189 3285 sw
tri 15189 3187 15287 3285 ne
rect 15287 3187 15641 3285
tri 15641 3187 15739 3285 sw
tri 15739 3187 15837 3285 ne
rect 15837 3187 16191 3285
tri 16191 3187 16289 3285 sw
tri 16289 3187 16387 3285 ne
rect 16387 3187 16741 3285
tri 16741 3187 16839 3285 sw
tri 16839 3187 16937 3285 ne
rect 16937 3187 17291 3285
tri 17291 3187 17389 3285 sw
tri 17389 3187 17487 3285 ne
rect 17487 3187 17841 3285
tri 17841 3187 17939 3285 sw
tri 17939 3187 18037 3285 ne
rect 18037 3187 18391 3285
tri 18391 3187 18489 3285 sw
tri 18489 3187 18587 3285 ne
rect 18587 3187 18941 3285
tri 18941 3187 19039 3285 sw
tri 19039 3187 19137 3285 ne
rect 19137 3187 19491 3285
tri 19491 3187 19589 3285 sw
tri 19589 3187 19687 3285 ne
rect 19687 3187 20300 3285
rect -2000 3089 339 3187
tri 339 3089 437 3187 sw
tri 437 3089 535 3187 ne
rect 535 3089 889 3187
tri 889 3089 987 3187 sw
tri 987 3089 1085 3187 ne
rect 1085 3089 1439 3187
tri 1439 3089 1537 3187 sw
tri 1537 3089 1635 3187 ne
rect 1635 3089 1989 3187
tri 1989 3089 2087 3187 sw
tri 2087 3089 2185 3187 ne
rect 2185 3089 2539 3187
tri 2539 3089 2637 3187 sw
tri 2637 3089 2735 3187 ne
rect 2735 3089 3089 3187
tri 3089 3089 3187 3187 sw
tri 3187 3089 3285 3187 ne
rect 3285 3089 3639 3187
tri 3639 3089 3737 3187 sw
tri 3737 3089 3835 3187 ne
rect 3835 3089 4189 3187
tri 4189 3089 4287 3187 sw
tri 4287 3089 4385 3187 ne
rect 4385 3089 4739 3187
tri 4739 3089 4837 3187 sw
tri 4837 3089 4935 3187 ne
rect 4935 3089 5289 3187
tri 5289 3089 5387 3187 sw
tri 5387 3089 5485 3187 ne
rect 5485 3089 5839 3187
tri 5839 3089 5937 3187 sw
tri 5937 3089 6035 3187 ne
rect 6035 3089 6389 3187
tri 6389 3089 6487 3187 sw
tri 6487 3089 6585 3187 ne
rect 6585 3089 6939 3187
tri 6939 3089 7037 3187 sw
tri 7037 3089 7135 3187 ne
rect 7135 3089 7489 3187
tri 7489 3089 7587 3187 sw
tri 7587 3089 7685 3187 ne
rect 7685 3089 8039 3187
tri 8039 3089 8137 3187 sw
tri 8137 3089 8235 3187 ne
rect 8235 3089 8589 3187
tri 8589 3089 8687 3187 sw
tri 8687 3089 8785 3187 ne
rect 8785 3089 9139 3187
tri 9139 3089 9237 3187 sw
tri 9237 3089 9335 3187 ne
rect 9335 3089 9689 3187
tri 9689 3089 9787 3187 sw
tri 9787 3089 9885 3187 ne
rect 9885 3089 10239 3187
tri 10239 3089 10337 3187 sw
tri 10337 3089 10435 3187 ne
rect 10435 3089 10789 3187
tri 10789 3089 10887 3187 sw
tri 10887 3089 10985 3187 ne
rect 10985 3089 11339 3187
tri 11339 3089 11437 3187 sw
tri 11437 3089 11535 3187 ne
rect 11535 3089 11889 3187
tri 11889 3089 11987 3187 sw
tri 11987 3089 12085 3187 ne
rect 12085 3089 12439 3187
tri 12439 3089 12537 3187 sw
tri 12537 3089 12635 3187 ne
rect 12635 3089 12989 3187
tri 12989 3089 13087 3187 sw
tri 13087 3089 13185 3187 ne
rect 13185 3089 13539 3187
tri 13539 3089 13637 3187 sw
tri 13637 3089 13735 3187 ne
rect 13735 3089 14089 3187
tri 14089 3089 14187 3187 sw
tri 14187 3089 14285 3187 ne
rect 14285 3089 14639 3187
tri 14639 3089 14737 3187 sw
tri 14737 3089 14835 3187 ne
rect 14835 3089 15189 3187
tri 15189 3089 15287 3187 sw
tri 15287 3089 15385 3187 ne
rect 15385 3089 15739 3187
tri 15739 3089 15837 3187 sw
tri 15837 3089 15935 3187 ne
rect 15935 3089 16289 3187
tri 16289 3089 16387 3187 sw
tri 16387 3089 16485 3187 ne
rect 16485 3089 16839 3187
tri 16839 3089 16937 3187 sw
tri 16937 3089 17035 3187 ne
rect 17035 3089 17389 3187
tri 17389 3089 17487 3187 sw
tri 17487 3089 17585 3187 ne
rect 17585 3089 17939 3187
tri 17939 3089 18037 3187 sw
tri 18037 3089 18135 3187 ne
rect 18135 3089 18489 3187
tri 18489 3089 18587 3187 sw
tri 18587 3089 18685 3187 ne
rect 18685 3089 19039 3187
tri 19039 3089 19137 3187 sw
tri 19137 3089 19235 3187 ne
rect 19235 3089 19589 3187
tri 19589 3089 19687 3187 sw
rect 20800 3089 21800 3737
rect -2000 3085 437 3089
rect -2000 2965 215 3085
rect 335 2991 437 3085
tri 437 2991 535 3089 sw
tri 535 2991 633 3089 ne
rect 633 3085 987 3089
rect 633 2991 765 3085
rect 335 2965 535 2991
rect -2000 2961 535 2965
rect -2000 2313 -1000 2961
tri 113 2863 211 2961 ne
rect 211 2913 535 2961
tri 535 2913 613 2991 sw
tri 633 2913 711 2991 ne
rect 711 2965 765 2991
rect 885 2991 987 3085
tri 987 2991 1085 3089 sw
tri 1085 2991 1183 3089 ne
rect 1183 3085 1537 3089
rect 1183 2991 1315 3085
rect 885 2965 1085 2991
rect 711 2913 1085 2965
tri 1085 2913 1163 2991 sw
tri 1183 2913 1261 2991 ne
rect 1261 2965 1315 2991
rect 1435 2991 1537 3085
tri 1537 2991 1635 3089 sw
tri 1635 2991 1733 3089 ne
rect 1733 3085 2087 3089
rect 1733 2991 1865 3085
rect 1435 2965 1635 2991
rect 1261 2913 1635 2965
tri 1635 2913 1713 2991 sw
tri 1733 2913 1811 2991 ne
rect 1811 2965 1865 2991
rect 1985 2991 2087 3085
tri 2087 2991 2185 3089 sw
tri 2185 2991 2283 3089 ne
rect 2283 3085 2637 3089
rect 2283 2991 2415 3085
rect 1985 2965 2185 2991
rect 1811 2913 2185 2965
tri 2185 2913 2263 2991 sw
tri 2283 2913 2361 2991 ne
rect 2361 2965 2415 2991
rect 2535 2991 2637 3085
tri 2637 2991 2735 3089 sw
tri 2735 2991 2833 3089 ne
rect 2833 3085 3187 3089
rect 2833 2991 2965 3085
rect 2535 2965 2735 2991
rect 2361 2913 2735 2965
tri 2735 2913 2813 2991 sw
tri 2833 2913 2911 2991 ne
rect 2911 2965 2965 2991
rect 3085 2991 3187 3085
tri 3187 2991 3285 3089 sw
tri 3285 2991 3383 3089 ne
rect 3383 3085 3737 3089
rect 3383 2991 3515 3085
rect 3085 2965 3285 2991
rect 2911 2913 3285 2965
tri 3285 2913 3363 2991 sw
tri 3383 2913 3461 2991 ne
rect 3461 2965 3515 2991
rect 3635 2991 3737 3085
tri 3737 2991 3835 3089 sw
tri 3835 2991 3933 3089 ne
rect 3933 3085 4287 3089
rect 3933 2991 4065 3085
rect 3635 2965 3835 2991
rect 3461 2913 3835 2965
tri 3835 2913 3913 2991 sw
tri 3933 2913 4011 2991 ne
rect 4011 2965 4065 2991
rect 4185 2991 4287 3085
tri 4287 2991 4385 3089 sw
tri 4385 2991 4483 3089 ne
rect 4483 3085 4837 3089
rect 4483 2991 4615 3085
rect 4185 2965 4385 2991
rect 4011 2913 4385 2965
tri 4385 2913 4463 2991 sw
tri 4483 2913 4561 2991 ne
rect 4561 2965 4615 2991
rect 4735 2991 4837 3085
tri 4837 2991 4935 3089 sw
tri 4935 2991 5033 3089 ne
rect 5033 3085 5387 3089
rect 5033 2991 5165 3085
rect 4735 2965 4935 2991
rect 4561 2913 4935 2965
tri 4935 2913 5013 2991 sw
tri 5033 2913 5111 2991 ne
rect 5111 2965 5165 2991
rect 5285 2991 5387 3085
tri 5387 2991 5485 3089 sw
tri 5485 2991 5583 3089 ne
rect 5583 3085 5937 3089
rect 5583 2991 5715 3085
rect 5285 2965 5485 2991
rect 5111 2913 5485 2965
tri 5485 2913 5563 2991 sw
tri 5583 2913 5661 2991 ne
rect 5661 2965 5715 2991
rect 5835 2991 5937 3085
tri 5937 2991 6035 3089 sw
tri 6035 2991 6133 3089 ne
rect 6133 3085 6487 3089
rect 6133 2991 6265 3085
rect 5835 2965 6035 2991
rect 5661 2913 6035 2965
tri 6035 2913 6113 2991 sw
tri 6133 2913 6211 2991 ne
rect 6211 2965 6265 2991
rect 6385 2991 6487 3085
tri 6487 2991 6585 3089 sw
tri 6585 2991 6683 3089 ne
rect 6683 3085 7037 3089
rect 6683 2991 6815 3085
rect 6385 2965 6585 2991
rect 6211 2913 6585 2965
tri 6585 2913 6663 2991 sw
tri 6683 2913 6761 2991 ne
rect 6761 2965 6815 2991
rect 6935 2991 7037 3085
tri 7037 2991 7135 3089 sw
tri 7135 2991 7233 3089 ne
rect 7233 3085 7587 3089
rect 7233 2991 7365 3085
rect 6935 2965 7135 2991
rect 6761 2913 7135 2965
tri 7135 2913 7213 2991 sw
tri 7233 2913 7311 2991 ne
rect 7311 2965 7365 2991
rect 7485 2991 7587 3085
tri 7587 2991 7685 3089 sw
tri 7685 2991 7783 3089 ne
rect 7783 3085 8137 3089
rect 7783 2991 7915 3085
rect 7485 2965 7685 2991
rect 7311 2913 7685 2965
tri 7685 2913 7763 2991 sw
tri 7783 2913 7861 2991 ne
rect 7861 2965 7915 2991
rect 8035 2991 8137 3085
tri 8137 2991 8235 3089 sw
tri 8235 2991 8333 3089 ne
rect 8333 3085 8687 3089
rect 8333 2991 8465 3085
rect 8035 2965 8235 2991
rect 7861 2913 8235 2965
tri 8235 2913 8313 2991 sw
tri 8333 2913 8411 2991 ne
rect 8411 2965 8465 2991
rect 8585 2991 8687 3085
tri 8687 2991 8785 3089 sw
tri 8785 2991 8883 3089 ne
rect 8883 3085 9237 3089
rect 8883 2991 9015 3085
rect 8585 2965 8785 2991
rect 8411 2913 8785 2965
tri 8785 2913 8863 2991 sw
tri 8883 2913 8961 2991 ne
rect 8961 2965 9015 2991
rect 9135 2991 9237 3085
tri 9237 2991 9335 3089 sw
tri 9335 2991 9433 3089 ne
rect 9433 3085 9787 3089
rect 9433 2991 9565 3085
rect 9135 2965 9335 2991
rect 8961 2913 9335 2965
tri 9335 2913 9413 2991 sw
tri 9433 2913 9511 2991 ne
rect 9511 2965 9565 2991
rect 9685 2991 9787 3085
tri 9787 2991 9885 3089 sw
tri 9885 2991 9983 3089 ne
rect 9983 3085 10337 3089
rect 9983 2991 10115 3085
rect 9685 2965 9885 2991
rect 9511 2913 9885 2965
tri 9885 2913 9963 2991 sw
tri 9983 2913 10061 2991 ne
rect 10061 2965 10115 2991
rect 10235 2991 10337 3085
tri 10337 2991 10435 3089 sw
tri 10435 2991 10533 3089 ne
rect 10533 3085 10887 3089
rect 10533 2991 10665 3085
rect 10235 2965 10435 2991
rect 10061 2913 10435 2965
tri 10435 2913 10513 2991 sw
tri 10533 2913 10611 2991 ne
rect 10611 2965 10665 2991
rect 10785 2991 10887 3085
tri 10887 2991 10985 3089 sw
tri 10985 2991 11083 3089 ne
rect 11083 3085 11437 3089
rect 11083 2991 11215 3085
rect 10785 2965 10985 2991
rect 10611 2913 10985 2965
tri 10985 2913 11063 2991 sw
tri 11083 2913 11161 2991 ne
rect 11161 2965 11215 2991
rect 11335 2991 11437 3085
tri 11437 2991 11535 3089 sw
tri 11535 2991 11633 3089 ne
rect 11633 3085 11987 3089
rect 11633 2991 11765 3085
rect 11335 2965 11535 2991
rect 11161 2913 11535 2965
tri 11535 2913 11613 2991 sw
tri 11633 2913 11711 2991 ne
rect 11711 2965 11765 2991
rect 11885 2991 11987 3085
tri 11987 2991 12085 3089 sw
tri 12085 2991 12183 3089 ne
rect 12183 3085 12537 3089
rect 12183 2991 12315 3085
rect 11885 2965 12085 2991
rect 11711 2913 12085 2965
tri 12085 2913 12163 2991 sw
tri 12183 2913 12261 2991 ne
rect 12261 2965 12315 2991
rect 12435 2991 12537 3085
tri 12537 2991 12635 3089 sw
tri 12635 2991 12733 3089 ne
rect 12733 3085 13087 3089
rect 12733 2991 12865 3085
rect 12435 2965 12635 2991
rect 12261 2913 12635 2965
tri 12635 2913 12713 2991 sw
tri 12733 2913 12811 2991 ne
rect 12811 2965 12865 2991
rect 12985 2991 13087 3085
tri 13087 2991 13185 3089 sw
tri 13185 2991 13283 3089 ne
rect 13283 3085 13637 3089
rect 13283 2991 13415 3085
rect 12985 2965 13185 2991
rect 12811 2913 13185 2965
tri 13185 2913 13263 2991 sw
tri 13283 2913 13361 2991 ne
rect 13361 2965 13415 2991
rect 13535 2991 13637 3085
tri 13637 2991 13735 3089 sw
tri 13735 2991 13833 3089 ne
rect 13833 3085 14187 3089
rect 13833 2991 13965 3085
rect 13535 2965 13735 2991
rect 13361 2913 13735 2965
tri 13735 2913 13813 2991 sw
tri 13833 2913 13911 2991 ne
rect 13911 2965 13965 2991
rect 14085 2991 14187 3085
tri 14187 2991 14285 3089 sw
tri 14285 2991 14383 3089 ne
rect 14383 3085 14737 3089
rect 14383 2991 14515 3085
rect 14085 2965 14285 2991
rect 13911 2913 14285 2965
tri 14285 2913 14363 2991 sw
tri 14383 2913 14461 2991 ne
rect 14461 2965 14515 2991
rect 14635 2991 14737 3085
tri 14737 2991 14835 3089 sw
tri 14835 2991 14933 3089 ne
rect 14933 3085 15287 3089
rect 14933 2991 15065 3085
rect 14635 2965 14835 2991
rect 14461 2913 14835 2965
tri 14835 2913 14913 2991 sw
tri 14933 2913 15011 2991 ne
rect 15011 2965 15065 2991
rect 15185 2991 15287 3085
tri 15287 2991 15385 3089 sw
tri 15385 2991 15483 3089 ne
rect 15483 3085 15837 3089
rect 15483 2991 15615 3085
rect 15185 2965 15385 2991
rect 15011 2913 15385 2965
tri 15385 2913 15463 2991 sw
tri 15483 2913 15561 2991 ne
rect 15561 2965 15615 2991
rect 15735 2991 15837 3085
tri 15837 2991 15935 3089 sw
tri 15935 2991 16033 3089 ne
rect 16033 3085 16387 3089
rect 16033 2991 16165 3085
rect 15735 2965 15935 2991
rect 15561 2913 15935 2965
tri 15935 2913 16013 2991 sw
tri 16033 2913 16111 2991 ne
rect 16111 2965 16165 2991
rect 16285 2991 16387 3085
tri 16387 2991 16485 3089 sw
tri 16485 2991 16583 3089 ne
rect 16583 3085 16937 3089
rect 16583 2991 16715 3085
rect 16285 2965 16485 2991
rect 16111 2913 16485 2965
tri 16485 2913 16563 2991 sw
tri 16583 2913 16661 2991 ne
rect 16661 2965 16715 2991
rect 16835 2991 16937 3085
tri 16937 2991 17035 3089 sw
tri 17035 2991 17133 3089 ne
rect 17133 3085 17487 3089
rect 17133 2991 17265 3085
rect 16835 2965 17035 2991
rect 16661 2913 17035 2965
tri 17035 2913 17113 2991 sw
tri 17133 2913 17211 2991 ne
rect 17211 2965 17265 2991
rect 17385 2991 17487 3085
tri 17487 2991 17585 3089 sw
tri 17585 2991 17683 3089 ne
rect 17683 3085 18037 3089
rect 17683 2991 17815 3085
rect 17385 2965 17585 2991
rect 17211 2913 17585 2965
tri 17585 2913 17663 2991 sw
tri 17683 2913 17761 2991 ne
rect 17761 2965 17815 2991
rect 17935 2991 18037 3085
tri 18037 2991 18135 3089 sw
tri 18135 2991 18233 3089 ne
rect 18233 3085 18587 3089
rect 18233 2991 18365 3085
rect 17935 2965 18135 2991
rect 17761 2913 18135 2965
tri 18135 2913 18213 2991 sw
tri 18233 2913 18311 2991 ne
rect 18311 2965 18365 2991
rect 18485 2991 18587 3085
tri 18587 2991 18685 3089 sw
tri 18685 2991 18783 3089 ne
rect 18783 3085 19137 3089
rect 18783 2991 18915 3085
rect 18485 2965 18685 2991
rect 18311 2913 18685 2965
tri 18685 2913 18763 2991 sw
tri 18783 2913 18861 2991 ne
rect 18861 2965 18915 2991
rect 19035 2991 19137 3085
tri 19137 2991 19235 3089 sw
tri 19235 2991 19333 3089 ne
rect 19333 3085 21800 3089
rect 19333 2991 19465 3085
rect 19035 2965 19235 2991
rect 18861 2913 19235 2965
tri 19235 2913 19313 2991 sw
tri 19333 2913 19411 2991 ne
rect 19411 2965 19465 2991
rect 19585 2965 21800 3085
rect 19411 2913 21800 2965
rect 211 2863 613 2913
rect -500 2813 113 2863
tri 113 2813 163 2863 sw
tri 211 2813 261 2863 ne
rect 261 2833 613 2863
tri 613 2833 693 2913 sw
tri 711 2833 791 2913 ne
rect 791 2833 1163 2913
tri 1163 2833 1243 2913 sw
tri 1261 2833 1341 2913 ne
rect 1341 2833 1713 2913
tri 1713 2833 1793 2913 sw
tri 1811 2833 1891 2913 ne
rect 1891 2833 2263 2913
tri 2263 2833 2343 2913 sw
tri 2361 2833 2441 2913 ne
rect 2441 2833 2813 2913
tri 2813 2833 2893 2913 sw
tri 2911 2833 2991 2913 ne
rect 2991 2833 3363 2913
tri 3363 2833 3443 2913 sw
tri 3461 2833 3541 2913 ne
rect 3541 2833 3913 2913
tri 3913 2833 3993 2913 sw
tri 4011 2833 4091 2913 ne
rect 4091 2833 4463 2913
tri 4463 2833 4543 2913 sw
tri 4561 2833 4641 2913 ne
rect 4641 2833 5013 2913
tri 5013 2833 5093 2913 sw
tri 5111 2833 5191 2913 ne
rect 5191 2833 5563 2913
tri 5563 2833 5643 2913 sw
tri 5661 2833 5741 2913 ne
rect 5741 2833 6113 2913
tri 6113 2833 6193 2913 sw
tri 6211 2833 6291 2913 ne
rect 6291 2833 6663 2913
tri 6663 2833 6743 2913 sw
tri 6761 2833 6841 2913 ne
rect 6841 2833 7213 2913
tri 7213 2833 7293 2913 sw
tri 7311 2833 7391 2913 ne
rect 7391 2833 7763 2913
tri 7763 2833 7843 2913 sw
tri 7861 2833 7941 2913 ne
rect 7941 2833 8313 2913
tri 8313 2833 8393 2913 sw
tri 8411 2833 8491 2913 ne
rect 8491 2833 8863 2913
tri 8863 2833 8943 2913 sw
tri 8961 2833 9041 2913 ne
rect 9041 2833 9413 2913
tri 9413 2833 9493 2913 sw
tri 9511 2833 9591 2913 ne
rect 9591 2833 9963 2913
tri 9963 2833 10043 2913 sw
tri 10061 2833 10141 2913 ne
rect 10141 2833 10513 2913
tri 10513 2833 10593 2913 sw
tri 10611 2833 10691 2913 ne
rect 10691 2833 11063 2913
tri 11063 2833 11143 2913 sw
tri 11161 2833 11241 2913 ne
rect 11241 2833 11613 2913
tri 11613 2833 11693 2913 sw
tri 11711 2833 11791 2913 ne
rect 11791 2833 12163 2913
tri 12163 2833 12243 2913 sw
tri 12261 2833 12341 2913 ne
rect 12341 2833 12713 2913
tri 12713 2833 12793 2913 sw
tri 12811 2833 12891 2913 ne
rect 12891 2833 13263 2913
tri 13263 2833 13343 2913 sw
tri 13361 2833 13441 2913 ne
rect 13441 2833 13813 2913
tri 13813 2833 13893 2913 sw
tri 13911 2833 13991 2913 ne
rect 13991 2833 14363 2913
tri 14363 2833 14443 2913 sw
tri 14461 2833 14541 2913 ne
rect 14541 2833 14913 2913
tri 14913 2833 14993 2913 sw
tri 15011 2833 15091 2913 ne
rect 15091 2833 15463 2913
tri 15463 2833 15543 2913 sw
tri 15561 2833 15641 2913 ne
rect 15641 2833 16013 2913
tri 16013 2833 16093 2913 sw
tri 16111 2833 16191 2913 ne
rect 16191 2833 16563 2913
tri 16563 2833 16643 2913 sw
tri 16661 2833 16741 2913 ne
rect 16741 2833 17113 2913
tri 17113 2833 17193 2913 sw
tri 17211 2833 17291 2913 ne
rect 17291 2833 17663 2913
tri 17663 2833 17743 2913 sw
tri 17761 2833 17841 2913 ne
rect 17841 2833 18213 2913
tri 18213 2833 18293 2913 sw
tri 18311 2833 18391 2913 ne
rect 18391 2833 18763 2913
tri 18763 2833 18843 2913 sw
tri 18861 2833 18941 2913 ne
rect 18941 2833 19313 2913
tri 19313 2833 19393 2913 sw
tri 19411 2833 19491 2913 ne
rect 19491 2833 20100 2913
rect 261 2813 693 2833
rect -500 2735 163 2813
tri 163 2735 241 2813 sw
tri 261 2735 339 2813 ne
rect 339 2735 693 2813
tri 693 2735 791 2833 sw
tri 791 2735 889 2833 ne
rect 889 2735 1243 2833
tri 1243 2735 1341 2833 sw
tri 1341 2735 1439 2833 ne
rect 1439 2735 1793 2833
tri 1793 2735 1891 2833 sw
tri 1891 2735 1989 2833 ne
rect 1989 2735 2343 2833
tri 2343 2735 2441 2833 sw
tri 2441 2735 2539 2833 ne
rect 2539 2735 2893 2833
tri 2893 2735 2991 2833 sw
tri 2991 2735 3089 2833 ne
rect 3089 2735 3443 2833
tri 3443 2735 3541 2833 sw
tri 3541 2735 3639 2833 ne
rect 3639 2735 3993 2833
tri 3993 2735 4091 2833 sw
tri 4091 2735 4189 2833 ne
rect 4189 2735 4543 2833
tri 4543 2735 4641 2833 sw
tri 4641 2735 4739 2833 ne
rect 4739 2735 5093 2833
tri 5093 2735 5191 2833 sw
tri 5191 2735 5289 2833 ne
rect 5289 2735 5643 2833
tri 5643 2735 5741 2833 sw
tri 5741 2735 5839 2833 ne
rect 5839 2735 6193 2833
tri 6193 2735 6291 2833 sw
tri 6291 2735 6389 2833 ne
rect 6389 2735 6743 2833
tri 6743 2735 6841 2833 sw
tri 6841 2735 6939 2833 ne
rect 6939 2735 7293 2833
tri 7293 2735 7391 2833 sw
tri 7391 2735 7489 2833 ne
rect 7489 2735 7843 2833
tri 7843 2735 7941 2833 sw
tri 7941 2735 8039 2833 ne
rect 8039 2735 8393 2833
tri 8393 2735 8491 2833 sw
tri 8491 2735 8589 2833 ne
rect 8589 2735 8943 2833
tri 8943 2735 9041 2833 sw
tri 9041 2735 9139 2833 ne
rect 9139 2735 9493 2833
tri 9493 2735 9591 2833 sw
tri 9591 2735 9689 2833 ne
rect 9689 2735 10043 2833
tri 10043 2735 10141 2833 sw
tri 10141 2735 10239 2833 ne
rect 10239 2735 10593 2833
tri 10593 2735 10691 2833 sw
tri 10691 2735 10789 2833 ne
rect 10789 2735 11143 2833
tri 11143 2735 11241 2833 sw
tri 11241 2735 11339 2833 ne
rect 11339 2735 11693 2833
tri 11693 2735 11791 2833 sw
tri 11791 2735 11889 2833 ne
rect 11889 2735 12243 2833
tri 12243 2735 12341 2833 sw
tri 12341 2735 12439 2833 ne
rect 12439 2735 12793 2833
tri 12793 2735 12891 2833 sw
tri 12891 2735 12989 2833 ne
rect 12989 2735 13343 2833
tri 13343 2735 13441 2833 sw
tri 13441 2735 13539 2833 ne
rect 13539 2735 13893 2833
tri 13893 2735 13991 2833 sw
tri 13991 2735 14089 2833 ne
rect 14089 2735 14443 2833
tri 14443 2735 14541 2833 sw
tri 14541 2735 14639 2833 ne
rect 14639 2735 14993 2833
tri 14993 2735 15091 2833 sw
tri 15091 2735 15189 2833 ne
rect 15189 2735 15543 2833
tri 15543 2735 15641 2833 sw
tri 15641 2735 15739 2833 ne
rect 15739 2735 16093 2833
tri 16093 2735 16191 2833 sw
tri 16191 2735 16289 2833 ne
rect 16289 2735 16643 2833
tri 16643 2735 16741 2833 sw
tri 16741 2735 16839 2833 ne
rect 16839 2735 17193 2833
tri 17193 2735 17291 2833 sw
tri 17291 2735 17389 2833 ne
rect 17389 2735 17743 2833
tri 17743 2735 17841 2833 sw
tri 17841 2735 17939 2833 ne
rect 17939 2735 18293 2833
tri 18293 2735 18391 2833 sw
tri 18391 2735 18489 2833 ne
rect 18489 2735 18843 2833
tri 18843 2735 18941 2833 sw
tri 18941 2735 19039 2833 ne
rect 19039 2735 19393 2833
tri 19393 2735 19491 2833 sw
tri 19491 2735 19589 2833 ne
rect 19589 2813 20100 2833
rect 20200 2813 21800 2913
rect 19589 2735 21800 2813
rect -500 2687 241 2735
rect -500 2587 -400 2687
rect -300 2637 241 2687
tri 241 2637 339 2735 sw
tri 339 2637 437 2735 ne
rect 437 2637 791 2735
tri 791 2637 889 2735 sw
tri 889 2637 987 2735 ne
rect 987 2637 1341 2735
tri 1341 2637 1439 2735 sw
tri 1439 2637 1537 2735 ne
rect 1537 2637 1891 2735
tri 1891 2637 1989 2735 sw
tri 1989 2637 2087 2735 ne
rect 2087 2637 2441 2735
tri 2441 2637 2539 2735 sw
tri 2539 2637 2637 2735 ne
rect 2637 2637 2991 2735
tri 2991 2637 3089 2735 sw
tri 3089 2637 3187 2735 ne
rect 3187 2637 3541 2735
tri 3541 2637 3639 2735 sw
tri 3639 2637 3737 2735 ne
rect 3737 2637 4091 2735
tri 4091 2637 4189 2735 sw
tri 4189 2637 4287 2735 ne
rect 4287 2637 4641 2735
tri 4641 2637 4739 2735 sw
tri 4739 2637 4837 2735 ne
rect 4837 2637 5191 2735
tri 5191 2637 5289 2735 sw
tri 5289 2637 5387 2735 ne
rect 5387 2637 5741 2735
tri 5741 2637 5839 2735 sw
tri 5839 2637 5937 2735 ne
rect 5937 2637 6291 2735
tri 6291 2637 6389 2735 sw
tri 6389 2637 6487 2735 ne
rect 6487 2637 6841 2735
tri 6841 2637 6939 2735 sw
tri 6939 2637 7037 2735 ne
rect 7037 2637 7391 2735
tri 7391 2637 7489 2735 sw
tri 7489 2637 7587 2735 ne
rect 7587 2637 7941 2735
tri 7941 2637 8039 2735 sw
tri 8039 2637 8137 2735 ne
rect 8137 2637 8491 2735
tri 8491 2637 8589 2735 sw
tri 8589 2637 8687 2735 ne
rect 8687 2637 9041 2735
tri 9041 2637 9139 2735 sw
tri 9139 2637 9237 2735 ne
rect 9237 2637 9591 2735
tri 9591 2637 9689 2735 sw
tri 9689 2637 9787 2735 ne
rect 9787 2637 10141 2735
tri 10141 2637 10239 2735 sw
tri 10239 2637 10337 2735 ne
rect 10337 2637 10691 2735
tri 10691 2637 10789 2735 sw
tri 10789 2637 10887 2735 ne
rect 10887 2637 11241 2735
tri 11241 2637 11339 2735 sw
tri 11339 2637 11437 2735 ne
rect 11437 2637 11791 2735
tri 11791 2637 11889 2735 sw
tri 11889 2637 11987 2735 ne
rect 11987 2637 12341 2735
tri 12341 2637 12439 2735 sw
tri 12439 2637 12537 2735 ne
rect 12537 2637 12891 2735
tri 12891 2637 12989 2735 sw
tri 12989 2637 13087 2735 ne
rect 13087 2637 13441 2735
tri 13441 2637 13539 2735 sw
tri 13539 2637 13637 2735 ne
rect 13637 2637 13991 2735
tri 13991 2637 14089 2735 sw
tri 14089 2637 14187 2735 ne
rect 14187 2637 14541 2735
tri 14541 2637 14639 2735 sw
tri 14639 2637 14737 2735 ne
rect 14737 2637 15091 2735
tri 15091 2637 15189 2735 sw
tri 15189 2637 15287 2735 ne
rect 15287 2637 15641 2735
tri 15641 2637 15739 2735 sw
tri 15739 2637 15837 2735 ne
rect 15837 2637 16191 2735
tri 16191 2637 16289 2735 sw
tri 16289 2637 16387 2735 ne
rect 16387 2637 16741 2735
tri 16741 2637 16839 2735 sw
tri 16839 2637 16937 2735 ne
rect 16937 2637 17291 2735
tri 17291 2637 17389 2735 sw
tri 17389 2637 17487 2735 ne
rect 17487 2637 17841 2735
tri 17841 2637 17939 2735 sw
tri 17939 2637 18037 2735 ne
rect 18037 2637 18391 2735
tri 18391 2637 18489 2735 sw
tri 18489 2637 18587 2735 ne
rect 18587 2637 18941 2735
tri 18941 2637 19039 2735 sw
tri 19039 2637 19137 2735 ne
rect 19137 2637 19491 2735
tri 19491 2637 19589 2735 sw
tri 19589 2637 19687 2735 ne
rect 19687 2637 21800 2735
rect -300 2587 339 2637
rect -500 2539 339 2587
tri 339 2539 437 2637 sw
tri 437 2539 535 2637 ne
rect 535 2539 889 2637
tri 889 2539 987 2637 sw
tri 987 2539 1085 2637 ne
rect 1085 2539 1439 2637
tri 1439 2539 1537 2637 sw
tri 1537 2539 1635 2637 ne
rect 1635 2539 1989 2637
tri 1989 2539 2087 2637 sw
tri 2087 2539 2185 2637 ne
rect 2185 2539 2539 2637
tri 2539 2539 2637 2637 sw
tri 2637 2539 2735 2637 ne
rect 2735 2539 3089 2637
tri 3089 2539 3187 2637 sw
tri 3187 2539 3285 2637 ne
rect 3285 2539 3639 2637
tri 3639 2539 3737 2637 sw
tri 3737 2539 3835 2637 ne
rect 3835 2539 4189 2637
tri 4189 2539 4287 2637 sw
tri 4287 2539 4385 2637 ne
rect 4385 2539 4739 2637
tri 4739 2539 4837 2637 sw
tri 4837 2539 4935 2637 ne
rect 4935 2539 5289 2637
tri 5289 2539 5387 2637 sw
tri 5387 2539 5485 2637 ne
rect 5485 2539 5839 2637
tri 5839 2539 5937 2637 sw
tri 5937 2539 6035 2637 ne
rect 6035 2539 6389 2637
tri 6389 2539 6487 2637 sw
tri 6487 2539 6585 2637 ne
rect 6585 2539 6939 2637
tri 6939 2539 7037 2637 sw
tri 7037 2539 7135 2637 ne
rect 7135 2539 7489 2637
tri 7489 2539 7587 2637 sw
tri 7587 2539 7685 2637 ne
rect 7685 2539 8039 2637
tri 8039 2539 8137 2637 sw
tri 8137 2539 8235 2637 ne
rect 8235 2539 8589 2637
tri 8589 2539 8687 2637 sw
tri 8687 2539 8785 2637 ne
rect 8785 2539 9139 2637
tri 9139 2539 9237 2637 sw
tri 9237 2539 9335 2637 ne
rect 9335 2539 9689 2637
tri 9689 2539 9787 2637 sw
tri 9787 2539 9885 2637 ne
rect 9885 2539 10239 2637
tri 10239 2539 10337 2637 sw
tri 10337 2539 10435 2637 ne
rect 10435 2539 10789 2637
tri 10789 2539 10887 2637 sw
tri 10887 2539 10985 2637 ne
rect 10985 2539 11339 2637
tri 11339 2539 11437 2637 sw
tri 11437 2539 11535 2637 ne
rect 11535 2539 11889 2637
tri 11889 2539 11987 2637 sw
tri 11987 2539 12085 2637 ne
rect 12085 2539 12439 2637
tri 12439 2539 12537 2637 sw
tri 12537 2539 12635 2637 ne
rect 12635 2539 12989 2637
tri 12989 2539 13087 2637 sw
tri 13087 2539 13185 2637 ne
rect 13185 2539 13539 2637
tri 13539 2539 13637 2637 sw
tri 13637 2539 13735 2637 ne
rect 13735 2539 14089 2637
tri 14089 2539 14187 2637 sw
tri 14187 2539 14285 2637 ne
rect 14285 2539 14639 2637
tri 14639 2539 14737 2637 sw
tri 14737 2539 14835 2637 ne
rect 14835 2539 15189 2637
tri 15189 2539 15287 2637 sw
tri 15287 2539 15385 2637 ne
rect 15385 2539 15739 2637
tri 15739 2539 15837 2637 sw
tri 15837 2539 15935 2637 ne
rect 15935 2539 16289 2637
tri 16289 2539 16387 2637 sw
tri 16387 2539 16485 2637 ne
rect 16485 2539 16839 2637
tri 16839 2539 16937 2637 sw
tri 16937 2539 17035 2637 ne
rect 17035 2539 17389 2637
tri 17389 2539 17487 2637 sw
tri 17487 2539 17585 2637 ne
rect 17585 2539 17939 2637
tri 17939 2539 18037 2637 sw
tri 18037 2539 18135 2637 ne
rect 18135 2539 18489 2637
tri 18489 2539 18587 2637 sw
tri 18587 2539 18685 2637 ne
rect 18685 2539 19039 2637
tri 19039 2539 19137 2637 sw
tri 19137 2539 19235 2637 ne
rect 19235 2539 19589 2637
tri 19589 2539 19687 2637 sw
rect -500 2535 437 2539
rect -500 2415 215 2535
rect 335 2441 437 2535
tri 437 2441 535 2539 sw
tri 535 2441 633 2539 ne
rect 633 2535 987 2539
rect 633 2441 765 2535
rect 335 2415 535 2441
rect -500 2411 535 2415
tri 535 2411 565 2441 sw
tri 633 2411 663 2441 ne
rect 663 2415 765 2441
rect 885 2441 987 2535
tri 987 2441 1085 2539 sw
tri 1085 2441 1183 2539 ne
rect 1183 2535 1537 2539
rect 1183 2441 1315 2535
rect 885 2415 1085 2441
rect 663 2411 1085 2415
tri 1085 2411 1115 2441 sw
tri 1183 2411 1213 2441 ne
rect 1213 2415 1315 2441
rect 1435 2441 1537 2535
tri 1537 2441 1635 2539 sw
tri 1635 2441 1733 2539 ne
rect 1733 2535 2087 2539
rect 1733 2441 1865 2535
rect 1435 2415 1635 2441
rect 1213 2411 1635 2415
tri 1635 2411 1665 2441 sw
tri 1733 2411 1763 2441 ne
rect 1763 2415 1865 2441
rect 1985 2441 2087 2535
tri 2087 2441 2185 2539 sw
tri 2185 2441 2283 2539 ne
rect 2283 2535 2637 2539
rect 2283 2441 2415 2535
rect 1985 2415 2185 2441
rect 1763 2411 2185 2415
tri 2185 2411 2215 2441 sw
tri 2283 2411 2313 2441 ne
rect 2313 2415 2415 2441
rect 2535 2441 2637 2535
tri 2637 2441 2735 2539 sw
tri 2735 2441 2833 2539 ne
rect 2833 2535 3187 2539
rect 2833 2441 2965 2535
rect 2535 2415 2735 2441
rect 2313 2411 2735 2415
tri 2735 2411 2765 2441 sw
tri 2833 2411 2863 2441 ne
rect 2863 2415 2965 2441
rect 3085 2441 3187 2535
tri 3187 2441 3285 2539 sw
tri 3285 2441 3383 2539 ne
rect 3383 2535 3737 2539
rect 3383 2441 3515 2535
rect 3085 2415 3285 2441
rect 2863 2411 3285 2415
tri 3285 2411 3315 2441 sw
tri 3383 2411 3413 2441 ne
rect 3413 2415 3515 2441
rect 3635 2441 3737 2535
tri 3737 2441 3835 2539 sw
tri 3835 2441 3933 2539 ne
rect 3933 2535 4287 2539
rect 3933 2441 4065 2535
rect 3635 2415 3835 2441
rect 3413 2411 3835 2415
tri 3835 2411 3865 2441 sw
tri 3933 2411 3963 2441 ne
rect 3963 2415 4065 2441
rect 4185 2441 4287 2535
tri 4287 2441 4385 2539 sw
tri 4385 2441 4483 2539 ne
rect 4483 2535 4837 2539
rect 4483 2441 4615 2535
rect 4185 2415 4385 2441
rect 3963 2411 4385 2415
tri 4385 2411 4415 2441 sw
tri 4483 2411 4513 2441 ne
rect 4513 2415 4615 2441
rect 4735 2441 4837 2535
tri 4837 2441 4935 2539 sw
tri 4935 2441 5033 2539 ne
rect 5033 2535 5387 2539
rect 5033 2441 5165 2535
rect 4735 2415 4935 2441
rect 4513 2411 4935 2415
tri 4935 2411 4965 2441 sw
tri 5033 2411 5063 2441 ne
rect 5063 2415 5165 2441
rect 5285 2441 5387 2535
tri 5387 2441 5485 2539 sw
tri 5485 2441 5583 2539 ne
rect 5583 2535 5937 2539
rect 5583 2441 5715 2535
rect 5285 2415 5485 2441
rect 5063 2411 5485 2415
tri 5485 2411 5515 2441 sw
tri 5583 2411 5613 2441 ne
rect 5613 2415 5715 2441
rect 5835 2441 5937 2535
tri 5937 2441 6035 2539 sw
tri 6035 2441 6133 2539 ne
rect 6133 2535 6487 2539
rect 6133 2441 6265 2535
rect 5835 2415 6035 2441
rect 5613 2411 6035 2415
tri 6035 2411 6065 2441 sw
tri 6133 2411 6163 2441 ne
rect 6163 2415 6265 2441
rect 6385 2441 6487 2535
tri 6487 2441 6585 2539 sw
tri 6585 2441 6683 2539 ne
rect 6683 2535 7037 2539
rect 6683 2441 6815 2535
rect 6385 2415 6585 2441
rect 6163 2411 6585 2415
tri 6585 2411 6615 2441 sw
tri 6683 2411 6713 2441 ne
rect 6713 2415 6815 2441
rect 6935 2441 7037 2535
tri 7037 2441 7135 2539 sw
tri 7135 2441 7233 2539 ne
rect 7233 2535 7587 2539
rect 7233 2441 7365 2535
rect 6935 2415 7135 2441
rect 6713 2411 7135 2415
tri 7135 2411 7165 2441 sw
tri 7233 2411 7263 2441 ne
rect 7263 2415 7365 2441
rect 7485 2441 7587 2535
tri 7587 2441 7685 2539 sw
tri 7685 2441 7783 2539 ne
rect 7783 2535 8137 2539
rect 7783 2441 7915 2535
rect 7485 2415 7685 2441
rect 7263 2411 7685 2415
tri 7685 2411 7715 2441 sw
tri 7783 2411 7813 2441 ne
rect 7813 2415 7915 2441
rect 8035 2441 8137 2535
tri 8137 2441 8235 2539 sw
tri 8235 2441 8333 2539 ne
rect 8333 2535 8687 2539
rect 8333 2441 8465 2535
rect 8035 2415 8235 2441
rect 7813 2411 8235 2415
tri 8235 2411 8265 2441 sw
tri 8333 2411 8363 2441 ne
rect 8363 2415 8465 2441
rect 8585 2441 8687 2535
tri 8687 2441 8785 2539 sw
tri 8785 2441 8883 2539 ne
rect 8883 2535 9237 2539
rect 8883 2441 9015 2535
rect 8585 2415 8785 2441
rect 8363 2411 8785 2415
tri 8785 2411 8815 2441 sw
tri 8883 2411 8913 2441 ne
rect 8913 2415 9015 2441
rect 9135 2441 9237 2535
tri 9237 2441 9335 2539 sw
tri 9335 2441 9433 2539 ne
rect 9433 2535 9787 2539
rect 9433 2441 9565 2535
rect 9135 2415 9335 2441
rect 8913 2411 9335 2415
tri 9335 2411 9365 2441 sw
tri 9433 2411 9463 2441 ne
rect 9463 2415 9565 2441
rect 9685 2441 9787 2535
tri 9787 2441 9885 2539 sw
tri 9885 2441 9983 2539 ne
rect 9983 2535 10337 2539
rect 9983 2441 10115 2535
rect 9685 2415 9885 2441
rect 9463 2411 9885 2415
tri 9885 2411 9915 2441 sw
tri 9983 2411 10013 2441 ne
rect 10013 2415 10115 2441
rect 10235 2441 10337 2535
tri 10337 2441 10435 2539 sw
tri 10435 2441 10533 2539 ne
rect 10533 2535 10887 2539
rect 10533 2441 10665 2535
rect 10235 2415 10435 2441
rect 10013 2411 10435 2415
tri 10435 2411 10465 2441 sw
tri 10533 2411 10563 2441 ne
rect 10563 2415 10665 2441
rect 10785 2441 10887 2535
tri 10887 2441 10985 2539 sw
tri 10985 2441 11083 2539 ne
rect 11083 2535 11437 2539
rect 11083 2441 11215 2535
rect 10785 2415 10985 2441
rect 10563 2411 10985 2415
tri 10985 2411 11015 2441 sw
tri 11083 2411 11113 2441 ne
rect 11113 2415 11215 2441
rect 11335 2441 11437 2535
tri 11437 2441 11535 2539 sw
tri 11535 2441 11633 2539 ne
rect 11633 2535 11987 2539
rect 11633 2441 11765 2535
rect 11335 2415 11535 2441
rect 11113 2411 11535 2415
tri 11535 2411 11565 2441 sw
tri 11633 2411 11663 2441 ne
rect 11663 2415 11765 2441
rect 11885 2441 11987 2535
tri 11987 2441 12085 2539 sw
tri 12085 2441 12183 2539 ne
rect 12183 2535 12537 2539
rect 12183 2441 12315 2535
rect 11885 2415 12085 2441
rect 11663 2411 12085 2415
tri 12085 2411 12115 2441 sw
tri 12183 2411 12213 2441 ne
rect 12213 2415 12315 2441
rect 12435 2441 12537 2535
tri 12537 2441 12635 2539 sw
tri 12635 2441 12733 2539 ne
rect 12733 2535 13087 2539
rect 12733 2441 12865 2535
rect 12435 2415 12635 2441
rect 12213 2411 12635 2415
tri 12635 2411 12665 2441 sw
tri 12733 2411 12763 2441 ne
rect 12763 2415 12865 2441
rect 12985 2441 13087 2535
tri 13087 2441 13185 2539 sw
tri 13185 2441 13283 2539 ne
rect 13283 2535 13637 2539
rect 13283 2441 13415 2535
rect 12985 2415 13185 2441
rect 12763 2411 13185 2415
tri 13185 2411 13215 2441 sw
tri 13283 2411 13313 2441 ne
rect 13313 2415 13415 2441
rect 13535 2441 13637 2535
tri 13637 2441 13735 2539 sw
tri 13735 2441 13833 2539 ne
rect 13833 2535 14187 2539
rect 13833 2441 13965 2535
rect 13535 2415 13735 2441
rect 13313 2411 13735 2415
tri 13735 2411 13765 2441 sw
tri 13833 2411 13863 2441 ne
rect 13863 2415 13965 2441
rect 14085 2441 14187 2535
tri 14187 2441 14285 2539 sw
tri 14285 2441 14383 2539 ne
rect 14383 2535 14737 2539
rect 14383 2441 14515 2535
rect 14085 2415 14285 2441
rect 13863 2411 14285 2415
tri 14285 2411 14315 2441 sw
tri 14383 2411 14413 2441 ne
rect 14413 2415 14515 2441
rect 14635 2441 14737 2535
tri 14737 2441 14835 2539 sw
tri 14835 2441 14933 2539 ne
rect 14933 2535 15287 2539
rect 14933 2441 15065 2535
rect 14635 2415 14835 2441
rect 14413 2411 14835 2415
tri 14835 2411 14865 2441 sw
tri 14933 2411 14963 2441 ne
rect 14963 2415 15065 2441
rect 15185 2441 15287 2535
tri 15287 2441 15385 2539 sw
tri 15385 2441 15483 2539 ne
rect 15483 2535 15837 2539
rect 15483 2441 15615 2535
rect 15185 2415 15385 2441
rect 14963 2411 15385 2415
tri 15385 2411 15415 2441 sw
tri 15483 2411 15513 2441 ne
rect 15513 2415 15615 2441
rect 15735 2441 15837 2535
tri 15837 2441 15935 2539 sw
tri 15935 2441 16033 2539 ne
rect 16033 2535 16387 2539
rect 16033 2441 16165 2535
rect 15735 2415 15935 2441
rect 15513 2411 15935 2415
tri 15935 2411 15965 2441 sw
tri 16033 2411 16063 2441 ne
rect 16063 2415 16165 2441
rect 16285 2441 16387 2535
tri 16387 2441 16485 2539 sw
tri 16485 2441 16583 2539 ne
rect 16583 2535 16937 2539
rect 16583 2441 16715 2535
rect 16285 2415 16485 2441
rect 16063 2411 16485 2415
tri 16485 2411 16515 2441 sw
tri 16583 2411 16613 2441 ne
rect 16613 2415 16715 2441
rect 16835 2441 16937 2535
tri 16937 2441 17035 2539 sw
tri 17035 2441 17133 2539 ne
rect 17133 2535 17487 2539
rect 17133 2441 17265 2535
rect 16835 2415 17035 2441
rect 16613 2411 17035 2415
tri 17035 2411 17065 2441 sw
tri 17133 2411 17163 2441 ne
rect 17163 2415 17265 2441
rect 17385 2441 17487 2535
tri 17487 2441 17585 2539 sw
tri 17585 2441 17683 2539 ne
rect 17683 2535 18037 2539
rect 17683 2441 17815 2535
rect 17385 2415 17585 2441
rect 17163 2411 17585 2415
tri 17585 2411 17615 2441 sw
tri 17683 2411 17713 2441 ne
rect 17713 2415 17815 2441
rect 17935 2441 18037 2535
tri 18037 2441 18135 2539 sw
tri 18135 2441 18233 2539 ne
rect 18233 2535 18587 2539
rect 18233 2441 18365 2535
rect 17935 2415 18135 2441
rect 17713 2411 18135 2415
tri 18135 2411 18165 2441 sw
tri 18233 2411 18263 2441 ne
rect 18263 2415 18365 2441
rect 18485 2441 18587 2535
tri 18587 2441 18685 2539 sw
tri 18685 2441 18783 2539 ne
rect 18783 2535 19137 2539
rect 18783 2441 18915 2535
rect 18485 2415 18685 2441
rect 18263 2411 18685 2415
tri 18685 2411 18715 2441 sw
tri 18783 2411 18813 2441 ne
rect 18813 2415 18915 2441
rect 19035 2441 19137 2535
tri 19137 2441 19235 2539 sw
tri 19235 2441 19333 2539 ne
rect 19333 2535 20300 2539
rect 19333 2441 19465 2535
rect 19035 2415 19235 2441
rect 18813 2411 19235 2415
tri 19235 2411 19265 2441 sw
tri 19333 2411 19363 2441 ne
rect 19363 2415 19465 2441
rect 19585 2415 20300 2535
rect 19363 2411 20300 2415
tri 113 2313 211 2411 ne
rect 211 2313 565 2411
tri 565 2313 663 2411 sw
tri 663 2313 761 2411 ne
rect 761 2313 1115 2411
tri 1115 2313 1213 2411 sw
tri 1213 2313 1311 2411 ne
rect 1311 2313 1665 2411
tri 1665 2313 1763 2411 sw
tri 1763 2313 1861 2411 ne
rect 1861 2313 2215 2411
tri 2215 2313 2313 2411 sw
tri 2313 2313 2411 2411 ne
rect 2411 2313 2765 2411
tri 2765 2313 2863 2411 sw
tri 2863 2313 2961 2411 ne
rect 2961 2313 3315 2411
tri 3315 2313 3413 2411 sw
tri 3413 2313 3511 2411 ne
rect 3511 2313 3865 2411
tri 3865 2313 3963 2411 sw
tri 3963 2313 4061 2411 ne
rect 4061 2313 4415 2411
tri 4415 2313 4513 2411 sw
tri 4513 2313 4611 2411 ne
rect 4611 2313 4965 2411
tri 4965 2313 5063 2411 sw
tri 5063 2313 5161 2411 ne
rect 5161 2313 5515 2411
tri 5515 2313 5613 2411 sw
tri 5613 2313 5711 2411 ne
rect 5711 2313 6065 2411
tri 6065 2313 6163 2411 sw
tri 6163 2313 6261 2411 ne
rect 6261 2313 6615 2411
tri 6615 2313 6713 2411 sw
tri 6713 2313 6811 2411 ne
rect 6811 2313 7165 2411
tri 7165 2313 7263 2411 sw
tri 7263 2313 7361 2411 ne
rect 7361 2313 7715 2411
tri 7715 2313 7813 2411 sw
tri 7813 2313 7911 2411 ne
rect 7911 2313 8265 2411
tri 8265 2313 8363 2411 sw
tri 8363 2313 8461 2411 ne
rect 8461 2313 8815 2411
tri 8815 2313 8913 2411 sw
tri 8913 2313 9011 2411 ne
rect 9011 2313 9365 2411
tri 9365 2313 9463 2411 sw
tri 9463 2313 9561 2411 ne
rect 9561 2313 9915 2411
tri 9915 2313 10013 2411 sw
tri 10013 2313 10111 2411 ne
rect 10111 2313 10465 2411
tri 10465 2313 10563 2411 sw
tri 10563 2313 10661 2411 ne
rect 10661 2313 11015 2411
tri 11015 2313 11113 2411 sw
tri 11113 2313 11211 2411 ne
rect 11211 2313 11565 2411
tri 11565 2313 11663 2411 sw
tri 11663 2313 11761 2411 ne
rect 11761 2313 12115 2411
tri 12115 2313 12213 2411 sw
tri 12213 2313 12311 2411 ne
rect 12311 2313 12665 2411
tri 12665 2313 12763 2411 sw
tri 12763 2313 12861 2411 ne
rect 12861 2313 13215 2411
tri 13215 2313 13313 2411 sw
tri 13313 2313 13411 2411 ne
rect 13411 2313 13765 2411
tri 13765 2313 13863 2411 sw
tri 13863 2313 13961 2411 ne
rect 13961 2313 14315 2411
tri 14315 2313 14413 2411 sw
tri 14413 2313 14511 2411 ne
rect 14511 2313 14865 2411
tri 14865 2313 14963 2411 sw
tri 14963 2313 15061 2411 ne
rect 15061 2313 15415 2411
tri 15415 2313 15513 2411 sw
tri 15513 2313 15611 2411 ne
rect 15611 2313 15965 2411
tri 15965 2313 16063 2411 sw
tri 16063 2313 16161 2411 ne
rect 16161 2313 16515 2411
tri 16515 2313 16613 2411 sw
tri 16613 2313 16711 2411 ne
rect 16711 2313 17065 2411
tri 17065 2313 17163 2411 sw
tri 17163 2313 17261 2411 ne
rect 17261 2313 17615 2411
tri 17615 2313 17713 2411 sw
tri 17713 2313 17811 2411 ne
rect 17811 2313 18165 2411
tri 18165 2313 18263 2411 sw
tri 18263 2313 18361 2411 ne
rect 18361 2313 18715 2411
tri 18715 2313 18813 2411 sw
tri 18813 2313 18911 2411 ne
rect 18911 2313 19265 2411
tri 19265 2313 19363 2411 sw
tri 19363 2313 19461 2411 ne
rect 19461 2313 20300 2411
rect -2000 2283 113 2313
tri 113 2283 143 2313 sw
tri 211 2283 241 2313 ne
rect 241 2283 663 2313
tri 663 2283 693 2313 sw
tri 761 2283 791 2313 ne
rect 791 2283 1213 2313
tri 1213 2283 1243 2313 sw
tri 1311 2283 1341 2313 ne
rect 1341 2283 1763 2313
tri 1763 2283 1793 2313 sw
tri 1861 2283 1891 2313 ne
rect 1891 2283 2313 2313
tri 2313 2283 2343 2313 sw
tri 2411 2283 2441 2313 ne
rect 2441 2283 2863 2313
tri 2863 2283 2893 2313 sw
tri 2961 2283 2991 2313 ne
rect 2991 2283 3413 2313
tri 3413 2283 3443 2313 sw
tri 3511 2283 3541 2313 ne
rect 3541 2283 3963 2313
tri 3963 2283 3993 2313 sw
tri 4061 2283 4091 2313 ne
rect 4091 2283 4513 2313
tri 4513 2283 4543 2313 sw
tri 4611 2283 4641 2313 ne
rect 4641 2283 5063 2313
tri 5063 2283 5093 2313 sw
tri 5161 2283 5191 2313 ne
rect 5191 2283 5613 2313
tri 5613 2283 5643 2313 sw
tri 5711 2283 5741 2313 ne
rect 5741 2283 6163 2313
tri 6163 2283 6193 2313 sw
tri 6261 2283 6291 2313 ne
rect 6291 2283 6713 2313
tri 6713 2283 6743 2313 sw
tri 6811 2283 6841 2313 ne
rect 6841 2283 7263 2313
tri 7263 2283 7293 2313 sw
tri 7361 2283 7391 2313 ne
rect 7391 2283 7813 2313
tri 7813 2283 7843 2313 sw
tri 7911 2283 7941 2313 ne
rect 7941 2283 8363 2313
tri 8363 2283 8393 2313 sw
tri 8461 2283 8491 2313 ne
rect 8491 2283 8913 2313
tri 8913 2283 8943 2313 sw
tri 9011 2283 9041 2313 ne
rect 9041 2283 9463 2313
tri 9463 2283 9493 2313 sw
tri 9561 2283 9591 2313 ne
rect 9591 2283 10013 2313
tri 10013 2283 10043 2313 sw
tri 10111 2283 10141 2313 ne
rect 10141 2283 10563 2313
tri 10563 2283 10593 2313 sw
tri 10661 2283 10691 2313 ne
rect 10691 2283 11113 2313
tri 11113 2283 11143 2313 sw
tri 11211 2283 11241 2313 ne
rect 11241 2283 11663 2313
tri 11663 2283 11693 2313 sw
tri 11761 2283 11791 2313 ne
rect 11791 2283 12213 2313
tri 12213 2283 12243 2313 sw
tri 12311 2283 12341 2313 ne
rect 12341 2283 12763 2313
tri 12763 2283 12793 2313 sw
tri 12861 2283 12891 2313 ne
rect 12891 2283 13313 2313
tri 13313 2283 13343 2313 sw
tri 13411 2283 13441 2313 ne
rect 13441 2283 13863 2313
tri 13863 2283 13893 2313 sw
tri 13961 2283 13991 2313 ne
rect 13991 2283 14413 2313
tri 14413 2283 14443 2313 sw
tri 14511 2283 14541 2313 ne
rect 14541 2283 14963 2313
tri 14963 2283 14993 2313 sw
tri 15061 2283 15091 2313 ne
rect 15091 2283 15513 2313
tri 15513 2283 15543 2313 sw
tri 15611 2283 15641 2313 ne
rect 15641 2283 16063 2313
tri 16063 2283 16093 2313 sw
tri 16161 2283 16191 2313 ne
rect 16191 2283 16613 2313
tri 16613 2283 16643 2313 sw
tri 16711 2283 16741 2313 ne
rect 16741 2283 17163 2313
tri 17163 2283 17193 2313 sw
tri 17261 2283 17291 2313 ne
rect 17291 2283 17713 2313
tri 17713 2283 17743 2313 sw
tri 17811 2283 17841 2313 ne
rect 17841 2283 18263 2313
tri 18263 2283 18293 2313 sw
tri 18361 2283 18391 2313 ne
rect 18391 2283 18813 2313
tri 18813 2283 18843 2313 sw
tri 18911 2283 18941 2313 ne
rect 18941 2283 19363 2313
tri 19363 2283 19393 2313 sw
tri 19461 2283 19491 2313 ne
rect 19491 2283 20300 2313
rect -2000 2185 143 2283
tri 143 2185 241 2283 sw
tri 241 2185 339 2283 ne
rect 339 2185 693 2283
tri 693 2185 791 2283 sw
tri 791 2185 889 2283 ne
rect 889 2185 1243 2283
tri 1243 2185 1341 2283 sw
tri 1341 2185 1439 2283 ne
rect 1439 2185 1793 2283
tri 1793 2185 1891 2283 sw
tri 1891 2185 1989 2283 ne
rect 1989 2185 2343 2283
tri 2343 2185 2441 2283 sw
tri 2441 2185 2539 2283 ne
rect 2539 2185 2893 2283
tri 2893 2185 2991 2283 sw
tri 2991 2185 3089 2283 ne
rect 3089 2185 3443 2283
tri 3443 2185 3541 2283 sw
tri 3541 2185 3639 2283 ne
rect 3639 2185 3993 2283
tri 3993 2185 4091 2283 sw
tri 4091 2185 4189 2283 ne
rect 4189 2185 4543 2283
tri 4543 2185 4641 2283 sw
tri 4641 2185 4739 2283 ne
rect 4739 2185 5093 2283
tri 5093 2185 5191 2283 sw
tri 5191 2185 5289 2283 ne
rect 5289 2185 5643 2283
tri 5643 2185 5741 2283 sw
tri 5741 2185 5839 2283 ne
rect 5839 2185 6193 2283
tri 6193 2185 6291 2283 sw
tri 6291 2185 6389 2283 ne
rect 6389 2185 6743 2283
tri 6743 2185 6841 2283 sw
tri 6841 2185 6939 2283 ne
rect 6939 2185 7293 2283
tri 7293 2185 7391 2283 sw
tri 7391 2185 7489 2283 ne
rect 7489 2185 7843 2283
tri 7843 2185 7941 2283 sw
tri 7941 2185 8039 2283 ne
rect 8039 2185 8393 2283
tri 8393 2185 8491 2283 sw
tri 8491 2185 8589 2283 ne
rect 8589 2185 8943 2283
tri 8943 2185 9041 2283 sw
tri 9041 2185 9139 2283 ne
rect 9139 2185 9493 2283
tri 9493 2185 9591 2283 sw
tri 9591 2185 9689 2283 ne
rect 9689 2185 10043 2283
tri 10043 2185 10141 2283 sw
tri 10141 2185 10239 2283 ne
rect 10239 2185 10593 2283
tri 10593 2185 10691 2283 sw
tri 10691 2185 10789 2283 ne
rect 10789 2185 11143 2283
tri 11143 2185 11241 2283 sw
tri 11241 2185 11339 2283 ne
rect 11339 2185 11693 2283
tri 11693 2185 11791 2283 sw
tri 11791 2185 11889 2283 ne
rect 11889 2185 12243 2283
tri 12243 2185 12341 2283 sw
tri 12341 2185 12439 2283 ne
rect 12439 2185 12793 2283
tri 12793 2185 12891 2283 sw
tri 12891 2185 12989 2283 ne
rect 12989 2185 13343 2283
tri 13343 2185 13441 2283 sw
tri 13441 2185 13539 2283 ne
rect 13539 2185 13893 2283
tri 13893 2185 13991 2283 sw
tri 13991 2185 14089 2283 ne
rect 14089 2185 14443 2283
tri 14443 2185 14541 2283 sw
tri 14541 2185 14639 2283 ne
rect 14639 2185 14993 2283
tri 14993 2185 15091 2283 sw
tri 15091 2185 15189 2283 ne
rect 15189 2185 15543 2283
tri 15543 2185 15641 2283 sw
tri 15641 2185 15739 2283 ne
rect 15739 2185 16093 2283
tri 16093 2185 16191 2283 sw
tri 16191 2185 16289 2283 ne
rect 16289 2185 16643 2283
tri 16643 2185 16741 2283 sw
tri 16741 2185 16839 2283 ne
rect 16839 2185 17193 2283
tri 17193 2185 17291 2283 sw
tri 17291 2185 17389 2283 ne
rect 17389 2185 17743 2283
tri 17743 2185 17841 2283 sw
tri 17841 2185 17939 2283 ne
rect 17939 2185 18293 2283
tri 18293 2185 18391 2283 sw
tri 18391 2185 18489 2283 ne
rect 18489 2185 18843 2283
tri 18843 2185 18941 2283 sw
tri 18941 2185 19039 2283 ne
rect 19039 2185 19393 2283
tri 19393 2185 19491 2283 sw
tri 19491 2185 19589 2283 ne
rect 19589 2185 20300 2283
rect -2000 2087 241 2185
tri 241 2087 339 2185 sw
tri 339 2087 437 2185 ne
rect 437 2087 791 2185
tri 791 2087 889 2185 sw
tri 889 2087 987 2185 ne
rect 987 2087 1341 2185
tri 1341 2087 1439 2185 sw
tri 1439 2087 1537 2185 ne
rect 1537 2087 1891 2185
tri 1891 2087 1989 2185 sw
tri 1989 2087 2087 2185 ne
rect 2087 2087 2441 2185
tri 2441 2087 2539 2185 sw
tri 2539 2087 2637 2185 ne
rect 2637 2087 2991 2185
tri 2991 2087 3089 2185 sw
tri 3089 2087 3187 2185 ne
rect 3187 2087 3541 2185
tri 3541 2087 3639 2185 sw
tri 3639 2087 3737 2185 ne
rect 3737 2087 4091 2185
tri 4091 2087 4189 2185 sw
tri 4189 2087 4287 2185 ne
rect 4287 2087 4641 2185
tri 4641 2087 4739 2185 sw
tri 4739 2087 4837 2185 ne
rect 4837 2087 5191 2185
tri 5191 2087 5289 2185 sw
tri 5289 2087 5387 2185 ne
rect 5387 2087 5741 2185
tri 5741 2087 5839 2185 sw
tri 5839 2087 5937 2185 ne
rect 5937 2087 6291 2185
tri 6291 2087 6389 2185 sw
tri 6389 2087 6487 2185 ne
rect 6487 2087 6841 2185
tri 6841 2087 6939 2185 sw
tri 6939 2087 7037 2185 ne
rect 7037 2087 7391 2185
tri 7391 2087 7489 2185 sw
tri 7489 2087 7587 2185 ne
rect 7587 2087 7941 2185
tri 7941 2087 8039 2185 sw
tri 8039 2087 8137 2185 ne
rect 8137 2087 8491 2185
tri 8491 2087 8589 2185 sw
tri 8589 2087 8687 2185 ne
rect 8687 2087 9041 2185
tri 9041 2087 9139 2185 sw
tri 9139 2087 9237 2185 ne
rect 9237 2087 9591 2185
tri 9591 2087 9689 2185 sw
tri 9689 2087 9787 2185 ne
rect 9787 2087 10141 2185
tri 10141 2087 10239 2185 sw
tri 10239 2087 10337 2185 ne
rect 10337 2087 10691 2185
tri 10691 2087 10789 2185 sw
tri 10789 2087 10887 2185 ne
rect 10887 2087 11241 2185
tri 11241 2087 11339 2185 sw
tri 11339 2087 11437 2185 ne
rect 11437 2087 11791 2185
tri 11791 2087 11889 2185 sw
tri 11889 2087 11987 2185 ne
rect 11987 2087 12341 2185
tri 12341 2087 12439 2185 sw
tri 12439 2087 12537 2185 ne
rect 12537 2087 12891 2185
tri 12891 2087 12989 2185 sw
tri 12989 2087 13087 2185 ne
rect 13087 2087 13441 2185
tri 13441 2087 13539 2185 sw
tri 13539 2087 13637 2185 ne
rect 13637 2087 13991 2185
tri 13991 2087 14089 2185 sw
tri 14089 2087 14187 2185 ne
rect 14187 2087 14541 2185
tri 14541 2087 14639 2185 sw
tri 14639 2087 14737 2185 ne
rect 14737 2087 15091 2185
tri 15091 2087 15189 2185 sw
tri 15189 2087 15287 2185 ne
rect 15287 2087 15641 2185
tri 15641 2087 15739 2185 sw
tri 15739 2087 15837 2185 ne
rect 15837 2087 16191 2185
tri 16191 2087 16289 2185 sw
tri 16289 2087 16387 2185 ne
rect 16387 2087 16741 2185
tri 16741 2087 16839 2185 sw
tri 16839 2087 16937 2185 ne
rect 16937 2087 17291 2185
tri 17291 2087 17389 2185 sw
tri 17389 2087 17487 2185 ne
rect 17487 2087 17841 2185
tri 17841 2087 17939 2185 sw
tri 17939 2087 18037 2185 ne
rect 18037 2087 18391 2185
tri 18391 2087 18489 2185 sw
tri 18489 2087 18587 2185 ne
rect 18587 2087 18941 2185
tri 18941 2087 19039 2185 sw
tri 19039 2087 19137 2185 ne
rect 19137 2087 19491 2185
tri 19491 2087 19589 2185 sw
tri 19589 2087 19687 2185 ne
rect 19687 2087 20300 2185
rect -2000 1989 339 2087
tri 339 1989 437 2087 sw
tri 437 1989 535 2087 ne
rect 535 1989 889 2087
tri 889 1989 987 2087 sw
tri 987 1989 1085 2087 ne
rect 1085 1989 1439 2087
tri 1439 1989 1537 2087 sw
tri 1537 1989 1635 2087 ne
rect 1635 1989 1989 2087
tri 1989 1989 2087 2087 sw
tri 2087 1989 2185 2087 ne
rect 2185 1989 2539 2087
tri 2539 1989 2637 2087 sw
tri 2637 1989 2735 2087 ne
rect 2735 1989 3089 2087
tri 3089 1989 3187 2087 sw
tri 3187 1989 3285 2087 ne
rect 3285 1989 3639 2087
tri 3639 1989 3737 2087 sw
tri 3737 1989 3835 2087 ne
rect 3835 1989 4189 2087
tri 4189 1989 4287 2087 sw
tri 4287 1989 4385 2087 ne
rect 4385 1989 4739 2087
tri 4739 1989 4837 2087 sw
tri 4837 1989 4935 2087 ne
rect 4935 1989 5289 2087
tri 5289 1989 5387 2087 sw
tri 5387 1989 5485 2087 ne
rect 5485 1989 5839 2087
tri 5839 1989 5937 2087 sw
tri 5937 1989 6035 2087 ne
rect 6035 1989 6389 2087
tri 6389 1989 6487 2087 sw
tri 6487 1989 6585 2087 ne
rect 6585 1989 6939 2087
tri 6939 1989 7037 2087 sw
tri 7037 1989 7135 2087 ne
rect 7135 1989 7489 2087
tri 7489 1989 7587 2087 sw
tri 7587 1989 7685 2087 ne
rect 7685 1989 8039 2087
tri 8039 1989 8137 2087 sw
tri 8137 1989 8235 2087 ne
rect 8235 1989 8589 2087
tri 8589 1989 8687 2087 sw
tri 8687 1989 8785 2087 ne
rect 8785 1989 9139 2087
tri 9139 1989 9237 2087 sw
tri 9237 1989 9335 2087 ne
rect 9335 1989 9689 2087
tri 9689 1989 9787 2087 sw
tri 9787 1989 9885 2087 ne
rect 9885 1989 10239 2087
tri 10239 1989 10337 2087 sw
tri 10337 1989 10435 2087 ne
rect 10435 1989 10789 2087
tri 10789 1989 10887 2087 sw
tri 10887 1989 10985 2087 ne
rect 10985 1989 11339 2087
tri 11339 1989 11437 2087 sw
tri 11437 1989 11535 2087 ne
rect 11535 1989 11889 2087
tri 11889 1989 11987 2087 sw
tri 11987 1989 12085 2087 ne
rect 12085 1989 12439 2087
tri 12439 1989 12537 2087 sw
tri 12537 1989 12635 2087 ne
rect 12635 1989 12989 2087
tri 12989 1989 13087 2087 sw
tri 13087 1989 13185 2087 ne
rect 13185 1989 13539 2087
tri 13539 1989 13637 2087 sw
tri 13637 1989 13735 2087 ne
rect 13735 1989 14089 2087
tri 14089 1989 14187 2087 sw
tri 14187 1989 14285 2087 ne
rect 14285 1989 14639 2087
tri 14639 1989 14737 2087 sw
tri 14737 1989 14835 2087 ne
rect 14835 1989 15189 2087
tri 15189 1989 15287 2087 sw
tri 15287 1989 15385 2087 ne
rect 15385 1989 15739 2087
tri 15739 1989 15837 2087 sw
tri 15837 1989 15935 2087 ne
rect 15935 1989 16289 2087
tri 16289 1989 16387 2087 sw
tri 16387 1989 16485 2087 ne
rect 16485 1989 16839 2087
tri 16839 1989 16937 2087 sw
tri 16937 1989 17035 2087 ne
rect 17035 1989 17389 2087
tri 17389 1989 17487 2087 sw
tri 17487 1989 17585 2087 ne
rect 17585 1989 17939 2087
tri 17939 1989 18037 2087 sw
tri 18037 1989 18135 2087 ne
rect 18135 1989 18489 2087
tri 18489 1989 18587 2087 sw
tri 18587 1989 18685 2087 ne
rect 18685 1989 19039 2087
tri 19039 1989 19137 2087 sw
tri 19137 1989 19235 2087 ne
rect 19235 1989 19589 2087
tri 19589 1989 19687 2087 sw
rect 20800 1989 21800 2637
rect -2000 1985 437 1989
rect -2000 1865 215 1985
rect 335 1891 437 1985
tri 437 1891 535 1989 sw
tri 535 1891 633 1989 ne
rect 633 1985 987 1989
rect 633 1891 765 1985
rect 335 1865 535 1891
rect -2000 1861 535 1865
rect -2000 1650 -1000 1861
tri 113 1763 211 1861 ne
rect 211 1813 535 1861
tri 535 1813 613 1891 sw
tri 633 1813 711 1891 ne
rect 711 1865 765 1891
rect 885 1891 987 1985
tri 987 1891 1085 1989 sw
tri 1085 1891 1183 1989 ne
rect 1183 1985 1537 1989
rect 1183 1891 1315 1985
rect 885 1865 1085 1891
rect 711 1813 1085 1865
tri 1085 1813 1163 1891 sw
tri 1183 1813 1261 1891 ne
rect 1261 1865 1315 1891
rect 1435 1891 1537 1985
tri 1537 1891 1635 1989 sw
tri 1635 1891 1733 1989 ne
rect 1733 1985 2087 1989
rect 1733 1891 1865 1985
rect 1435 1865 1635 1891
rect 1261 1813 1635 1865
tri 1635 1813 1713 1891 sw
tri 1733 1813 1811 1891 ne
rect 1811 1865 1865 1891
rect 1985 1891 2087 1985
tri 2087 1891 2185 1989 sw
tri 2185 1891 2283 1989 ne
rect 2283 1985 2637 1989
rect 2283 1891 2415 1985
rect 1985 1865 2185 1891
rect 1811 1813 2185 1865
tri 2185 1813 2263 1891 sw
tri 2283 1813 2361 1891 ne
rect 2361 1865 2415 1891
rect 2535 1891 2637 1985
tri 2637 1891 2735 1989 sw
tri 2735 1891 2833 1989 ne
rect 2833 1985 3187 1989
rect 2833 1891 2965 1985
rect 2535 1865 2735 1891
rect 2361 1813 2735 1865
tri 2735 1813 2813 1891 sw
tri 2833 1813 2911 1891 ne
rect 2911 1865 2965 1891
rect 3085 1891 3187 1985
tri 3187 1891 3285 1989 sw
tri 3285 1891 3383 1989 ne
rect 3383 1985 3737 1989
rect 3383 1891 3515 1985
rect 3085 1865 3285 1891
rect 2911 1813 3285 1865
tri 3285 1813 3363 1891 sw
tri 3383 1813 3461 1891 ne
rect 3461 1865 3515 1891
rect 3635 1891 3737 1985
tri 3737 1891 3835 1989 sw
tri 3835 1891 3933 1989 ne
rect 3933 1985 4287 1989
rect 3933 1891 4065 1985
rect 3635 1865 3835 1891
rect 3461 1813 3835 1865
tri 3835 1813 3913 1891 sw
tri 3933 1813 4011 1891 ne
rect 4011 1865 4065 1891
rect 4185 1891 4287 1985
tri 4287 1891 4385 1989 sw
tri 4385 1891 4483 1989 ne
rect 4483 1985 4837 1989
rect 4483 1891 4615 1985
rect 4185 1865 4385 1891
rect 4011 1813 4385 1865
tri 4385 1813 4463 1891 sw
tri 4483 1813 4561 1891 ne
rect 4561 1865 4615 1891
rect 4735 1891 4837 1985
tri 4837 1891 4935 1989 sw
tri 4935 1891 5033 1989 ne
rect 5033 1985 5387 1989
rect 5033 1891 5165 1985
rect 4735 1865 4935 1891
rect 4561 1813 4935 1865
tri 4935 1813 5013 1891 sw
tri 5033 1813 5111 1891 ne
rect 5111 1865 5165 1891
rect 5285 1891 5387 1985
tri 5387 1891 5485 1989 sw
tri 5485 1891 5583 1989 ne
rect 5583 1985 5937 1989
rect 5583 1891 5715 1985
rect 5285 1865 5485 1891
rect 5111 1813 5485 1865
tri 5485 1813 5563 1891 sw
tri 5583 1813 5661 1891 ne
rect 5661 1865 5715 1891
rect 5835 1891 5937 1985
tri 5937 1891 6035 1989 sw
tri 6035 1891 6133 1989 ne
rect 6133 1985 6487 1989
rect 6133 1891 6265 1985
rect 5835 1865 6035 1891
rect 5661 1813 6035 1865
tri 6035 1813 6113 1891 sw
tri 6133 1813 6211 1891 ne
rect 6211 1865 6265 1891
rect 6385 1891 6487 1985
tri 6487 1891 6585 1989 sw
tri 6585 1891 6683 1989 ne
rect 6683 1985 7037 1989
rect 6683 1891 6815 1985
rect 6385 1865 6585 1891
rect 6211 1813 6585 1865
tri 6585 1813 6663 1891 sw
tri 6683 1813 6761 1891 ne
rect 6761 1865 6815 1891
rect 6935 1891 7037 1985
tri 7037 1891 7135 1989 sw
tri 7135 1891 7233 1989 ne
rect 7233 1985 7587 1989
rect 7233 1891 7365 1985
rect 6935 1865 7135 1891
rect 6761 1813 7135 1865
tri 7135 1813 7213 1891 sw
tri 7233 1813 7311 1891 ne
rect 7311 1865 7365 1891
rect 7485 1891 7587 1985
tri 7587 1891 7685 1989 sw
tri 7685 1891 7783 1989 ne
rect 7783 1985 8137 1989
rect 7783 1891 7915 1985
rect 7485 1865 7685 1891
rect 7311 1813 7685 1865
tri 7685 1813 7763 1891 sw
tri 7783 1813 7861 1891 ne
rect 7861 1865 7915 1891
rect 8035 1891 8137 1985
tri 8137 1891 8235 1989 sw
tri 8235 1891 8333 1989 ne
rect 8333 1985 8687 1989
rect 8333 1891 8465 1985
rect 8035 1865 8235 1891
rect 7861 1813 8235 1865
tri 8235 1813 8313 1891 sw
tri 8333 1813 8411 1891 ne
rect 8411 1865 8465 1891
rect 8585 1891 8687 1985
tri 8687 1891 8785 1989 sw
tri 8785 1891 8883 1989 ne
rect 8883 1985 9237 1989
rect 8883 1891 9015 1985
rect 8585 1865 8785 1891
rect 8411 1813 8785 1865
tri 8785 1813 8863 1891 sw
tri 8883 1813 8961 1891 ne
rect 8961 1865 9015 1891
rect 9135 1891 9237 1985
tri 9237 1891 9335 1989 sw
tri 9335 1891 9433 1989 ne
rect 9433 1985 9787 1989
rect 9433 1891 9565 1985
rect 9135 1865 9335 1891
rect 8961 1813 9335 1865
tri 9335 1813 9413 1891 sw
tri 9433 1813 9511 1891 ne
rect 9511 1865 9565 1891
rect 9685 1891 9787 1985
tri 9787 1891 9885 1989 sw
tri 9885 1891 9983 1989 ne
rect 9983 1985 10337 1989
rect 9983 1891 10115 1985
rect 9685 1865 9885 1891
rect 9511 1813 9885 1865
tri 9885 1813 9963 1891 sw
tri 9983 1813 10061 1891 ne
rect 10061 1865 10115 1891
rect 10235 1891 10337 1985
tri 10337 1891 10435 1989 sw
tri 10435 1891 10533 1989 ne
rect 10533 1985 10887 1989
rect 10533 1891 10665 1985
rect 10235 1865 10435 1891
rect 10061 1813 10435 1865
tri 10435 1813 10513 1891 sw
tri 10533 1813 10611 1891 ne
rect 10611 1865 10665 1891
rect 10785 1891 10887 1985
tri 10887 1891 10985 1989 sw
tri 10985 1891 11083 1989 ne
rect 11083 1985 11437 1989
rect 11083 1891 11215 1985
rect 10785 1865 10985 1891
rect 10611 1813 10985 1865
tri 10985 1813 11063 1891 sw
tri 11083 1813 11161 1891 ne
rect 11161 1865 11215 1891
rect 11335 1891 11437 1985
tri 11437 1891 11535 1989 sw
tri 11535 1891 11633 1989 ne
rect 11633 1985 11987 1989
rect 11633 1891 11765 1985
rect 11335 1865 11535 1891
rect 11161 1813 11535 1865
tri 11535 1813 11613 1891 sw
tri 11633 1813 11711 1891 ne
rect 11711 1865 11765 1891
rect 11885 1891 11987 1985
tri 11987 1891 12085 1989 sw
tri 12085 1891 12183 1989 ne
rect 12183 1985 12537 1989
rect 12183 1891 12315 1985
rect 11885 1865 12085 1891
rect 11711 1813 12085 1865
tri 12085 1813 12163 1891 sw
tri 12183 1813 12261 1891 ne
rect 12261 1865 12315 1891
rect 12435 1891 12537 1985
tri 12537 1891 12635 1989 sw
tri 12635 1891 12733 1989 ne
rect 12733 1985 13087 1989
rect 12733 1891 12865 1985
rect 12435 1865 12635 1891
rect 12261 1813 12635 1865
tri 12635 1813 12713 1891 sw
tri 12733 1813 12811 1891 ne
rect 12811 1865 12865 1891
rect 12985 1891 13087 1985
tri 13087 1891 13185 1989 sw
tri 13185 1891 13283 1989 ne
rect 13283 1985 13637 1989
rect 13283 1891 13415 1985
rect 12985 1865 13185 1891
rect 12811 1813 13185 1865
tri 13185 1813 13263 1891 sw
tri 13283 1813 13361 1891 ne
rect 13361 1865 13415 1891
rect 13535 1891 13637 1985
tri 13637 1891 13735 1989 sw
tri 13735 1891 13833 1989 ne
rect 13833 1985 14187 1989
rect 13833 1891 13965 1985
rect 13535 1865 13735 1891
rect 13361 1813 13735 1865
tri 13735 1813 13813 1891 sw
tri 13833 1813 13911 1891 ne
rect 13911 1865 13965 1891
rect 14085 1891 14187 1985
tri 14187 1891 14285 1989 sw
tri 14285 1891 14383 1989 ne
rect 14383 1985 14737 1989
rect 14383 1891 14515 1985
rect 14085 1865 14285 1891
rect 13911 1813 14285 1865
tri 14285 1813 14363 1891 sw
tri 14383 1813 14461 1891 ne
rect 14461 1865 14515 1891
rect 14635 1891 14737 1985
tri 14737 1891 14835 1989 sw
tri 14835 1891 14933 1989 ne
rect 14933 1985 15287 1989
rect 14933 1891 15065 1985
rect 14635 1865 14835 1891
rect 14461 1813 14835 1865
tri 14835 1813 14913 1891 sw
tri 14933 1813 15011 1891 ne
rect 15011 1865 15065 1891
rect 15185 1891 15287 1985
tri 15287 1891 15385 1989 sw
tri 15385 1891 15483 1989 ne
rect 15483 1985 15837 1989
rect 15483 1891 15615 1985
rect 15185 1865 15385 1891
rect 15011 1813 15385 1865
tri 15385 1813 15463 1891 sw
tri 15483 1813 15561 1891 ne
rect 15561 1865 15615 1891
rect 15735 1891 15837 1985
tri 15837 1891 15935 1989 sw
tri 15935 1891 16033 1989 ne
rect 16033 1985 16387 1989
rect 16033 1891 16165 1985
rect 15735 1865 15935 1891
rect 15561 1813 15935 1865
tri 15935 1813 16013 1891 sw
tri 16033 1813 16111 1891 ne
rect 16111 1865 16165 1891
rect 16285 1891 16387 1985
tri 16387 1891 16485 1989 sw
tri 16485 1891 16583 1989 ne
rect 16583 1985 16937 1989
rect 16583 1891 16715 1985
rect 16285 1865 16485 1891
rect 16111 1813 16485 1865
tri 16485 1813 16563 1891 sw
tri 16583 1813 16661 1891 ne
rect 16661 1865 16715 1891
rect 16835 1891 16937 1985
tri 16937 1891 17035 1989 sw
tri 17035 1891 17133 1989 ne
rect 17133 1985 17487 1989
rect 17133 1891 17265 1985
rect 16835 1865 17035 1891
rect 16661 1813 17035 1865
tri 17035 1813 17113 1891 sw
tri 17133 1813 17211 1891 ne
rect 17211 1865 17265 1891
rect 17385 1891 17487 1985
tri 17487 1891 17585 1989 sw
tri 17585 1891 17683 1989 ne
rect 17683 1985 18037 1989
rect 17683 1891 17815 1985
rect 17385 1865 17585 1891
rect 17211 1813 17585 1865
tri 17585 1813 17663 1891 sw
tri 17683 1813 17761 1891 ne
rect 17761 1865 17815 1891
rect 17935 1891 18037 1985
tri 18037 1891 18135 1989 sw
tri 18135 1891 18233 1989 ne
rect 18233 1985 18587 1989
rect 18233 1891 18365 1985
rect 17935 1865 18135 1891
rect 17761 1813 18135 1865
tri 18135 1813 18213 1891 sw
tri 18233 1813 18311 1891 ne
rect 18311 1865 18365 1891
rect 18485 1891 18587 1985
tri 18587 1891 18685 1989 sw
tri 18685 1891 18783 1989 ne
rect 18783 1985 19137 1989
rect 18783 1891 18915 1985
rect 18485 1865 18685 1891
rect 18311 1813 18685 1865
tri 18685 1813 18763 1891 sw
tri 18783 1813 18861 1891 ne
rect 18861 1865 18915 1891
rect 19035 1891 19137 1985
tri 19137 1891 19235 1989 sw
tri 19235 1891 19333 1989 ne
rect 19333 1985 21800 1989
rect 19333 1891 19465 1985
rect 19035 1865 19235 1891
rect 18861 1813 19235 1865
tri 19235 1813 19313 1891 sw
tri 19333 1813 19411 1891 ne
rect 19411 1865 19465 1891
rect 19585 1865 21800 1985
rect 19411 1813 21800 1865
rect 211 1763 613 1813
rect -500 1713 113 1763
tri 113 1713 163 1763 sw
tri 211 1713 261 1763 ne
rect 261 1733 613 1763
tri 613 1733 693 1813 sw
tri 711 1733 791 1813 ne
rect 791 1733 1163 1813
tri 1163 1733 1243 1813 sw
tri 1261 1733 1341 1813 ne
rect 1341 1733 1713 1813
tri 1713 1733 1793 1813 sw
tri 1811 1733 1891 1813 ne
rect 1891 1733 2263 1813
tri 2263 1733 2343 1813 sw
tri 2361 1733 2441 1813 ne
rect 2441 1733 2813 1813
tri 2813 1733 2893 1813 sw
tri 2911 1733 2991 1813 ne
rect 2991 1733 3363 1813
tri 3363 1733 3443 1813 sw
tri 3461 1733 3541 1813 ne
rect 3541 1733 3913 1813
tri 3913 1733 3993 1813 sw
tri 4011 1733 4091 1813 ne
rect 4091 1733 4463 1813
tri 4463 1733 4543 1813 sw
tri 4561 1733 4641 1813 ne
rect 4641 1733 5013 1813
tri 5013 1733 5093 1813 sw
tri 5111 1733 5191 1813 ne
rect 5191 1733 5563 1813
tri 5563 1733 5643 1813 sw
tri 5661 1733 5741 1813 ne
rect 5741 1733 6113 1813
tri 6113 1733 6193 1813 sw
tri 6211 1733 6291 1813 ne
rect 6291 1733 6663 1813
tri 6663 1733 6743 1813 sw
tri 6761 1733 6841 1813 ne
rect 6841 1733 7213 1813
tri 7213 1733 7293 1813 sw
tri 7311 1733 7391 1813 ne
rect 7391 1733 7763 1813
tri 7763 1733 7843 1813 sw
tri 7861 1733 7941 1813 ne
rect 7941 1733 8313 1813
tri 8313 1733 8393 1813 sw
tri 8411 1733 8491 1813 ne
rect 8491 1733 8863 1813
tri 8863 1733 8943 1813 sw
tri 8961 1733 9041 1813 ne
rect 9041 1733 9413 1813
tri 9413 1733 9493 1813 sw
tri 9511 1733 9591 1813 ne
rect 9591 1733 9963 1813
tri 9963 1733 10043 1813 sw
tri 10061 1733 10141 1813 ne
rect 10141 1733 10513 1813
tri 10513 1733 10593 1813 sw
tri 10611 1733 10691 1813 ne
rect 10691 1733 11063 1813
tri 11063 1733 11143 1813 sw
tri 11161 1733 11241 1813 ne
rect 11241 1733 11613 1813
tri 11613 1733 11693 1813 sw
tri 11711 1733 11791 1813 ne
rect 11791 1733 12163 1813
tri 12163 1733 12243 1813 sw
tri 12261 1733 12341 1813 ne
rect 12341 1733 12713 1813
tri 12713 1733 12793 1813 sw
tri 12811 1733 12891 1813 ne
rect 12891 1733 13263 1813
tri 13263 1733 13343 1813 sw
tri 13361 1733 13441 1813 ne
rect 13441 1733 13813 1813
tri 13813 1733 13893 1813 sw
tri 13911 1733 13991 1813 ne
rect 13991 1733 14363 1813
tri 14363 1733 14443 1813 sw
tri 14461 1733 14541 1813 ne
rect 14541 1733 14913 1813
tri 14913 1733 14993 1813 sw
tri 15011 1733 15091 1813 ne
rect 15091 1733 15463 1813
tri 15463 1733 15543 1813 sw
tri 15561 1733 15641 1813 ne
rect 15641 1733 16013 1813
tri 16013 1733 16093 1813 sw
tri 16111 1733 16191 1813 ne
rect 16191 1733 16563 1813
tri 16563 1733 16643 1813 sw
tri 16661 1733 16741 1813 ne
rect 16741 1733 17113 1813
tri 17113 1733 17193 1813 sw
tri 17211 1733 17291 1813 ne
rect 17291 1733 17663 1813
tri 17663 1733 17743 1813 sw
tri 17761 1733 17841 1813 ne
rect 17841 1733 18213 1813
tri 18213 1733 18293 1813 sw
tri 18311 1733 18391 1813 ne
rect 18391 1733 18763 1813
tri 18763 1733 18843 1813 sw
tri 18861 1733 18941 1813 ne
rect 18941 1733 19313 1813
tri 19313 1733 19393 1813 sw
tri 19411 1733 19491 1813 ne
rect 19491 1733 20100 1813
rect 261 1713 693 1733
rect -500 1635 163 1713
tri 163 1635 241 1713 sw
tri 261 1635 339 1713 ne
rect 339 1635 693 1713
tri 693 1635 791 1733 sw
tri 791 1635 889 1733 ne
rect 889 1635 1243 1733
tri 1243 1635 1341 1733 sw
tri 1341 1635 1439 1733 ne
rect 1439 1635 1793 1733
tri 1793 1635 1891 1733 sw
tri 1891 1635 1989 1733 ne
rect 1989 1635 2343 1733
tri 2343 1635 2441 1733 sw
tri 2441 1635 2539 1733 ne
rect 2539 1635 2893 1733
tri 2893 1635 2991 1733 sw
tri 2991 1635 3089 1733 ne
rect 3089 1635 3443 1733
tri 3443 1635 3541 1733 sw
tri 3541 1635 3639 1733 ne
rect 3639 1635 3993 1733
tri 3993 1635 4091 1733 sw
tri 4091 1635 4189 1733 ne
rect 4189 1635 4543 1733
tri 4543 1635 4641 1733 sw
tri 4641 1635 4739 1733 ne
rect 4739 1635 5093 1733
tri 5093 1635 5191 1733 sw
tri 5191 1635 5289 1733 ne
rect 5289 1635 5643 1733
tri 5643 1635 5741 1733 sw
tri 5741 1635 5839 1733 ne
rect 5839 1635 6193 1733
tri 6193 1635 6291 1733 sw
tri 6291 1635 6389 1733 ne
rect 6389 1635 6743 1733
tri 6743 1635 6841 1733 sw
tri 6841 1635 6939 1733 ne
rect 6939 1635 7293 1733
tri 7293 1635 7391 1733 sw
tri 7391 1635 7489 1733 ne
rect 7489 1635 7843 1733
tri 7843 1635 7941 1733 sw
tri 7941 1635 8039 1733 ne
rect 8039 1635 8393 1733
tri 8393 1635 8491 1733 sw
tri 8491 1635 8589 1733 ne
rect 8589 1635 8943 1733
tri 8943 1635 9041 1733 sw
tri 9041 1635 9139 1733 ne
rect 9139 1635 9493 1733
tri 9493 1635 9591 1733 sw
tri 9591 1635 9689 1733 ne
rect 9689 1635 10043 1733
tri 10043 1635 10141 1733 sw
tri 10141 1635 10239 1733 ne
rect 10239 1635 10593 1733
tri 10593 1635 10691 1733 sw
tri 10691 1635 10789 1733 ne
rect 10789 1635 11143 1733
tri 11143 1635 11241 1733 sw
tri 11241 1635 11339 1733 ne
rect 11339 1635 11693 1733
tri 11693 1635 11791 1733 sw
tri 11791 1635 11889 1733 ne
rect 11889 1635 12243 1733
tri 12243 1635 12341 1733 sw
tri 12341 1635 12439 1733 ne
rect 12439 1635 12793 1733
tri 12793 1635 12891 1733 sw
tri 12891 1635 12989 1733 ne
rect 12989 1635 13343 1733
tri 13343 1635 13441 1733 sw
tri 13441 1635 13539 1733 ne
rect 13539 1635 13893 1733
tri 13893 1635 13991 1733 sw
tri 13991 1635 14089 1733 ne
rect 14089 1635 14443 1733
tri 14443 1635 14541 1733 sw
tri 14541 1635 14639 1733 ne
rect 14639 1635 14993 1733
tri 14993 1635 15091 1733 sw
tri 15091 1635 15189 1733 ne
rect 15189 1635 15543 1733
tri 15543 1635 15641 1733 sw
tri 15641 1635 15739 1733 ne
rect 15739 1635 16093 1733
tri 16093 1635 16191 1733 sw
tri 16191 1635 16289 1733 ne
rect 16289 1635 16643 1733
tri 16643 1635 16741 1733 sw
tri 16741 1635 16839 1733 ne
rect 16839 1635 17193 1733
tri 17193 1635 17291 1733 sw
tri 17291 1635 17389 1733 ne
rect 17389 1635 17743 1733
tri 17743 1635 17841 1733 sw
tri 17841 1635 17939 1733 ne
rect 17939 1635 18293 1733
tri 18293 1635 18391 1733 sw
tri 18391 1635 18489 1733 ne
rect 18489 1635 18843 1733
tri 18843 1635 18941 1733 sw
tri 18941 1635 19039 1733 ne
rect 19039 1635 19393 1733
tri 19393 1635 19491 1733 sw
tri 19491 1635 19589 1733 ne
rect 19589 1713 20100 1733
rect 20200 1713 21800 1813
rect 19589 1635 21800 1713
rect -500 1587 241 1635
rect -500 1487 -400 1587
rect -300 1537 241 1587
tri 241 1537 339 1635 sw
tri 339 1537 437 1635 ne
rect 437 1537 791 1635
tri 791 1537 889 1635 sw
tri 889 1537 987 1635 ne
rect 987 1537 1341 1635
tri 1341 1537 1439 1635 sw
tri 1439 1537 1537 1635 ne
rect 1537 1537 1891 1635
tri 1891 1537 1989 1635 sw
tri 1989 1537 2087 1635 ne
rect 2087 1537 2441 1635
tri 2441 1537 2539 1635 sw
tri 2539 1537 2637 1635 ne
rect 2637 1537 2991 1635
tri 2991 1537 3089 1635 sw
tri 3089 1537 3187 1635 ne
rect 3187 1537 3541 1635
tri 3541 1537 3639 1635 sw
tri 3639 1537 3737 1635 ne
rect 3737 1537 4091 1635
tri 4091 1537 4189 1635 sw
tri 4189 1537 4287 1635 ne
rect 4287 1537 4641 1635
tri 4641 1537 4739 1635 sw
tri 4739 1537 4837 1635 ne
rect 4837 1537 5191 1635
tri 5191 1537 5289 1635 sw
tri 5289 1537 5387 1635 ne
rect 5387 1537 5741 1635
tri 5741 1537 5839 1635 sw
tri 5839 1537 5937 1635 ne
rect 5937 1537 6291 1635
tri 6291 1537 6389 1635 sw
tri 6389 1537 6487 1635 ne
rect 6487 1537 6841 1635
tri 6841 1537 6939 1635 sw
tri 6939 1537 7037 1635 ne
rect 7037 1537 7391 1635
tri 7391 1537 7489 1635 sw
tri 7489 1537 7587 1635 ne
rect 7587 1537 7941 1635
tri 7941 1537 8039 1635 sw
tri 8039 1537 8137 1635 ne
rect 8137 1537 8491 1635
tri 8491 1537 8589 1635 sw
tri 8589 1537 8687 1635 ne
rect 8687 1537 9041 1635
tri 9041 1537 9139 1635 sw
tri 9139 1537 9237 1635 ne
rect 9237 1537 9591 1635
tri 9591 1537 9689 1635 sw
tri 9689 1537 9787 1635 ne
rect 9787 1537 10141 1635
tri 10141 1537 10239 1635 sw
tri 10239 1537 10337 1635 ne
rect 10337 1537 10691 1635
tri 10691 1537 10789 1635 sw
tri 10789 1537 10887 1635 ne
rect 10887 1537 11241 1635
tri 11241 1537 11339 1635 sw
tri 11339 1537 11437 1635 ne
rect 11437 1537 11791 1635
tri 11791 1537 11889 1635 sw
tri 11889 1537 11987 1635 ne
rect 11987 1537 12341 1635
tri 12341 1537 12439 1635 sw
tri 12439 1537 12537 1635 ne
rect 12537 1537 12891 1635
tri 12891 1537 12989 1635 sw
tri 12989 1537 13087 1635 ne
rect 13087 1537 13441 1635
tri 13441 1537 13539 1635 sw
tri 13539 1537 13637 1635 ne
rect 13637 1537 13991 1635
tri 13991 1537 14089 1635 sw
tri 14089 1537 14187 1635 ne
rect 14187 1537 14541 1635
tri 14541 1537 14639 1635 sw
tri 14639 1537 14737 1635 ne
rect 14737 1537 15091 1635
tri 15091 1537 15189 1635 sw
tri 15189 1537 15287 1635 ne
rect 15287 1537 15641 1635
tri 15641 1537 15739 1635 sw
tri 15739 1537 15837 1635 ne
rect 15837 1537 16191 1635
tri 16191 1537 16289 1635 sw
tri 16289 1537 16387 1635 ne
rect 16387 1537 16741 1635
tri 16741 1537 16839 1635 sw
tri 16839 1537 16937 1635 ne
rect 16937 1537 17291 1635
tri 17291 1537 17389 1635 sw
tri 17389 1537 17487 1635 ne
rect 17487 1537 17841 1635
tri 17841 1537 17939 1635 sw
tri 17939 1537 18037 1635 ne
rect 18037 1537 18391 1635
tri 18391 1537 18489 1635 sw
tri 18489 1537 18587 1635 ne
rect 18587 1537 18941 1635
tri 18941 1537 19039 1635 sw
tri 19039 1537 19137 1635 ne
rect 19137 1537 19491 1635
tri 19491 1537 19589 1635 sw
tri 19589 1537 19687 1635 ne
rect 19687 1537 21800 1635
rect -300 1487 339 1537
rect -500 1439 339 1487
tri 339 1439 437 1537 sw
tri 437 1439 535 1537 ne
rect 535 1439 889 1537
tri 889 1439 987 1537 sw
tri 987 1439 1085 1537 ne
rect 1085 1439 1439 1537
tri 1439 1439 1537 1537 sw
tri 1537 1439 1635 1537 ne
rect 1635 1439 1989 1537
tri 1989 1439 2087 1537 sw
tri 2087 1439 2185 1537 ne
rect 2185 1439 2539 1537
tri 2539 1439 2637 1537 sw
tri 2637 1439 2735 1537 ne
rect 2735 1439 3089 1537
tri 3089 1439 3187 1537 sw
tri 3187 1439 3285 1537 ne
rect 3285 1439 3639 1537
tri 3639 1439 3737 1537 sw
tri 3737 1439 3835 1537 ne
rect 3835 1439 4189 1537
tri 4189 1439 4287 1537 sw
tri 4287 1439 4385 1537 ne
rect 4385 1439 4739 1537
tri 4739 1439 4837 1537 sw
tri 4837 1439 4935 1537 ne
rect 4935 1439 5289 1537
tri 5289 1439 5387 1537 sw
tri 5387 1439 5485 1537 ne
rect 5485 1439 5839 1537
tri 5839 1439 5937 1537 sw
tri 5937 1439 6035 1537 ne
rect 6035 1439 6389 1537
tri 6389 1439 6487 1537 sw
tri 6487 1439 6585 1537 ne
rect 6585 1439 6939 1537
tri 6939 1439 7037 1537 sw
tri 7037 1439 7135 1537 ne
rect 7135 1439 7489 1537
tri 7489 1439 7587 1537 sw
tri 7587 1439 7685 1537 ne
rect 7685 1439 8039 1537
tri 8039 1439 8137 1537 sw
tri 8137 1439 8235 1537 ne
rect 8235 1439 8589 1537
tri 8589 1439 8687 1537 sw
tri 8687 1439 8785 1537 ne
rect 8785 1439 9139 1537
tri 9139 1439 9237 1537 sw
tri 9237 1439 9335 1537 ne
rect 9335 1439 9689 1537
tri 9689 1439 9787 1537 sw
tri 9787 1439 9885 1537 ne
rect 9885 1439 10239 1537
tri 10239 1439 10337 1537 sw
tri 10337 1439 10435 1537 ne
rect 10435 1439 10789 1537
tri 10789 1439 10887 1537 sw
tri 10887 1439 10985 1537 ne
rect 10985 1439 11339 1537
tri 11339 1439 11437 1537 sw
tri 11437 1439 11535 1537 ne
rect 11535 1439 11889 1537
tri 11889 1439 11987 1537 sw
tri 11987 1439 12085 1537 ne
rect 12085 1439 12439 1537
tri 12439 1439 12537 1537 sw
tri 12537 1439 12635 1537 ne
rect 12635 1439 12989 1537
tri 12989 1439 13087 1537 sw
tri 13087 1439 13185 1537 ne
rect 13185 1439 13539 1537
tri 13539 1439 13637 1537 sw
tri 13637 1439 13735 1537 ne
rect 13735 1439 14089 1537
tri 14089 1439 14187 1537 sw
tri 14187 1439 14285 1537 ne
rect 14285 1439 14639 1537
tri 14639 1439 14737 1537 sw
tri 14737 1439 14835 1537 ne
rect 14835 1439 15189 1537
tri 15189 1439 15287 1537 sw
tri 15287 1439 15385 1537 ne
rect 15385 1439 15739 1537
tri 15739 1439 15837 1537 sw
tri 15837 1439 15935 1537 ne
rect 15935 1439 16289 1537
tri 16289 1439 16387 1537 sw
tri 16387 1439 16485 1537 ne
rect 16485 1439 16839 1537
tri 16839 1439 16937 1537 sw
tri 16937 1439 17035 1537 ne
rect 17035 1439 17389 1537
tri 17389 1439 17487 1537 sw
tri 17487 1439 17585 1537 ne
rect 17585 1439 17939 1537
tri 17939 1439 18037 1537 sw
tri 18037 1439 18135 1537 ne
rect 18135 1439 18489 1537
tri 18489 1439 18587 1537 sw
tri 18587 1439 18685 1537 ne
rect 18685 1439 19039 1537
tri 19039 1439 19137 1537 sw
tri 19137 1439 19235 1537 ne
rect 19235 1439 19589 1537
tri 19589 1439 19687 1537 sw
rect -500 1435 437 1439
rect -500 1315 215 1435
rect 335 1341 437 1435
tri 437 1341 535 1439 sw
tri 535 1341 633 1439 ne
rect 633 1435 987 1439
rect 633 1341 765 1435
rect 335 1315 535 1341
rect -500 1311 535 1315
tri 535 1311 565 1341 sw
tri 633 1311 663 1341 ne
rect 663 1315 765 1341
rect 885 1341 987 1435
tri 987 1341 1085 1439 sw
tri 1085 1341 1183 1439 ne
rect 1183 1435 1537 1439
rect 1183 1341 1315 1435
rect 885 1315 1085 1341
rect 663 1311 1085 1315
tri 1085 1311 1115 1341 sw
tri 1183 1311 1213 1341 ne
rect 1213 1315 1315 1341
rect 1435 1341 1537 1435
tri 1537 1341 1635 1439 sw
tri 1635 1341 1733 1439 ne
rect 1733 1435 2087 1439
rect 1733 1341 1865 1435
rect 1435 1315 1635 1341
rect 1213 1311 1635 1315
tri 1635 1311 1665 1341 sw
tri 1733 1311 1763 1341 ne
rect 1763 1315 1865 1341
rect 1985 1341 2087 1435
tri 2087 1341 2185 1439 sw
tri 2185 1341 2283 1439 ne
rect 2283 1435 2637 1439
rect 2283 1341 2415 1435
rect 1985 1315 2185 1341
rect 1763 1311 2185 1315
tri 2185 1311 2215 1341 sw
tri 2283 1311 2313 1341 ne
rect 2313 1315 2415 1341
rect 2535 1341 2637 1435
tri 2637 1341 2735 1439 sw
tri 2735 1341 2833 1439 ne
rect 2833 1435 3187 1439
rect 2833 1341 2965 1435
rect 2535 1315 2735 1341
rect 2313 1311 2735 1315
tri 2735 1311 2765 1341 sw
tri 2833 1311 2863 1341 ne
rect 2863 1315 2965 1341
rect 3085 1341 3187 1435
tri 3187 1341 3285 1439 sw
tri 3285 1341 3383 1439 ne
rect 3383 1435 3737 1439
rect 3383 1341 3515 1435
rect 3085 1315 3285 1341
rect 2863 1311 3285 1315
tri 3285 1311 3315 1341 sw
tri 3383 1311 3413 1341 ne
rect 3413 1315 3515 1341
rect 3635 1341 3737 1435
tri 3737 1341 3835 1439 sw
tri 3835 1341 3933 1439 ne
rect 3933 1435 4287 1439
rect 3933 1341 4065 1435
rect 3635 1315 3835 1341
rect 3413 1311 3835 1315
tri 3835 1311 3865 1341 sw
tri 3933 1311 3963 1341 ne
rect 3963 1315 4065 1341
rect 4185 1341 4287 1435
tri 4287 1341 4385 1439 sw
tri 4385 1341 4483 1439 ne
rect 4483 1435 4837 1439
rect 4483 1341 4615 1435
rect 4185 1315 4385 1341
rect 3963 1311 4385 1315
tri 4385 1311 4415 1341 sw
tri 4483 1311 4513 1341 ne
rect 4513 1315 4615 1341
rect 4735 1341 4837 1435
tri 4837 1341 4935 1439 sw
tri 4935 1341 5033 1439 ne
rect 5033 1435 5387 1439
rect 5033 1341 5165 1435
rect 4735 1315 4935 1341
rect 4513 1311 4935 1315
tri 4935 1311 4965 1341 sw
tri 5033 1311 5063 1341 ne
rect 5063 1315 5165 1341
rect 5285 1341 5387 1435
tri 5387 1341 5485 1439 sw
tri 5485 1341 5583 1439 ne
rect 5583 1435 5937 1439
rect 5583 1341 5715 1435
rect 5285 1315 5485 1341
rect 5063 1311 5485 1315
tri 5485 1311 5515 1341 sw
tri 5583 1311 5613 1341 ne
rect 5613 1315 5715 1341
rect 5835 1341 5937 1435
tri 5937 1341 6035 1439 sw
tri 6035 1341 6133 1439 ne
rect 6133 1435 6487 1439
rect 6133 1341 6265 1435
rect 5835 1315 6035 1341
rect 5613 1311 6035 1315
tri 6035 1311 6065 1341 sw
tri 6133 1311 6163 1341 ne
rect 6163 1315 6265 1341
rect 6385 1341 6487 1435
tri 6487 1341 6585 1439 sw
tri 6585 1341 6683 1439 ne
rect 6683 1435 7037 1439
rect 6683 1341 6815 1435
rect 6385 1315 6585 1341
rect 6163 1311 6585 1315
tri 6585 1311 6615 1341 sw
tri 6683 1311 6713 1341 ne
rect 6713 1315 6815 1341
rect 6935 1341 7037 1435
tri 7037 1341 7135 1439 sw
tri 7135 1341 7233 1439 ne
rect 7233 1435 7587 1439
rect 7233 1341 7365 1435
rect 6935 1315 7135 1341
rect 6713 1311 7135 1315
tri 7135 1311 7165 1341 sw
tri 7233 1311 7263 1341 ne
rect 7263 1315 7365 1341
rect 7485 1341 7587 1435
tri 7587 1341 7685 1439 sw
tri 7685 1341 7783 1439 ne
rect 7783 1435 8137 1439
rect 7783 1341 7915 1435
rect 7485 1315 7685 1341
rect 7263 1311 7685 1315
tri 7685 1311 7715 1341 sw
tri 7783 1311 7813 1341 ne
rect 7813 1315 7915 1341
rect 8035 1341 8137 1435
tri 8137 1341 8235 1439 sw
tri 8235 1341 8333 1439 ne
rect 8333 1435 8687 1439
rect 8333 1341 8465 1435
rect 8035 1315 8235 1341
rect 7813 1311 8235 1315
tri 8235 1311 8265 1341 sw
tri 8333 1311 8363 1341 ne
rect 8363 1315 8465 1341
rect 8585 1341 8687 1435
tri 8687 1341 8785 1439 sw
tri 8785 1341 8883 1439 ne
rect 8883 1435 9237 1439
rect 8883 1341 9015 1435
rect 8585 1315 8785 1341
rect 8363 1311 8785 1315
tri 8785 1311 8815 1341 sw
tri 8883 1311 8913 1341 ne
rect 8913 1315 9015 1341
rect 9135 1341 9237 1435
tri 9237 1341 9335 1439 sw
tri 9335 1341 9433 1439 ne
rect 9433 1435 9787 1439
rect 9433 1341 9565 1435
rect 9135 1315 9335 1341
rect 8913 1311 9335 1315
tri 9335 1311 9365 1341 sw
tri 9433 1311 9463 1341 ne
rect 9463 1315 9565 1341
rect 9685 1341 9787 1435
tri 9787 1341 9885 1439 sw
tri 9885 1341 9983 1439 ne
rect 9983 1435 10337 1439
rect 9983 1341 10115 1435
rect 9685 1315 9885 1341
rect 9463 1311 9885 1315
tri 9885 1311 9915 1341 sw
tri 9983 1311 10013 1341 ne
rect 10013 1315 10115 1341
rect 10235 1341 10337 1435
tri 10337 1341 10435 1439 sw
tri 10435 1341 10533 1439 ne
rect 10533 1435 10887 1439
rect 10533 1341 10665 1435
rect 10235 1315 10435 1341
rect 10013 1311 10435 1315
tri 10435 1311 10465 1341 sw
tri 10533 1311 10563 1341 ne
rect 10563 1315 10665 1341
rect 10785 1341 10887 1435
tri 10887 1341 10985 1439 sw
tri 10985 1341 11083 1439 ne
rect 11083 1435 11437 1439
rect 11083 1341 11215 1435
rect 10785 1315 10985 1341
rect 10563 1311 10985 1315
tri 10985 1311 11015 1341 sw
tri 11083 1311 11113 1341 ne
rect 11113 1315 11215 1341
rect 11335 1341 11437 1435
tri 11437 1341 11535 1439 sw
tri 11535 1341 11633 1439 ne
rect 11633 1435 11987 1439
rect 11633 1341 11765 1435
rect 11335 1315 11535 1341
rect 11113 1311 11535 1315
tri 11535 1311 11565 1341 sw
tri 11633 1311 11663 1341 ne
rect 11663 1315 11765 1341
rect 11885 1341 11987 1435
tri 11987 1341 12085 1439 sw
tri 12085 1341 12183 1439 ne
rect 12183 1435 12537 1439
rect 12183 1341 12315 1435
rect 11885 1315 12085 1341
rect 11663 1311 12085 1315
tri 12085 1311 12115 1341 sw
tri 12183 1311 12213 1341 ne
rect 12213 1315 12315 1341
rect 12435 1341 12537 1435
tri 12537 1341 12635 1439 sw
tri 12635 1341 12733 1439 ne
rect 12733 1435 13087 1439
rect 12733 1341 12865 1435
rect 12435 1315 12635 1341
rect 12213 1311 12635 1315
tri 12635 1311 12665 1341 sw
tri 12733 1311 12763 1341 ne
rect 12763 1315 12865 1341
rect 12985 1341 13087 1435
tri 13087 1341 13185 1439 sw
tri 13185 1341 13283 1439 ne
rect 13283 1435 13637 1439
rect 13283 1341 13415 1435
rect 12985 1315 13185 1341
rect 12763 1311 13185 1315
tri 13185 1311 13215 1341 sw
tri 13283 1311 13313 1341 ne
rect 13313 1315 13415 1341
rect 13535 1341 13637 1435
tri 13637 1341 13735 1439 sw
tri 13735 1341 13833 1439 ne
rect 13833 1435 14187 1439
rect 13833 1341 13965 1435
rect 13535 1315 13735 1341
rect 13313 1311 13735 1315
tri 13735 1311 13765 1341 sw
tri 13833 1311 13863 1341 ne
rect 13863 1315 13965 1341
rect 14085 1341 14187 1435
tri 14187 1341 14285 1439 sw
tri 14285 1341 14383 1439 ne
rect 14383 1435 14737 1439
rect 14383 1341 14515 1435
rect 14085 1315 14285 1341
rect 13863 1311 14285 1315
tri 14285 1311 14315 1341 sw
tri 14383 1311 14413 1341 ne
rect 14413 1315 14515 1341
rect 14635 1341 14737 1435
tri 14737 1341 14835 1439 sw
tri 14835 1341 14933 1439 ne
rect 14933 1435 15287 1439
rect 14933 1341 15065 1435
rect 14635 1315 14835 1341
rect 14413 1311 14835 1315
tri 14835 1311 14865 1341 sw
tri 14933 1311 14963 1341 ne
rect 14963 1315 15065 1341
rect 15185 1341 15287 1435
tri 15287 1341 15385 1439 sw
tri 15385 1341 15483 1439 ne
rect 15483 1435 15837 1439
rect 15483 1341 15615 1435
rect 15185 1315 15385 1341
rect 14963 1311 15385 1315
tri 15385 1311 15415 1341 sw
tri 15483 1311 15513 1341 ne
rect 15513 1315 15615 1341
rect 15735 1341 15837 1435
tri 15837 1341 15935 1439 sw
tri 15935 1341 16033 1439 ne
rect 16033 1435 16387 1439
rect 16033 1341 16165 1435
rect 15735 1315 15935 1341
rect 15513 1311 15935 1315
tri 15935 1311 15965 1341 sw
tri 16033 1311 16063 1341 ne
rect 16063 1315 16165 1341
rect 16285 1341 16387 1435
tri 16387 1341 16485 1439 sw
tri 16485 1341 16583 1439 ne
rect 16583 1435 16937 1439
rect 16583 1341 16715 1435
rect 16285 1315 16485 1341
rect 16063 1311 16485 1315
tri 16485 1311 16515 1341 sw
tri 16583 1311 16613 1341 ne
rect 16613 1315 16715 1341
rect 16835 1341 16937 1435
tri 16937 1341 17035 1439 sw
tri 17035 1341 17133 1439 ne
rect 17133 1435 17487 1439
rect 17133 1341 17265 1435
rect 16835 1315 17035 1341
rect 16613 1311 17035 1315
tri 17035 1311 17065 1341 sw
tri 17133 1311 17163 1341 ne
rect 17163 1315 17265 1341
rect 17385 1341 17487 1435
tri 17487 1341 17585 1439 sw
tri 17585 1341 17683 1439 ne
rect 17683 1435 18037 1439
rect 17683 1341 17815 1435
rect 17385 1315 17585 1341
rect 17163 1311 17585 1315
tri 17585 1311 17615 1341 sw
tri 17683 1311 17713 1341 ne
rect 17713 1315 17815 1341
rect 17935 1341 18037 1435
tri 18037 1341 18135 1439 sw
tri 18135 1341 18233 1439 ne
rect 18233 1435 18587 1439
rect 18233 1341 18365 1435
rect 17935 1315 18135 1341
rect 17713 1311 18135 1315
tri 18135 1311 18165 1341 sw
tri 18233 1311 18263 1341 ne
rect 18263 1315 18365 1341
rect 18485 1341 18587 1435
tri 18587 1341 18685 1439 sw
tri 18685 1341 18783 1439 ne
rect 18783 1435 19137 1439
rect 18783 1341 18915 1435
rect 18485 1315 18685 1341
rect 18263 1311 18685 1315
tri 18685 1311 18715 1341 sw
tri 18783 1311 18813 1341 ne
rect 18813 1315 18915 1341
rect 19035 1341 19137 1435
tri 19137 1341 19235 1439 sw
tri 19235 1341 19333 1439 ne
rect 19333 1435 20300 1439
rect 19333 1341 19465 1435
rect 19035 1315 19235 1341
rect 18813 1311 19235 1315
tri 19235 1311 19265 1341 sw
tri 19333 1311 19363 1341 ne
rect 19363 1315 19465 1341
rect 19585 1315 20300 1435
rect 19363 1311 20300 1315
tri 113 1213 211 1311 ne
rect 211 1213 565 1311
tri 565 1213 663 1311 sw
tri 663 1213 761 1311 ne
rect 761 1213 1115 1311
tri 1115 1213 1213 1311 sw
tri 1213 1213 1311 1311 ne
rect 1311 1213 1665 1311
tri 1665 1213 1763 1311 sw
tri 1763 1213 1861 1311 ne
rect 1861 1213 2215 1311
tri 2215 1213 2313 1311 sw
tri 2313 1213 2411 1311 ne
rect 2411 1213 2765 1311
tri 2765 1213 2863 1311 sw
tri 2863 1213 2961 1311 ne
rect 2961 1213 3315 1311
tri 3315 1213 3413 1311 sw
tri 3413 1213 3511 1311 ne
rect 3511 1213 3865 1311
tri 3865 1213 3963 1311 sw
tri 3963 1213 4061 1311 ne
rect 4061 1213 4415 1311
tri 4415 1213 4513 1311 sw
tri 4513 1213 4611 1311 ne
rect 4611 1213 4965 1311
tri 4965 1213 5063 1311 sw
tri 5063 1213 5161 1311 ne
rect 5161 1213 5515 1311
tri 5515 1213 5613 1311 sw
tri 5613 1213 5711 1311 ne
rect 5711 1213 6065 1311
tri 6065 1213 6163 1311 sw
tri 6163 1213 6261 1311 ne
rect 6261 1213 6615 1311
tri 6615 1213 6713 1311 sw
tri 6713 1213 6811 1311 ne
rect 6811 1213 7165 1311
tri 7165 1213 7263 1311 sw
tri 7263 1213 7361 1311 ne
rect 7361 1213 7715 1311
tri 7715 1213 7813 1311 sw
tri 7813 1213 7911 1311 ne
rect 7911 1213 8265 1311
tri 8265 1213 8363 1311 sw
tri 8363 1213 8461 1311 ne
rect 8461 1213 8815 1311
tri 8815 1213 8913 1311 sw
tri 8913 1213 9011 1311 ne
rect 9011 1213 9365 1311
tri 9365 1213 9463 1311 sw
tri 9463 1213 9561 1311 ne
rect 9561 1213 9915 1311
tri 9915 1213 10013 1311 sw
tri 10013 1213 10111 1311 ne
rect 10111 1213 10465 1311
tri 10465 1213 10563 1311 sw
tri 10563 1213 10661 1311 ne
rect 10661 1213 11015 1311
tri 11015 1213 11113 1311 sw
tri 11113 1213 11211 1311 ne
rect 11211 1213 11565 1311
tri 11565 1213 11663 1311 sw
tri 11663 1213 11761 1311 ne
rect 11761 1213 12115 1311
tri 12115 1213 12213 1311 sw
tri 12213 1213 12311 1311 ne
rect 12311 1213 12665 1311
tri 12665 1213 12763 1311 sw
tri 12763 1213 12861 1311 ne
rect 12861 1213 13215 1311
tri 13215 1213 13313 1311 sw
tri 13313 1213 13411 1311 ne
rect 13411 1213 13765 1311
tri 13765 1213 13863 1311 sw
tri 13863 1213 13961 1311 ne
rect 13961 1213 14315 1311
tri 14315 1213 14413 1311 sw
tri 14413 1213 14511 1311 ne
rect 14511 1213 14865 1311
tri 14865 1213 14963 1311 sw
tri 14963 1213 15061 1311 ne
rect 15061 1213 15415 1311
tri 15415 1213 15513 1311 sw
tri 15513 1213 15611 1311 ne
rect 15611 1213 15965 1311
tri 15965 1213 16063 1311 sw
tri 16063 1213 16161 1311 ne
rect 16161 1213 16515 1311
tri 16515 1213 16613 1311 sw
tri 16613 1213 16711 1311 ne
rect 16711 1213 17065 1311
tri 17065 1213 17163 1311 sw
tri 17163 1213 17261 1311 ne
rect 17261 1213 17615 1311
tri 17615 1213 17713 1311 sw
tri 17713 1213 17811 1311 ne
rect 17811 1213 18165 1311
tri 18165 1213 18263 1311 sw
tri 18263 1213 18361 1311 ne
rect 18361 1213 18715 1311
tri 18715 1213 18813 1311 sw
tri 18813 1213 18911 1311 ne
rect 18911 1213 19265 1311
tri 19265 1213 19363 1311 sw
tri 19363 1213 19461 1311 ne
rect 19461 1213 20300 1311
rect -1000 1183 113 1213
tri 113 1183 143 1213 sw
tri 211 1183 241 1213 ne
rect 241 1183 663 1213
tri 663 1183 693 1213 sw
tri 761 1183 791 1213 ne
rect 791 1183 1213 1213
tri 1213 1183 1243 1213 sw
tri 1311 1183 1341 1213 ne
rect 1341 1183 1763 1213
tri 1763 1183 1793 1213 sw
tri 1861 1183 1891 1213 ne
rect 1891 1183 2313 1213
tri 2313 1183 2343 1213 sw
tri 2411 1183 2441 1213 ne
rect 2441 1183 2863 1213
tri 2863 1183 2893 1213 sw
tri 2961 1183 2991 1213 ne
rect 2991 1183 3413 1213
tri 3413 1183 3443 1213 sw
tri 3511 1183 3541 1213 ne
rect 3541 1183 3963 1213
tri 3963 1183 3993 1213 sw
tri 4061 1183 4091 1213 ne
rect 4091 1183 4513 1213
tri 4513 1183 4543 1213 sw
tri 4611 1183 4641 1213 ne
rect 4641 1183 5063 1213
tri 5063 1183 5093 1213 sw
tri 5161 1183 5191 1213 ne
rect 5191 1183 5613 1213
tri 5613 1183 5643 1213 sw
tri 5711 1183 5741 1213 ne
rect 5741 1183 6163 1213
tri 6163 1183 6193 1213 sw
tri 6261 1183 6291 1213 ne
rect 6291 1183 6713 1213
tri 6713 1183 6743 1213 sw
tri 6811 1183 6841 1213 ne
rect 6841 1183 7263 1213
tri 7263 1183 7293 1213 sw
tri 7361 1183 7391 1213 ne
rect 7391 1183 7813 1213
tri 7813 1183 7843 1213 sw
tri 7911 1183 7941 1213 ne
rect 7941 1183 8363 1213
tri 8363 1183 8393 1213 sw
tri 8461 1183 8491 1213 ne
rect 8491 1183 8913 1213
tri 8913 1183 8943 1213 sw
tri 9011 1183 9041 1213 ne
rect 9041 1183 9463 1213
tri 9463 1183 9493 1213 sw
tri 9561 1183 9591 1213 ne
rect 9591 1183 10013 1213
tri 10013 1183 10043 1213 sw
tri 10111 1183 10141 1213 ne
rect 10141 1183 10563 1213
tri 10563 1183 10593 1213 sw
tri 10661 1183 10691 1213 ne
rect 10691 1183 11113 1213
tri 11113 1183 11143 1213 sw
tri 11211 1183 11241 1213 ne
rect 11241 1183 11663 1213
tri 11663 1183 11693 1213 sw
tri 11761 1183 11791 1213 ne
rect 11791 1183 12213 1213
tri 12213 1183 12243 1213 sw
tri 12311 1183 12341 1213 ne
rect 12341 1183 12763 1213
tri 12763 1183 12793 1213 sw
tri 12861 1183 12891 1213 ne
rect 12891 1183 13313 1213
tri 13313 1183 13343 1213 sw
tri 13411 1183 13441 1213 ne
rect 13441 1183 13863 1213
tri 13863 1183 13893 1213 sw
tri 13961 1183 13991 1213 ne
rect 13991 1183 14413 1213
tri 14413 1183 14443 1213 sw
tri 14511 1183 14541 1213 ne
rect 14541 1183 14963 1213
tri 14963 1183 14993 1213 sw
tri 15061 1183 15091 1213 ne
rect 15091 1183 15513 1213
tri 15513 1183 15543 1213 sw
tri 15611 1183 15641 1213 ne
rect 15641 1183 16063 1213
tri 16063 1183 16093 1213 sw
tri 16161 1183 16191 1213 ne
rect 16191 1183 16613 1213
tri 16613 1183 16643 1213 sw
tri 16711 1183 16741 1213 ne
rect 16741 1183 17163 1213
tri 17163 1183 17193 1213 sw
tri 17261 1183 17291 1213 ne
rect 17291 1183 17713 1213
tri 17713 1183 17743 1213 sw
tri 17811 1183 17841 1213 ne
rect 17841 1183 18263 1213
tri 18263 1183 18293 1213 sw
tri 18361 1183 18391 1213 ne
rect 18391 1183 18813 1213
tri 18813 1183 18843 1213 sw
tri 18911 1183 18941 1213 ne
rect 18941 1183 19363 1213
tri 19363 1183 19393 1213 sw
tri 19461 1183 19491 1213 ne
rect 19491 1183 20300 1213
rect -1000 1085 143 1183
tri 143 1085 241 1183 sw
tri 241 1085 339 1183 ne
rect 339 1085 693 1183
tri 693 1085 791 1183 sw
tri 791 1085 889 1183 ne
rect 889 1085 1243 1183
tri 1243 1085 1341 1183 sw
tri 1341 1085 1439 1183 ne
rect 1439 1085 1793 1183
tri 1793 1085 1891 1183 sw
tri 1891 1085 1989 1183 ne
rect 1989 1085 2343 1183
tri 2343 1085 2441 1183 sw
tri 2441 1085 2539 1183 ne
rect 2539 1085 2893 1183
tri 2893 1085 2991 1183 sw
tri 2991 1085 3089 1183 ne
rect 3089 1085 3443 1183
tri 3443 1085 3541 1183 sw
tri 3541 1085 3639 1183 ne
rect 3639 1085 3993 1183
tri 3993 1085 4091 1183 sw
tri 4091 1085 4189 1183 ne
rect 4189 1085 4543 1183
tri 4543 1085 4641 1183 sw
tri 4641 1085 4739 1183 ne
rect 4739 1085 5093 1183
tri 5093 1085 5191 1183 sw
tri 5191 1085 5289 1183 ne
rect 5289 1085 5643 1183
tri 5643 1085 5741 1183 sw
tri 5741 1085 5839 1183 ne
rect 5839 1085 6193 1183
tri 6193 1085 6291 1183 sw
tri 6291 1085 6389 1183 ne
rect 6389 1085 6743 1183
tri 6743 1085 6841 1183 sw
tri 6841 1085 6939 1183 ne
rect 6939 1085 7293 1183
tri 7293 1085 7391 1183 sw
tri 7391 1085 7489 1183 ne
rect 7489 1085 7843 1183
tri 7843 1085 7941 1183 sw
tri 7941 1085 8039 1183 ne
rect 8039 1085 8393 1183
tri 8393 1085 8491 1183 sw
tri 8491 1085 8589 1183 ne
rect 8589 1085 8943 1183
tri 8943 1085 9041 1183 sw
tri 9041 1085 9139 1183 ne
rect 9139 1085 9493 1183
tri 9493 1085 9591 1183 sw
tri 9591 1085 9689 1183 ne
rect 9689 1085 10043 1183
tri 10043 1085 10141 1183 sw
tri 10141 1085 10239 1183 ne
rect 10239 1085 10593 1183
tri 10593 1085 10691 1183 sw
tri 10691 1085 10789 1183 ne
rect 10789 1085 11143 1183
tri 11143 1085 11241 1183 sw
tri 11241 1085 11339 1183 ne
rect 11339 1085 11693 1183
tri 11693 1085 11791 1183 sw
tri 11791 1085 11889 1183 ne
rect 11889 1085 12243 1183
tri 12243 1085 12341 1183 sw
tri 12341 1085 12439 1183 ne
rect 12439 1085 12793 1183
tri 12793 1085 12891 1183 sw
tri 12891 1085 12989 1183 ne
rect 12989 1085 13343 1183
tri 13343 1085 13441 1183 sw
tri 13441 1085 13539 1183 ne
rect 13539 1085 13893 1183
tri 13893 1085 13991 1183 sw
tri 13991 1085 14089 1183 ne
rect 14089 1085 14443 1183
tri 14443 1085 14541 1183 sw
tri 14541 1085 14639 1183 ne
rect 14639 1085 14993 1183
tri 14993 1085 15091 1183 sw
tri 15091 1085 15189 1183 ne
rect 15189 1085 15543 1183
tri 15543 1085 15641 1183 sw
tri 15641 1085 15739 1183 ne
rect 15739 1085 16093 1183
tri 16093 1085 16191 1183 sw
tri 16191 1085 16289 1183 ne
rect 16289 1085 16643 1183
tri 16643 1085 16741 1183 sw
tri 16741 1085 16839 1183 ne
rect 16839 1085 17193 1183
tri 17193 1085 17291 1183 sw
tri 17291 1085 17389 1183 ne
rect 17389 1085 17743 1183
tri 17743 1085 17841 1183 sw
tri 17841 1085 17939 1183 ne
rect 17939 1085 18293 1183
tri 18293 1085 18391 1183 sw
tri 18391 1085 18489 1183 ne
rect 18489 1085 18843 1183
tri 18843 1085 18941 1183 sw
tri 18941 1085 19039 1183 ne
rect 19039 1085 19393 1183
tri 19393 1085 19491 1183 sw
tri 19491 1085 19589 1183 ne
rect 19589 1085 20300 1183
rect -1000 987 241 1085
tri 241 987 339 1085 sw
tri 339 987 437 1085 ne
rect 437 987 791 1085
tri 791 987 889 1085 sw
tri 889 987 987 1085 ne
rect 987 987 1341 1085
tri 1341 987 1439 1085 sw
tri 1439 987 1537 1085 ne
rect 1537 987 1891 1085
tri 1891 987 1989 1085 sw
tri 1989 987 2087 1085 ne
rect 2087 987 2441 1085
tri 2441 987 2539 1085 sw
tri 2539 987 2637 1085 ne
rect 2637 987 2991 1085
tri 2991 987 3089 1085 sw
tri 3089 987 3187 1085 ne
rect 3187 987 3541 1085
tri 3541 987 3639 1085 sw
tri 3639 987 3737 1085 ne
rect 3737 987 4091 1085
tri 4091 987 4189 1085 sw
tri 4189 987 4287 1085 ne
rect 4287 987 4641 1085
tri 4641 987 4739 1085 sw
tri 4739 987 4837 1085 ne
rect 4837 987 5191 1085
tri 5191 987 5289 1085 sw
tri 5289 987 5387 1085 ne
rect 5387 987 5741 1085
tri 5741 987 5839 1085 sw
tri 5839 987 5937 1085 ne
rect 5937 987 6291 1085
tri 6291 987 6389 1085 sw
tri 6389 987 6487 1085 ne
rect 6487 987 6841 1085
tri 6841 987 6939 1085 sw
tri 6939 987 7037 1085 ne
rect 7037 987 7391 1085
tri 7391 987 7489 1085 sw
tri 7489 987 7587 1085 ne
rect 7587 987 7941 1085
tri 7941 987 8039 1085 sw
tri 8039 987 8137 1085 ne
rect 8137 987 8491 1085
tri 8491 987 8589 1085 sw
tri 8589 987 8687 1085 ne
rect 8687 987 9041 1085
tri 9041 987 9139 1085 sw
tri 9139 987 9237 1085 ne
rect 9237 987 9591 1085
tri 9591 987 9689 1085 sw
tri 9689 987 9787 1085 ne
rect 9787 987 10141 1085
tri 10141 987 10239 1085 sw
tri 10239 987 10337 1085 ne
rect 10337 987 10691 1085
tri 10691 987 10789 1085 sw
tri 10789 987 10887 1085 ne
rect 10887 987 11241 1085
tri 11241 987 11339 1085 sw
tri 11339 987 11437 1085 ne
rect 11437 987 11791 1085
tri 11791 987 11889 1085 sw
tri 11889 987 11987 1085 ne
rect 11987 987 12341 1085
tri 12341 987 12439 1085 sw
tri 12439 987 12537 1085 ne
rect 12537 987 12891 1085
tri 12891 987 12989 1085 sw
tri 12989 987 13087 1085 ne
rect 13087 987 13441 1085
tri 13441 987 13539 1085 sw
tri 13539 987 13637 1085 ne
rect 13637 987 13991 1085
tri 13991 987 14089 1085 sw
tri 14089 987 14187 1085 ne
rect 14187 987 14541 1085
tri 14541 987 14639 1085 sw
tri 14639 987 14737 1085 ne
rect 14737 987 15091 1085
tri 15091 987 15189 1085 sw
tri 15189 987 15287 1085 ne
rect 15287 987 15641 1085
tri 15641 987 15739 1085 sw
tri 15739 987 15837 1085 ne
rect 15837 987 16191 1085
tri 16191 987 16289 1085 sw
tri 16289 987 16387 1085 ne
rect 16387 987 16741 1085
tri 16741 987 16839 1085 sw
tri 16839 987 16937 1085 ne
rect 16937 987 17291 1085
tri 17291 987 17389 1085 sw
tri 17389 987 17487 1085 ne
rect 17487 987 17841 1085
tri 17841 987 17939 1085 sw
tri 17939 987 18037 1085 ne
rect 18037 987 18391 1085
tri 18391 987 18489 1085 sw
tri 18489 987 18587 1085 ne
rect 18587 987 18941 1085
tri 18941 987 19039 1085 sw
tri 19039 987 19137 1085 ne
rect 19137 987 19491 1085
tri 19491 987 19589 1085 sw
tri 19589 987 19687 1085 ne
rect 19687 987 20300 1085
rect -1000 889 339 987
tri 339 889 437 987 sw
tri 437 889 535 987 ne
rect 535 889 889 987
tri 889 889 987 987 sw
tri 987 889 1085 987 ne
rect 1085 889 1439 987
tri 1439 889 1537 987 sw
tri 1537 889 1635 987 ne
rect 1635 889 1989 987
tri 1989 889 2087 987 sw
tri 2087 889 2185 987 ne
rect 2185 889 2539 987
tri 2539 889 2637 987 sw
tri 2637 889 2735 987 ne
rect 2735 889 3089 987
tri 3089 889 3187 987 sw
tri 3187 889 3285 987 ne
rect 3285 889 3639 987
tri 3639 889 3737 987 sw
tri 3737 889 3835 987 ne
rect 3835 889 4189 987
tri 4189 889 4287 987 sw
tri 4287 889 4385 987 ne
rect 4385 889 4739 987
tri 4739 889 4837 987 sw
tri 4837 889 4935 987 ne
rect 4935 889 5289 987
tri 5289 889 5387 987 sw
tri 5387 889 5485 987 ne
rect 5485 889 5839 987
tri 5839 889 5937 987 sw
tri 5937 889 6035 987 ne
rect 6035 889 6389 987
tri 6389 889 6487 987 sw
tri 6487 889 6585 987 ne
rect 6585 889 6939 987
tri 6939 889 7037 987 sw
tri 7037 889 7135 987 ne
rect 7135 889 7489 987
tri 7489 889 7587 987 sw
tri 7587 889 7685 987 ne
rect 7685 889 8039 987
tri 8039 889 8137 987 sw
tri 8137 889 8235 987 ne
rect 8235 889 8589 987
tri 8589 889 8687 987 sw
tri 8687 889 8785 987 ne
rect 8785 889 9139 987
tri 9139 889 9237 987 sw
tri 9237 889 9335 987 ne
rect 9335 889 9689 987
tri 9689 889 9787 987 sw
tri 9787 889 9885 987 ne
rect 9885 889 10239 987
tri 10239 889 10337 987 sw
tri 10337 889 10435 987 ne
rect 10435 889 10789 987
tri 10789 889 10887 987 sw
tri 10887 889 10985 987 ne
rect 10985 889 11339 987
tri 11339 889 11437 987 sw
tri 11437 889 11535 987 ne
rect 11535 889 11889 987
tri 11889 889 11987 987 sw
tri 11987 889 12085 987 ne
rect 12085 889 12439 987
tri 12439 889 12537 987 sw
tri 12537 889 12635 987 ne
rect 12635 889 12989 987
tri 12989 889 13087 987 sw
tri 13087 889 13185 987 ne
rect 13185 889 13539 987
tri 13539 889 13637 987 sw
tri 13637 889 13735 987 ne
rect 13735 889 14089 987
tri 14089 889 14187 987 sw
tri 14187 889 14285 987 ne
rect 14285 889 14639 987
tri 14639 889 14737 987 sw
tri 14737 889 14835 987 ne
rect 14835 889 15189 987
tri 15189 889 15287 987 sw
tri 15287 889 15385 987 ne
rect 15385 889 15739 987
tri 15739 889 15837 987 sw
tri 15837 889 15935 987 ne
rect 15935 889 16289 987
tri 16289 889 16387 987 sw
tri 16387 889 16485 987 ne
rect 16485 889 16839 987
tri 16839 889 16937 987 sw
tri 16937 889 17035 987 ne
rect 17035 889 17389 987
tri 17389 889 17487 987 sw
tri 17487 889 17585 987 ne
rect 17585 889 17939 987
tri 17939 889 18037 987 sw
tri 18037 889 18135 987 ne
rect 18135 889 18489 987
tri 18489 889 18587 987 sw
tri 18587 889 18685 987 ne
rect 18685 889 19039 987
tri 19039 889 19137 987 sw
tri 19137 889 19235 987 ne
rect 19235 889 19589 987
tri 19589 889 19687 987 sw
rect 20800 889 21800 1537
rect -1000 885 437 889
rect -1000 765 215 885
rect 335 791 437 885
tri 437 791 535 889 sw
tri 535 791 633 889 ne
rect 633 885 987 889
rect 633 791 765 885
rect 335 765 535 791
rect -1000 761 535 765
tri 113 663 211 761 ne
rect 211 713 535 761
tri 535 713 613 791 sw
tri 633 713 711 791 ne
rect 711 765 765 791
rect 885 791 987 885
tri 987 791 1085 889 sw
tri 1085 791 1183 889 ne
rect 1183 885 1537 889
rect 1183 791 1315 885
rect 885 765 1085 791
rect 711 713 1085 765
tri 1085 713 1163 791 sw
tri 1183 713 1261 791 ne
rect 1261 765 1315 791
rect 1435 791 1537 885
tri 1537 791 1635 889 sw
tri 1635 791 1733 889 ne
rect 1733 885 2087 889
rect 1733 791 1865 885
rect 1435 765 1635 791
rect 1261 713 1635 765
tri 1635 713 1713 791 sw
tri 1733 713 1811 791 ne
rect 1811 765 1865 791
rect 1985 791 2087 885
tri 2087 791 2185 889 sw
tri 2185 791 2283 889 ne
rect 2283 885 2637 889
rect 2283 791 2415 885
rect 1985 765 2185 791
rect 1811 713 2185 765
tri 2185 713 2263 791 sw
tri 2283 713 2361 791 ne
rect 2361 765 2415 791
rect 2535 791 2637 885
tri 2637 791 2735 889 sw
tri 2735 791 2833 889 ne
rect 2833 885 3187 889
rect 2833 791 2965 885
rect 2535 765 2735 791
rect 2361 713 2735 765
tri 2735 713 2813 791 sw
tri 2833 713 2911 791 ne
rect 2911 765 2965 791
rect 3085 791 3187 885
tri 3187 791 3285 889 sw
tri 3285 791 3383 889 ne
rect 3383 885 3737 889
rect 3383 791 3515 885
rect 3085 765 3285 791
rect 2911 713 3285 765
tri 3285 713 3363 791 sw
tri 3383 713 3461 791 ne
rect 3461 765 3515 791
rect 3635 791 3737 885
tri 3737 791 3835 889 sw
tri 3835 791 3933 889 ne
rect 3933 885 4287 889
rect 3933 791 4065 885
rect 3635 765 3835 791
rect 3461 713 3835 765
tri 3835 713 3913 791 sw
tri 3933 713 4011 791 ne
rect 4011 765 4065 791
rect 4185 791 4287 885
tri 4287 791 4385 889 sw
tri 4385 791 4483 889 ne
rect 4483 885 4837 889
rect 4483 791 4615 885
rect 4185 765 4385 791
rect 4011 713 4385 765
tri 4385 713 4463 791 sw
tri 4483 713 4561 791 ne
rect 4561 765 4615 791
rect 4735 791 4837 885
tri 4837 791 4935 889 sw
tri 4935 791 5033 889 ne
rect 5033 885 5387 889
rect 5033 791 5165 885
rect 4735 765 4935 791
rect 4561 713 4935 765
tri 4935 713 5013 791 sw
tri 5033 713 5111 791 ne
rect 5111 765 5165 791
rect 5285 791 5387 885
tri 5387 791 5485 889 sw
tri 5485 791 5583 889 ne
rect 5583 885 5937 889
rect 5583 791 5715 885
rect 5285 765 5485 791
rect 5111 713 5485 765
tri 5485 713 5563 791 sw
tri 5583 713 5661 791 ne
rect 5661 765 5715 791
rect 5835 791 5937 885
tri 5937 791 6035 889 sw
tri 6035 791 6133 889 ne
rect 6133 885 6487 889
rect 6133 791 6265 885
rect 5835 765 6035 791
rect 5661 713 6035 765
tri 6035 713 6113 791 sw
tri 6133 713 6211 791 ne
rect 6211 765 6265 791
rect 6385 791 6487 885
tri 6487 791 6585 889 sw
tri 6585 791 6683 889 ne
rect 6683 885 7037 889
rect 6683 791 6815 885
rect 6385 765 6585 791
rect 6211 713 6585 765
tri 6585 713 6663 791 sw
tri 6683 713 6761 791 ne
rect 6761 765 6815 791
rect 6935 791 7037 885
tri 7037 791 7135 889 sw
tri 7135 791 7233 889 ne
rect 7233 885 7587 889
rect 7233 791 7365 885
rect 6935 765 7135 791
rect 6761 713 7135 765
tri 7135 713 7213 791 sw
tri 7233 713 7311 791 ne
rect 7311 765 7365 791
rect 7485 791 7587 885
tri 7587 791 7685 889 sw
tri 7685 791 7783 889 ne
rect 7783 885 8137 889
rect 7783 791 7915 885
rect 7485 765 7685 791
rect 7311 713 7685 765
tri 7685 713 7763 791 sw
tri 7783 713 7861 791 ne
rect 7861 765 7915 791
rect 8035 791 8137 885
tri 8137 791 8235 889 sw
tri 8235 791 8333 889 ne
rect 8333 885 8687 889
rect 8333 791 8465 885
rect 8035 765 8235 791
rect 7861 713 8235 765
tri 8235 713 8313 791 sw
tri 8333 713 8411 791 ne
rect 8411 765 8465 791
rect 8585 791 8687 885
tri 8687 791 8785 889 sw
tri 8785 791 8883 889 ne
rect 8883 885 9237 889
rect 8883 791 9015 885
rect 8585 765 8785 791
rect 8411 713 8785 765
tri 8785 713 8863 791 sw
tri 8883 713 8961 791 ne
rect 8961 765 9015 791
rect 9135 791 9237 885
tri 9237 791 9335 889 sw
tri 9335 791 9433 889 ne
rect 9433 885 9787 889
rect 9433 791 9565 885
rect 9135 765 9335 791
rect 8961 713 9335 765
tri 9335 713 9413 791 sw
tri 9433 713 9511 791 ne
rect 9511 765 9565 791
rect 9685 791 9787 885
tri 9787 791 9885 889 sw
tri 9885 791 9983 889 ne
rect 9983 885 10337 889
rect 9983 791 10115 885
rect 9685 765 9885 791
rect 9511 713 9885 765
tri 9885 713 9963 791 sw
tri 9983 713 10061 791 ne
rect 10061 765 10115 791
rect 10235 791 10337 885
tri 10337 791 10435 889 sw
tri 10435 791 10533 889 ne
rect 10533 885 10887 889
rect 10533 791 10665 885
rect 10235 765 10435 791
rect 10061 713 10435 765
tri 10435 713 10513 791 sw
tri 10533 713 10611 791 ne
rect 10611 765 10665 791
rect 10785 791 10887 885
tri 10887 791 10985 889 sw
tri 10985 791 11083 889 ne
rect 11083 885 11437 889
rect 11083 791 11215 885
rect 10785 765 10985 791
rect 10611 713 10985 765
tri 10985 713 11063 791 sw
tri 11083 713 11161 791 ne
rect 11161 765 11215 791
rect 11335 791 11437 885
tri 11437 791 11535 889 sw
tri 11535 791 11633 889 ne
rect 11633 885 11987 889
rect 11633 791 11765 885
rect 11335 765 11535 791
rect 11161 713 11535 765
tri 11535 713 11613 791 sw
tri 11633 713 11711 791 ne
rect 11711 765 11765 791
rect 11885 791 11987 885
tri 11987 791 12085 889 sw
tri 12085 791 12183 889 ne
rect 12183 885 12537 889
rect 12183 791 12315 885
rect 11885 765 12085 791
rect 11711 713 12085 765
tri 12085 713 12163 791 sw
tri 12183 713 12261 791 ne
rect 12261 765 12315 791
rect 12435 791 12537 885
tri 12537 791 12635 889 sw
tri 12635 791 12733 889 ne
rect 12733 885 13087 889
rect 12733 791 12865 885
rect 12435 765 12635 791
rect 12261 713 12635 765
tri 12635 713 12713 791 sw
tri 12733 713 12811 791 ne
rect 12811 765 12865 791
rect 12985 791 13087 885
tri 13087 791 13185 889 sw
tri 13185 791 13283 889 ne
rect 13283 885 13637 889
rect 13283 791 13415 885
rect 12985 765 13185 791
rect 12811 713 13185 765
tri 13185 713 13263 791 sw
tri 13283 713 13361 791 ne
rect 13361 765 13415 791
rect 13535 791 13637 885
tri 13637 791 13735 889 sw
tri 13735 791 13833 889 ne
rect 13833 885 14187 889
rect 13833 791 13965 885
rect 13535 765 13735 791
rect 13361 713 13735 765
tri 13735 713 13813 791 sw
tri 13833 713 13911 791 ne
rect 13911 765 13965 791
rect 14085 791 14187 885
tri 14187 791 14285 889 sw
tri 14285 791 14383 889 ne
rect 14383 885 14737 889
rect 14383 791 14515 885
rect 14085 765 14285 791
rect 13911 713 14285 765
tri 14285 713 14363 791 sw
tri 14383 713 14461 791 ne
rect 14461 765 14515 791
rect 14635 791 14737 885
tri 14737 791 14835 889 sw
tri 14835 791 14933 889 ne
rect 14933 885 15287 889
rect 14933 791 15065 885
rect 14635 765 14835 791
rect 14461 713 14835 765
tri 14835 713 14913 791 sw
tri 14933 713 15011 791 ne
rect 15011 765 15065 791
rect 15185 791 15287 885
tri 15287 791 15385 889 sw
tri 15385 791 15483 889 ne
rect 15483 885 15837 889
rect 15483 791 15615 885
rect 15185 765 15385 791
rect 15011 713 15385 765
tri 15385 713 15463 791 sw
tri 15483 713 15561 791 ne
rect 15561 765 15615 791
rect 15735 791 15837 885
tri 15837 791 15935 889 sw
tri 15935 791 16033 889 ne
rect 16033 885 16387 889
rect 16033 791 16165 885
rect 15735 765 15935 791
rect 15561 713 15935 765
tri 15935 713 16013 791 sw
tri 16033 713 16111 791 ne
rect 16111 765 16165 791
rect 16285 791 16387 885
tri 16387 791 16485 889 sw
tri 16485 791 16583 889 ne
rect 16583 885 16937 889
rect 16583 791 16715 885
rect 16285 765 16485 791
rect 16111 713 16485 765
tri 16485 713 16563 791 sw
tri 16583 713 16661 791 ne
rect 16661 765 16715 791
rect 16835 791 16937 885
tri 16937 791 17035 889 sw
tri 17035 791 17133 889 ne
rect 17133 885 17487 889
rect 17133 791 17265 885
rect 16835 765 17035 791
rect 16661 713 17035 765
tri 17035 713 17113 791 sw
tri 17133 713 17211 791 ne
rect 17211 765 17265 791
rect 17385 791 17487 885
tri 17487 791 17585 889 sw
tri 17585 791 17683 889 ne
rect 17683 885 18037 889
rect 17683 791 17815 885
rect 17385 765 17585 791
rect 17211 713 17585 765
tri 17585 713 17663 791 sw
tri 17683 713 17761 791 ne
rect 17761 765 17815 791
rect 17935 791 18037 885
tri 18037 791 18135 889 sw
tri 18135 791 18233 889 ne
rect 18233 885 18587 889
rect 18233 791 18365 885
rect 17935 765 18135 791
rect 17761 713 18135 765
tri 18135 713 18213 791 sw
tri 18233 713 18311 791 ne
rect 18311 765 18365 791
rect 18485 791 18587 885
tri 18587 791 18685 889 sw
tri 18685 791 18783 889 ne
rect 18783 885 19137 889
rect 18783 791 18915 885
rect 18485 765 18685 791
rect 18311 713 18685 765
tri 18685 713 18763 791 sw
tri 18783 713 18861 791 ne
rect 18861 765 18915 791
rect 19035 791 19137 885
tri 19137 791 19235 889 sw
tri 19235 791 19333 889 ne
rect 19333 885 21800 889
rect 19333 791 19465 885
rect 19035 765 19235 791
rect 18861 713 19235 765
tri 19235 713 19313 791 sw
tri 19333 713 19411 791 ne
rect 19411 765 19465 791
rect 19585 765 21800 885
rect 19411 713 21800 765
rect 211 663 613 713
rect -500 613 113 663
tri 113 613 163 663 sw
tri 211 613 261 663 ne
rect 261 633 613 663
tri 613 633 693 713 sw
tri 711 633 791 713 ne
rect 791 633 1163 713
tri 1163 633 1243 713 sw
tri 1261 633 1341 713 ne
rect 1341 633 1713 713
tri 1713 633 1793 713 sw
tri 1811 633 1891 713 ne
rect 1891 633 2263 713
tri 2263 633 2343 713 sw
tri 2361 633 2441 713 ne
rect 2441 633 2813 713
tri 2813 633 2893 713 sw
tri 2911 633 2991 713 ne
rect 2991 633 3363 713
tri 3363 633 3443 713 sw
tri 3461 633 3541 713 ne
rect 3541 633 3913 713
tri 3913 633 3993 713 sw
tri 4011 633 4091 713 ne
rect 4091 633 4463 713
tri 4463 633 4543 713 sw
tri 4561 633 4641 713 ne
rect 4641 633 5013 713
tri 5013 633 5093 713 sw
tri 5111 633 5191 713 ne
rect 5191 633 5563 713
tri 5563 633 5643 713 sw
tri 5661 633 5741 713 ne
rect 5741 633 6113 713
tri 6113 633 6193 713 sw
tri 6211 633 6291 713 ne
rect 6291 633 6663 713
tri 6663 633 6743 713 sw
tri 6761 633 6841 713 ne
rect 6841 633 7213 713
tri 7213 633 7293 713 sw
tri 7311 633 7391 713 ne
rect 7391 633 7763 713
tri 7763 633 7843 713 sw
tri 7861 633 7941 713 ne
rect 7941 633 8313 713
tri 8313 633 8393 713 sw
tri 8411 633 8491 713 ne
rect 8491 633 8863 713
tri 8863 633 8943 713 sw
tri 8961 633 9041 713 ne
rect 9041 633 9413 713
tri 9413 633 9493 713 sw
tri 9511 633 9591 713 ne
rect 9591 633 9963 713
tri 9963 633 10043 713 sw
tri 10061 633 10141 713 ne
rect 10141 633 10513 713
tri 10513 633 10593 713 sw
tri 10611 633 10691 713 ne
rect 10691 633 11063 713
tri 11063 633 11143 713 sw
tri 11161 633 11241 713 ne
rect 11241 633 11613 713
tri 11613 633 11693 713 sw
tri 11711 633 11791 713 ne
rect 11791 633 12163 713
tri 12163 633 12243 713 sw
tri 12261 633 12341 713 ne
rect 12341 633 12713 713
tri 12713 633 12793 713 sw
tri 12811 633 12891 713 ne
rect 12891 633 13263 713
tri 13263 633 13343 713 sw
tri 13361 633 13441 713 ne
rect 13441 633 13813 713
tri 13813 633 13893 713 sw
tri 13911 633 13991 713 ne
rect 13991 633 14363 713
tri 14363 633 14443 713 sw
tri 14461 633 14541 713 ne
rect 14541 633 14913 713
tri 14913 633 14993 713 sw
tri 15011 633 15091 713 ne
rect 15091 633 15463 713
tri 15463 633 15543 713 sw
tri 15561 633 15641 713 ne
rect 15641 633 16013 713
tri 16013 633 16093 713 sw
tri 16111 633 16191 713 ne
rect 16191 633 16563 713
tri 16563 633 16643 713 sw
tri 16661 633 16741 713 ne
rect 16741 633 17113 713
tri 17113 633 17193 713 sw
tri 17211 633 17291 713 ne
rect 17291 633 17663 713
tri 17663 633 17743 713 sw
tri 17761 633 17841 713 ne
rect 17841 633 18213 713
tri 18213 633 18293 713 sw
tri 18311 633 18391 713 ne
rect 18391 633 18763 713
tri 18763 633 18843 713 sw
tri 18861 633 18941 713 ne
rect 18941 633 19313 713
tri 19313 633 19393 713 sw
tri 19411 633 19491 713 ne
rect 19491 633 20100 713
rect 261 613 693 633
rect -500 535 163 613
tri 163 535 241 613 sw
tri 261 535 339 613 ne
rect 339 535 693 613
tri 693 535 791 633 sw
tri 791 535 889 633 ne
rect 889 535 1243 633
tri 1243 535 1341 633 sw
tri 1341 535 1439 633 ne
rect 1439 535 1793 633
tri 1793 535 1891 633 sw
tri 1891 535 1989 633 ne
rect 1989 535 2343 633
tri 2343 535 2441 633 sw
tri 2441 535 2539 633 ne
rect 2539 535 2893 633
tri 2893 535 2991 633 sw
tri 2991 535 3089 633 ne
rect 3089 535 3443 633
tri 3443 535 3541 633 sw
tri 3541 535 3639 633 ne
rect 3639 535 3993 633
tri 3993 535 4091 633 sw
tri 4091 535 4189 633 ne
rect 4189 535 4543 633
tri 4543 535 4641 633 sw
tri 4641 535 4739 633 ne
rect 4739 535 5093 633
tri 5093 535 5191 633 sw
tri 5191 535 5289 633 ne
rect 5289 535 5643 633
tri 5643 535 5741 633 sw
tri 5741 535 5839 633 ne
rect 5839 535 6193 633
tri 6193 535 6291 633 sw
tri 6291 535 6389 633 ne
rect 6389 535 6743 633
tri 6743 535 6841 633 sw
tri 6841 535 6939 633 ne
rect 6939 535 7293 633
tri 7293 535 7391 633 sw
tri 7391 535 7489 633 ne
rect 7489 535 7843 633
tri 7843 535 7941 633 sw
tri 7941 535 8039 633 ne
rect 8039 535 8393 633
tri 8393 535 8491 633 sw
tri 8491 535 8589 633 ne
rect 8589 535 8943 633
tri 8943 535 9041 633 sw
tri 9041 535 9139 633 ne
rect 9139 535 9493 633
tri 9493 535 9591 633 sw
tri 9591 535 9689 633 ne
rect 9689 535 10043 633
tri 10043 535 10141 633 sw
tri 10141 535 10239 633 ne
rect 10239 535 10593 633
tri 10593 535 10691 633 sw
tri 10691 535 10789 633 ne
rect 10789 535 11143 633
tri 11143 535 11241 633 sw
tri 11241 535 11339 633 ne
rect 11339 535 11693 633
tri 11693 535 11791 633 sw
tri 11791 535 11889 633 ne
rect 11889 535 12243 633
tri 12243 535 12341 633 sw
tri 12341 535 12439 633 ne
rect 12439 535 12793 633
tri 12793 535 12891 633 sw
tri 12891 535 12989 633 ne
rect 12989 535 13343 633
tri 13343 535 13441 633 sw
tri 13441 535 13539 633 ne
rect 13539 535 13893 633
tri 13893 535 13991 633 sw
tri 13991 535 14089 633 ne
rect 14089 535 14443 633
tri 14443 535 14541 633 sw
tri 14541 535 14639 633 ne
rect 14639 535 14993 633
tri 14993 535 15091 633 sw
tri 15091 535 15189 633 ne
rect 15189 535 15543 633
tri 15543 535 15641 633 sw
tri 15641 535 15739 633 ne
rect 15739 535 16093 633
tri 16093 535 16191 633 sw
tri 16191 535 16289 633 ne
rect 16289 535 16643 633
tri 16643 535 16741 633 sw
tri 16741 535 16839 633 ne
rect 16839 535 17193 633
tri 17193 535 17291 633 sw
tri 17291 535 17389 633 ne
rect 17389 535 17743 633
tri 17743 535 17841 633 sw
tri 17841 535 17939 633 ne
rect 17939 535 18293 633
tri 18293 535 18391 633 sw
tri 18391 535 18489 633 ne
rect 18489 535 18843 633
tri 18843 535 18941 633 sw
tri 18941 535 19039 633 ne
rect 19039 535 19393 633
tri 19393 535 19491 633 sw
tri 19491 535 19589 633 ne
rect 19589 613 20100 633
rect 20200 613 21800 713
rect 19589 535 21800 613
rect -500 487 241 535
rect -500 387 -400 487
rect -300 437 241 487
tri 241 437 339 535 sw
tri 339 437 437 535 ne
rect 437 437 791 535
tri 791 437 889 535 sw
tri 889 437 987 535 ne
rect 987 437 1341 535
tri 1341 437 1439 535 sw
tri 1439 437 1537 535 ne
rect 1537 437 1891 535
tri 1891 437 1989 535 sw
tri 1989 437 2087 535 ne
rect 2087 437 2441 535
tri 2441 437 2539 535 sw
tri 2539 437 2637 535 ne
rect 2637 437 2991 535
tri 2991 437 3089 535 sw
tri 3089 437 3187 535 ne
rect 3187 437 3541 535
tri 3541 437 3639 535 sw
tri 3639 437 3737 535 ne
rect 3737 437 4091 535
tri 4091 437 4189 535 sw
tri 4189 437 4287 535 ne
rect 4287 437 4641 535
tri 4641 437 4739 535 sw
tri 4739 437 4837 535 ne
rect 4837 437 5191 535
tri 5191 437 5289 535 sw
tri 5289 437 5387 535 ne
rect 5387 437 5741 535
tri 5741 437 5839 535 sw
tri 5839 437 5937 535 ne
rect 5937 437 6291 535
tri 6291 437 6389 535 sw
tri 6389 437 6487 535 ne
rect 6487 437 6841 535
tri 6841 437 6939 535 sw
tri 6939 437 7037 535 ne
rect 7037 437 7391 535
tri 7391 437 7489 535 sw
tri 7489 437 7587 535 ne
rect 7587 437 7941 535
tri 7941 437 8039 535 sw
tri 8039 437 8137 535 ne
rect 8137 437 8491 535
tri 8491 437 8589 535 sw
tri 8589 437 8687 535 ne
rect 8687 437 9041 535
tri 9041 437 9139 535 sw
tri 9139 437 9237 535 ne
rect 9237 437 9591 535
tri 9591 437 9689 535 sw
tri 9689 437 9787 535 ne
rect 9787 437 10141 535
tri 10141 437 10239 535 sw
tri 10239 437 10337 535 ne
rect 10337 437 10691 535
tri 10691 437 10789 535 sw
tri 10789 437 10887 535 ne
rect 10887 437 11241 535
tri 11241 437 11339 535 sw
tri 11339 437 11437 535 ne
rect 11437 437 11791 535
tri 11791 437 11889 535 sw
tri 11889 437 11987 535 ne
rect 11987 437 12341 535
tri 12341 437 12439 535 sw
tri 12439 437 12537 535 ne
rect 12537 437 12891 535
tri 12891 437 12989 535 sw
tri 12989 437 13087 535 ne
rect 13087 437 13441 535
tri 13441 437 13539 535 sw
tri 13539 437 13637 535 ne
rect 13637 437 13991 535
tri 13991 437 14089 535 sw
tri 14089 437 14187 535 ne
rect 14187 437 14541 535
tri 14541 437 14639 535 sw
tri 14639 437 14737 535 ne
rect 14737 437 15091 535
tri 15091 437 15189 535 sw
tri 15189 437 15287 535 ne
rect 15287 437 15641 535
tri 15641 437 15739 535 sw
tri 15739 437 15837 535 ne
rect 15837 437 16191 535
tri 16191 437 16289 535 sw
tri 16289 437 16387 535 ne
rect 16387 437 16741 535
tri 16741 437 16839 535 sw
tri 16839 437 16937 535 ne
rect 16937 437 17291 535
tri 17291 437 17389 535 sw
tri 17389 437 17487 535 ne
rect 17487 437 17841 535
tri 17841 437 17939 535 sw
tri 17939 437 18037 535 ne
rect 18037 437 18391 535
tri 18391 437 18489 535 sw
tri 18489 437 18587 535 ne
rect 18587 437 18941 535
tri 18941 437 19039 535 sw
tri 19039 437 19137 535 ne
rect 19137 437 19491 535
tri 19491 437 19589 535 sw
tri 19589 437 19687 535 ne
rect 19687 437 21800 535
rect -300 387 339 437
rect -500 339 339 387
tri 339 339 437 437 sw
tri 437 339 535 437 ne
rect 535 339 889 437
tri 889 339 987 437 sw
tri 987 339 1085 437 ne
rect 1085 339 1439 437
tri 1439 339 1537 437 sw
tri 1537 339 1635 437 ne
rect 1635 339 1989 437
tri 1989 339 2087 437 sw
tri 2087 339 2185 437 ne
rect 2185 339 2539 437
tri 2539 339 2637 437 sw
tri 2637 339 2735 437 ne
rect 2735 339 3089 437
tri 3089 339 3187 437 sw
tri 3187 339 3285 437 ne
rect 3285 339 3639 437
tri 3639 339 3737 437 sw
tri 3737 339 3835 437 ne
rect 3835 339 4189 437
tri 4189 339 4287 437 sw
tri 4287 339 4385 437 ne
rect 4385 339 4739 437
tri 4739 339 4837 437 sw
tri 4837 339 4935 437 ne
rect 4935 339 5289 437
tri 5289 339 5387 437 sw
tri 5387 339 5485 437 ne
rect 5485 339 5839 437
tri 5839 339 5937 437 sw
tri 5937 339 6035 437 ne
rect 6035 339 6389 437
tri 6389 339 6487 437 sw
tri 6487 339 6585 437 ne
rect 6585 339 6939 437
tri 6939 339 7037 437 sw
tri 7037 339 7135 437 ne
rect 7135 339 7489 437
tri 7489 339 7587 437 sw
tri 7587 339 7685 437 ne
rect 7685 339 8039 437
tri 8039 339 8137 437 sw
tri 8137 339 8235 437 ne
rect 8235 339 8589 437
tri 8589 339 8687 437 sw
tri 8687 339 8785 437 ne
rect 8785 339 9139 437
tri 9139 339 9237 437 sw
tri 9237 339 9335 437 ne
rect 9335 339 9689 437
tri 9689 339 9787 437 sw
tri 9787 339 9885 437 ne
rect 9885 339 10239 437
tri 10239 339 10337 437 sw
tri 10337 339 10435 437 ne
rect 10435 339 10789 437
tri 10789 339 10887 437 sw
tri 10887 339 10985 437 ne
rect 10985 339 11339 437
tri 11339 339 11437 437 sw
tri 11437 339 11535 437 ne
rect 11535 339 11889 437
tri 11889 339 11987 437 sw
tri 11987 339 12085 437 ne
rect 12085 339 12439 437
tri 12439 339 12537 437 sw
tri 12537 339 12635 437 ne
rect 12635 339 12989 437
tri 12989 339 13087 437 sw
tri 13087 339 13185 437 ne
rect 13185 339 13539 437
tri 13539 339 13637 437 sw
tri 13637 339 13735 437 ne
rect 13735 339 14089 437
tri 14089 339 14187 437 sw
tri 14187 339 14285 437 ne
rect 14285 339 14639 437
tri 14639 339 14737 437 sw
tri 14737 339 14835 437 ne
rect 14835 339 15189 437
tri 15189 339 15287 437 sw
tri 15287 339 15385 437 ne
rect 15385 339 15739 437
tri 15739 339 15837 437 sw
tri 15837 339 15935 437 ne
rect 15935 339 16289 437
tri 16289 339 16387 437 sw
tri 16387 339 16485 437 ne
rect 16485 339 16839 437
tri 16839 339 16937 437 sw
tri 16937 339 17035 437 ne
rect 17035 339 17389 437
tri 17389 339 17487 437 sw
tri 17487 339 17585 437 ne
rect 17585 339 17939 437
tri 17939 339 18037 437 sw
tri 18037 339 18135 437 ne
rect 18135 339 18489 437
tri 18489 339 18587 437 sw
tri 18587 339 18685 437 ne
rect 18685 339 19039 437
tri 19039 339 19137 437 sw
tri 19137 339 19235 437 ne
rect 19235 339 19589 437
tri 19589 339 19687 437 sw
rect -500 335 437 339
rect -500 215 215 335
rect 335 241 437 335
tri 437 241 535 339 sw
tri 535 241 633 339 ne
rect 633 335 987 339
rect 633 241 765 335
rect 335 215 535 241
rect -500 211 535 215
tri 535 211 565 241 sw
tri 633 211 663 241 ne
rect 663 215 765 241
rect 885 241 987 335
tri 987 241 1085 339 sw
tri 1085 241 1183 339 ne
rect 1183 335 1537 339
rect 1183 241 1315 335
rect 885 215 1085 241
rect 663 211 1085 215
tri 1085 211 1115 241 sw
tri 1183 211 1213 241 ne
rect 1213 215 1315 241
rect 1435 241 1537 335
tri 1537 241 1635 339 sw
tri 1635 241 1733 339 ne
rect 1733 335 2087 339
rect 1733 241 1865 335
rect 1435 215 1635 241
rect 1213 211 1635 215
tri 1635 211 1665 241 sw
tri 1733 211 1763 241 ne
rect 1763 215 1865 241
rect 1985 241 2087 335
tri 2087 241 2185 339 sw
tri 2185 241 2283 339 ne
rect 2283 335 2637 339
rect 2283 241 2415 335
rect 1985 215 2185 241
rect 1763 211 2185 215
tri 2185 211 2215 241 sw
tri 2283 211 2313 241 ne
rect 2313 215 2415 241
rect 2535 241 2637 335
tri 2637 241 2735 339 sw
tri 2735 241 2833 339 ne
rect 2833 335 3187 339
rect 2833 241 2965 335
rect 2535 215 2735 241
rect 2313 211 2735 215
tri 2735 211 2765 241 sw
tri 2833 211 2863 241 ne
rect 2863 215 2965 241
rect 3085 241 3187 335
tri 3187 241 3285 339 sw
tri 3285 241 3383 339 ne
rect 3383 335 3737 339
rect 3383 241 3515 335
rect 3085 215 3285 241
rect 2863 211 3285 215
tri 3285 211 3315 241 sw
tri 3383 211 3413 241 ne
rect 3413 215 3515 241
rect 3635 241 3737 335
tri 3737 241 3835 339 sw
tri 3835 241 3933 339 ne
rect 3933 335 4287 339
rect 3933 241 4065 335
rect 3635 215 3835 241
rect 3413 211 3835 215
tri 3835 211 3865 241 sw
tri 3933 211 3963 241 ne
rect 3963 215 4065 241
rect 4185 241 4287 335
tri 4287 241 4385 339 sw
tri 4385 241 4483 339 ne
rect 4483 335 4837 339
rect 4483 241 4615 335
rect 4185 215 4385 241
rect 3963 211 4385 215
tri 4385 211 4415 241 sw
tri 4483 211 4513 241 ne
rect 4513 215 4615 241
rect 4735 241 4837 335
tri 4837 241 4935 339 sw
tri 4935 241 5033 339 ne
rect 5033 335 5387 339
rect 5033 241 5165 335
rect 4735 215 4935 241
rect 4513 211 4935 215
tri 4935 211 4965 241 sw
tri 5033 211 5063 241 ne
rect 5063 215 5165 241
rect 5285 241 5387 335
tri 5387 241 5485 339 sw
tri 5485 241 5583 339 ne
rect 5583 335 5937 339
rect 5583 241 5715 335
rect 5285 215 5485 241
rect 5063 211 5485 215
tri 5485 211 5515 241 sw
tri 5583 211 5613 241 ne
rect 5613 215 5715 241
rect 5835 241 5937 335
tri 5937 241 6035 339 sw
tri 6035 241 6133 339 ne
rect 6133 335 6487 339
rect 6133 241 6265 335
rect 5835 215 6035 241
rect 5613 211 6035 215
tri 6035 211 6065 241 sw
tri 6133 211 6163 241 ne
rect 6163 215 6265 241
rect 6385 241 6487 335
tri 6487 241 6585 339 sw
tri 6585 241 6683 339 ne
rect 6683 335 7037 339
rect 6683 241 6815 335
rect 6385 215 6585 241
rect 6163 211 6585 215
tri 6585 211 6615 241 sw
tri 6683 211 6713 241 ne
rect 6713 215 6815 241
rect 6935 241 7037 335
tri 7037 241 7135 339 sw
tri 7135 241 7233 339 ne
rect 7233 335 7587 339
rect 7233 241 7365 335
rect 6935 215 7135 241
rect 6713 211 7135 215
tri 7135 211 7165 241 sw
tri 7233 211 7263 241 ne
rect 7263 215 7365 241
rect 7485 241 7587 335
tri 7587 241 7685 339 sw
tri 7685 241 7783 339 ne
rect 7783 335 8137 339
rect 7783 241 7915 335
rect 7485 215 7685 241
rect 7263 211 7685 215
tri 7685 211 7715 241 sw
tri 7783 211 7813 241 ne
rect 7813 215 7915 241
rect 8035 241 8137 335
tri 8137 241 8235 339 sw
tri 8235 241 8333 339 ne
rect 8333 335 8687 339
rect 8333 241 8465 335
rect 8035 215 8235 241
rect 7813 211 8235 215
tri 8235 211 8265 241 sw
tri 8333 211 8363 241 ne
rect 8363 215 8465 241
rect 8585 241 8687 335
tri 8687 241 8785 339 sw
tri 8785 241 8883 339 ne
rect 8883 335 9237 339
rect 8883 241 9015 335
rect 8585 215 8785 241
rect 8363 211 8785 215
tri 8785 211 8815 241 sw
tri 8883 211 8913 241 ne
rect 8913 215 9015 241
rect 9135 241 9237 335
tri 9237 241 9335 339 sw
tri 9335 241 9433 339 ne
rect 9433 335 9787 339
rect 9433 241 9565 335
rect 9135 215 9335 241
rect 8913 211 9335 215
tri 9335 211 9365 241 sw
tri 9433 211 9463 241 ne
rect 9463 215 9565 241
rect 9685 241 9787 335
tri 9787 241 9885 339 sw
tri 9885 241 9983 339 ne
rect 9983 335 10337 339
rect 9983 241 10115 335
rect 9685 215 9885 241
rect 9463 211 9885 215
tri 9885 211 9915 241 sw
tri 9983 211 10013 241 ne
rect 10013 215 10115 241
rect 10235 241 10337 335
tri 10337 241 10435 339 sw
tri 10435 241 10533 339 ne
rect 10533 335 10887 339
rect 10533 241 10665 335
rect 10235 215 10435 241
rect 10013 211 10435 215
tri 10435 211 10465 241 sw
tri 10533 211 10563 241 ne
rect 10563 215 10665 241
rect 10785 241 10887 335
tri 10887 241 10985 339 sw
tri 10985 241 11083 339 ne
rect 11083 335 11437 339
rect 11083 241 11215 335
rect 10785 215 10985 241
rect 10563 211 10985 215
tri 10985 211 11015 241 sw
tri 11083 211 11113 241 ne
rect 11113 215 11215 241
rect 11335 241 11437 335
tri 11437 241 11535 339 sw
tri 11535 241 11633 339 ne
rect 11633 335 11987 339
rect 11633 241 11765 335
rect 11335 215 11535 241
rect 11113 211 11535 215
tri 11535 211 11565 241 sw
tri 11633 211 11663 241 ne
rect 11663 215 11765 241
rect 11885 241 11987 335
tri 11987 241 12085 339 sw
tri 12085 241 12183 339 ne
rect 12183 335 12537 339
rect 12183 241 12315 335
rect 11885 215 12085 241
rect 11663 211 12085 215
tri 12085 211 12115 241 sw
tri 12183 211 12213 241 ne
rect 12213 215 12315 241
rect 12435 241 12537 335
tri 12537 241 12635 339 sw
tri 12635 241 12733 339 ne
rect 12733 335 13087 339
rect 12733 241 12865 335
rect 12435 215 12635 241
rect 12213 211 12635 215
tri 12635 211 12665 241 sw
tri 12733 211 12763 241 ne
rect 12763 215 12865 241
rect 12985 241 13087 335
tri 13087 241 13185 339 sw
tri 13185 241 13283 339 ne
rect 13283 335 13637 339
rect 13283 241 13415 335
rect 12985 215 13185 241
rect 12763 211 13185 215
tri 13185 211 13215 241 sw
tri 13283 211 13313 241 ne
rect 13313 215 13415 241
rect 13535 241 13637 335
tri 13637 241 13735 339 sw
tri 13735 241 13833 339 ne
rect 13833 335 14187 339
rect 13833 241 13965 335
rect 13535 215 13735 241
rect 13313 211 13735 215
tri 13735 211 13765 241 sw
tri 13833 211 13863 241 ne
rect 13863 215 13965 241
rect 14085 241 14187 335
tri 14187 241 14285 339 sw
tri 14285 241 14383 339 ne
rect 14383 335 14737 339
rect 14383 241 14515 335
rect 14085 215 14285 241
rect 13863 211 14285 215
tri 14285 211 14315 241 sw
tri 14383 211 14413 241 ne
rect 14413 215 14515 241
rect 14635 241 14737 335
tri 14737 241 14835 339 sw
tri 14835 241 14933 339 ne
rect 14933 335 15287 339
rect 14933 241 15065 335
rect 14635 215 14835 241
rect 14413 211 14835 215
tri 14835 211 14865 241 sw
tri 14933 211 14963 241 ne
rect 14963 215 15065 241
rect 15185 241 15287 335
tri 15287 241 15385 339 sw
tri 15385 241 15483 339 ne
rect 15483 335 15837 339
rect 15483 241 15615 335
rect 15185 215 15385 241
rect 14963 211 15385 215
tri 15385 211 15415 241 sw
tri 15483 211 15513 241 ne
rect 15513 215 15615 241
rect 15735 241 15837 335
tri 15837 241 15935 339 sw
tri 15935 241 16033 339 ne
rect 16033 335 16387 339
rect 16033 241 16165 335
rect 15735 215 15935 241
rect 15513 211 15935 215
tri 15935 211 15965 241 sw
tri 16033 211 16063 241 ne
rect 16063 215 16165 241
rect 16285 241 16387 335
tri 16387 241 16485 339 sw
tri 16485 241 16583 339 ne
rect 16583 335 16937 339
rect 16583 241 16715 335
rect 16285 215 16485 241
rect 16063 211 16485 215
tri 16485 211 16515 241 sw
tri 16583 211 16613 241 ne
rect 16613 215 16715 241
rect 16835 241 16937 335
tri 16937 241 17035 339 sw
tri 17035 241 17133 339 ne
rect 17133 335 17487 339
rect 17133 241 17265 335
rect 16835 215 17035 241
rect 16613 211 17035 215
tri 17035 211 17065 241 sw
tri 17133 211 17163 241 ne
rect 17163 215 17265 241
rect 17385 241 17487 335
tri 17487 241 17585 339 sw
tri 17585 241 17683 339 ne
rect 17683 335 18037 339
rect 17683 241 17815 335
rect 17385 215 17585 241
rect 17163 211 17585 215
tri 17585 211 17615 241 sw
tri 17683 211 17713 241 ne
rect 17713 215 17815 241
rect 17935 241 18037 335
tri 18037 241 18135 339 sw
tri 18135 241 18233 339 ne
rect 18233 335 18587 339
rect 18233 241 18365 335
rect 17935 215 18135 241
rect 17713 211 18135 215
tri 18135 211 18165 241 sw
tri 18233 211 18263 241 ne
rect 18263 215 18365 241
rect 18485 241 18587 335
tri 18587 241 18685 339 sw
tri 18685 241 18783 339 ne
rect 18783 335 19137 339
rect 18783 241 18915 335
rect 18485 215 18685 241
rect 18263 211 18685 215
tri 18685 211 18715 241 sw
tri 18783 211 18813 241 ne
rect 18813 215 18915 241
rect 19035 241 19137 335
tri 19137 241 19235 339 sw
tri 19235 241 19333 339 ne
rect 19333 335 20300 339
rect 19333 241 19465 335
rect 19035 215 19235 241
rect 18813 211 19235 215
tri 19235 211 19265 241 sw
tri 19333 211 19363 241 ne
rect 19363 215 19465 241
rect 19585 215 20300 335
rect 19363 211 20300 215
tri 113 113 211 211 ne
rect 211 113 565 211
tri 565 113 663 211 sw
tri 663 113 761 211 ne
rect 761 113 1115 211
tri 1115 113 1213 211 sw
tri 1213 113 1311 211 ne
rect 1311 113 1665 211
tri 1665 113 1763 211 sw
tri 1763 113 1861 211 ne
rect 1861 113 2215 211
tri 2215 113 2313 211 sw
tri 2313 113 2411 211 ne
rect 2411 113 2765 211
tri 2765 113 2863 211 sw
tri 2863 113 2961 211 ne
rect 2961 113 3315 211
tri 3315 113 3413 211 sw
tri 3413 113 3511 211 ne
rect 3511 113 3865 211
tri 3865 113 3963 211 sw
tri 3963 113 4061 211 ne
rect 4061 113 4415 211
tri 4415 113 4513 211 sw
tri 4513 113 4611 211 ne
rect 4611 113 4965 211
tri 4965 113 5063 211 sw
tri 5063 113 5161 211 ne
rect 5161 113 5515 211
tri 5515 113 5613 211 sw
tri 5613 113 5711 211 ne
rect 5711 113 6065 211
tri 6065 113 6163 211 sw
tri 6163 113 6261 211 ne
rect 6261 113 6615 211
tri 6615 113 6713 211 sw
tri 6713 113 6811 211 ne
rect 6811 113 7165 211
tri 7165 113 7263 211 sw
tri 7263 113 7361 211 ne
rect 7361 113 7715 211
tri 7715 113 7813 211 sw
tri 7813 113 7911 211 ne
rect 7911 113 8265 211
tri 8265 113 8363 211 sw
tri 8363 113 8461 211 ne
rect 8461 113 8815 211
tri 8815 113 8913 211 sw
tri 8913 113 9011 211 ne
rect 9011 113 9365 211
tri 9365 113 9463 211 sw
tri 9463 113 9561 211 ne
rect 9561 113 9915 211
tri 9915 113 10013 211 sw
tri 10013 113 10111 211 ne
rect 10111 113 10465 211
tri 10465 113 10563 211 sw
tri 10563 113 10661 211 ne
rect 10661 113 11015 211
tri 11015 113 11113 211 sw
tri 11113 113 11211 211 ne
rect 11211 113 11565 211
tri 11565 113 11663 211 sw
tri 11663 113 11761 211 ne
rect 11761 113 12115 211
tri 12115 113 12213 211 sw
tri 12213 113 12311 211 ne
rect 12311 113 12665 211
tri 12665 113 12763 211 sw
tri 12763 113 12861 211 ne
rect 12861 113 13215 211
tri 13215 113 13313 211 sw
tri 13313 113 13411 211 ne
rect 13411 113 13765 211
tri 13765 113 13863 211 sw
tri 13863 113 13961 211 ne
rect 13961 113 14315 211
tri 14315 113 14413 211 sw
tri 14413 113 14511 211 ne
rect 14511 113 14865 211
tri 14865 113 14963 211 sw
tri 14963 113 15061 211 ne
rect 15061 113 15415 211
tri 15415 113 15513 211 sw
tri 15513 113 15611 211 ne
rect 15611 113 15965 211
tri 15965 113 16063 211 sw
tri 16063 113 16161 211 ne
rect 16161 113 16515 211
tri 16515 113 16613 211 sw
tri 16613 113 16711 211 ne
rect 16711 113 17065 211
tri 17065 113 17163 211 sw
tri 17163 113 17261 211 ne
rect 17261 113 17615 211
tri 17615 113 17713 211 sw
tri 17713 113 17811 211 ne
rect 17811 113 18165 211
tri 18165 113 18263 211 sw
tri 18263 113 18361 211 ne
rect 18361 113 18715 211
tri 18715 113 18813 211 sw
tri 18813 113 18911 211 ne
rect 18911 113 19265 211
tri 19265 113 19363 211 sw
tri 19363 113 19461 211 ne
rect 211 -300 663 113
rect 211 -400 387 -300
rect 487 -400 663 -300
rect 211 -1000 663 -400
rect 761 -500 1213 113
rect 1311 -300 1763 113
rect 1311 -400 1487 -300
rect 1587 -400 1763 -300
rect 1311 -1000 1763 -400
rect 1861 -500 2313 113
rect 2411 -300 2863 113
rect 2411 -400 2587 -300
rect 2687 -400 2863 -300
rect 2411 -1000 2863 -400
rect 2961 -500 3413 113
rect 3511 -300 3963 113
rect 3511 -400 3687 -300
rect 3787 -400 3963 -300
rect 3511 -1000 3963 -400
rect 4061 -500 4513 113
rect 4611 -300 5063 113
rect 4611 -400 4787 -300
rect 4887 -400 5063 -300
rect 4611 -1000 5063 -400
rect 5161 -500 5613 113
rect 5711 -300 6163 113
rect 5711 -400 5887 -300
rect 5987 -400 6163 -300
rect 5711 -1000 6163 -400
rect 6261 -500 6713 113
rect 6811 -300 7263 113
rect 6811 -400 6987 -300
rect 7087 -400 7263 -300
rect 6811 -1000 7263 -400
rect 7361 -500 7813 113
rect 7911 -300 8363 113
rect 7911 -400 8087 -300
rect 8187 -400 8363 -300
rect 7911 -1000 8363 -400
rect 8461 -500 8913 113
rect 9011 -300 9463 113
rect 9011 -400 9187 -300
rect 9287 -400 9463 -300
rect 9011 -1000 9463 -400
rect 9561 -500 10013 113
rect 10111 -300 10563 113
rect 10111 -400 10287 -300
rect 10387 -400 10563 -300
rect 10111 -1000 10563 -400
rect 10661 -500 11113 113
rect 11211 -300 11663 113
rect 11211 -400 11387 -300
rect 11487 -400 11663 -300
rect 11211 -1000 11663 -400
rect 11761 -500 12213 113
rect 12311 -300 12763 113
rect 12311 -400 12487 -300
rect 12587 -400 12763 -300
rect 12311 -1000 12763 -400
rect 12861 -500 13313 113
rect 13411 -300 13863 113
rect 13411 -400 13587 -300
rect 13687 -400 13863 -300
rect 13411 -1000 13863 -400
rect 13961 -500 14413 113
rect 14511 -300 14963 113
rect 14511 -400 14687 -300
rect 14787 -400 14963 -300
rect 14511 -1000 14963 -400
rect 15061 -500 15513 113
rect 15611 -300 16063 113
rect 15611 -400 15787 -300
rect 15887 -400 16063 -300
rect 15611 -1000 16063 -400
rect 16161 -500 16613 113
rect 16711 -300 17163 113
rect 16711 -400 16887 -300
rect 16987 -400 17163 -300
rect 16711 -1000 17163 -400
rect 17261 -500 17713 113
rect 17811 -300 18263 113
rect 17811 -400 17987 -300
rect 18087 -400 18263 -300
rect 17811 -1000 18263 -400
rect 18361 -500 18813 113
rect 18911 -300 19363 113
rect 18911 -400 19087 -300
rect 19187 -400 19363 -300
rect 18911 -1000 19363 -400
rect 19461 -113 20300 211
rect 19461 -500 19913 -113
rect 20800 -1000 21800 437
rect 0 -2000 21800 -1000
<< via3 >>
rect 613 20100 713 20200
rect 1713 20100 1813 20200
rect 2813 20100 2913 20200
rect 3913 20100 4013 20200
rect 5013 20100 5113 20200
rect 6113 20100 6213 20200
rect 7213 20100 7313 20200
rect 8313 20100 8413 20200
rect 9413 20100 9513 20200
rect 10513 20100 10613 20200
rect 11613 20100 11713 20200
rect 12713 20100 12813 20200
rect 13813 20100 13913 20200
rect 14913 20100 15013 20200
rect 16013 20100 16113 20200
rect 17113 20100 17213 20200
rect 18213 20100 18313 20200
rect 19313 20100 19413 20200
rect 215 19465 335 19585
rect 765 19465 885 19585
rect 1315 19465 1435 19585
rect 1865 19465 1985 19585
rect 2415 19465 2535 19585
rect 2965 19465 3085 19585
rect 3515 19465 3635 19585
rect 4065 19465 4185 19585
rect 4615 19465 4735 19585
rect 5165 19465 5285 19585
rect 5715 19465 5835 19585
rect 6265 19465 6385 19585
rect 6815 19465 6935 19585
rect 7365 19465 7485 19585
rect 7915 19465 8035 19585
rect 8465 19465 8585 19585
rect 9015 19465 9135 19585
rect 9565 19465 9685 19585
rect 10115 19465 10235 19585
rect 10665 19465 10785 19585
rect 11215 19465 11335 19585
rect 11765 19465 11885 19585
rect 12315 19465 12435 19585
rect 12865 19465 12985 19585
rect 13415 19465 13535 19585
rect 13965 19465 14085 19585
rect 14515 19465 14635 19585
rect 15065 19465 15185 19585
rect 15615 19465 15735 19585
rect 16165 19465 16285 19585
rect 16715 19465 16835 19585
rect 17265 19465 17385 19585
rect 17815 19465 17935 19585
rect 18365 19465 18485 19585
rect 18915 19465 19035 19585
rect 19465 19465 19585 19585
rect 20100 19313 20200 19413
rect -400 19087 -300 19187
rect 215 18915 335 19035
rect 19465 18915 19585 19035
rect 215 18365 335 18485
rect 19465 18365 19585 18485
rect 20100 18213 20200 18313
rect -400 17987 -300 18087
rect 215 17815 335 17935
rect 19465 17815 19585 17935
rect 215 17265 335 17385
rect 19465 17265 19585 17385
rect 20100 17113 20200 17213
rect -400 16887 -300 16987
rect 215 16715 335 16835
rect 19465 16715 19585 16835
rect 215 16165 335 16285
rect 19465 16165 19585 16285
rect 20100 16013 20200 16113
rect -400 15787 -300 15887
rect 215 15615 335 15735
rect 19465 15615 19585 15735
rect 215 15065 335 15185
rect 19465 15065 19585 15185
rect 20100 14913 20200 15013
rect -400 14687 -300 14787
rect 215 14515 335 14635
rect 19465 14515 19585 14635
rect 215 13965 335 14085
rect 19465 13965 19585 14085
rect 20100 13813 20200 13913
rect -400 13587 -300 13687
rect 215 13415 335 13535
rect 19465 13415 19585 13535
rect 215 12865 335 12985
rect 19465 12865 19585 12985
rect 20100 12713 20200 12813
rect -400 12487 -300 12587
rect 215 12315 335 12435
rect 19465 12315 19585 12435
rect 215 11765 335 11885
rect 19465 11765 19585 11885
rect 20100 11613 20200 11713
rect -400 11387 -300 11487
rect 215 11215 335 11335
rect 19465 11215 19585 11335
rect 215 10665 335 10785
rect 19465 10665 19585 10785
rect 20100 10513 20200 10613
rect -400 10287 -300 10387
rect 215 10115 335 10235
rect 19465 10115 19585 10235
rect 215 9565 335 9685
rect 19465 9565 19585 9685
rect 20100 9413 20200 9513
rect -400 9187 -300 9287
rect 215 9015 335 9135
rect 19465 9015 19585 9135
rect 215 8465 335 8585
rect 19465 8465 19585 8585
rect 20100 8313 20200 8413
rect -400 8087 -300 8187
rect 215 7915 335 8035
rect 19465 7915 19585 8035
rect 215 7365 335 7485
rect 19465 7365 19585 7485
rect 20100 7213 20200 7313
rect -400 6987 -300 7087
rect 215 6815 335 6935
rect 19465 6815 19585 6935
rect 215 6265 335 6385
rect 19465 6265 19585 6385
rect 20100 6113 20200 6213
rect -400 5887 -300 5987
rect 215 5715 335 5835
rect 19465 5715 19585 5835
rect 215 5165 335 5285
rect 19465 5165 19585 5285
rect 20100 5013 20200 5113
rect -400 4787 -300 4887
rect 215 4615 335 4735
rect 19465 4615 19585 4735
rect 215 4065 335 4185
rect 19465 4065 19585 4185
rect 20100 3913 20200 4013
rect -400 3687 -300 3787
rect 215 3515 335 3635
rect 19465 3515 19585 3635
rect 215 2965 335 3085
rect 19465 2965 19585 3085
rect 20100 2813 20200 2913
rect -400 2587 -300 2687
rect 215 2415 335 2535
rect 19465 2415 19585 2535
rect 215 1865 335 1985
rect 19465 1865 19585 1985
rect 20100 1713 20200 1813
rect -400 1487 -300 1587
rect 215 1315 335 1435
rect 19465 1315 19585 1435
rect 215 765 335 885
rect 19465 765 19585 885
rect 20100 613 20200 713
rect -400 387 -300 487
rect 215 215 335 335
rect 765 215 885 335
rect 1315 215 1435 335
rect 1865 215 1985 335
rect 2415 215 2535 335
rect 2965 215 3085 335
rect 3515 215 3635 335
rect 4065 215 4185 335
rect 4615 215 4735 335
rect 5165 215 5285 335
rect 5715 215 5835 335
rect 6265 215 6385 335
rect 6815 215 6935 335
rect 7365 215 7485 335
rect 7915 215 8035 335
rect 8465 215 8585 335
rect 9015 215 9135 335
rect 9565 215 9685 335
rect 10115 215 10235 335
rect 10665 215 10785 335
rect 11215 215 11335 335
rect 11765 215 11885 335
rect 12315 215 12435 335
rect 12865 215 12985 335
rect 13415 215 13535 335
rect 13965 215 14085 335
rect 14515 215 14635 335
rect 15065 215 15185 335
rect 15615 215 15735 335
rect 16165 215 16285 335
rect 16715 215 16835 335
rect 17265 215 17385 335
rect 17815 215 17935 335
rect 18365 215 18485 335
rect 18915 215 19035 335
rect 19465 215 19585 335
rect 387 -400 487 -300
rect 1487 -400 1587 -300
rect 2587 -400 2687 -300
rect 3687 -400 3787 -300
rect 4787 -400 4887 -300
rect 5887 -400 5987 -300
rect 6987 -400 7087 -300
rect 8087 -400 8187 -300
rect 9187 -400 9287 -300
rect 10287 -400 10387 -300
rect 11387 -400 11487 -300
rect 12487 -400 12587 -300
rect 13587 -400 13687 -300
rect 14687 -400 14787 -300
rect 15787 -400 15887 -300
rect 16887 -400 16987 -300
rect 17987 -400 18087 -300
rect 19087 -400 19187 -300
<< metal4 >>
rect -2000 20800 19800 21800
rect -2000 19913 -1000 20800
rect -113 19913 339 20800
rect -2000 19589 339 19913
rect 437 20200 889 20300
rect 437 20100 613 20200
rect 713 20100 889 20200
rect 437 19687 889 20100
rect 987 19687 1439 20800
rect 1537 20200 1989 20300
rect 1537 20100 1713 20200
rect 1813 20100 1989 20200
rect 1537 19687 1989 20100
rect 2087 19687 2539 20800
rect 2637 20200 3089 20300
rect 2637 20100 2813 20200
rect 2913 20100 3089 20200
rect 2637 19687 3089 20100
rect 3187 19687 3639 20800
rect 3737 20200 4189 20300
rect 3737 20100 3913 20200
rect 4013 20100 4189 20200
rect 3737 19687 4189 20100
rect 4287 19687 4739 20800
rect 4837 20200 5289 20300
rect 4837 20100 5013 20200
rect 5113 20100 5289 20200
rect 4837 19687 5289 20100
rect 5387 19687 5839 20800
rect 5937 20200 6389 20300
rect 5937 20100 6113 20200
rect 6213 20100 6389 20200
rect 5937 19687 6389 20100
rect 6487 19687 6939 20800
rect 7037 20200 7489 20300
rect 7037 20100 7213 20200
rect 7313 20100 7489 20200
rect 7037 19687 7489 20100
rect 7587 19687 8039 20800
rect 8137 20200 8589 20300
rect 8137 20100 8313 20200
rect 8413 20100 8589 20200
rect 8137 19687 8589 20100
rect 8687 19687 9139 20800
rect 9237 20200 9689 20300
rect 9237 20100 9413 20200
rect 9513 20100 9689 20200
rect 9237 19687 9689 20100
rect 9787 19687 10239 20800
rect 10337 20200 10789 20300
rect 10337 20100 10513 20200
rect 10613 20100 10789 20200
rect 10337 19687 10789 20100
rect 10887 19687 11339 20800
rect 11437 20200 11889 20300
rect 11437 20100 11613 20200
rect 11713 20100 11889 20200
rect 11437 19687 11889 20100
rect 11987 19687 12439 20800
rect 12537 20200 12989 20300
rect 12537 20100 12713 20200
rect 12813 20100 12989 20200
rect 12537 19687 12989 20100
rect 13087 19687 13539 20800
rect 13637 20200 14089 20300
rect 13637 20100 13813 20200
rect 13913 20100 14089 20200
rect 13637 19687 14089 20100
rect 14187 19687 14639 20800
rect 14737 20200 15189 20300
rect 14737 20100 14913 20200
rect 15013 20100 15189 20200
rect 14737 19687 15189 20100
rect 15287 19687 15739 20800
rect 15837 20200 16289 20300
rect 15837 20100 16013 20200
rect 16113 20100 16289 20200
rect 15837 19687 16289 20100
rect 16387 19687 16839 20800
rect 16937 20200 17389 20300
rect 16937 20100 17113 20200
rect 17213 20100 17389 20200
rect 16937 19687 17389 20100
rect 17487 19687 17939 20800
rect 18037 20200 18489 20300
rect 18037 20100 18213 20200
rect 18313 20100 18489 20200
rect 18037 19687 18489 20100
rect 18587 19687 19039 20800
rect 19137 20200 19589 20300
rect 19137 20100 19313 20200
rect 19413 20100 19589 20200
rect 19137 19687 19589 20100
tri 339 19589 437 19687 sw
tri 437 19589 535 19687 ne
rect 535 19589 889 19687
tri 889 19589 987 19687 sw
tri 987 19589 1085 19687 ne
rect 1085 19589 1439 19687
tri 1439 19589 1537 19687 sw
tri 1537 19589 1635 19687 ne
rect 1635 19589 1989 19687
tri 1989 19589 2087 19687 sw
tri 2087 19589 2185 19687 ne
rect 2185 19589 2539 19687
tri 2539 19589 2637 19687 sw
tri 2637 19589 2735 19687 ne
rect 2735 19589 3089 19687
tri 3089 19589 3187 19687 sw
tri 3187 19589 3285 19687 ne
rect 3285 19589 3639 19687
tri 3639 19589 3737 19687 sw
tri 3737 19589 3835 19687 ne
rect 3835 19589 4189 19687
tri 4189 19589 4287 19687 sw
tri 4287 19589 4385 19687 ne
rect 4385 19589 4739 19687
tri 4739 19589 4837 19687 sw
tri 4837 19589 4935 19687 ne
rect 4935 19589 5289 19687
tri 5289 19589 5387 19687 sw
tri 5387 19589 5485 19687 ne
rect 5485 19589 5839 19687
tri 5839 19589 5937 19687 sw
tri 5937 19589 6035 19687 ne
rect 6035 19589 6389 19687
tri 6389 19589 6487 19687 sw
tri 6487 19589 6585 19687 ne
rect 6585 19589 6939 19687
tri 6939 19589 7037 19687 sw
tri 7037 19589 7135 19687 ne
rect 7135 19589 7489 19687
tri 7489 19589 7587 19687 sw
tri 7587 19589 7685 19687 ne
rect 7685 19589 8039 19687
tri 8039 19589 8137 19687 sw
tri 8137 19589 8235 19687 ne
rect 8235 19589 8589 19687
tri 8589 19589 8687 19687 sw
tri 8687 19589 8785 19687 ne
rect 8785 19589 9139 19687
tri 9139 19589 9237 19687 sw
tri 9237 19589 9335 19687 ne
rect 9335 19589 9689 19687
tri 9689 19589 9787 19687 sw
tri 9787 19589 9885 19687 ne
rect 9885 19589 10239 19687
tri 10239 19589 10337 19687 sw
tri 10337 19589 10435 19687 ne
rect 10435 19589 10789 19687
tri 10789 19589 10887 19687 sw
tri 10887 19589 10985 19687 ne
rect 10985 19589 11339 19687
tri 11339 19589 11437 19687 sw
tri 11437 19589 11535 19687 ne
rect 11535 19589 11889 19687
tri 11889 19589 11987 19687 sw
tri 11987 19589 12085 19687 ne
rect 12085 19589 12439 19687
tri 12439 19589 12537 19687 sw
tri 12537 19589 12635 19687 ne
rect 12635 19589 12989 19687
tri 12989 19589 13087 19687 sw
tri 13087 19589 13185 19687 ne
rect 13185 19589 13539 19687
tri 13539 19589 13637 19687 sw
tri 13637 19589 13735 19687 ne
rect 13735 19589 14089 19687
tri 14089 19589 14187 19687 sw
tri 14187 19589 14285 19687 ne
rect 14285 19589 14639 19687
tri 14639 19589 14737 19687 sw
tri 14737 19589 14835 19687 ne
rect 14835 19589 15189 19687
tri 15189 19589 15287 19687 sw
tri 15287 19589 15385 19687 ne
rect 15385 19589 15739 19687
tri 15739 19589 15837 19687 sw
tri 15837 19589 15935 19687 ne
rect 15935 19589 16289 19687
tri 16289 19589 16387 19687 sw
tri 16387 19589 16485 19687 ne
rect 16485 19589 16839 19687
tri 16839 19589 16937 19687 sw
tri 16937 19589 17035 19687 ne
rect 17035 19589 17389 19687
tri 17389 19589 17487 19687 sw
tri 17487 19589 17585 19687 ne
rect 17585 19589 17939 19687
tri 17939 19589 18037 19687 sw
tri 18037 19589 18135 19687 ne
rect 18135 19589 18489 19687
tri 18489 19589 18587 19687 sw
tri 18587 19589 18685 19687 ne
rect 18685 19589 19039 19687
tri 19039 19589 19137 19687 sw
tri 19137 19589 19235 19687 ne
rect 19235 19589 19589 19687
tri 19589 19589 19687 19687 sw
rect 20800 19589 21800 19800
rect -2000 19585 437 19589
rect -2000 19465 215 19585
rect 335 19491 437 19585
tri 437 19491 535 19589 sw
tri 535 19491 633 19589 ne
rect 633 19585 987 19589
rect 633 19491 765 19585
rect 335 19465 535 19491
rect -2000 19461 535 19465
rect -2000 18813 -1000 19461
tri 113 19363 211 19461 ne
rect 211 19413 535 19461
tri 535 19413 613 19491 sw
tri 633 19413 711 19491 ne
rect 711 19465 765 19491
rect 885 19491 987 19585
tri 987 19491 1085 19589 sw
tri 1085 19491 1183 19589 ne
rect 1183 19585 1537 19589
rect 1183 19491 1315 19585
rect 885 19465 1085 19491
rect 711 19413 1085 19465
tri 1085 19413 1163 19491 sw
tri 1183 19413 1261 19491 ne
rect 1261 19465 1315 19491
rect 1435 19491 1537 19585
tri 1537 19491 1635 19589 sw
tri 1635 19491 1733 19589 ne
rect 1733 19585 2087 19589
rect 1733 19491 1865 19585
rect 1435 19465 1635 19491
rect 1261 19413 1635 19465
tri 1635 19413 1713 19491 sw
tri 1733 19413 1811 19491 ne
rect 1811 19465 1865 19491
rect 1985 19491 2087 19585
tri 2087 19491 2185 19589 sw
tri 2185 19491 2283 19589 ne
rect 2283 19585 2637 19589
rect 2283 19491 2415 19585
rect 1985 19465 2185 19491
rect 1811 19413 2185 19465
tri 2185 19413 2263 19491 sw
tri 2283 19413 2361 19491 ne
rect 2361 19465 2415 19491
rect 2535 19491 2637 19585
tri 2637 19491 2735 19589 sw
tri 2735 19491 2833 19589 ne
rect 2833 19585 3187 19589
rect 2833 19491 2965 19585
rect 2535 19465 2735 19491
rect 2361 19413 2735 19465
tri 2735 19413 2813 19491 sw
tri 2833 19413 2911 19491 ne
rect 2911 19465 2965 19491
rect 3085 19491 3187 19585
tri 3187 19491 3285 19589 sw
tri 3285 19491 3383 19589 ne
rect 3383 19585 3737 19589
rect 3383 19491 3515 19585
rect 3085 19465 3285 19491
rect 2911 19413 3285 19465
tri 3285 19413 3363 19491 sw
tri 3383 19413 3461 19491 ne
rect 3461 19465 3515 19491
rect 3635 19491 3737 19585
tri 3737 19491 3835 19589 sw
tri 3835 19491 3933 19589 ne
rect 3933 19585 4287 19589
rect 3933 19491 4065 19585
rect 3635 19465 3835 19491
rect 3461 19413 3835 19465
tri 3835 19413 3913 19491 sw
tri 3933 19413 4011 19491 ne
rect 4011 19465 4065 19491
rect 4185 19491 4287 19585
tri 4287 19491 4385 19589 sw
tri 4385 19491 4483 19589 ne
rect 4483 19585 4837 19589
rect 4483 19491 4615 19585
rect 4185 19465 4385 19491
rect 4011 19413 4385 19465
tri 4385 19413 4463 19491 sw
tri 4483 19413 4561 19491 ne
rect 4561 19465 4615 19491
rect 4735 19491 4837 19585
tri 4837 19491 4935 19589 sw
tri 4935 19491 5033 19589 ne
rect 5033 19585 5387 19589
rect 5033 19491 5165 19585
rect 4735 19465 4935 19491
rect 4561 19413 4935 19465
tri 4935 19413 5013 19491 sw
tri 5033 19413 5111 19491 ne
rect 5111 19465 5165 19491
rect 5285 19491 5387 19585
tri 5387 19491 5485 19589 sw
tri 5485 19491 5583 19589 ne
rect 5583 19585 5937 19589
rect 5583 19491 5715 19585
rect 5285 19465 5485 19491
rect 5111 19413 5485 19465
tri 5485 19413 5563 19491 sw
tri 5583 19413 5661 19491 ne
rect 5661 19465 5715 19491
rect 5835 19491 5937 19585
tri 5937 19491 6035 19589 sw
tri 6035 19491 6133 19589 ne
rect 6133 19585 6487 19589
rect 6133 19491 6265 19585
rect 5835 19465 6035 19491
rect 5661 19413 6035 19465
tri 6035 19413 6113 19491 sw
tri 6133 19413 6211 19491 ne
rect 6211 19465 6265 19491
rect 6385 19491 6487 19585
tri 6487 19491 6585 19589 sw
tri 6585 19491 6683 19589 ne
rect 6683 19585 7037 19589
rect 6683 19491 6815 19585
rect 6385 19465 6585 19491
rect 6211 19413 6585 19465
tri 6585 19413 6663 19491 sw
tri 6683 19413 6761 19491 ne
rect 6761 19465 6815 19491
rect 6935 19491 7037 19585
tri 7037 19491 7135 19589 sw
tri 7135 19491 7233 19589 ne
rect 7233 19585 7587 19589
rect 7233 19491 7365 19585
rect 6935 19465 7135 19491
rect 6761 19413 7135 19465
tri 7135 19413 7213 19491 sw
tri 7233 19413 7311 19491 ne
rect 7311 19465 7365 19491
rect 7485 19491 7587 19585
tri 7587 19491 7685 19589 sw
tri 7685 19491 7783 19589 ne
rect 7783 19585 8137 19589
rect 7783 19491 7915 19585
rect 7485 19465 7685 19491
rect 7311 19413 7685 19465
tri 7685 19413 7763 19491 sw
tri 7783 19413 7861 19491 ne
rect 7861 19465 7915 19491
rect 8035 19491 8137 19585
tri 8137 19491 8235 19589 sw
tri 8235 19491 8333 19589 ne
rect 8333 19585 8687 19589
rect 8333 19491 8465 19585
rect 8035 19465 8235 19491
rect 7861 19413 8235 19465
tri 8235 19413 8313 19491 sw
tri 8333 19413 8411 19491 ne
rect 8411 19465 8465 19491
rect 8585 19491 8687 19585
tri 8687 19491 8785 19589 sw
tri 8785 19491 8883 19589 ne
rect 8883 19585 9237 19589
rect 8883 19491 9015 19585
rect 8585 19465 8785 19491
rect 8411 19413 8785 19465
tri 8785 19413 8863 19491 sw
tri 8883 19413 8961 19491 ne
rect 8961 19465 9015 19491
rect 9135 19491 9237 19585
tri 9237 19491 9335 19589 sw
tri 9335 19491 9433 19589 ne
rect 9433 19585 9787 19589
rect 9433 19491 9565 19585
rect 9135 19465 9335 19491
rect 8961 19413 9335 19465
tri 9335 19413 9413 19491 sw
tri 9433 19413 9511 19491 ne
rect 9511 19465 9565 19491
rect 9685 19491 9787 19585
tri 9787 19491 9885 19589 sw
tri 9885 19491 9983 19589 ne
rect 9983 19585 10337 19589
rect 9983 19491 10115 19585
rect 9685 19465 9885 19491
rect 9511 19413 9885 19465
tri 9885 19413 9963 19491 sw
tri 9983 19413 10061 19491 ne
rect 10061 19465 10115 19491
rect 10235 19491 10337 19585
tri 10337 19491 10435 19589 sw
tri 10435 19491 10533 19589 ne
rect 10533 19585 10887 19589
rect 10533 19491 10665 19585
rect 10235 19465 10435 19491
rect 10061 19413 10435 19465
tri 10435 19413 10513 19491 sw
tri 10533 19413 10611 19491 ne
rect 10611 19465 10665 19491
rect 10785 19491 10887 19585
tri 10887 19491 10985 19589 sw
tri 10985 19491 11083 19589 ne
rect 11083 19585 11437 19589
rect 11083 19491 11215 19585
rect 10785 19465 10985 19491
rect 10611 19413 10985 19465
tri 10985 19413 11063 19491 sw
tri 11083 19413 11161 19491 ne
rect 11161 19465 11215 19491
rect 11335 19491 11437 19585
tri 11437 19491 11535 19589 sw
tri 11535 19491 11633 19589 ne
rect 11633 19585 11987 19589
rect 11633 19491 11765 19585
rect 11335 19465 11535 19491
rect 11161 19413 11535 19465
tri 11535 19413 11613 19491 sw
tri 11633 19413 11711 19491 ne
rect 11711 19465 11765 19491
rect 11885 19491 11987 19585
tri 11987 19491 12085 19589 sw
tri 12085 19491 12183 19589 ne
rect 12183 19585 12537 19589
rect 12183 19491 12315 19585
rect 11885 19465 12085 19491
rect 11711 19413 12085 19465
tri 12085 19413 12163 19491 sw
tri 12183 19413 12261 19491 ne
rect 12261 19465 12315 19491
rect 12435 19491 12537 19585
tri 12537 19491 12635 19589 sw
tri 12635 19491 12733 19589 ne
rect 12733 19585 13087 19589
rect 12733 19491 12865 19585
rect 12435 19465 12635 19491
rect 12261 19413 12635 19465
tri 12635 19413 12713 19491 sw
tri 12733 19413 12811 19491 ne
rect 12811 19465 12865 19491
rect 12985 19491 13087 19585
tri 13087 19491 13185 19589 sw
tri 13185 19491 13283 19589 ne
rect 13283 19585 13637 19589
rect 13283 19491 13415 19585
rect 12985 19465 13185 19491
rect 12811 19413 13185 19465
tri 13185 19413 13263 19491 sw
tri 13283 19413 13361 19491 ne
rect 13361 19465 13415 19491
rect 13535 19491 13637 19585
tri 13637 19491 13735 19589 sw
tri 13735 19491 13833 19589 ne
rect 13833 19585 14187 19589
rect 13833 19491 13965 19585
rect 13535 19465 13735 19491
rect 13361 19413 13735 19465
tri 13735 19413 13813 19491 sw
tri 13833 19413 13911 19491 ne
rect 13911 19465 13965 19491
rect 14085 19491 14187 19585
tri 14187 19491 14285 19589 sw
tri 14285 19491 14383 19589 ne
rect 14383 19585 14737 19589
rect 14383 19491 14515 19585
rect 14085 19465 14285 19491
rect 13911 19413 14285 19465
tri 14285 19413 14363 19491 sw
tri 14383 19413 14461 19491 ne
rect 14461 19465 14515 19491
rect 14635 19491 14737 19585
tri 14737 19491 14835 19589 sw
tri 14835 19491 14933 19589 ne
rect 14933 19585 15287 19589
rect 14933 19491 15065 19585
rect 14635 19465 14835 19491
rect 14461 19413 14835 19465
tri 14835 19413 14913 19491 sw
tri 14933 19413 15011 19491 ne
rect 15011 19465 15065 19491
rect 15185 19491 15287 19585
tri 15287 19491 15385 19589 sw
tri 15385 19491 15483 19589 ne
rect 15483 19585 15837 19589
rect 15483 19491 15615 19585
rect 15185 19465 15385 19491
rect 15011 19413 15385 19465
tri 15385 19413 15463 19491 sw
tri 15483 19413 15561 19491 ne
rect 15561 19465 15615 19491
rect 15735 19491 15837 19585
tri 15837 19491 15935 19589 sw
tri 15935 19491 16033 19589 ne
rect 16033 19585 16387 19589
rect 16033 19491 16165 19585
rect 15735 19465 15935 19491
rect 15561 19413 15935 19465
tri 15935 19413 16013 19491 sw
tri 16033 19413 16111 19491 ne
rect 16111 19465 16165 19491
rect 16285 19491 16387 19585
tri 16387 19491 16485 19589 sw
tri 16485 19491 16583 19589 ne
rect 16583 19585 16937 19589
rect 16583 19491 16715 19585
rect 16285 19465 16485 19491
rect 16111 19413 16485 19465
tri 16485 19413 16563 19491 sw
tri 16583 19413 16661 19491 ne
rect 16661 19465 16715 19491
rect 16835 19491 16937 19585
tri 16937 19491 17035 19589 sw
tri 17035 19491 17133 19589 ne
rect 17133 19585 17487 19589
rect 17133 19491 17265 19585
rect 16835 19465 17035 19491
rect 16661 19413 17035 19465
tri 17035 19413 17113 19491 sw
tri 17133 19413 17211 19491 ne
rect 17211 19465 17265 19491
rect 17385 19491 17487 19585
tri 17487 19491 17585 19589 sw
tri 17585 19491 17683 19589 ne
rect 17683 19585 18037 19589
rect 17683 19491 17815 19585
rect 17385 19465 17585 19491
rect 17211 19413 17585 19465
tri 17585 19413 17663 19491 sw
tri 17683 19413 17761 19491 ne
rect 17761 19465 17815 19491
rect 17935 19491 18037 19585
tri 18037 19491 18135 19589 sw
tri 18135 19491 18233 19589 ne
rect 18233 19585 18587 19589
rect 18233 19491 18365 19585
rect 17935 19465 18135 19491
rect 17761 19413 18135 19465
tri 18135 19413 18213 19491 sw
tri 18233 19413 18311 19491 ne
rect 18311 19465 18365 19491
rect 18485 19491 18587 19585
tri 18587 19491 18685 19589 sw
tri 18685 19491 18783 19589 ne
rect 18783 19585 19137 19589
rect 18783 19491 18915 19585
rect 18485 19465 18685 19491
rect 18311 19413 18685 19465
tri 18685 19413 18763 19491 sw
tri 18783 19413 18861 19491 ne
rect 18861 19465 18915 19491
rect 19035 19491 19137 19585
tri 19137 19491 19235 19589 sw
tri 19235 19491 19333 19589 ne
rect 19333 19585 21800 19589
rect 19333 19491 19465 19585
rect 19035 19465 19235 19491
rect 18861 19413 19235 19465
tri 19235 19413 19313 19491 sw
tri 19333 19413 19411 19491 ne
rect 19411 19465 19465 19491
rect 19585 19465 21800 19585
rect 19411 19413 21800 19465
rect 211 19363 613 19413
rect -500 19313 113 19363
tri 113 19313 163 19363 sw
tri 211 19313 261 19363 ne
rect 261 19333 613 19363
tri 613 19333 693 19413 sw
tri 711 19333 791 19413 ne
rect 791 19333 1163 19413
tri 1163 19333 1243 19413 sw
tri 1261 19333 1341 19413 ne
rect 1341 19333 1713 19413
tri 1713 19333 1793 19413 sw
tri 1811 19333 1891 19413 ne
rect 1891 19333 2263 19413
tri 2263 19333 2343 19413 sw
tri 2361 19333 2441 19413 ne
rect 2441 19333 2813 19413
tri 2813 19333 2893 19413 sw
tri 2911 19333 2991 19413 ne
rect 2991 19333 3363 19413
tri 3363 19333 3443 19413 sw
tri 3461 19333 3541 19413 ne
rect 3541 19333 3913 19413
tri 3913 19333 3993 19413 sw
tri 4011 19333 4091 19413 ne
rect 4091 19333 4463 19413
tri 4463 19333 4543 19413 sw
tri 4561 19333 4641 19413 ne
rect 4641 19333 5013 19413
tri 5013 19333 5093 19413 sw
tri 5111 19333 5191 19413 ne
rect 5191 19333 5563 19413
tri 5563 19333 5643 19413 sw
tri 5661 19333 5741 19413 ne
rect 5741 19333 6113 19413
tri 6113 19333 6193 19413 sw
tri 6211 19333 6291 19413 ne
rect 6291 19333 6663 19413
tri 6663 19333 6743 19413 sw
tri 6761 19333 6841 19413 ne
rect 6841 19333 7213 19413
tri 7213 19333 7293 19413 sw
tri 7311 19333 7391 19413 ne
rect 7391 19333 7763 19413
tri 7763 19333 7843 19413 sw
tri 7861 19333 7941 19413 ne
rect 7941 19333 8313 19413
tri 8313 19333 8393 19413 sw
tri 8411 19333 8491 19413 ne
rect 8491 19333 8863 19413
tri 8863 19333 8943 19413 sw
tri 8961 19333 9041 19413 ne
rect 9041 19333 9413 19413
tri 9413 19333 9493 19413 sw
tri 9511 19333 9591 19413 ne
rect 9591 19333 9963 19413
tri 9963 19333 10043 19413 sw
tri 10061 19333 10141 19413 ne
rect 10141 19333 10513 19413
tri 10513 19333 10593 19413 sw
tri 10611 19333 10691 19413 ne
rect 10691 19333 11063 19413
tri 11063 19333 11143 19413 sw
tri 11161 19333 11241 19413 ne
rect 11241 19333 11613 19413
tri 11613 19333 11693 19413 sw
tri 11711 19333 11791 19413 ne
rect 11791 19333 12163 19413
tri 12163 19333 12243 19413 sw
tri 12261 19333 12341 19413 ne
rect 12341 19333 12713 19413
tri 12713 19333 12793 19413 sw
tri 12811 19333 12891 19413 ne
rect 12891 19333 13263 19413
tri 13263 19333 13343 19413 sw
tri 13361 19333 13441 19413 ne
rect 13441 19333 13813 19413
tri 13813 19333 13893 19413 sw
tri 13911 19333 13991 19413 ne
rect 13991 19333 14363 19413
tri 14363 19333 14443 19413 sw
tri 14461 19333 14541 19413 ne
rect 14541 19333 14913 19413
tri 14913 19333 14993 19413 sw
tri 15011 19333 15091 19413 ne
rect 15091 19333 15463 19413
tri 15463 19333 15543 19413 sw
tri 15561 19333 15641 19413 ne
rect 15641 19333 16013 19413
tri 16013 19333 16093 19413 sw
tri 16111 19333 16191 19413 ne
rect 16191 19333 16563 19413
tri 16563 19333 16643 19413 sw
tri 16661 19333 16741 19413 ne
rect 16741 19333 17113 19413
tri 17113 19333 17193 19413 sw
tri 17211 19333 17291 19413 ne
rect 17291 19333 17663 19413
tri 17663 19333 17743 19413 sw
tri 17761 19333 17841 19413 ne
rect 17841 19333 18213 19413
tri 18213 19333 18293 19413 sw
tri 18311 19333 18391 19413 ne
rect 18391 19333 18763 19413
tri 18763 19333 18843 19413 sw
tri 18861 19333 18941 19413 ne
rect 18941 19333 19313 19413
tri 19313 19333 19393 19413 sw
tri 19411 19333 19491 19413 ne
rect 19491 19333 20100 19413
rect 261 19313 693 19333
rect -500 19235 163 19313
tri 163 19235 241 19313 sw
tri 261 19235 339 19313 ne
rect 339 19235 693 19313
tri 693 19235 791 19333 sw
tri 791 19235 889 19333 ne
rect 889 19235 1243 19333
tri 1243 19235 1341 19333 sw
tri 1341 19235 1439 19333 ne
rect 1439 19235 1793 19333
tri 1793 19235 1891 19333 sw
tri 1891 19235 1989 19333 ne
rect 1989 19235 2343 19333
tri 2343 19235 2441 19333 sw
tri 2441 19235 2539 19333 ne
rect 2539 19235 2893 19333
tri 2893 19235 2991 19333 sw
tri 2991 19235 3089 19333 ne
rect 3089 19235 3443 19333
tri 3443 19235 3541 19333 sw
tri 3541 19235 3639 19333 ne
rect 3639 19235 3993 19333
tri 3993 19235 4091 19333 sw
tri 4091 19235 4189 19333 ne
rect 4189 19235 4543 19333
tri 4543 19235 4641 19333 sw
tri 4641 19235 4739 19333 ne
rect 4739 19235 5093 19333
tri 5093 19235 5191 19333 sw
tri 5191 19235 5289 19333 ne
rect 5289 19235 5643 19333
tri 5643 19235 5741 19333 sw
tri 5741 19235 5839 19333 ne
rect 5839 19235 6193 19333
tri 6193 19235 6291 19333 sw
tri 6291 19235 6389 19333 ne
rect 6389 19235 6743 19333
tri 6743 19235 6841 19333 sw
tri 6841 19235 6939 19333 ne
rect 6939 19235 7293 19333
tri 7293 19235 7391 19333 sw
tri 7391 19235 7489 19333 ne
rect 7489 19235 7843 19333
tri 7843 19235 7941 19333 sw
tri 7941 19235 8039 19333 ne
rect 8039 19235 8393 19333
tri 8393 19235 8491 19333 sw
tri 8491 19235 8589 19333 ne
rect 8589 19235 8943 19333
tri 8943 19235 9041 19333 sw
tri 9041 19235 9139 19333 ne
rect 9139 19235 9493 19333
tri 9493 19235 9591 19333 sw
tri 9591 19235 9689 19333 ne
rect 9689 19235 10043 19333
tri 10043 19235 10141 19333 sw
tri 10141 19235 10239 19333 ne
rect 10239 19235 10593 19333
tri 10593 19235 10691 19333 sw
tri 10691 19235 10789 19333 ne
rect 10789 19235 11143 19333
tri 11143 19235 11241 19333 sw
tri 11241 19235 11339 19333 ne
rect 11339 19235 11693 19333
tri 11693 19235 11791 19333 sw
tri 11791 19235 11889 19333 ne
rect 11889 19235 12243 19333
tri 12243 19235 12341 19333 sw
tri 12341 19235 12439 19333 ne
rect 12439 19235 12793 19333
tri 12793 19235 12891 19333 sw
tri 12891 19235 12989 19333 ne
rect 12989 19235 13343 19333
tri 13343 19235 13441 19333 sw
tri 13441 19235 13539 19333 ne
rect 13539 19235 13893 19333
tri 13893 19235 13991 19333 sw
tri 13991 19235 14089 19333 ne
rect 14089 19235 14443 19333
tri 14443 19235 14541 19333 sw
tri 14541 19235 14639 19333 ne
rect 14639 19235 14993 19333
tri 14993 19235 15091 19333 sw
tri 15091 19235 15189 19333 ne
rect 15189 19235 15543 19333
tri 15543 19235 15641 19333 sw
tri 15641 19235 15739 19333 ne
rect 15739 19235 16093 19333
tri 16093 19235 16191 19333 sw
tri 16191 19235 16289 19333 ne
rect 16289 19235 16643 19333
tri 16643 19235 16741 19333 sw
tri 16741 19235 16839 19333 ne
rect 16839 19235 17193 19333
tri 17193 19235 17291 19333 sw
tri 17291 19235 17389 19333 ne
rect 17389 19235 17743 19333
tri 17743 19235 17841 19333 sw
tri 17841 19235 17939 19333 ne
rect 17939 19235 18293 19333
tri 18293 19235 18391 19333 sw
tri 18391 19235 18489 19333 ne
rect 18489 19235 18843 19333
tri 18843 19235 18941 19333 sw
tri 18941 19235 19039 19333 ne
rect 19039 19235 19393 19333
tri 19393 19235 19491 19333 sw
tri 19491 19235 19589 19333 ne
rect 19589 19313 20100 19333
rect 20200 19313 21800 19413
rect 19589 19235 21800 19313
rect -500 19187 241 19235
rect -500 19087 -400 19187
rect -300 19137 241 19187
tri 241 19137 339 19235 sw
tri 339 19137 437 19235 ne
rect 437 19137 791 19235
tri 791 19137 889 19235 sw
tri 889 19137 987 19235 ne
rect 987 19137 1341 19235
tri 1341 19137 1439 19235 sw
tri 1439 19137 1537 19235 ne
rect 1537 19137 1891 19235
tri 1891 19137 1989 19235 sw
tri 1989 19137 2087 19235 ne
rect 2087 19137 2441 19235
tri 2441 19137 2539 19235 sw
tri 2539 19137 2637 19235 ne
rect 2637 19137 2991 19235
tri 2991 19137 3089 19235 sw
tri 3089 19137 3187 19235 ne
rect 3187 19137 3541 19235
tri 3541 19137 3639 19235 sw
tri 3639 19137 3737 19235 ne
rect 3737 19137 4091 19235
tri 4091 19137 4189 19235 sw
tri 4189 19137 4287 19235 ne
rect 4287 19137 4641 19235
tri 4641 19137 4739 19235 sw
tri 4739 19137 4837 19235 ne
rect 4837 19137 5191 19235
tri 5191 19137 5289 19235 sw
tri 5289 19137 5387 19235 ne
rect 5387 19137 5741 19235
tri 5741 19137 5839 19235 sw
tri 5839 19137 5937 19235 ne
rect 5937 19137 6291 19235
tri 6291 19137 6389 19235 sw
tri 6389 19137 6487 19235 ne
rect 6487 19137 6841 19235
tri 6841 19137 6939 19235 sw
tri 6939 19137 7037 19235 ne
rect 7037 19137 7391 19235
tri 7391 19137 7489 19235 sw
tri 7489 19137 7587 19235 ne
rect 7587 19137 7941 19235
tri 7941 19137 8039 19235 sw
tri 8039 19137 8137 19235 ne
rect 8137 19137 8491 19235
tri 8491 19137 8589 19235 sw
tri 8589 19137 8687 19235 ne
rect 8687 19137 9041 19235
tri 9041 19137 9139 19235 sw
tri 9139 19137 9237 19235 ne
rect 9237 19137 9591 19235
tri 9591 19137 9689 19235 sw
tri 9689 19137 9787 19235 ne
rect 9787 19137 10141 19235
tri 10141 19137 10239 19235 sw
tri 10239 19137 10337 19235 ne
rect 10337 19137 10691 19235
tri 10691 19137 10789 19235 sw
tri 10789 19137 10887 19235 ne
rect 10887 19137 11241 19235
tri 11241 19137 11339 19235 sw
tri 11339 19137 11437 19235 ne
rect 11437 19137 11791 19235
tri 11791 19137 11889 19235 sw
tri 11889 19137 11987 19235 ne
rect 11987 19137 12341 19235
tri 12341 19137 12439 19235 sw
tri 12439 19137 12537 19235 ne
rect 12537 19137 12891 19235
tri 12891 19137 12989 19235 sw
tri 12989 19137 13087 19235 ne
rect 13087 19137 13441 19235
tri 13441 19137 13539 19235 sw
tri 13539 19137 13637 19235 ne
rect 13637 19137 13991 19235
tri 13991 19137 14089 19235 sw
tri 14089 19137 14187 19235 ne
rect 14187 19137 14541 19235
tri 14541 19137 14639 19235 sw
tri 14639 19137 14737 19235 ne
rect 14737 19137 15091 19235
tri 15091 19137 15189 19235 sw
tri 15189 19137 15287 19235 ne
rect 15287 19137 15641 19235
tri 15641 19137 15739 19235 sw
tri 15739 19137 15837 19235 ne
rect 15837 19137 16191 19235
tri 16191 19137 16289 19235 sw
tri 16289 19137 16387 19235 ne
rect 16387 19137 16741 19235
tri 16741 19137 16839 19235 sw
tri 16839 19137 16937 19235 ne
rect 16937 19137 17291 19235
tri 17291 19137 17389 19235 sw
tri 17389 19137 17487 19235 ne
rect 17487 19137 17841 19235
tri 17841 19137 17939 19235 sw
tri 17939 19137 18037 19235 ne
rect 18037 19137 18391 19235
tri 18391 19137 18489 19235 sw
tri 18489 19137 18587 19235 ne
rect 18587 19137 18941 19235
tri 18941 19137 19039 19235 sw
tri 19039 19137 19137 19235 ne
rect 19137 19137 19491 19235
tri 19491 19137 19589 19235 sw
tri 19589 19137 19687 19235 ne
rect 19687 19137 21800 19235
rect -300 19087 339 19137
rect -500 19039 339 19087
tri 339 19039 437 19137 sw
tri 437 19039 535 19137 ne
rect 535 19039 889 19137
tri 889 19039 987 19137 sw
tri 987 19039 1085 19137 ne
rect 1085 19039 1439 19137
tri 1439 19039 1537 19137 sw
tri 1537 19039 1635 19137 ne
rect 1635 19039 1989 19137
tri 1989 19039 2087 19137 sw
tri 2087 19039 2185 19137 ne
rect 2185 19039 2539 19137
tri 2539 19039 2637 19137 sw
tri 2637 19039 2735 19137 ne
rect 2735 19039 3089 19137
tri 3089 19039 3187 19137 sw
tri 3187 19039 3285 19137 ne
rect 3285 19039 3639 19137
tri 3639 19039 3737 19137 sw
tri 3737 19039 3835 19137 ne
rect 3835 19039 4189 19137
tri 4189 19039 4287 19137 sw
tri 4287 19039 4385 19137 ne
rect 4385 19039 4739 19137
tri 4739 19039 4837 19137 sw
tri 4837 19039 4935 19137 ne
rect 4935 19039 5289 19137
tri 5289 19039 5387 19137 sw
tri 5387 19039 5485 19137 ne
rect 5485 19039 5839 19137
tri 5839 19039 5937 19137 sw
tri 5937 19039 6035 19137 ne
rect 6035 19039 6389 19137
tri 6389 19039 6487 19137 sw
tri 6487 19039 6585 19137 ne
rect 6585 19039 6939 19137
tri 6939 19039 7037 19137 sw
tri 7037 19039 7135 19137 ne
rect 7135 19039 7489 19137
tri 7489 19039 7587 19137 sw
tri 7587 19039 7685 19137 ne
rect 7685 19039 8039 19137
tri 8039 19039 8137 19137 sw
tri 8137 19039 8235 19137 ne
rect 8235 19039 8589 19137
tri 8589 19039 8687 19137 sw
tri 8687 19039 8785 19137 ne
rect 8785 19039 9139 19137
tri 9139 19039 9237 19137 sw
tri 9237 19039 9335 19137 ne
rect 9335 19039 9689 19137
tri 9689 19039 9787 19137 sw
tri 9787 19039 9885 19137 ne
rect 9885 19039 10239 19137
tri 10239 19039 10337 19137 sw
tri 10337 19039 10435 19137 ne
rect 10435 19039 10789 19137
tri 10789 19039 10887 19137 sw
tri 10887 19039 10985 19137 ne
rect 10985 19039 11339 19137
tri 11339 19039 11437 19137 sw
tri 11437 19039 11535 19137 ne
rect 11535 19039 11889 19137
tri 11889 19039 11987 19137 sw
tri 11987 19039 12085 19137 ne
rect 12085 19039 12439 19137
tri 12439 19039 12537 19137 sw
tri 12537 19039 12635 19137 ne
rect 12635 19039 12989 19137
tri 12989 19039 13087 19137 sw
tri 13087 19039 13185 19137 ne
rect 13185 19039 13539 19137
tri 13539 19039 13637 19137 sw
tri 13637 19039 13735 19137 ne
rect 13735 19039 14089 19137
tri 14089 19039 14187 19137 sw
tri 14187 19039 14285 19137 ne
rect 14285 19039 14639 19137
tri 14639 19039 14737 19137 sw
tri 14737 19039 14835 19137 ne
rect 14835 19039 15189 19137
tri 15189 19039 15287 19137 sw
tri 15287 19039 15385 19137 ne
rect 15385 19039 15739 19137
tri 15739 19039 15837 19137 sw
tri 15837 19039 15935 19137 ne
rect 15935 19039 16289 19137
tri 16289 19039 16387 19137 sw
tri 16387 19039 16485 19137 ne
rect 16485 19039 16839 19137
tri 16839 19039 16937 19137 sw
tri 16937 19039 17035 19137 ne
rect 17035 19039 17389 19137
tri 17389 19039 17487 19137 sw
tri 17487 19039 17585 19137 ne
rect 17585 19039 17939 19137
tri 17939 19039 18037 19137 sw
tri 18037 19039 18135 19137 ne
rect 18135 19039 18489 19137
tri 18489 19039 18587 19137 sw
tri 18587 19039 18685 19137 ne
rect 18685 19039 19039 19137
tri 19039 19039 19137 19137 sw
tri 19137 19039 19235 19137 ne
rect 19235 19039 19589 19137
tri 19589 19039 19687 19137 sw
rect -500 19035 437 19039
rect -500 18915 215 19035
rect 335 18941 437 19035
tri 437 18941 535 19039 sw
tri 535 18941 633 19039 ne
rect 633 19035 987 19039
rect 633 18941 765 19035
rect 335 18915 535 18941
rect -500 18911 535 18915
tri 535 18911 565 18941 sw
tri 633 18911 663 18941 ne
rect 663 18915 765 18941
rect 885 18941 987 19035
tri 987 18941 1085 19039 sw
tri 1085 18941 1183 19039 ne
rect 1183 19035 1537 19039
rect 1183 18941 1315 19035
rect 885 18915 1085 18941
rect 663 18911 1085 18915
tri 1085 18911 1115 18941 sw
tri 1183 18911 1213 18941 ne
rect 1213 18915 1315 18941
rect 1435 18941 1537 19035
tri 1537 18941 1635 19039 sw
tri 1635 18941 1733 19039 ne
rect 1733 19035 2087 19039
rect 1733 18941 1865 19035
rect 1435 18915 1635 18941
rect 1213 18911 1635 18915
tri 1635 18911 1665 18941 sw
tri 1733 18911 1763 18941 ne
rect 1763 18915 1865 18941
rect 1985 18941 2087 19035
tri 2087 18941 2185 19039 sw
tri 2185 18941 2283 19039 ne
rect 2283 19035 2637 19039
rect 2283 18941 2415 19035
rect 1985 18915 2185 18941
rect 1763 18911 2185 18915
tri 2185 18911 2215 18941 sw
tri 2283 18911 2313 18941 ne
rect 2313 18915 2415 18941
rect 2535 18941 2637 19035
tri 2637 18941 2735 19039 sw
tri 2735 18941 2833 19039 ne
rect 2833 19035 3187 19039
rect 2833 18941 2965 19035
rect 2535 18915 2735 18941
rect 2313 18911 2735 18915
tri 2735 18911 2765 18941 sw
tri 2833 18911 2863 18941 ne
rect 2863 18915 2965 18941
rect 3085 18941 3187 19035
tri 3187 18941 3285 19039 sw
tri 3285 18941 3383 19039 ne
rect 3383 19035 3737 19039
rect 3383 18941 3515 19035
rect 3085 18915 3285 18941
rect 2863 18911 3285 18915
tri 3285 18911 3315 18941 sw
tri 3383 18911 3413 18941 ne
rect 3413 18915 3515 18941
rect 3635 18941 3737 19035
tri 3737 18941 3835 19039 sw
tri 3835 18941 3933 19039 ne
rect 3933 19035 4287 19039
rect 3933 18941 4065 19035
rect 3635 18915 3835 18941
rect 3413 18911 3835 18915
tri 3835 18911 3865 18941 sw
tri 3933 18911 3963 18941 ne
rect 3963 18915 4065 18941
rect 4185 18941 4287 19035
tri 4287 18941 4385 19039 sw
tri 4385 18941 4483 19039 ne
rect 4483 19035 4837 19039
rect 4483 18941 4615 19035
rect 4185 18915 4385 18941
rect 3963 18911 4385 18915
tri 4385 18911 4415 18941 sw
tri 4483 18911 4513 18941 ne
rect 4513 18915 4615 18941
rect 4735 18941 4837 19035
tri 4837 18941 4935 19039 sw
tri 4935 18941 5033 19039 ne
rect 5033 19035 5387 19039
rect 5033 18941 5165 19035
rect 4735 18915 4935 18941
rect 4513 18911 4935 18915
tri 4935 18911 4965 18941 sw
tri 5033 18911 5063 18941 ne
rect 5063 18915 5165 18941
rect 5285 18941 5387 19035
tri 5387 18941 5485 19039 sw
tri 5485 18941 5583 19039 ne
rect 5583 19035 5937 19039
rect 5583 18941 5715 19035
rect 5285 18915 5485 18941
rect 5063 18911 5485 18915
tri 5485 18911 5515 18941 sw
tri 5583 18911 5613 18941 ne
rect 5613 18915 5715 18941
rect 5835 18941 5937 19035
tri 5937 18941 6035 19039 sw
tri 6035 18941 6133 19039 ne
rect 6133 19035 6487 19039
rect 6133 18941 6265 19035
rect 5835 18915 6035 18941
rect 5613 18911 6035 18915
tri 6035 18911 6065 18941 sw
tri 6133 18911 6163 18941 ne
rect 6163 18915 6265 18941
rect 6385 18941 6487 19035
tri 6487 18941 6585 19039 sw
tri 6585 18941 6683 19039 ne
rect 6683 19035 7037 19039
rect 6683 18941 6815 19035
rect 6385 18915 6585 18941
rect 6163 18911 6585 18915
tri 6585 18911 6615 18941 sw
tri 6683 18911 6713 18941 ne
rect 6713 18915 6815 18941
rect 6935 18941 7037 19035
tri 7037 18941 7135 19039 sw
tri 7135 18941 7233 19039 ne
rect 7233 19035 7587 19039
rect 7233 18941 7365 19035
rect 6935 18915 7135 18941
rect 6713 18911 7135 18915
tri 7135 18911 7165 18941 sw
tri 7233 18911 7263 18941 ne
rect 7263 18915 7365 18941
rect 7485 18941 7587 19035
tri 7587 18941 7685 19039 sw
tri 7685 18941 7783 19039 ne
rect 7783 19035 8137 19039
rect 7783 18941 7915 19035
rect 7485 18915 7685 18941
rect 7263 18911 7685 18915
tri 7685 18911 7715 18941 sw
tri 7783 18911 7813 18941 ne
rect 7813 18915 7915 18941
rect 8035 18941 8137 19035
tri 8137 18941 8235 19039 sw
tri 8235 18941 8333 19039 ne
rect 8333 19035 8687 19039
rect 8333 18941 8465 19035
rect 8035 18915 8235 18941
rect 7813 18911 8235 18915
tri 8235 18911 8265 18941 sw
tri 8333 18911 8363 18941 ne
rect 8363 18915 8465 18941
rect 8585 18941 8687 19035
tri 8687 18941 8785 19039 sw
tri 8785 18941 8883 19039 ne
rect 8883 19035 9237 19039
rect 8883 18941 9015 19035
rect 8585 18915 8785 18941
rect 8363 18911 8785 18915
tri 8785 18911 8815 18941 sw
tri 8883 18911 8913 18941 ne
rect 8913 18915 9015 18941
rect 9135 18941 9237 19035
tri 9237 18941 9335 19039 sw
tri 9335 18941 9433 19039 ne
rect 9433 19035 9787 19039
rect 9433 18941 9565 19035
rect 9135 18915 9335 18941
rect 8913 18911 9335 18915
tri 9335 18911 9365 18941 sw
tri 9433 18911 9463 18941 ne
rect 9463 18915 9565 18941
rect 9685 18941 9787 19035
tri 9787 18941 9885 19039 sw
tri 9885 18941 9983 19039 ne
rect 9983 19035 10337 19039
rect 9983 18941 10115 19035
rect 9685 18915 9885 18941
rect 9463 18911 9885 18915
tri 9885 18911 9915 18941 sw
tri 9983 18911 10013 18941 ne
rect 10013 18915 10115 18941
rect 10235 18941 10337 19035
tri 10337 18941 10435 19039 sw
tri 10435 18941 10533 19039 ne
rect 10533 19035 10887 19039
rect 10533 18941 10665 19035
rect 10235 18915 10435 18941
rect 10013 18911 10435 18915
tri 10435 18911 10465 18941 sw
tri 10533 18911 10563 18941 ne
rect 10563 18915 10665 18941
rect 10785 18941 10887 19035
tri 10887 18941 10985 19039 sw
tri 10985 18941 11083 19039 ne
rect 11083 19035 11437 19039
rect 11083 18941 11215 19035
rect 10785 18915 10985 18941
rect 10563 18911 10985 18915
tri 10985 18911 11015 18941 sw
tri 11083 18911 11113 18941 ne
rect 11113 18915 11215 18941
rect 11335 18941 11437 19035
tri 11437 18941 11535 19039 sw
tri 11535 18941 11633 19039 ne
rect 11633 19035 11987 19039
rect 11633 18941 11765 19035
rect 11335 18915 11535 18941
rect 11113 18911 11535 18915
tri 11535 18911 11565 18941 sw
tri 11633 18911 11663 18941 ne
rect 11663 18915 11765 18941
rect 11885 18941 11987 19035
tri 11987 18941 12085 19039 sw
tri 12085 18941 12183 19039 ne
rect 12183 19035 12537 19039
rect 12183 18941 12315 19035
rect 11885 18915 12085 18941
rect 11663 18911 12085 18915
tri 12085 18911 12115 18941 sw
tri 12183 18911 12213 18941 ne
rect 12213 18915 12315 18941
rect 12435 18941 12537 19035
tri 12537 18941 12635 19039 sw
tri 12635 18941 12733 19039 ne
rect 12733 19035 13087 19039
rect 12733 18941 12865 19035
rect 12435 18915 12635 18941
rect 12213 18911 12635 18915
tri 12635 18911 12665 18941 sw
tri 12733 18911 12763 18941 ne
rect 12763 18915 12865 18941
rect 12985 18941 13087 19035
tri 13087 18941 13185 19039 sw
tri 13185 18941 13283 19039 ne
rect 13283 19035 13637 19039
rect 13283 18941 13415 19035
rect 12985 18915 13185 18941
rect 12763 18911 13185 18915
tri 13185 18911 13215 18941 sw
tri 13283 18911 13313 18941 ne
rect 13313 18915 13415 18941
rect 13535 18941 13637 19035
tri 13637 18941 13735 19039 sw
tri 13735 18941 13833 19039 ne
rect 13833 19035 14187 19039
rect 13833 18941 13965 19035
rect 13535 18915 13735 18941
rect 13313 18911 13735 18915
tri 13735 18911 13765 18941 sw
tri 13833 18911 13863 18941 ne
rect 13863 18915 13965 18941
rect 14085 18941 14187 19035
tri 14187 18941 14285 19039 sw
tri 14285 18941 14383 19039 ne
rect 14383 19035 14737 19039
rect 14383 18941 14515 19035
rect 14085 18915 14285 18941
rect 13863 18911 14285 18915
tri 14285 18911 14315 18941 sw
tri 14383 18911 14413 18941 ne
rect 14413 18915 14515 18941
rect 14635 18941 14737 19035
tri 14737 18941 14835 19039 sw
tri 14835 18941 14933 19039 ne
rect 14933 19035 15287 19039
rect 14933 18941 15065 19035
rect 14635 18915 14835 18941
rect 14413 18911 14835 18915
tri 14835 18911 14865 18941 sw
tri 14933 18911 14963 18941 ne
rect 14963 18915 15065 18941
rect 15185 18941 15287 19035
tri 15287 18941 15385 19039 sw
tri 15385 18941 15483 19039 ne
rect 15483 19035 15837 19039
rect 15483 18941 15615 19035
rect 15185 18915 15385 18941
rect 14963 18911 15385 18915
tri 15385 18911 15415 18941 sw
tri 15483 18911 15513 18941 ne
rect 15513 18915 15615 18941
rect 15735 18941 15837 19035
tri 15837 18941 15935 19039 sw
tri 15935 18941 16033 19039 ne
rect 16033 19035 16387 19039
rect 16033 18941 16165 19035
rect 15735 18915 15935 18941
rect 15513 18911 15935 18915
tri 15935 18911 15965 18941 sw
tri 16033 18911 16063 18941 ne
rect 16063 18915 16165 18941
rect 16285 18941 16387 19035
tri 16387 18941 16485 19039 sw
tri 16485 18941 16583 19039 ne
rect 16583 19035 16937 19039
rect 16583 18941 16715 19035
rect 16285 18915 16485 18941
rect 16063 18911 16485 18915
tri 16485 18911 16515 18941 sw
tri 16583 18911 16613 18941 ne
rect 16613 18915 16715 18941
rect 16835 18941 16937 19035
tri 16937 18941 17035 19039 sw
tri 17035 18941 17133 19039 ne
rect 17133 19035 17487 19039
rect 17133 18941 17265 19035
rect 16835 18915 17035 18941
rect 16613 18911 17035 18915
tri 17035 18911 17065 18941 sw
tri 17133 18911 17163 18941 ne
rect 17163 18915 17265 18941
rect 17385 18941 17487 19035
tri 17487 18941 17585 19039 sw
tri 17585 18941 17683 19039 ne
rect 17683 19035 18037 19039
rect 17683 18941 17815 19035
rect 17385 18915 17585 18941
rect 17163 18911 17585 18915
tri 17585 18911 17615 18941 sw
tri 17683 18911 17713 18941 ne
rect 17713 18915 17815 18941
rect 17935 18941 18037 19035
tri 18037 18941 18135 19039 sw
tri 18135 18941 18233 19039 ne
rect 18233 19035 18587 19039
rect 18233 18941 18365 19035
rect 17935 18915 18135 18941
rect 17713 18911 18135 18915
tri 18135 18911 18165 18941 sw
tri 18233 18911 18263 18941 ne
rect 18263 18915 18365 18941
rect 18485 18941 18587 19035
tri 18587 18941 18685 19039 sw
tri 18685 18941 18783 19039 ne
rect 18783 19035 19137 19039
rect 18783 18941 18915 19035
rect 18485 18915 18685 18941
rect 18263 18911 18685 18915
tri 18685 18911 18715 18941 sw
tri 18783 18911 18813 18941 ne
rect 18813 18915 18915 18941
rect 19035 18941 19137 19035
tri 19137 18941 19235 19039 sw
tri 19235 18941 19333 19039 ne
rect 19333 19035 20300 19039
rect 19333 18941 19465 19035
rect 19035 18915 19235 18941
rect 18813 18911 19235 18915
tri 19235 18911 19265 18941 sw
tri 19333 18911 19363 18941 ne
rect 19363 18915 19465 18941
rect 19585 18915 20300 19035
rect 19363 18911 20300 18915
tri 113 18813 211 18911 ne
rect 211 18813 565 18911
tri 565 18813 663 18911 sw
tri 663 18813 761 18911 ne
rect 761 18813 1115 18911
tri 1115 18813 1213 18911 sw
tri 1213 18813 1311 18911 ne
rect 1311 18813 1665 18911
tri 1665 18813 1763 18911 sw
tri 1763 18813 1861 18911 ne
rect 1861 18813 2215 18911
tri 2215 18813 2313 18911 sw
tri 2313 18813 2411 18911 ne
rect 2411 18813 2765 18911
tri 2765 18813 2863 18911 sw
tri 2863 18813 2961 18911 ne
rect 2961 18813 3315 18911
tri 3315 18813 3413 18911 sw
tri 3413 18813 3511 18911 ne
rect 3511 18813 3865 18911
tri 3865 18813 3963 18911 sw
tri 3963 18813 4061 18911 ne
rect 4061 18813 4415 18911
tri 4415 18813 4513 18911 sw
tri 4513 18813 4611 18911 ne
rect 4611 18813 4965 18911
tri 4965 18813 5063 18911 sw
tri 5063 18813 5161 18911 ne
rect 5161 18813 5515 18911
tri 5515 18813 5613 18911 sw
tri 5613 18813 5711 18911 ne
rect 5711 18813 6065 18911
tri 6065 18813 6163 18911 sw
tri 6163 18813 6261 18911 ne
rect 6261 18813 6615 18911
tri 6615 18813 6713 18911 sw
tri 6713 18813 6811 18911 ne
rect 6811 18813 7165 18911
tri 7165 18813 7263 18911 sw
tri 7263 18813 7361 18911 ne
rect 7361 18813 7715 18911
tri 7715 18813 7813 18911 sw
tri 7813 18813 7911 18911 ne
rect 7911 18813 8265 18911
tri 8265 18813 8363 18911 sw
tri 8363 18813 8461 18911 ne
rect 8461 18813 8815 18911
tri 8815 18813 8913 18911 sw
tri 8913 18813 9011 18911 ne
rect 9011 18813 9365 18911
tri 9365 18813 9463 18911 sw
tri 9463 18813 9561 18911 ne
rect 9561 18813 9915 18911
tri 9915 18813 10013 18911 sw
tri 10013 18813 10111 18911 ne
rect 10111 18813 10465 18911
tri 10465 18813 10563 18911 sw
tri 10563 18813 10661 18911 ne
rect 10661 18813 11015 18911
tri 11015 18813 11113 18911 sw
tri 11113 18813 11211 18911 ne
rect 11211 18813 11565 18911
tri 11565 18813 11663 18911 sw
tri 11663 18813 11761 18911 ne
rect 11761 18813 12115 18911
tri 12115 18813 12213 18911 sw
tri 12213 18813 12311 18911 ne
rect 12311 18813 12665 18911
tri 12665 18813 12763 18911 sw
tri 12763 18813 12861 18911 ne
rect 12861 18813 13215 18911
tri 13215 18813 13313 18911 sw
tri 13313 18813 13411 18911 ne
rect 13411 18813 13765 18911
tri 13765 18813 13863 18911 sw
tri 13863 18813 13961 18911 ne
rect 13961 18813 14315 18911
tri 14315 18813 14413 18911 sw
tri 14413 18813 14511 18911 ne
rect 14511 18813 14865 18911
tri 14865 18813 14963 18911 sw
tri 14963 18813 15061 18911 ne
rect 15061 18813 15415 18911
tri 15415 18813 15513 18911 sw
tri 15513 18813 15611 18911 ne
rect 15611 18813 15965 18911
tri 15965 18813 16063 18911 sw
tri 16063 18813 16161 18911 ne
rect 16161 18813 16515 18911
tri 16515 18813 16613 18911 sw
tri 16613 18813 16711 18911 ne
rect 16711 18813 17065 18911
tri 17065 18813 17163 18911 sw
tri 17163 18813 17261 18911 ne
rect 17261 18813 17615 18911
tri 17615 18813 17713 18911 sw
tri 17713 18813 17811 18911 ne
rect 17811 18813 18165 18911
tri 18165 18813 18263 18911 sw
tri 18263 18813 18361 18911 ne
rect 18361 18813 18715 18911
tri 18715 18813 18813 18911 sw
tri 18813 18813 18911 18911 ne
rect 18911 18813 19265 18911
tri 19265 18813 19363 18911 sw
tri 19363 18813 19461 18911 ne
rect 19461 18813 20300 18911
rect -2000 18783 113 18813
tri 113 18783 143 18813 sw
tri 211 18783 241 18813 ne
rect 241 18783 663 18813
tri 663 18783 693 18813 sw
tri 761 18783 791 18813 ne
rect 791 18783 1213 18813
tri 1213 18783 1243 18813 sw
tri 1311 18783 1341 18813 ne
rect 1341 18783 1763 18813
tri 1763 18783 1793 18813 sw
tri 1861 18783 1891 18813 ne
rect 1891 18783 2313 18813
tri 2313 18783 2343 18813 sw
tri 2411 18783 2441 18813 ne
rect 2441 18783 2863 18813
tri 2863 18783 2893 18813 sw
tri 2961 18783 2991 18813 ne
rect 2991 18783 3413 18813
tri 3413 18783 3443 18813 sw
tri 3511 18783 3541 18813 ne
rect 3541 18783 3963 18813
tri 3963 18783 3993 18813 sw
tri 4061 18783 4091 18813 ne
rect 4091 18783 4513 18813
tri 4513 18783 4543 18813 sw
tri 4611 18783 4641 18813 ne
rect 4641 18783 5063 18813
tri 5063 18783 5093 18813 sw
tri 5161 18783 5191 18813 ne
rect 5191 18783 5613 18813
tri 5613 18783 5643 18813 sw
tri 5711 18783 5741 18813 ne
rect 5741 18783 6163 18813
tri 6163 18783 6193 18813 sw
tri 6261 18783 6291 18813 ne
rect 6291 18783 6713 18813
tri 6713 18783 6743 18813 sw
tri 6811 18783 6841 18813 ne
rect 6841 18783 7263 18813
tri 7263 18783 7293 18813 sw
tri 7361 18783 7391 18813 ne
rect 7391 18783 7813 18813
tri 7813 18783 7843 18813 sw
tri 7911 18783 7941 18813 ne
rect 7941 18783 8363 18813
tri 8363 18783 8393 18813 sw
tri 8461 18783 8491 18813 ne
rect 8491 18783 8913 18813
tri 8913 18783 8943 18813 sw
tri 9011 18783 9041 18813 ne
rect 9041 18783 9463 18813
tri 9463 18783 9493 18813 sw
tri 9561 18783 9591 18813 ne
rect 9591 18783 10013 18813
tri 10013 18783 10043 18813 sw
tri 10111 18783 10141 18813 ne
rect 10141 18783 10563 18813
tri 10563 18783 10593 18813 sw
tri 10661 18783 10691 18813 ne
rect 10691 18783 11113 18813
tri 11113 18783 11143 18813 sw
tri 11211 18783 11241 18813 ne
rect 11241 18783 11663 18813
tri 11663 18783 11693 18813 sw
tri 11761 18783 11791 18813 ne
rect 11791 18783 12213 18813
tri 12213 18783 12243 18813 sw
tri 12311 18783 12341 18813 ne
rect 12341 18783 12763 18813
tri 12763 18783 12793 18813 sw
tri 12861 18783 12891 18813 ne
rect 12891 18783 13313 18813
tri 13313 18783 13343 18813 sw
tri 13411 18783 13441 18813 ne
rect 13441 18783 13863 18813
tri 13863 18783 13893 18813 sw
tri 13961 18783 13991 18813 ne
rect 13991 18783 14413 18813
tri 14413 18783 14443 18813 sw
tri 14511 18783 14541 18813 ne
rect 14541 18783 14963 18813
tri 14963 18783 14993 18813 sw
tri 15061 18783 15091 18813 ne
rect 15091 18783 15513 18813
tri 15513 18783 15543 18813 sw
tri 15611 18783 15641 18813 ne
rect 15641 18783 16063 18813
tri 16063 18783 16093 18813 sw
tri 16161 18783 16191 18813 ne
rect 16191 18783 16613 18813
tri 16613 18783 16643 18813 sw
tri 16711 18783 16741 18813 ne
rect 16741 18783 17163 18813
tri 17163 18783 17193 18813 sw
tri 17261 18783 17291 18813 ne
rect 17291 18783 17713 18813
tri 17713 18783 17743 18813 sw
tri 17811 18783 17841 18813 ne
rect 17841 18783 18263 18813
tri 18263 18783 18293 18813 sw
tri 18361 18783 18391 18813 ne
rect 18391 18783 18813 18813
tri 18813 18783 18843 18813 sw
tri 18911 18783 18941 18813 ne
rect 18941 18783 19363 18813
tri 19363 18783 19393 18813 sw
tri 19461 18783 19491 18813 ne
rect 19491 18783 20300 18813
rect -2000 18685 143 18783
tri 143 18685 241 18783 sw
tri 241 18685 339 18783 ne
rect 339 18685 693 18783
tri 693 18685 791 18783 sw
tri 791 18685 889 18783 ne
rect 889 18685 1243 18783
tri 1243 18685 1341 18783 sw
tri 1341 18685 1439 18783 ne
rect 1439 18685 1793 18783
tri 1793 18685 1891 18783 sw
tri 1891 18685 1989 18783 ne
rect 1989 18685 2343 18783
tri 2343 18685 2441 18783 sw
tri 2441 18685 2539 18783 ne
rect 2539 18685 2893 18783
tri 2893 18685 2991 18783 sw
tri 2991 18685 3089 18783 ne
rect 3089 18685 3443 18783
tri 3443 18685 3541 18783 sw
tri 3541 18685 3639 18783 ne
rect 3639 18685 3993 18783
tri 3993 18685 4091 18783 sw
tri 4091 18685 4189 18783 ne
rect 4189 18685 4543 18783
tri 4543 18685 4641 18783 sw
tri 4641 18685 4739 18783 ne
rect 4739 18685 5093 18783
tri 5093 18685 5191 18783 sw
tri 5191 18685 5289 18783 ne
rect 5289 18685 5643 18783
tri 5643 18685 5741 18783 sw
tri 5741 18685 5839 18783 ne
rect 5839 18685 6193 18783
tri 6193 18685 6291 18783 sw
tri 6291 18685 6389 18783 ne
rect 6389 18685 6743 18783
tri 6743 18685 6841 18783 sw
tri 6841 18685 6939 18783 ne
rect 6939 18685 7293 18783
tri 7293 18685 7391 18783 sw
tri 7391 18685 7489 18783 ne
rect 7489 18685 7843 18783
tri 7843 18685 7941 18783 sw
tri 7941 18685 8039 18783 ne
rect 8039 18685 8393 18783
tri 8393 18685 8491 18783 sw
tri 8491 18685 8589 18783 ne
rect 8589 18685 8943 18783
tri 8943 18685 9041 18783 sw
tri 9041 18685 9139 18783 ne
rect 9139 18685 9493 18783
tri 9493 18685 9591 18783 sw
tri 9591 18685 9689 18783 ne
rect 9689 18685 10043 18783
tri 10043 18685 10141 18783 sw
tri 10141 18685 10239 18783 ne
rect 10239 18685 10593 18783
tri 10593 18685 10691 18783 sw
tri 10691 18685 10789 18783 ne
rect 10789 18685 11143 18783
tri 11143 18685 11241 18783 sw
tri 11241 18685 11339 18783 ne
rect 11339 18685 11693 18783
tri 11693 18685 11791 18783 sw
tri 11791 18685 11889 18783 ne
rect 11889 18685 12243 18783
tri 12243 18685 12341 18783 sw
tri 12341 18685 12439 18783 ne
rect 12439 18685 12793 18783
tri 12793 18685 12891 18783 sw
tri 12891 18685 12989 18783 ne
rect 12989 18685 13343 18783
tri 13343 18685 13441 18783 sw
tri 13441 18685 13539 18783 ne
rect 13539 18685 13893 18783
tri 13893 18685 13991 18783 sw
tri 13991 18685 14089 18783 ne
rect 14089 18685 14443 18783
tri 14443 18685 14541 18783 sw
tri 14541 18685 14639 18783 ne
rect 14639 18685 14993 18783
tri 14993 18685 15091 18783 sw
tri 15091 18685 15189 18783 ne
rect 15189 18685 15543 18783
tri 15543 18685 15641 18783 sw
tri 15641 18685 15739 18783 ne
rect 15739 18685 16093 18783
tri 16093 18685 16191 18783 sw
tri 16191 18685 16289 18783 ne
rect 16289 18685 16643 18783
tri 16643 18685 16741 18783 sw
tri 16741 18685 16839 18783 ne
rect 16839 18685 17193 18783
tri 17193 18685 17291 18783 sw
tri 17291 18685 17389 18783 ne
rect 17389 18685 17743 18783
tri 17743 18685 17841 18783 sw
tri 17841 18685 17939 18783 ne
rect 17939 18685 18293 18783
tri 18293 18685 18391 18783 sw
tri 18391 18685 18489 18783 ne
rect 18489 18685 18843 18783
tri 18843 18685 18941 18783 sw
tri 18941 18685 19039 18783 ne
rect 19039 18685 19393 18783
tri 19393 18685 19491 18783 sw
tri 19491 18685 19589 18783 ne
rect 19589 18685 20300 18783
rect -2000 18587 241 18685
tri 241 18587 339 18685 sw
tri 339 18587 437 18685 ne
rect 437 18587 791 18685
tri 791 18587 889 18685 sw
tri 889 18587 987 18685 ne
rect 987 18587 1341 18685
tri 1341 18587 1439 18685 sw
tri 1439 18587 1537 18685 ne
rect 1537 18587 1891 18685
tri 1891 18587 1989 18685 sw
tri 1989 18587 2087 18685 ne
rect 2087 18587 2441 18685
tri 2441 18587 2539 18685 sw
tri 2539 18587 2637 18685 ne
rect 2637 18587 2991 18685
tri 2991 18587 3089 18685 sw
tri 3089 18587 3187 18685 ne
rect 3187 18587 3541 18685
tri 3541 18587 3639 18685 sw
tri 3639 18587 3737 18685 ne
rect 3737 18587 4091 18685
tri 4091 18587 4189 18685 sw
tri 4189 18587 4287 18685 ne
rect 4287 18587 4641 18685
tri 4641 18587 4739 18685 sw
tri 4739 18587 4837 18685 ne
rect 4837 18587 5191 18685
tri 5191 18587 5289 18685 sw
tri 5289 18587 5387 18685 ne
rect 5387 18587 5741 18685
tri 5741 18587 5839 18685 sw
tri 5839 18587 5937 18685 ne
rect 5937 18587 6291 18685
tri 6291 18587 6389 18685 sw
tri 6389 18587 6487 18685 ne
rect 6487 18587 6841 18685
tri 6841 18587 6939 18685 sw
tri 6939 18587 7037 18685 ne
rect 7037 18587 7391 18685
tri 7391 18587 7489 18685 sw
tri 7489 18587 7587 18685 ne
rect 7587 18587 7941 18685
tri 7941 18587 8039 18685 sw
tri 8039 18587 8137 18685 ne
rect 8137 18587 8491 18685
tri 8491 18587 8589 18685 sw
tri 8589 18587 8687 18685 ne
rect 8687 18587 9041 18685
tri 9041 18587 9139 18685 sw
tri 9139 18587 9237 18685 ne
rect 9237 18587 9591 18685
tri 9591 18587 9689 18685 sw
tri 9689 18587 9787 18685 ne
rect 9787 18587 10141 18685
tri 10141 18587 10239 18685 sw
tri 10239 18587 10337 18685 ne
rect 10337 18587 10691 18685
tri 10691 18587 10789 18685 sw
tri 10789 18587 10887 18685 ne
rect 10887 18587 11241 18685
tri 11241 18587 11339 18685 sw
tri 11339 18587 11437 18685 ne
rect 11437 18587 11791 18685
tri 11791 18587 11889 18685 sw
tri 11889 18587 11987 18685 ne
rect 11987 18587 12341 18685
tri 12341 18587 12439 18685 sw
tri 12439 18587 12537 18685 ne
rect 12537 18587 12891 18685
tri 12891 18587 12989 18685 sw
tri 12989 18587 13087 18685 ne
rect 13087 18587 13441 18685
tri 13441 18587 13539 18685 sw
tri 13539 18587 13637 18685 ne
rect 13637 18587 13991 18685
tri 13991 18587 14089 18685 sw
tri 14089 18587 14187 18685 ne
rect 14187 18587 14541 18685
tri 14541 18587 14639 18685 sw
tri 14639 18587 14737 18685 ne
rect 14737 18587 15091 18685
tri 15091 18587 15189 18685 sw
tri 15189 18587 15287 18685 ne
rect 15287 18587 15641 18685
tri 15641 18587 15739 18685 sw
tri 15739 18587 15837 18685 ne
rect 15837 18587 16191 18685
tri 16191 18587 16289 18685 sw
tri 16289 18587 16387 18685 ne
rect 16387 18587 16741 18685
tri 16741 18587 16839 18685 sw
tri 16839 18587 16937 18685 ne
rect 16937 18587 17291 18685
tri 17291 18587 17389 18685 sw
tri 17389 18587 17487 18685 ne
rect 17487 18587 17841 18685
tri 17841 18587 17939 18685 sw
tri 17939 18587 18037 18685 ne
rect 18037 18587 18391 18685
tri 18391 18587 18489 18685 sw
tri 18489 18587 18587 18685 ne
rect 18587 18587 18941 18685
tri 18941 18587 19039 18685 sw
tri 19039 18587 19137 18685 ne
rect 19137 18587 19491 18685
tri 19491 18587 19589 18685 sw
tri 19589 18587 19687 18685 ne
rect 19687 18587 20300 18685
rect -2000 18489 339 18587
tri 339 18489 437 18587 sw
tri 437 18489 535 18587 ne
rect 535 18489 889 18587
tri 889 18489 987 18587 sw
tri 987 18489 1085 18587 ne
rect 1085 18489 1439 18587
tri 1439 18489 1537 18587 sw
tri 1537 18489 1635 18587 ne
rect 1635 18489 1989 18587
tri 1989 18489 2087 18587 sw
tri 2087 18489 2185 18587 ne
rect 2185 18489 2539 18587
tri 2539 18489 2637 18587 sw
tri 2637 18489 2735 18587 ne
rect 2735 18489 3089 18587
tri 3089 18489 3187 18587 sw
tri 3187 18489 3285 18587 ne
rect 3285 18489 3639 18587
tri 3639 18489 3737 18587 sw
tri 3737 18489 3835 18587 ne
rect 3835 18489 4189 18587
tri 4189 18489 4287 18587 sw
tri 4287 18489 4385 18587 ne
rect 4385 18489 4739 18587
tri 4739 18489 4837 18587 sw
tri 4837 18489 4935 18587 ne
rect 4935 18489 5289 18587
tri 5289 18489 5387 18587 sw
tri 5387 18489 5485 18587 ne
rect 5485 18489 5839 18587
tri 5839 18489 5937 18587 sw
tri 5937 18489 6035 18587 ne
rect 6035 18489 6389 18587
tri 6389 18489 6487 18587 sw
tri 6487 18489 6585 18587 ne
rect 6585 18489 6939 18587
tri 6939 18489 7037 18587 sw
tri 7037 18489 7135 18587 ne
rect 7135 18489 7489 18587
tri 7489 18489 7587 18587 sw
tri 7587 18489 7685 18587 ne
rect 7685 18489 8039 18587
tri 8039 18489 8137 18587 sw
tri 8137 18489 8235 18587 ne
rect 8235 18489 8589 18587
tri 8589 18489 8687 18587 sw
tri 8687 18489 8785 18587 ne
rect 8785 18489 9139 18587
tri 9139 18489 9237 18587 sw
tri 9237 18489 9335 18587 ne
rect 9335 18489 9689 18587
tri 9689 18489 9787 18587 sw
tri 9787 18489 9885 18587 ne
rect 9885 18489 10239 18587
tri 10239 18489 10337 18587 sw
tri 10337 18489 10435 18587 ne
rect 10435 18489 10789 18587
tri 10789 18489 10887 18587 sw
tri 10887 18489 10985 18587 ne
rect 10985 18489 11339 18587
tri 11339 18489 11437 18587 sw
tri 11437 18489 11535 18587 ne
rect 11535 18489 11889 18587
tri 11889 18489 11987 18587 sw
tri 11987 18489 12085 18587 ne
rect 12085 18489 12439 18587
tri 12439 18489 12537 18587 sw
tri 12537 18489 12635 18587 ne
rect 12635 18489 12989 18587
tri 12989 18489 13087 18587 sw
tri 13087 18489 13185 18587 ne
rect 13185 18489 13539 18587
tri 13539 18489 13637 18587 sw
tri 13637 18489 13735 18587 ne
rect 13735 18489 14089 18587
tri 14089 18489 14187 18587 sw
tri 14187 18489 14285 18587 ne
rect 14285 18489 14639 18587
tri 14639 18489 14737 18587 sw
tri 14737 18489 14835 18587 ne
rect 14835 18489 15189 18587
tri 15189 18489 15287 18587 sw
tri 15287 18489 15385 18587 ne
rect 15385 18489 15739 18587
tri 15739 18489 15837 18587 sw
tri 15837 18489 15935 18587 ne
rect 15935 18489 16289 18587
tri 16289 18489 16387 18587 sw
tri 16387 18489 16485 18587 ne
rect 16485 18489 16839 18587
tri 16839 18489 16937 18587 sw
tri 16937 18489 17035 18587 ne
rect 17035 18489 17389 18587
tri 17389 18489 17487 18587 sw
tri 17487 18489 17585 18587 ne
rect 17585 18489 17939 18587
tri 17939 18489 18037 18587 sw
tri 18037 18489 18135 18587 ne
rect 18135 18489 18489 18587
tri 18489 18489 18587 18587 sw
tri 18587 18489 18685 18587 ne
rect 18685 18489 19039 18587
tri 19039 18489 19137 18587 sw
tri 19137 18489 19235 18587 ne
rect 19235 18489 19589 18587
tri 19589 18489 19687 18587 sw
rect 20800 18489 21800 19137
rect -2000 18485 437 18489
rect -2000 18365 215 18485
rect 335 18391 437 18485
tri 437 18391 535 18489 sw
tri 535 18391 633 18489 ne
rect 633 18485 987 18489
rect 633 18391 765 18485
rect 335 18365 535 18391
rect -2000 18361 535 18365
rect -2000 17713 -1000 18361
tri 113 18263 211 18361 ne
rect 211 18313 535 18361
tri 535 18313 613 18391 sw
tri 633 18313 711 18391 ne
rect 711 18365 765 18391
rect 885 18391 987 18485
tri 987 18391 1085 18489 sw
tri 1085 18391 1183 18489 ne
rect 1183 18485 1537 18489
rect 1183 18391 1315 18485
rect 885 18365 1085 18391
rect 711 18313 1085 18365
tri 1085 18313 1163 18391 sw
tri 1183 18313 1261 18391 ne
rect 1261 18365 1315 18391
rect 1435 18391 1537 18485
tri 1537 18391 1635 18489 sw
tri 1635 18391 1733 18489 ne
rect 1733 18485 2087 18489
rect 1733 18391 1865 18485
rect 1435 18365 1635 18391
rect 1261 18313 1635 18365
tri 1635 18313 1713 18391 sw
tri 1733 18313 1811 18391 ne
rect 1811 18365 1865 18391
rect 1985 18391 2087 18485
tri 2087 18391 2185 18489 sw
tri 2185 18391 2283 18489 ne
rect 2283 18485 2637 18489
rect 2283 18391 2415 18485
rect 1985 18365 2185 18391
rect 1811 18313 2185 18365
tri 2185 18313 2263 18391 sw
tri 2283 18313 2361 18391 ne
rect 2361 18365 2415 18391
rect 2535 18391 2637 18485
tri 2637 18391 2735 18489 sw
tri 2735 18391 2833 18489 ne
rect 2833 18485 3187 18489
rect 2833 18391 2965 18485
rect 2535 18365 2735 18391
rect 2361 18313 2735 18365
tri 2735 18313 2813 18391 sw
tri 2833 18313 2911 18391 ne
rect 2911 18365 2965 18391
rect 3085 18391 3187 18485
tri 3187 18391 3285 18489 sw
tri 3285 18391 3383 18489 ne
rect 3383 18485 3737 18489
rect 3383 18391 3515 18485
rect 3085 18365 3285 18391
rect 2911 18313 3285 18365
tri 3285 18313 3363 18391 sw
tri 3383 18313 3461 18391 ne
rect 3461 18365 3515 18391
rect 3635 18391 3737 18485
tri 3737 18391 3835 18489 sw
tri 3835 18391 3933 18489 ne
rect 3933 18485 4287 18489
rect 3933 18391 4065 18485
rect 3635 18365 3835 18391
rect 3461 18313 3835 18365
tri 3835 18313 3913 18391 sw
tri 3933 18313 4011 18391 ne
rect 4011 18365 4065 18391
rect 4185 18391 4287 18485
tri 4287 18391 4385 18489 sw
tri 4385 18391 4483 18489 ne
rect 4483 18485 4837 18489
rect 4483 18391 4615 18485
rect 4185 18365 4385 18391
rect 4011 18313 4385 18365
tri 4385 18313 4463 18391 sw
tri 4483 18313 4561 18391 ne
rect 4561 18365 4615 18391
rect 4735 18391 4837 18485
tri 4837 18391 4935 18489 sw
tri 4935 18391 5033 18489 ne
rect 5033 18485 5387 18489
rect 5033 18391 5165 18485
rect 4735 18365 4935 18391
rect 4561 18313 4935 18365
tri 4935 18313 5013 18391 sw
tri 5033 18313 5111 18391 ne
rect 5111 18365 5165 18391
rect 5285 18391 5387 18485
tri 5387 18391 5485 18489 sw
tri 5485 18391 5583 18489 ne
rect 5583 18485 5937 18489
rect 5583 18391 5715 18485
rect 5285 18365 5485 18391
rect 5111 18313 5485 18365
tri 5485 18313 5563 18391 sw
tri 5583 18313 5661 18391 ne
rect 5661 18365 5715 18391
rect 5835 18391 5937 18485
tri 5937 18391 6035 18489 sw
tri 6035 18391 6133 18489 ne
rect 6133 18485 6487 18489
rect 6133 18391 6265 18485
rect 5835 18365 6035 18391
rect 5661 18313 6035 18365
tri 6035 18313 6113 18391 sw
tri 6133 18313 6211 18391 ne
rect 6211 18365 6265 18391
rect 6385 18391 6487 18485
tri 6487 18391 6585 18489 sw
tri 6585 18391 6683 18489 ne
rect 6683 18485 7037 18489
rect 6683 18391 6815 18485
rect 6385 18365 6585 18391
rect 6211 18313 6585 18365
tri 6585 18313 6663 18391 sw
tri 6683 18313 6761 18391 ne
rect 6761 18365 6815 18391
rect 6935 18391 7037 18485
tri 7037 18391 7135 18489 sw
tri 7135 18391 7233 18489 ne
rect 7233 18485 7587 18489
rect 7233 18391 7365 18485
rect 6935 18365 7135 18391
rect 6761 18313 7135 18365
tri 7135 18313 7213 18391 sw
tri 7233 18313 7311 18391 ne
rect 7311 18365 7365 18391
rect 7485 18391 7587 18485
tri 7587 18391 7685 18489 sw
tri 7685 18391 7783 18489 ne
rect 7783 18485 8137 18489
rect 7783 18391 7915 18485
rect 7485 18365 7685 18391
rect 7311 18313 7685 18365
tri 7685 18313 7763 18391 sw
tri 7783 18313 7861 18391 ne
rect 7861 18365 7915 18391
rect 8035 18391 8137 18485
tri 8137 18391 8235 18489 sw
tri 8235 18391 8333 18489 ne
rect 8333 18485 8687 18489
rect 8333 18391 8465 18485
rect 8035 18365 8235 18391
rect 7861 18313 8235 18365
tri 8235 18313 8313 18391 sw
tri 8333 18313 8411 18391 ne
rect 8411 18365 8465 18391
rect 8585 18391 8687 18485
tri 8687 18391 8785 18489 sw
tri 8785 18391 8883 18489 ne
rect 8883 18485 9237 18489
rect 8883 18391 9015 18485
rect 8585 18365 8785 18391
rect 8411 18313 8785 18365
tri 8785 18313 8863 18391 sw
tri 8883 18313 8961 18391 ne
rect 8961 18365 9015 18391
rect 9135 18391 9237 18485
tri 9237 18391 9335 18489 sw
tri 9335 18391 9433 18489 ne
rect 9433 18485 9787 18489
rect 9433 18391 9565 18485
rect 9135 18365 9335 18391
rect 8961 18313 9335 18365
tri 9335 18313 9413 18391 sw
tri 9433 18313 9511 18391 ne
rect 9511 18365 9565 18391
rect 9685 18391 9787 18485
tri 9787 18391 9885 18489 sw
tri 9885 18391 9983 18489 ne
rect 9983 18485 10337 18489
rect 9983 18391 10115 18485
rect 9685 18365 9885 18391
rect 9511 18313 9885 18365
tri 9885 18313 9963 18391 sw
tri 9983 18313 10061 18391 ne
rect 10061 18365 10115 18391
rect 10235 18391 10337 18485
tri 10337 18391 10435 18489 sw
tri 10435 18391 10533 18489 ne
rect 10533 18485 10887 18489
rect 10533 18391 10665 18485
rect 10235 18365 10435 18391
rect 10061 18313 10435 18365
tri 10435 18313 10513 18391 sw
tri 10533 18313 10611 18391 ne
rect 10611 18365 10665 18391
rect 10785 18391 10887 18485
tri 10887 18391 10985 18489 sw
tri 10985 18391 11083 18489 ne
rect 11083 18485 11437 18489
rect 11083 18391 11215 18485
rect 10785 18365 10985 18391
rect 10611 18313 10985 18365
tri 10985 18313 11063 18391 sw
tri 11083 18313 11161 18391 ne
rect 11161 18365 11215 18391
rect 11335 18391 11437 18485
tri 11437 18391 11535 18489 sw
tri 11535 18391 11633 18489 ne
rect 11633 18485 11987 18489
rect 11633 18391 11765 18485
rect 11335 18365 11535 18391
rect 11161 18313 11535 18365
tri 11535 18313 11613 18391 sw
tri 11633 18313 11711 18391 ne
rect 11711 18365 11765 18391
rect 11885 18391 11987 18485
tri 11987 18391 12085 18489 sw
tri 12085 18391 12183 18489 ne
rect 12183 18485 12537 18489
rect 12183 18391 12315 18485
rect 11885 18365 12085 18391
rect 11711 18313 12085 18365
tri 12085 18313 12163 18391 sw
tri 12183 18313 12261 18391 ne
rect 12261 18365 12315 18391
rect 12435 18391 12537 18485
tri 12537 18391 12635 18489 sw
tri 12635 18391 12733 18489 ne
rect 12733 18485 13087 18489
rect 12733 18391 12865 18485
rect 12435 18365 12635 18391
rect 12261 18313 12635 18365
tri 12635 18313 12713 18391 sw
tri 12733 18313 12811 18391 ne
rect 12811 18365 12865 18391
rect 12985 18391 13087 18485
tri 13087 18391 13185 18489 sw
tri 13185 18391 13283 18489 ne
rect 13283 18485 13637 18489
rect 13283 18391 13415 18485
rect 12985 18365 13185 18391
rect 12811 18313 13185 18365
tri 13185 18313 13263 18391 sw
tri 13283 18313 13361 18391 ne
rect 13361 18365 13415 18391
rect 13535 18391 13637 18485
tri 13637 18391 13735 18489 sw
tri 13735 18391 13833 18489 ne
rect 13833 18485 14187 18489
rect 13833 18391 13965 18485
rect 13535 18365 13735 18391
rect 13361 18313 13735 18365
tri 13735 18313 13813 18391 sw
tri 13833 18313 13911 18391 ne
rect 13911 18365 13965 18391
rect 14085 18391 14187 18485
tri 14187 18391 14285 18489 sw
tri 14285 18391 14383 18489 ne
rect 14383 18485 14737 18489
rect 14383 18391 14515 18485
rect 14085 18365 14285 18391
rect 13911 18313 14285 18365
tri 14285 18313 14363 18391 sw
tri 14383 18313 14461 18391 ne
rect 14461 18365 14515 18391
rect 14635 18391 14737 18485
tri 14737 18391 14835 18489 sw
tri 14835 18391 14933 18489 ne
rect 14933 18485 15287 18489
rect 14933 18391 15065 18485
rect 14635 18365 14835 18391
rect 14461 18313 14835 18365
tri 14835 18313 14913 18391 sw
tri 14933 18313 15011 18391 ne
rect 15011 18365 15065 18391
rect 15185 18391 15287 18485
tri 15287 18391 15385 18489 sw
tri 15385 18391 15483 18489 ne
rect 15483 18485 15837 18489
rect 15483 18391 15615 18485
rect 15185 18365 15385 18391
rect 15011 18313 15385 18365
tri 15385 18313 15463 18391 sw
tri 15483 18313 15561 18391 ne
rect 15561 18365 15615 18391
rect 15735 18391 15837 18485
tri 15837 18391 15935 18489 sw
tri 15935 18391 16033 18489 ne
rect 16033 18485 16387 18489
rect 16033 18391 16165 18485
rect 15735 18365 15935 18391
rect 15561 18313 15935 18365
tri 15935 18313 16013 18391 sw
tri 16033 18313 16111 18391 ne
rect 16111 18365 16165 18391
rect 16285 18391 16387 18485
tri 16387 18391 16485 18489 sw
tri 16485 18391 16583 18489 ne
rect 16583 18485 16937 18489
rect 16583 18391 16715 18485
rect 16285 18365 16485 18391
rect 16111 18313 16485 18365
tri 16485 18313 16563 18391 sw
tri 16583 18313 16661 18391 ne
rect 16661 18365 16715 18391
rect 16835 18391 16937 18485
tri 16937 18391 17035 18489 sw
tri 17035 18391 17133 18489 ne
rect 17133 18485 17487 18489
rect 17133 18391 17265 18485
rect 16835 18365 17035 18391
rect 16661 18313 17035 18365
tri 17035 18313 17113 18391 sw
tri 17133 18313 17211 18391 ne
rect 17211 18365 17265 18391
rect 17385 18391 17487 18485
tri 17487 18391 17585 18489 sw
tri 17585 18391 17683 18489 ne
rect 17683 18485 18037 18489
rect 17683 18391 17815 18485
rect 17385 18365 17585 18391
rect 17211 18313 17585 18365
tri 17585 18313 17663 18391 sw
tri 17683 18313 17761 18391 ne
rect 17761 18365 17815 18391
rect 17935 18391 18037 18485
tri 18037 18391 18135 18489 sw
tri 18135 18391 18233 18489 ne
rect 18233 18485 18587 18489
rect 18233 18391 18365 18485
rect 17935 18365 18135 18391
rect 17761 18313 18135 18365
tri 18135 18313 18213 18391 sw
tri 18233 18313 18311 18391 ne
rect 18311 18365 18365 18391
rect 18485 18391 18587 18485
tri 18587 18391 18685 18489 sw
tri 18685 18391 18783 18489 ne
rect 18783 18485 19137 18489
rect 18783 18391 18915 18485
rect 18485 18365 18685 18391
rect 18311 18313 18685 18365
tri 18685 18313 18763 18391 sw
tri 18783 18313 18861 18391 ne
rect 18861 18365 18915 18391
rect 19035 18391 19137 18485
tri 19137 18391 19235 18489 sw
tri 19235 18391 19333 18489 ne
rect 19333 18485 21800 18489
rect 19333 18391 19465 18485
rect 19035 18365 19235 18391
rect 18861 18313 19235 18365
tri 19235 18313 19313 18391 sw
tri 19333 18313 19411 18391 ne
rect 19411 18365 19465 18391
rect 19585 18365 21800 18485
rect 19411 18313 21800 18365
rect 211 18263 613 18313
rect -500 18213 113 18263
tri 113 18213 163 18263 sw
tri 211 18213 261 18263 ne
rect 261 18233 613 18263
tri 613 18233 693 18313 sw
tri 711 18233 791 18313 ne
rect 791 18233 1163 18313
tri 1163 18233 1243 18313 sw
tri 1261 18233 1341 18313 ne
rect 1341 18233 1713 18313
tri 1713 18233 1793 18313 sw
tri 1811 18233 1891 18313 ne
rect 1891 18233 2263 18313
tri 2263 18233 2343 18313 sw
tri 2361 18233 2441 18313 ne
rect 2441 18233 2813 18313
tri 2813 18233 2893 18313 sw
tri 2911 18233 2991 18313 ne
rect 2991 18233 3363 18313
tri 3363 18233 3443 18313 sw
tri 3461 18233 3541 18313 ne
rect 3541 18233 3913 18313
tri 3913 18233 3993 18313 sw
tri 4011 18233 4091 18313 ne
rect 4091 18233 4463 18313
tri 4463 18233 4543 18313 sw
tri 4561 18233 4641 18313 ne
rect 4641 18233 5013 18313
tri 5013 18233 5093 18313 sw
tri 5111 18233 5191 18313 ne
rect 5191 18233 5563 18313
tri 5563 18233 5643 18313 sw
tri 5661 18233 5741 18313 ne
rect 5741 18233 6113 18313
tri 6113 18233 6193 18313 sw
tri 6211 18233 6291 18313 ne
rect 6291 18233 6663 18313
tri 6663 18233 6743 18313 sw
tri 6761 18233 6841 18313 ne
rect 6841 18233 7213 18313
tri 7213 18233 7293 18313 sw
tri 7311 18233 7391 18313 ne
rect 7391 18233 7763 18313
tri 7763 18233 7843 18313 sw
tri 7861 18233 7941 18313 ne
rect 7941 18233 8313 18313
tri 8313 18233 8393 18313 sw
tri 8411 18233 8491 18313 ne
rect 8491 18233 8863 18313
tri 8863 18233 8943 18313 sw
tri 8961 18233 9041 18313 ne
rect 9041 18233 9413 18313
tri 9413 18233 9493 18313 sw
tri 9511 18233 9591 18313 ne
rect 9591 18233 9963 18313
tri 9963 18233 10043 18313 sw
tri 10061 18233 10141 18313 ne
rect 10141 18233 10513 18313
tri 10513 18233 10593 18313 sw
tri 10611 18233 10691 18313 ne
rect 10691 18233 11063 18313
tri 11063 18233 11143 18313 sw
tri 11161 18233 11241 18313 ne
rect 11241 18233 11613 18313
tri 11613 18233 11693 18313 sw
tri 11711 18233 11791 18313 ne
rect 11791 18233 12163 18313
tri 12163 18233 12243 18313 sw
tri 12261 18233 12341 18313 ne
rect 12341 18233 12713 18313
tri 12713 18233 12793 18313 sw
tri 12811 18233 12891 18313 ne
rect 12891 18233 13263 18313
tri 13263 18233 13343 18313 sw
tri 13361 18233 13441 18313 ne
rect 13441 18233 13813 18313
tri 13813 18233 13893 18313 sw
tri 13911 18233 13991 18313 ne
rect 13991 18233 14363 18313
tri 14363 18233 14443 18313 sw
tri 14461 18233 14541 18313 ne
rect 14541 18233 14913 18313
tri 14913 18233 14993 18313 sw
tri 15011 18233 15091 18313 ne
rect 15091 18233 15463 18313
tri 15463 18233 15543 18313 sw
tri 15561 18233 15641 18313 ne
rect 15641 18233 16013 18313
tri 16013 18233 16093 18313 sw
tri 16111 18233 16191 18313 ne
rect 16191 18233 16563 18313
tri 16563 18233 16643 18313 sw
tri 16661 18233 16741 18313 ne
rect 16741 18233 17113 18313
tri 17113 18233 17193 18313 sw
tri 17211 18233 17291 18313 ne
rect 17291 18233 17663 18313
tri 17663 18233 17743 18313 sw
tri 17761 18233 17841 18313 ne
rect 17841 18233 18213 18313
tri 18213 18233 18293 18313 sw
tri 18311 18233 18391 18313 ne
rect 18391 18233 18763 18313
tri 18763 18233 18843 18313 sw
tri 18861 18233 18941 18313 ne
rect 18941 18233 19313 18313
tri 19313 18233 19393 18313 sw
tri 19411 18233 19491 18313 ne
rect 19491 18233 20100 18313
rect 261 18213 693 18233
rect -500 18135 163 18213
tri 163 18135 241 18213 sw
tri 261 18135 339 18213 ne
rect 339 18135 693 18213
tri 693 18135 791 18233 sw
tri 791 18135 889 18233 ne
rect 889 18135 1243 18233
tri 1243 18135 1341 18233 sw
tri 1341 18135 1439 18233 ne
rect 1439 18135 1793 18233
tri 1793 18135 1891 18233 sw
tri 1891 18135 1989 18233 ne
rect 1989 18135 2343 18233
tri 2343 18135 2441 18233 sw
tri 2441 18135 2539 18233 ne
rect 2539 18135 2893 18233
tri 2893 18135 2991 18233 sw
tri 2991 18135 3089 18233 ne
rect 3089 18135 3443 18233
tri 3443 18135 3541 18233 sw
tri 3541 18135 3639 18233 ne
rect 3639 18135 3993 18233
tri 3993 18135 4091 18233 sw
tri 4091 18135 4189 18233 ne
rect 4189 18135 4543 18233
tri 4543 18135 4641 18233 sw
tri 4641 18135 4739 18233 ne
rect 4739 18135 5093 18233
tri 5093 18135 5191 18233 sw
tri 5191 18135 5289 18233 ne
rect 5289 18135 5643 18233
tri 5643 18135 5741 18233 sw
tri 5741 18135 5839 18233 ne
rect 5839 18135 6193 18233
tri 6193 18135 6291 18233 sw
tri 6291 18135 6389 18233 ne
rect 6389 18135 6743 18233
tri 6743 18135 6841 18233 sw
tri 6841 18135 6939 18233 ne
rect 6939 18135 7293 18233
tri 7293 18135 7391 18233 sw
tri 7391 18135 7489 18233 ne
rect 7489 18135 7843 18233
tri 7843 18135 7941 18233 sw
tri 7941 18135 8039 18233 ne
rect 8039 18135 8393 18233
tri 8393 18135 8491 18233 sw
tri 8491 18135 8589 18233 ne
rect 8589 18135 8943 18233
tri 8943 18135 9041 18233 sw
tri 9041 18135 9139 18233 ne
rect 9139 18135 9493 18233
tri 9493 18135 9591 18233 sw
tri 9591 18135 9689 18233 ne
rect 9689 18135 10043 18233
tri 10043 18135 10141 18233 sw
tri 10141 18135 10239 18233 ne
rect 10239 18135 10593 18233
tri 10593 18135 10691 18233 sw
tri 10691 18135 10789 18233 ne
rect 10789 18135 11143 18233
tri 11143 18135 11241 18233 sw
tri 11241 18135 11339 18233 ne
rect 11339 18135 11693 18233
tri 11693 18135 11791 18233 sw
tri 11791 18135 11889 18233 ne
rect 11889 18135 12243 18233
tri 12243 18135 12341 18233 sw
tri 12341 18135 12439 18233 ne
rect 12439 18135 12793 18233
tri 12793 18135 12891 18233 sw
tri 12891 18135 12989 18233 ne
rect 12989 18135 13343 18233
tri 13343 18135 13441 18233 sw
tri 13441 18135 13539 18233 ne
rect 13539 18135 13893 18233
tri 13893 18135 13991 18233 sw
tri 13991 18135 14089 18233 ne
rect 14089 18135 14443 18233
tri 14443 18135 14541 18233 sw
tri 14541 18135 14639 18233 ne
rect 14639 18135 14993 18233
tri 14993 18135 15091 18233 sw
tri 15091 18135 15189 18233 ne
rect 15189 18135 15543 18233
tri 15543 18135 15641 18233 sw
tri 15641 18135 15739 18233 ne
rect 15739 18135 16093 18233
tri 16093 18135 16191 18233 sw
tri 16191 18135 16289 18233 ne
rect 16289 18135 16643 18233
tri 16643 18135 16741 18233 sw
tri 16741 18135 16839 18233 ne
rect 16839 18135 17193 18233
tri 17193 18135 17291 18233 sw
tri 17291 18135 17389 18233 ne
rect 17389 18135 17743 18233
tri 17743 18135 17841 18233 sw
tri 17841 18135 17939 18233 ne
rect 17939 18135 18293 18233
tri 18293 18135 18391 18233 sw
tri 18391 18135 18489 18233 ne
rect 18489 18135 18843 18233
tri 18843 18135 18941 18233 sw
tri 18941 18135 19039 18233 ne
rect 19039 18135 19393 18233
tri 19393 18135 19491 18233 sw
tri 19491 18135 19589 18233 ne
rect 19589 18213 20100 18233
rect 20200 18213 21800 18313
rect 19589 18135 21800 18213
rect -500 18087 241 18135
rect -500 17987 -400 18087
rect -300 18037 241 18087
tri 241 18037 339 18135 sw
tri 339 18037 437 18135 ne
rect 437 18037 791 18135
tri 791 18037 889 18135 sw
tri 889 18037 987 18135 ne
rect 987 18037 1341 18135
tri 1341 18037 1439 18135 sw
tri 1439 18037 1537 18135 ne
rect 1537 18037 1891 18135
tri 1891 18037 1989 18135 sw
tri 1989 18037 2087 18135 ne
rect 2087 18037 2441 18135
tri 2441 18037 2539 18135 sw
tri 2539 18037 2637 18135 ne
rect 2637 18037 2991 18135
tri 2991 18037 3089 18135 sw
tri 3089 18037 3187 18135 ne
rect 3187 18037 3541 18135
tri 3541 18037 3639 18135 sw
tri 3639 18037 3737 18135 ne
rect 3737 18037 4091 18135
tri 4091 18037 4189 18135 sw
tri 4189 18037 4287 18135 ne
rect 4287 18037 4641 18135
tri 4641 18037 4739 18135 sw
tri 4739 18037 4837 18135 ne
rect 4837 18037 5191 18135
tri 5191 18037 5289 18135 sw
tri 5289 18037 5387 18135 ne
rect 5387 18037 5741 18135
tri 5741 18037 5839 18135 sw
tri 5839 18037 5937 18135 ne
rect 5937 18037 6291 18135
tri 6291 18037 6389 18135 sw
tri 6389 18037 6487 18135 ne
rect 6487 18037 6841 18135
tri 6841 18037 6939 18135 sw
tri 6939 18037 7037 18135 ne
rect 7037 18037 7391 18135
tri 7391 18037 7489 18135 sw
tri 7489 18037 7587 18135 ne
rect 7587 18037 7941 18135
tri 7941 18037 8039 18135 sw
tri 8039 18037 8137 18135 ne
rect 8137 18037 8491 18135
tri 8491 18037 8589 18135 sw
tri 8589 18037 8687 18135 ne
rect 8687 18037 9041 18135
tri 9041 18037 9139 18135 sw
tri 9139 18037 9237 18135 ne
rect 9237 18037 9591 18135
tri 9591 18037 9689 18135 sw
tri 9689 18037 9787 18135 ne
rect 9787 18037 10141 18135
tri 10141 18037 10239 18135 sw
tri 10239 18037 10337 18135 ne
rect 10337 18037 10691 18135
tri 10691 18037 10789 18135 sw
tri 10789 18037 10887 18135 ne
rect 10887 18037 11241 18135
tri 11241 18037 11339 18135 sw
tri 11339 18037 11437 18135 ne
rect 11437 18037 11791 18135
tri 11791 18037 11889 18135 sw
tri 11889 18037 11987 18135 ne
rect 11987 18037 12341 18135
tri 12341 18037 12439 18135 sw
tri 12439 18037 12537 18135 ne
rect 12537 18037 12891 18135
tri 12891 18037 12989 18135 sw
tri 12989 18037 13087 18135 ne
rect 13087 18037 13441 18135
tri 13441 18037 13539 18135 sw
tri 13539 18037 13637 18135 ne
rect 13637 18037 13991 18135
tri 13991 18037 14089 18135 sw
tri 14089 18037 14187 18135 ne
rect 14187 18037 14541 18135
tri 14541 18037 14639 18135 sw
tri 14639 18037 14737 18135 ne
rect 14737 18037 15091 18135
tri 15091 18037 15189 18135 sw
tri 15189 18037 15287 18135 ne
rect 15287 18037 15641 18135
tri 15641 18037 15739 18135 sw
tri 15739 18037 15837 18135 ne
rect 15837 18037 16191 18135
tri 16191 18037 16289 18135 sw
tri 16289 18037 16387 18135 ne
rect 16387 18037 16741 18135
tri 16741 18037 16839 18135 sw
tri 16839 18037 16937 18135 ne
rect 16937 18037 17291 18135
tri 17291 18037 17389 18135 sw
tri 17389 18037 17487 18135 ne
rect 17487 18037 17841 18135
tri 17841 18037 17939 18135 sw
tri 17939 18037 18037 18135 ne
rect 18037 18037 18391 18135
tri 18391 18037 18489 18135 sw
tri 18489 18037 18587 18135 ne
rect 18587 18037 18941 18135
tri 18941 18037 19039 18135 sw
tri 19039 18037 19137 18135 ne
rect 19137 18037 19491 18135
tri 19491 18037 19589 18135 sw
tri 19589 18037 19687 18135 ne
rect 19687 18037 21800 18135
rect -300 17987 339 18037
rect -500 17939 339 17987
tri 339 17939 437 18037 sw
tri 437 17939 535 18037 ne
rect 535 17939 889 18037
tri 889 17939 987 18037 sw
tri 987 17939 1085 18037 ne
rect 1085 17939 1439 18037
tri 1439 17939 1537 18037 sw
tri 1537 17939 1635 18037 ne
rect 1635 17939 1989 18037
tri 1989 17939 2087 18037 sw
tri 2087 17939 2185 18037 ne
rect 2185 17939 2539 18037
tri 2539 17939 2637 18037 sw
tri 2637 17939 2735 18037 ne
rect 2735 17939 3089 18037
tri 3089 17939 3187 18037 sw
tri 3187 17939 3285 18037 ne
rect 3285 17939 3639 18037
tri 3639 17939 3737 18037 sw
tri 3737 17939 3835 18037 ne
rect 3835 17939 4189 18037
tri 4189 17939 4287 18037 sw
tri 4287 17939 4385 18037 ne
rect 4385 17939 4739 18037
tri 4739 17939 4837 18037 sw
tri 4837 17939 4935 18037 ne
rect 4935 17939 5289 18037
tri 5289 17939 5387 18037 sw
tri 5387 17939 5485 18037 ne
rect 5485 17939 5839 18037
tri 5839 17939 5937 18037 sw
tri 5937 17939 6035 18037 ne
rect 6035 17939 6389 18037
tri 6389 17939 6487 18037 sw
tri 6487 17939 6585 18037 ne
rect 6585 17939 6939 18037
tri 6939 17939 7037 18037 sw
tri 7037 17939 7135 18037 ne
rect 7135 17939 7489 18037
tri 7489 17939 7587 18037 sw
tri 7587 17939 7685 18037 ne
rect 7685 17939 8039 18037
tri 8039 17939 8137 18037 sw
tri 8137 17939 8235 18037 ne
rect 8235 17939 8589 18037
tri 8589 17939 8687 18037 sw
tri 8687 17939 8785 18037 ne
rect 8785 17939 9139 18037
tri 9139 17939 9237 18037 sw
tri 9237 17939 9335 18037 ne
rect 9335 17939 9689 18037
tri 9689 17939 9787 18037 sw
tri 9787 17939 9885 18037 ne
rect 9885 17939 10239 18037
tri 10239 17939 10337 18037 sw
tri 10337 17939 10435 18037 ne
rect 10435 17939 10789 18037
tri 10789 17939 10887 18037 sw
tri 10887 17939 10985 18037 ne
rect 10985 17939 11339 18037
tri 11339 17939 11437 18037 sw
tri 11437 17939 11535 18037 ne
rect 11535 17939 11889 18037
tri 11889 17939 11987 18037 sw
tri 11987 17939 12085 18037 ne
rect 12085 17939 12439 18037
tri 12439 17939 12537 18037 sw
tri 12537 17939 12635 18037 ne
rect 12635 17939 12989 18037
tri 12989 17939 13087 18037 sw
tri 13087 17939 13185 18037 ne
rect 13185 17939 13539 18037
tri 13539 17939 13637 18037 sw
tri 13637 17939 13735 18037 ne
rect 13735 17939 14089 18037
tri 14089 17939 14187 18037 sw
tri 14187 17939 14285 18037 ne
rect 14285 17939 14639 18037
tri 14639 17939 14737 18037 sw
tri 14737 17939 14835 18037 ne
rect 14835 17939 15189 18037
tri 15189 17939 15287 18037 sw
tri 15287 17939 15385 18037 ne
rect 15385 17939 15739 18037
tri 15739 17939 15837 18037 sw
tri 15837 17939 15935 18037 ne
rect 15935 17939 16289 18037
tri 16289 17939 16387 18037 sw
tri 16387 17939 16485 18037 ne
rect 16485 17939 16839 18037
tri 16839 17939 16937 18037 sw
tri 16937 17939 17035 18037 ne
rect 17035 17939 17389 18037
tri 17389 17939 17487 18037 sw
tri 17487 17939 17585 18037 ne
rect 17585 17939 17939 18037
tri 17939 17939 18037 18037 sw
tri 18037 17939 18135 18037 ne
rect 18135 17939 18489 18037
tri 18489 17939 18587 18037 sw
tri 18587 17939 18685 18037 ne
rect 18685 17939 19039 18037
tri 19039 17939 19137 18037 sw
tri 19137 17939 19235 18037 ne
rect 19235 17939 19589 18037
tri 19589 17939 19687 18037 sw
rect -500 17935 437 17939
rect -500 17815 215 17935
rect 335 17841 437 17935
tri 437 17841 535 17939 sw
tri 535 17841 633 17939 ne
rect 633 17935 987 17939
rect 633 17841 765 17935
rect 335 17815 535 17841
rect -500 17811 535 17815
tri 535 17811 565 17841 sw
tri 633 17811 663 17841 ne
rect 663 17815 765 17841
rect 885 17841 987 17935
tri 987 17841 1085 17939 sw
tri 1085 17841 1183 17939 ne
rect 1183 17935 1537 17939
rect 1183 17841 1315 17935
rect 885 17815 1085 17841
rect 663 17811 1085 17815
tri 1085 17811 1115 17841 sw
tri 1183 17811 1213 17841 ne
rect 1213 17815 1315 17841
rect 1435 17841 1537 17935
tri 1537 17841 1635 17939 sw
tri 1635 17841 1733 17939 ne
rect 1733 17935 2087 17939
rect 1733 17841 1865 17935
rect 1435 17815 1635 17841
rect 1213 17811 1635 17815
tri 1635 17811 1665 17841 sw
tri 1733 17811 1763 17841 ne
rect 1763 17815 1865 17841
rect 1985 17841 2087 17935
tri 2087 17841 2185 17939 sw
tri 2185 17841 2283 17939 ne
rect 2283 17935 2637 17939
rect 2283 17841 2415 17935
rect 1985 17815 2185 17841
rect 1763 17811 2185 17815
tri 2185 17811 2215 17841 sw
tri 2283 17811 2313 17841 ne
rect 2313 17815 2415 17841
rect 2535 17841 2637 17935
tri 2637 17841 2735 17939 sw
tri 2735 17841 2833 17939 ne
rect 2833 17935 3187 17939
rect 2833 17841 2965 17935
rect 2535 17815 2735 17841
rect 2313 17811 2735 17815
tri 2735 17811 2765 17841 sw
tri 2833 17811 2863 17841 ne
rect 2863 17815 2965 17841
rect 3085 17841 3187 17935
tri 3187 17841 3285 17939 sw
tri 3285 17841 3383 17939 ne
rect 3383 17935 3737 17939
rect 3383 17841 3515 17935
rect 3085 17815 3285 17841
rect 2863 17811 3285 17815
tri 3285 17811 3315 17841 sw
tri 3383 17811 3413 17841 ne
rect 3413 17815 3515 17841
rect 3635 17841 3737 17935
tri 3737 17841 3835 17939 sw
tri 3835 17841 3933 17939 ne
rect 3933 17935 4287 17939
rect 3933 17841 4065 17935
rect 3635 17815 3835 17841
rect 3413 17811 3835 17815
tri 3835 17811 3865 17841 sw
tri 3933 17811 3963 17841 ne
rect 3963 17815 4065 17841
rect 4185 17841 4287 17935
tri 4287 17841 4385 17939 sw
tri 4385 17841 4483 17939 ne
rect 4483 17935 4837 17939
rect 4483 17841 4615 17935
rect 4185 17815 4385 17841
rect 3963 17811 4385 17815
tri 4385 17811 4415 17841 sw
tri 4483 17811 4513 17841 ne
rect 4513 17815 4615 17841
rect 4735 17841 4837 17935
tri 4837 17841 4935 17939 sw
tri 4935 17841 5033 17939 ne
rect 5033 17935 5387 17939
rect 5033 17841 5165 17935
rect 4735 17815 4935 17841
rect 4513 17811 4935 17815
tri 4935 17811 4965 17841 sw
tri 5033 17811 5063 17841 ne
rect 5063 17815 5165 17841
rect 5285 17841 5387 17935
tri 5387 17841 5485 17939 sw
tri 5485 17841 5583 17939 ne
rect 5583 17935 5937 17939
rect 5583 17841 5715 17935
rect 5285 17815 5485 17841
rect 5063 17811 5485 17815
tri 5485 17811 5515 17841 sw
tri 5583 17811 5613 17841 ne
rect 5613 17815 5715 17841
rect 5835 17841 5937 17935
tri 5937 17841 6035 17939 sw
tri 6035 17841 6133 17939 ne
rect 6133 17935 6487 17939
rect 6133 17841 6265 17935
rect 5835 17815 6035 17841
rect 5613 17811 6035 17815
tri 6035 17811 6065 17841 sw
tri 6133 17811 6163 17841 ne
rect 6163 17815 6265 17841
rect 6385 17841 6487 17935
tri 6487 17841 6585 17939 sw
tri 6585 17841 6683 17939 ne
rect 6683 17935 7037 17939
rect 6683 17841 6815 17935
rect 6385 17815 6585 17841
rect 6163 17811 6585 17815
tri 6585 17811 6615 17841 sw
tri 6683 17811 6713 17841 ne
rect 6713 17815 6815 17841
rect 6935 17841 7037 17935
tri 7037 17841 7135 17939 sw
tri 7135 17841 7233 17939 ne
rect 7233 17935 7587 17939
rect 7233 17841 7365 17935
rect 6935 17815 7135 17841
rect 6713 17811 7135 17815
tri 7135 17811 7165 17841 sw
tri 7233 17811 7263 17841 ne
rect 7263 17815 7365 17841
rect 7485 17841 7587 17935
tri 7587 17841 7685 17939 sw
tri 7685 17841 7783 17939 ne
rect 7783 17935 8137 17939
rect 7783 17841 7915 17935
rect 7485 17815 7685 17841
rect 7263 17811 7685 17815
tri 7685 17811 7715 17841 sw
tri 7783 17811 7813 17841 ne
rect 7813 17815 7915 17841
rect 8035 17841 8137 17935
tri 8137 17841 8235 17939 sw
tri 8235 17841 8333 17939 ne
rect 8333 17935 8687 17939
rect 8333 17841 8465 17935
rect 8035 17815 8235 17841
rect 7813 17811 8235 17815
tri 8235 17811 8265 17841 sw
tri 8333 17811 8363 17841 ne
rect 8363 17815 8465 17841
rect 8585 17841 8687 17935
tri 8687 17841 8785 17939 sw
tri 8785 17841 8883 17939 ne
rect 8883 17935 9237 17939
rect 8883 17841 9015 17935
rect 8585 17815 8785 17841
rect 8363 17811 8785 17815
tri 8785 17811 8815 17841 sw
tri 8883 17811 8913 17841 ne
rect 8913 17815 9015 17841
rect 9135 17841 9237 17935
tri 9237 17841 9335 17939 sw
tri 9335 17841 9433 17939 ne
rect 9433 17935 9787 17939
rect 9433 17841 9565 17935
rect 9135 17815 9335 17841
rect 8913 17811 9335 17815
tri 9335 17811 9365 17841 sw
tri 9433 17811 9463 17841 ne
rect 9463 17815 9565 17841
rect 9685 17841 9787 17935
tri 9787 17841 9885 17939 sw
tri 9885 17841 9983 17939 ne
rect 9983 17935 10337 17939
rect 9983 17841 10115 17935
rect 9685 17815 9885 17841
rect 9463 17811 9885 17815
tri 9885 17811 9915 17841 sw
tri 9983 17811 10013 17841 ne
rect 10013 17815 10115 17841
rect 10235 17841 10337 17935
tri 10337 17841 10435 17939 sw
tri 10435 17841 10533 17939 ne
rect 10533 17935 10887 17939
rect 10533 17841 10665 17935
rect 10235 17815 10435 17841
rect 10013 17811 10435 17815
tri 10435 17811 10465 17841 sw
tri 10533 17811 10563 17841 ne
rect 10563 17815 10665 17841
rect 10785 17841 10887 17935
tri 10887 17841 10985 17939 sw
tri 10985 17841 11083 17939 ne
rect 11083 17935 11437 17939
rect 11083 17841 11215 17935
rect 10785 17815 10985 17841
rect 10563 17811 10985 17815
tri 10985 17811 11015 17841 sw
tri 11083 17811 11113 17841 ne
rect 11113 17815 11215 17841
rect 11335 17841 11437 17935
tri 11437 17841 11535 17939 sw
tri 11535 17841 11633 17939 ne
rect 11633 17935 11987 17939
rect 11633 17841 11765 17935
rect 11335 17815 11535 17841
rect 11113 17811 11535 17815
tri 11535 17811 11565 17841 sw
tri 11633 17811 11663 17841 ne
rect 11663 17815 11765 17841
rect 11885 17841 11987 17935
tri 11987 17841 12085 17939 sw
tri 12085 17841 12183 17939 ne
rect 12183 17935 12537 17939
rect 12183 17841 12315 17935
rect 11885 17815 12085 17841
rect 11663 17811 12085 17815
tri 12085 17811 12115 17841 sw
tri 12183 17811 12213 17841 ne
rect 12213 17815 12315 17841
rect 12435 17841 12537 17935
tri 12537 17841 12635 17939 sw
tri 12635 17841 12733 17939 ne
rect 12733 17935 13087 17939
rect 12733 17841 12865 17935
rect 12435 17815 12635 17841
rect 12213 17811 12635 17815
tri 12635 17811 12665 17841 sw
tri 12733 17811 12763 17841 ne
rect 12763 17815 12865 17841
rect 12985 17841 13087 17935
tri 13087 17841 13185 17939 sw
tri 13185 17841 13283 17939 ne
rect 13283 17935 13637 17939
rect 13283 17841 13415 17935
rect 12985 17815 13185 17841
rect 12763 17811 13185 17815
tri 13185 17811 13215 17841 sw
tri 13283 17811 13313 17841 ne
rect 13313 17815 13415 17841
rect 13535 17841 13637 17935
tri 13637 17841 13735 17939 sw
tri 13735 17841 13833 17939 ne
rect 13833 17935 14187 17939
rect 13833 17841 13965 17935
rect 13535 17815 13735 17841
rect 13313 17811 13735 17815
tri 13735 17811 13765 17841 sw
tri 13833 17811 13863 17841 ne
rect 13863 17815 13965 17841
rect 14085 17841 14187 17935
tri 14187 17841 14285 17939 sw
tri 14285 17841 14383 17939 ne
rect 14383 17935 14737 17939
rect 14383 17841 14515 17935
rect 14085 17815 14285 17841
rect 13863 17811 14285 17815
tri 14285 17811 14315 17841 sw
tri 14383 17811 14413 17841 ne
rect 14413 17815 14515 17841
rect 14635 17841 14737 17935
tri 14737 17841 14835 17939 sw
tri 14835 17841 14933 17939 ne
rect 14933 17935 15287 17939
rect 14933 17841 15065 17935
rect 14635 17815 14835 17841
rect 14413 17811 14835 17815
tri 14835 17811 14865 17841 sw
tri 14933 17811 14963 17841 ne
rect 14963 17815 15065 17841
rect 15185 17841 15287 17935
tri 15287 17841 15385 17939 sw
tri 15385 17841 15483 17939 ne
rect 15483 17935 15837 17939
rect 15483 17841 15615 17935
rect 15185 17815 15385 17841
rect 14963 17811 15385 17815
tri 15385 17811 15415 17841 sw
tri 15483 17811 15513 17841 ne
rect 15513 17815 15615 17841
rect 15735 17841 15837 17935
tri 15837 17841 15935 17939 sw
tri 15935 17841 16033 17939 ne
rect 16033 17935 16387 17939
rect 16033 17841 16165 17935
rect 15735 17815 15935 17841
rect 15513 17811 15935 17815
tri 15935 17811 15965 17841 sw
tri 16033 17811 16063 17841 ne
rect 16063 17815 16165 17841
rect 16285 17841 16387 17935
tri 16387 17841 16485 17939 sw
tri 16485 17841 16583 17939 ne
rect 16583 17935 16937 17939
rect 16583 17841 16715 17935
rect 16285 17815 16485 17841
rect 16063 17811 16485 17815
tri 16485 17811 16515 17841 sw
tri 16583 17811 16613 17841 ne
rect 16613 17815 16715 17841
rect 16835 17841 16937 17935
tri 16937 17841 17035 17939 sw
tri 17035 17841 17133 17939 ne
rect 17133 17935 17487 17939
rect 17133 17841 17265 17935
rect 16835 17815 17035 17841
rect 16613 17811 17035 17815
tri 17035 17811 17065 17841 sw
tri 17133 17811 17163 17841 ne
rect 17163 17815 17265 17841
rect 17385 17841 17487 17935
tri 17487 17841 17585 17939 sw
tri 17585 17841 17683 17939 ne
rect 17683 17935 18037 17939
rect 17683 17841 17815 17935
rect 17385 17815 17585 17841
rect 17163 17811 17585 17815
tri 17585 17811 17615 17841 sw
tri 17683 17811 17713 17841 ne
rect 17713 17815 17815 17841
rect 17935 17841 18037 17935
tri 18037 17841 18135 17939 sw
tri 18135 17841 18233 17939 ne
rect 18233 17935 18587 17939
rect 18233 17841 18365 17935
rect 17935 17815 18135 17841
rect 17713 17811 18135 17815
tri 18135 17811 18165 17841 sw
tri 18233 17811 18263 17841 ne
rect 18263 17815 18365 17841
rect 18485 17841 18587 17935
tri 18587 17841 18685 17939 sw
tri 18685 17841 18783 17939 ne
rect 18783 17935 19137 17939
rect 18783 17841 18915 17935
rect 18485 17815 18685 17841
rect 18263 17811 18685 17815
tri 18685 17811 18715 17841 sw
tri 18783 17811 18813 17841 ne
rect 18813 17815 18915 17841
rect 19035 17841 19137 17935
tri 19137 17841 19235 17939 sw
tri 19235 17841 19333 17939 ne
rect 19333 17935 20300 17939
rect 19333 17841 19465 17935
rect 19035 17815 19235 17841
rect 18813 17811 19235 17815
tri 19235 17811 19265 17841 sw
tri 19333 17811 19363 17841 ne
rect 19363 17815 19465 17841
rect 19585 17815 20300 17935
rect 19363 17811 20300 17815
tri 113 17713 211 17811 ne
rect 211 17713 565 17811
tri 565 17713 663 17811 sw
tri 663 17713 761 17811 ne
rect 761 17713 1115 17811
tri 1115 17713 1213 17811 sw
tri 1213 17713 1311 17811 ne
rect 1311 17713 1665 17811
tri 1665 17713 1763 17811 sw
tri 1763 17713 1861 17811 ne
rect 1861 17713 2215 17811
tri 2215 17713 2313 17811 sw
tri 2313 17713 2411 17811 ne
rect 2411 17713 2765 17811
tri 2765 17713 2863 17811 sw
tri 2863 17713 2961 17811 ne
rect 2961 17713 3315 17811
tri 3315 17713 3413 17811 sw
tri 3413 17713 3511 17811 ne
rect 3511 17713 3865 17811
tri 3865 17713 3963 17811 sw
tri 3963 17713 4061 17811 ne
rect 4061 17713 4415 17811
tri 4415 17713 4513 17811 sw
tri 4513 17713 4611 17811 ne
rect 4611 17713 4965 17811
tri 4965 17713 5063 17811 sw
tri 5063 17713 5161 17811 ne
rect 5161 17713 5515 17811
tri 5515 17713 5613 17811 sw
tri 5613 17713 5711 17811 ne
rect 5711 17713 6065 17811
tri 6065 17713 6163 17811 sw
tri 6163 17713 6261 17811 ne
rect 6261 17713 6615 17811
tri 6615 17713 6713 17811 sw
tri 6713 17713 6811 17811 ne
rect 6811 17713 7165 17811
tri 7165 17713 7263 17811 sw
tri 7263 17713 7361 17811 ne
rect 7361 17713 7715 17811
tri 7715 17713 7813 17811 sw
tri 7813 17713 7911 17811 ne
rect 7911 17713 8265 17811
tri 8265 17713 8363 17811 sw
tri 8363 17713 8461 17811 ne
rect 8461 17713 8815 17811
tri 8815 17713 8913 17811 sw
tri 8913 17713 9011 17811 ne
rect 9011 17713 9365 17811
tri 9365 17713 9463 17811 sw
tri 9463 17713 9561 17811 ne
rect 9561 17713 9915 17811
tri 9915 17713 10013 17811 sw
tri 10013 17713 10111 17811 ne
rect 10111 17713 10465 17811
tri 10465 17713 10563 17811 sw
tri 10563 17713 10661 17811 ne
rect 10661 17713 11015 17811
tri 11015 17713 11113 17811 sw
tri 11113 17713 11211 17811 ne
rect 11211 17713 11565 17811
tri 11565 17713 11663 17811 sw
tri 11663 17713 11761 17811 ne
rect 11761 17713 12115 17811
tri 12115 17713 12213 17811 sw
tri 12213 17713 12311 17811 ne
rect 12311 17713 12665 17811
tri 12665 17713 12763 17811 sw
tri 12763 17713 12861 17811 ne
rect 12861 17713 13215 17811
tri 13215 17713 13313 17811 sw
tri 13313 17713 13411 17811 ne
rect 13411 17713 13765 17811
tri 13765 17713 13863 17811 sw
tri 13863 17713 13961 17811 ne
rect 13961 17713 14315 17811
tri 14315 17713 14413 17811 sw
tri 14413 17713 14511 17811 ne
rect 14511 17713 14865 17811
tri 14865 17713 14963 17811 sw
tri 14963 17713 15061 17811 ne
rect 15061 17713 15415 17811
tri 15415 17713 15513 17811 sw
tri 15513 17713 15611 17811 ne
rect 15611 17713 15965 17811
tri 15965 17713 16063 17811 sw
tri 16063 17713 16161 17811 ne
rect 16161 17713 16515 17811
tri 16515 17713 16613 17811 sw
tri 16613 17713 16711 17811 ne
rect 16711 17713 17065 17811
tri 17065 17713 17163 17811 sw
tri 17163 17713 17261 17811 ne
rect 17261 17713 17615 17811
tri 17615 17713 17713 17811 sw
tri 17713 17713 17811 17811 ne
rect 17811 17713 18165 17811
tri 18165 17713 18263 17811 sw
tri 18263 17713 18361 17811 ne
rect 18361 17713 18715 17811
tri 18715 17713 18813 17811 sw
tri 18813 17713 18911 17811 ne
rect 18911 17713 19265 17811
tri 19265 17713 19363 17811 sw
tri 19363 17713 19461 17811 ne
rect 19461 17713 20300 17811
rect -2000 17683 113 17713
tri 113 17683 143 17713 sw
tri 211 17683 241 17713 ne
rect 241 17683 663 17713
tri 663 17683 693 17713 sw
tri 761 17683 791 17713 ne
rect 791 17683 1213 17713
tri 1213 17683 1243 17713 sw
tri 1311 17683 1341 17713 ne
rect 1341 17683 1763 17713
tri 1763 17683 1793 17713 sw
tri 1861 17683 1891 17713 ne
rect 1891 17683 2313 17713
tri 2313 17683 2343 17713 sw
tri 2411 17683 2441 17713 ne
rect 2441 17683 2863 17713
tri 2863 17683 2893 17713 sw
tri 2961 17683 2991 17713 ne
rect 2991 17683 3413 17713
tri 3413 17683 3443 17713 sw
tri 3511 17683 3541 17713 ne
rect 3541 17683 3963 17713
tri 3963 17683 3993 17713 sw
tri 4061 17683 4091 17713 ne
rect 4091 17683 4513 17713
tri 4513 17683 4543 17713 sw
tri 4611 17683 4641 17713 ne
rect 4641 17683 5063 17713
tri 5063 17683 5093 17713 sw
tri 5161 17683 5191 17713 ne
rect 5191 17683 5613 17713
tri 5613 17683 5643 17713 sw
tri 5711 17683 5741 17713 ne
rect 5741 17683 6163 17713
tri 6163 17683 6193 17713 sw
tri 6261 17683 6291 17713 ne
rect 6291 17683 6713 17713
tri 6713 17683 6743 17713 sw
tri 6811 17683 6841 17713 ne
rect 6841 17683 7263 17713
tri 7263 17683 7293 17713 sw
tri 7361 17683 7391 17713 ne
rect 7391 17683 7813 17713
tri 7813 17683 7843 17713 sw
tri 7911 17683 7941 17713 ne
rect 7941 17683 8363 17713
tri 8363 17683 8393 17713 sw
tri 8461 17683 8491 17713 ne
rect 8491 17683 8913 17713
tri 8913 17683 8943 17713 sw
tri 9011 17683 9041 17713 ne
rect 9041 17683 9463 17713
tri 9463 17683 9493 17713 sw
tri 9561 17683 9591 17713 ne
rect 9591 17683 10013 17713
tri 10013 17683 10043 17713 sw
tri 10111 17683 10141 17713 ne
rect 10141 17683 10563 17713
tri 10563 17683 10593 17713 sw
tri 10661 17683 10691 17713 ne
rect 10691 17683 11113 17713
tri 11113 17683 11143 17713 sw
tri 11211 17683 11241 17713 ne
rect 11241 17683 11663 17713
tri 11663 17683 11693 17713 sw
tri 11761 17683 11791 17713 ne
rect 11791 17683 12213 17713
tri 12213 17683 12243 17713 sw
tri 12311 17683 12341 17713 ne
rect 12341 17683 12763 17713
tri 12763 17683 12793 17713 sw
tri 12861 17683 12891 17713 ne
rect 12891 17683 13313 17713
tri 13313 17683 13343 17713 sw
tri 13411 17683 13441 17713 ne
rect 13441 17683 13863 17713
tri 13863 17683 13893 17713 sw
tri 13961 17683 13991 17713 ne
rect 13991 17683 14413 17713
tri 14413 17683 14443 17713 sw
tri 14511 17683 14541 17713 ne
rect 14541 17683 14963 17713
tri 14963 17683 14993 17713 sw
tri 15061 17683 15091 17713 ne
rect 15091 17683 15513 17713
tri 15513 17683 15543 17713 sw
tri 15611 17683 15641 17713 ne
rect 15641 17683 16063 17713
tri 16063 17683 16093 17713 sw
tri 16161 17683 16191 17713 ne
rect 16191 17683 16613 17713
tri 16613 17683 16643 17713 sw
tri 16711 17683 16741 17713 ne
rect 16741 17683 17163 17713
tri 17163 17683 17193 17713 sw
tri 17261 17683 17291 17713 ne
rect 17291 17683 17713 17713
tri 17713 17683 17743 17713 sw
tri 17811 17683 17841 17713 ne
rect 17841 17683 18263 17713
tri 18263 17683 18293 17713 sw
tri 18361 17683 18391 17713 ne
rect 18391 17683 18813 17713
tri 18813 17683 18843 17713 sw
tri 18911 17683 18941 17713 ne
rect 18941 17683 19363 17713
tri 19363 17683 19393 17713 sw
tri 19461 17683 19491 17713 ne
rect 19491 17683 20300 17713
rect -2000 17585 143 17683
tri 143 17585 241 17683 sw
tri 241 17585 339 17683 ne
rect 339 17585 693 17683
tri 693 17585 791 17683 sw
tri 791 17585 889 17683 ne
rect 889 17585 1243 17683
tri 1243 17585 1341 17683 sw
tri 1341 17585 1439 17683 ne
rect 1439 17585 1793 17683
tri 1793 17585 1891 17683 sw
tri 1891 17585 1989 17683 ne
rect 1989 17585 2343 17683
tri 2343 17585 2441 17683 sw
tri 2441 17585 2539 17683 ne
rect 2539 17585 2893 17683
tri 2893 17585 2991 17683 sw
tri 2991 17585 3089 17683 ne
rect 3089 17585 3443 17683
tri 3443 17585 3541 17683 sw
tri 3541 17585 3639 17683 ne
rect 3639 17585 3993 17683
tri 3993 17585 4091 17683 sw
tri 4091 17585 4189 17683 ne
rect 4189 17585 4543 17683
tri 4543 17585 4641 17683 sw
tri 4641 17585 4739 17683 ne
rect 4739 17585 5093 17683
tri 5093 17585 5191 17683 sw
tri 5191 17585 5289 17683 ne
rect 5289 17585 5643 17683
tri 5643 17585 5741 17683 sw
tri 5741 17585 5839 17683 ne
rect 5839 17585 6193 17683
tri 6193 17585 6291 17683 sw
tri 6291 17585 6389 17683 ne
rect 6389 17585 6743 17683
tri 6743 17585 6841 17683 sw
tri 6841 17585 6939 17683 ne
rect 6939 17585 7293 17683
tri 7293 17585 7391 17683 sw
tri 7391 17585 7489 17683 ne
rect 7489 17585 7843 17683
tri 7843 17585 7941 17683 sw
tri 7941 17585 8039 17683 ne
rect 8039 17585 8393 17683
tri 8393 17585 8491 17683 sw
tri 8491 17585 8589 17683 ne
rect 8589 17585 8943 17683
tri 8943 17585 9041 17683 sw
tri 9041 17585 9139 17683 ne
rect 9139 17585 9493 17683
tri 9493 17585 9591 17683 sw
tri 9591 17585 9689 17683 ne
rect 9689 17585 10043 17683
tri 10043 17585 10141 17683 sw
tri 10141 17585 10239 17683 ne
rect 10239 17585 10593 17683
tri 10593 17585 10691 17683 sw
tri 10691 17585 10789 17683 ne
rect 10789 17585 11143 17683
tri 11143 17585 11241 17683 sw
tri 11241 17585 11339 17683 ne
rect 11339 17585 11693 17683
tri 11693 17585 11791 17683 sw
tri 11791 17585 11889 17683 ne
rect 11889 17585 12243 17683
tri 12243 17585 12341 17683 sw
tri 12341 17585 12439 17683 ne
rect 12439 17585 12793 17683
tri 12793 17585 12891 17683 sw
tri 12891 17585 12989 17683 ne
rect 12989 17585 13343 17683
tri 13343 17585 13441 17683 sw
tri 13441 17585 13539 17683 ne
rect 13539 17585 13893 17683
tri 13893 17585 13991 17683 sw
tri 13991 17585 14089 17683 ne
rect 14089 17585 14443 17683
tri 14443 17585 14541 17683 sw
tri 14541 17585 14639 17683 ne
rect 14639 17585 14993 17683
tri 14993 17585 15091 17683 sw
tri 15091 17585 15189 17683 ne
rect 15189 17585 15543 17683
tri 15543 17585 15641 17683 sw
tri 15641 17585 15739 17683 ne
rect 15739 17585 16093 17683
tri 16093 17585 16191 17683 sw
tri 16191 17585 16289 17683 ne
rect 16289 17585 16643 17683
tri 16643 17585 16741 17683 sw
tri 16741 17585 16839 17683 ne
rect 16839 17585 17193 17683
tri 17193 17585 17291 17683 sw
tri 17291 17585 17389 17683 ne
rect 17389 17585 17743 17683
tri 17743 17585 17841 17683 sw
tri 17841 17585 17939 17683 ne
rect 17939 17585 18293 17683
tri 18293 17585 18391 17683 sw
tri 18391 17585 18489 17683 ne
rect 18489 17585 18843 17683
tri 18843 17585 18941 17683 sw
tri 18941 17585 19039 17683 ne
rect 19039 17585 19393 17683
tri 19393 17585 19491 17683 sw
tri 19491 17585 19589 17683 ne
rect 19589 17585 20300 17683
rect -2000 17487 241 17585
tri 241 17487 339 17585 sw
tri 339 17487 437 17585 ne
rect 437 17487 791 17585
tri 791 17487 889 17585 sw
tri 889 17487 987 17585 ne
rect 987 17487 1341 17585
tri 1341 17487 1439 17585 sw
tri 1439 17487 1537 17585 ne
rect 1537 17487 1891 17585
tri 1891 17487 1989 17585 sw
tri 1989 17487 2087 17585 ne
rect 2087 17487 2441 17585
tri 2441 17487 2539 17585 sw
tri 2539 17487 2637 17585 ne
rect 2637 17487 2991 17585
tri 2991 17487 3089 17585 sw
tri 3089 17487 3187 17585 ne
rect 3187 17487 3541 17585
tri 3541 17487 3639 17585 sw
tri 3639 17487 3737 17585 ne
rect 3737 17487 4091 17585
tri 4091 17487 4189 17585 sw
tri 4189 17487 4287 17585 ne
rect 4287 17487 4641 17585
tri 4641 17487 4739 17585 sw
tri 4739 17487 4837 17585 ne
rect 4837 17487 5191 17585
tri 5191 17487 5289 17585 sw
tri 5289 17487 5387 17585 ne
rect 5387 17487 5741 17585
tri 5741 17487 5839 17585 sw
tri 5839 17487 5937 17585 ne
rect 5937 17487 6291 17585
tri 6291 17487 6389 17585 sw
tri 6389 17487 6487 17585 ne
rect 6487 17487 6841 17585
tri 6841 17487 6939 17585 sw
tri 6939 17487 7037 17585 ne
rect 7037 17487 7391 17585
tri 7391 17487 7489 17585 sw
tri 7489 17487 7587 17585 ne
rect 7587 17487 7941 17585
tri 7941 17487 8039 17585 sw
tri 8039 17487 8137 17585 ne
rect 8137 17487 8491 17585
tri 8491 17487 8589 17585 sw
tri 8589 17487 8687 17585 ne
rect 8687 17487 9041 17585
tri 9041 17487 9139 17585 sw
tri 9139 17487 9237 17585 ne
rect 9237 17487 9591 17585
tri 9591 17487 9689 17585 sw
tri 9689 17487 9787 17585 ne
rect 9787 17487 10141 17585
tri 10141 17487 10239 17585 sw
tri 10239 17487 10337 17585 ne
rect 10337 17487 10691 17585
tri 10691 17487 10789 17585 sw
tri 10789 17487 10887 17585 ne
rect 10887 17487 11241 17585
tri 11241 17487 11339 17585 sw
tri 11339 17487 11437 17585 ne
rect 11437 17487 11791 17585
tri 11791 17487 11889 17585 sw
tri 11889 17487 11987 17585 ne
rect 11987 17487 12341 17585
tri 12341 17487 12439 17585 sw
tri 12439 17487 12537 17585 ne
rect 12537 17487 12891 17585
tri 12891 17487 12989 17585 sw
tri 12989 17487 13087 17585 ne
rect 13087 17487 13441 17585
tri 13441 17487 13539 17585 sw
tri 13539 17487 13637 17585 ne
rect 13637 17487 13991 17585
tri 13991 17487 14089 17585 sw
tri 14089 17487 14187 17585 ne
rect 14187 17487 14541 17585
tri 14541 17487 14639 17585 sw
tri 14639 17487 14737 17585 ne
rect 14737 17487 15091 17585
tri 15091 17487 15189 17585 sw
tri 15189 17487 15287 17585 ne
rect 15287 17487 15641 17585
tri 15641 17487 15739 17585 sw
tri 15739 17487 15837 17585 ne
rect 15837 17487 16191 17585
tri 16191 17487 16289 17585 sw
tri 16289 17487 16387 17585 ne
rect 16387 17487 16741 17585
tri 16741 17487 16839 17585 sw
tri 16839 17487 16937 17585 ne
rect 16937 17487 17291 17585
tri 17291 17487 17389 17585 sw
tri 17389 17487 17487 17585 ne
rect 17487 17487 17841 17585
tri 17841 17487 17939 17585 sw
tri 17939 17487 18037 17585 ne
rect 18037 17487 18391 17585
tri 18391 17487 18489 17585 sw
tri 18489 17487 18587 17585 ne
rect 18587 17487 18941 17585
tri 18941 17487 19039 17585 sw
tri 19039 17487 19137 17585 ne
rect 19137 17487 19491 17585
tri 19491 17487 19589 17585 sw
tri 19589 17487 19687 17585 ne
rect 19687 17487 20300 17585
rect -2000 17389 339 17487
tri 339 17389 437 17487 sw
tri 437 17389 535 17487 ne
rect 535 17389 889 17487
tri 889 17389 987 17487 sw
tri 987 17389 1085 17487 ne
rect 1085 17389 1439 17487
tri 1439 17389 1537 17487 sw
tri 1537 17389 1635 17487 ne
rect 1635 17389 1989 17487
tri 1989 17389 2087 17487 sw
tri 2087 17389 2185 17487 ne
rect 2185 17389 2539 17487
tri 2539 17389 2637 17487 sw
tri 2637 17389 2735 17487 ne
rect 2735 17389 3089 17487
tri 3089 17389 3187 17487 sw
tri 3187 17389 3285 17487 ne
rect 3285 17389 3639 17487
tri 3639 17389 3737 17487 sw
tri 3737 17389 3835 17487 ne
rect 3835 17389 4189 17487
tri 4189 17389 4287 17487 sw
tri 4287 17389 4385 17487 ne
rect 4385 17389 4739 17487
tri 4739 17389 4837 17487 sw
tri 4837 17389 4935 17487 ne
rect 4935 17389 5289 17487
tri 5289 17389 5387 17487 sw
tri 5387 17389 5485 17487 ne
rect 5485 17389 5839 17487
tri 5839 17389 5937 17487 sw
tri 5937 17389 6035 17487 ne
rect 6035 17389 6389 17487
tri 6389 17389 6487 17487 sw
tri 6487 17389 6585 17487 ne
rect 6585 17389 6939 17487
tri 6939 17389 7037 17487 sw
tri 7037 17389 7135 17487 ne
rect 7135 17389 7489 17487
tri 7489 17389 7587 17487 sw
tri 7587 17389 7685 17487 ne
rect 7685 17389 8039 17487
tri 8039 17389 8137 17487 sw
tri 8137 17389 8235 17487 ne
rect 8235 17389 8589 17487
tri 8589 17389 8687 17487 sw
tri 8687 17389 8785 17487 ne
rect 8785 17389 9139 17487
tri 9139 17389 9237 17487 sw
tri 9237 17389 9335 17487 ne
rect 9335 17389 9689 17487
tri 9689 17389 9787 17487 sw
tri 9787 17389 9885 17487 ne
rect 9885 17389 10239 17487
tri 10239 17389 10337 17487 sw
tri 10337 17389 10435 17487 ne
rect 10435 17389 10789 17487
tri 10789 17389 10887 17487 sw
tri 10887 17389 10985 17487 ne
rect 10985 17389 11339 17487
tri 11339 17389 11437 17487 sw
tri 11437 17389 11535 17487 ne
rect 11535 17389 11889 17487
tri 11889 17389 11987 17487 sw
tri 11987 17389 12085 17487 ne
rect 12085 17389 12439 17487
tri 12439 17389 12537 17487 sw
tri 12537 17389 12635 17487 ne
rect 12635 17389 12989 17487
tri 12989 17389 13087 17487 sw
tri 13087 17389 13185 17487 ne
rect 13185 17389 13539 17487
tri 13539 17389 13637 17487 sw
tri 13637 17389 13735 17487 ne
rect 13735 17389 14089 17487
tri 14089 17389 14187 17487 sw
tri 14187 17389 14285 17487 ne
rect 14285 17389 14639 17487
tri 14639 17389 14737 17487 sw
tri 14737 17389 14835 17487 ne
rect 14835 17389 15189 17487
tri 15189 17389 15287 17487 sw
tri 15287 17389 15385 17487 ne
rect 15385 17389 15739 17487
tri 15739 17389 15837 17487 sw
tri 15837 17389 15935 17487 ne
rect 15935 17389 16289 17487
tri 16289 17389 16387 17487 sw
tri 16387 17389 16485 17487 ne
rect 16485 17389 16839 17487
tri 16839 17389 16937 17487 sw
tri 16937 17389 17035 17487 ne
rect 17035 17389 17389 17487
tri 17389 17389 17487 17487 sw
tri 17487 17389 17585 17487 ne
rect 17585 17389 17939 17487
tri 17939 17389 18037 17487 sw
tri 18037 17389 18135 17487 ne
rect 18135 17389 18489 17487
tri 18489 17389 18587 17487 sw
tri 18587 17389 18685 17487 ne
rect 18685 17389 19039 17487
tri 19039 17389 19137 17487 sw
tri 19137 17389 19235 17487 ne
rect 19235 17389 19589 17487
tri 19589 17389 19687 17487 sw
rect 20800 17389 21800 18037
rect -2000 17385 437 17389
rect -2000 17265 215 17385
rect 335 17291 437 17385
tri 437 17291 535 17389 sw
tri 535 17291 633 17389 ne
rect 633 17385 987 17389
rect 633 17291 765 17385
rect 335 17265 535 17291
rect -2000 17261 535 17265
rect -2000 16613 -1000 17261
tri 113 17163 211 17261 ne
rect 211 17213 535 17261
tri 535 17213 613 17291 sw
tri 633 17213 711 17291 ne
rect 711 17265 765 17291
rect 885 17291 987 17385
tri 987 17291 1085 17389 sw
tri 1085 17291 1183 17389 ne
rect 1183 17385 1537 17389
rect 1183 17291 1315 17385
rect 885 17265 1085 17291
rect 711 17213 1085 17265
tri 1085 17213 1163 17291 sw
tri 1183 17213 1261 17291 ne
rect 1261 17265 1315 17291
rect 1435 17291 1537 17385
tri 1537 17291 1635 17389 sw
tri 1635 17291 1733 17389 ne
rect 1733 17385 2087 17389
rect 1733 17291 1865 17385
rect 1435 17265 1635 17291
rect 1261 17213 1635 17265
tri 1635 17213 1713 17291 sw
tri 1733 17213 1811 17291 ne
rect 1811 17265 1865 17291
rect 1985 17291 2087 17385
tri 2087 17291 2185 17389 sw
tri 2185 17291 2283 17389 ne
rect 2283 17385 2637 17389
rect 2283 17291 2415 17385
rect 1985 17265 2185 17291
rect 1811 17213 2185 17265
tri 2185 17213 2263 17291 sw
tri 2283 17213 2361 17291 ne
rect 2361 17265 2415 17291
rect 2535 17291 2637 17385
tri 2637 17291 2735 17389 sw
tri 2735 17291 2833 17389 ne
rect 2833 17385 3187 17389
rect 2833 17291 2965 17385
rect 2535 17265 2735 17291
rect 2361 17213 2735 17265
tri 2735 17213 2813 17291 sw
tri 2833 17213 2911 17291 ne
rect 2911 17265 2965 17291
rect 3085 17291 3187 17385
tri 3187 17291 3285 17389 sw
tri 3285 17291 3383 17389 ne
rect 3383 17385 3737 17389
rect 3383 17291 3515 17385
rect 3085 17265 3285 17291
rect 2911 17213 3285 17265
tri 3285 17213 3363 17291 sw
tri 3383 17213 3461 17291 ne
rect 3461 17265 3515 17291
rect 3635 17291 3737 17385
tri 3737 17291 3835 17389 sw
tri 3835 17291 3933 17389 ne
rect 3933 17385 4287 17389
rect 3933 17291 4065 17385
rect 3635 17265 3835 17291
rect 3461 17213 3835 17265
tri 3835 17213 3913 17291 sw
tri 3933 17213 4011 17291 ne
rect 4011 17265 4065 17291
rect 4185 17291 4287 17385
tri 4287 17291 4385 17389 sw
tri 4385 17291 4483 17389 ne
rect 4483 17385 4837 17389
rect 4483 17291 4615 17385
rect 4185 17265 4385 17291
rect 4011 17213 4385 17265
tri 4385 17213 4463 17291 sw
tri 4483 17213 4561 17291 ne
rect 4561 17265 4615 17291
rect 4735 17291 4837 17385
tri 4837 17291 4935 17389 sw
tri 4935 17291 5033 17389 ne
rect 5033 17385 5387 17389
rect 5033 17291 5165 17385
rect 4735 17265 4935 17291
rect 4561 17213 4935 17265
tri 4935 17213 5013 17291 sw
tri 5033 17213 5111 17291 ne
rect 5111 17265 5165 17291
rect 5285 17291 5387 17385
tri 5387 17291 5485 17389 sw
tri 5485 17291 5583 17389 ne
rect 5583 17385 5937 17389
rect 5583 17291 5715 17385
rect 5285 17265 5485 17291
rect 5111 17213 5485 17265
tri 5485 17213 5563 17291 sw
tri 5583 17213 5661 17291 ne
rect 5661 17265 5715 17291
rect 5835 17291 5937 17385
tri 5937 17291 6035 17389 sw
tri 6035 17291 6133 17389 ne
rect 6133 17385 6487 17389
rect 6133 17291 6265 17385
rect 5835 17265 6035 17291
rect 5661 17213 6035 17265
tri 6035 17213 6113 17291 sw
tri 6133 17213 6211 17291 ne
rect 6211 17265 6265 17291
rect 6385 17291 6487 17385
tri 6487 17291 6585 17389 sw
tri 6585 17291 6683 17389 ne
rect 6683 17385 7037 17389
rect 6683 17291 6815 17385
rect 6385 17265 6585 17291
rect 6211 17213 6585 17265
tri 6585 17213 6663 17291 sw
tri 6683 17213 6761 17291 ne
rect 6761 17265 6815 17291
rect 6935 17291 7037 17385
tri 7037 17291 7135 17389 sw
tri 7135 17291 7233 17389 ne
rect 7233 17385 7587 17389
rect 7233 17291 7365 17385
rect 6935 17265 7135 17291
rect 6761 17213 7135 17265
tri 7135 17213 7213 17291 sw
tri 7233 17213 7311 17291 ne
rect 7311 17265 7365 17291
rect 7485 17291 7587 17385
tri 7587 17291 7685 17389 sw
tri 7685 17291 7783 17389 ne
rect 7783 17385 8137 17389
rect 7783 17291 7915 17385
rect 7485 17265 7685 17291
rect 7311 17213 7685 17265
tri 7685 17213 7763 17291 sw
tri 7783 17213 7861 17291 ne
rect 7861 17265 7915 17291
rect 8035 17291 8137 17385
tri 8137 17291 8235 17389 sw
tri 8235 17291 8333 17389 ne
rect 8333 17385 8687 17389
rect 8333 17291 8465 17385
rect 8035 17265 8235 17291
rect 7861 17213 8235 17265
tri 8235 17213 8313 17291 sw
tri 8333 17213 8411 17291 ne
rect 8411 17265 8465 17291
rect 8585 17291 8687 17385
tri 8687 17291 8785 17389 sw
tri 8785 17291 8883 17389 ne
rect 8883 17385 9237 17389
rect 8883 17291 9015 17385
rect 8585 17265 8785 17291
rect 8411 17213 8785 17265
tri 8785 17213 8863 17291 sw
tri 8883 17213 8961 17291 ne
rect 8961 17265 9015 17291
rect 9135 17291 9237 17385
tri 9237 17291 9335 17389 sw
tri 9335 17291 9433 17389 ne
rect 9433 17385 9787 17389
rect 9433 17291 9565 17385
rect 9135 17265 9335 17291
rect 8961 17213 9335 17265
tri 9335 17213 9413 17291 sw
tri 9433 17213 9511 17291 ne
rect 9511 17265 9565 17291
rect 9685 17291 9787 17385
tri 9787 17291 9885 17389 sw
tri 9885 17291 9983 17389 ne
rect 9983 17385 10337 17389
rect 9983 17291 10115 17385
rect 9685 17265 9885 17291
rect 9511 17213 9885 17265
tri 9885 17213 9963 17291 sw
tri 9983 17213 10061 17291 ne
rect 10061 17265 10115 17291
rect 10235 17291 10337 17385
tri 10337 17291 10435 17389 sw
tri 10435 17291 10533 17389 ne
rect 10533 17385 10887 17389
rect 10533 17291 10665 17385
rect 10235 17265 10435 17291
rect 10061 17213 10435 17265
tri 10435 17213 10513 17291 sw
tri 10533 17213 10611 17291 ne
rect 10611 17265 10665 17291
rect 10785 17291 10887 17385
tri 10887 17291 10985 17389 sw
tri 10985 17291 11083 17389 ne
rect 11083 17385 11437 17389
rect 11083 17291 11215 17385
rect 10785 17265 10985 17291
rect 10611 17213 10985 17265
tri 10985 17213 11063 17291 sw
tri 11083 17213 11161 17291 ne
rect 11161 17265 11215 17291
rect 11335 17291 11437 17385
tri 11437 17291 11535 17389 sw
tri 11535 17291 11633 17389 ne
rect 11633 17385 11987 17389
rect 11633 17291 11765 17385
rect 11335 17265 11535 17291
rect 11161 17213 11535 17265
tri 11535 17213 11613 17291 sw
tri 11633 17213 11711 17291 ne
rect 11711 17265 11765 17291
rect 11885 17291 11987 17385
tri 11987 17291 12085 17389 sw
tri 12085 17291 12183 17389 ne
rect 12183 17385 12537 17389
rect 12183 17291 12315 17385
rect 11885 17265 12085 17291
rect 11711 17213 12085 17265
tri 12085 17213 12163 17291 sw
tri 12183 17213 12261 17291 ne
rect 12261 17265 12315 17291
rect 12435 17291 12537 17385
tri 12537 17291 12635 17389 sw
tri 12635 17291 12733 17389 ne
rect 12733 17385 13087 17389
rect 12733 17291 12865 17385
rect 12435 17265 12635 17291
rect 12261 17213 12635 17265
tri 12635 17213 12713 17291 sw
tri 12733 17213 12811 17291 ne
rect 12811 17265 12865 17291
rect 12985 17291 13087 17385
tri 13087 17291 13185 17389 sw
tri 13185 17291 13283 17389 ne
rect 13283 17385 13637 17389
rect 13283 17291 13415 17385
rect 12985 17265 13185 17291
rect 12811 17213 13185 17265
tri 13185 17213 13263 17291 sw
tri 13283 17213 13361 17291 ne
rect 13361 17265 13415 17291
rect 13535 17291 13637 17385
tri 13637 17291 13735 17389 sw
tri 13735 17291 13833 17389 ne
rect 13833 17385 14187 17389
rect 13833 17291 13965 17385
rect 13535 17265 13735 17291
rect 13361 17213 13735 17265
tri 13735 17213 13813 17291 sw
tri 13833 17213 13911 17291 ne
rect 13911 17265 13965 17291
rect 14085 17291 14187 17385
tri 14187 17291 14285 17389 sw
tri 14285 17291 14383 17389 ne
rect 14383 17385 14737 17389
rect 14383 17291 14515 17385
rect 14085 17265 14285 17291
rect 13911 17213 14285 17265
tri 14285 17213 14363 17291 sw
tri 14383 17213 14461 17291 ne
rect 14461 17265 14515 17291
rect 14635 17291 14737 17385
tri 14737 17291 14835 17389 sw
tri 14835 17291 14933 17389 ne
rect 14933 17385 15287 17389
rect 14933 17291 15065 17385
rect 14635 17265 14835 17291
rect 14461 17213 14835 17265
tri 14835 17213 14913 17291 sw
tri 14933 17213 15011 17291 ne
rect 15011 17265 15065 17291
rect 15185 17291 15287 17385
tri 15287 17291 15385 17389 sw
tri 15385 17291 15483 17389 ne
rect 15483 17385 15837 17389
rect 15483 17291 15615 17385
rect 15185 17265 15385 17291
rect 15011 17213 15385 17265
tri 15385 17213 15463 17291 sw
tri 15483 17213 15561 17291 ne
rect 15561 17265 15615 17291
rect 15735 17291 15837 17385
tri 15837 17291 15935 17389 sw
tri 15935 17291 16033 17389 ne
rect 16033 17385 16387 17389
rect 16033 17291 16165 17385
rect 15735 17265 15935 17291
rect 15561 17213 15935 17265
tri 15935 17213 16013 17291 sw
tri 16033 17213 16111 17291 ne
rect 16111 17265 16165 17291
rect 16285 17291 16387 17385
tri 16387 17291 16485 17389 sw
tri 16485 17291 16583 17389 ne
rect 16583 17385 16937 17389
rect 16583 17291 16715 17385
rect 16285 17265 16485 17291
rect 16111 17213 16485 17265
tri 16485 17213 16563 17291 sw
tri 16583 17213 16661 17291 ne
rect 16661 17265 16715 17291
rect 16835 17291 16937 17385
tri 16937 17291 17035 17389 sw
tri 17035 17291 17133 17389 ne
rect 17133 17385 17487 17389
rect 17133 17291 17265 17385
rect 16835 17265 17035 17291
rect 16661 17213 17035 17265
tri 17035 17213 17113 17291 sw
tri 17133 17213 17211 17291 ne
rect 17211 17265 17265 17291
rect 17385 17291 17487 17385
tri 17487 17291 17585 17389 sw
tri 17585 17291 17683 17389 ne
rect 17683 17385 18037 17389
rect 17683 17291 17815 17385
rect 17385 17265 17585 17291
rect 17211 17213 17585 17265
tri 17585 17213 17663 17291 sw
tri 17683 17213 17761 17291 ne
rect 17761 17265 17815 17291
rect 17935 17291 18037 17385
tri 18037 17291 18135 17389 sw
tri 18135 17291 18233 17389 ne
rect 18233 17385 18587 17389
rect 18233 17291 18365 17385
rect 17935 17265 18135 17291
rect 17761 17213 18135 17265
tri 18135 17213 18213 17291 sw
tri 18233 17213 18311 17291 ne
rect 18311 17265 18365 17291
rect 18485 17291 18587 17385
tri 18587 17291 18685 17389 sw
tri 18685 17291 18783 17389 ne
rect 18783 17385 19137 17389
rect 18783 17291 18915 17385
rect 18485 17265 18685 17291
rect 18311 17213 18685 17265
tri 18685 17213 18763 17291 sw
tri 18783 17213 18861 17291 ne
rect 18861 17265 18915 17291
rect 19035 17291 19137 17385
tri 19137 17291 19235 17389 sw
tri 19235 17291 19333 17389 ne
rect 19333 17385 21800 17389
rect 19333 17291 19465 17385
rect 19035 17265 19235 17291
rect 18861 17213 19235 17265
tri 19235 17213 19313 17291 sw
tri 19333 17213 19411 17291 ne
rect 19411 17265 19465 17291
rect 19585 17265 21800 17385
rect 19411 17213 21800 17265
rect 211 17163 613 17213
rect -500 17113 113 17163
tri 113 17113 163 17163 sw
tri 211 17113 261 17163 ne
rect 261 17133 613 17163
tri 613 17133 693 17213 sw
tri 711 17133 791 17213 ne
rect 791 17133 1163 17213
tri 1163 17133 1243 17213 sw
tri 1261 17133 1341 17213 ne
rect 1341 17133 1713 17213
tri 1713 17133 1793 17213 sw
tri 1811 17133 1891 17213 ne
rect 1891 17133 2263 17213
tri 2263 17133 2343 17213 sw
tri 2361 17133 2441 17213 ne
rect 2441 17133 2813 17213
tri 2813 17133 2893 17213 sw
tri 2911 17133 2991 17213 ne
rect 2991 17133 3363 17213
tri 3363 17133 3443 17213 sw
tri 3461 17133 3541 17213 ne
rect 3541 17133 3913 17213
tri 3913 17133 3993 17213 sw
tri 4011 17133 4091 17213 ne
rect 4091 17133 4463 17213
tri 4463 17133 4543 17213 sw
tri 4561 17133 4641 17213 ne
rect 4641 17133 5013 17213
tri 5013 17133 5093 17213 sw
tri 5111 17133 5191 17213 ne
rect 5191 17133 5563 17213
tri 5563 17133 5643 17213 sw
tri 5661 17133 5741 17213 ne
rect 5741 17133 6113 17213
tri 6113 17133 6193 17213 sw
tri 6211 17133 6291 17213 ne
rect 6291 17133 6663 17213
tri 6663 17133 6743 17213 sw
tri 6761 17133 6841 17213 ne
rect 6841 17133 7213 17213
tri 7213 17133 7293 17213 sw
tri 7311 17133 7391 17213 ne
rect 7391 17133 7763 17213
tri 7763 17133 7843 17213 sw
tri 7861 17133 7941 17213 ne
rect 7941 17133 8313 17213
tri 8313 17133 8393 17213 sw
tri 8411 17133 8491 17213 ne
rect 8491 17133 8863 17213
tri 8863 17133 8943 17213 sw
tri 8961 17133 9041 17213 ne
rect 9041 17133 9413 17213
tri 9413 17133 9493 17213 sw
tri 9511 17133 9591 17213 ne
rect 9591 17133 9963 17213
tri 9963 17133 10043 17213 sw
tri 10061 17133 10141 17213 ne
rect 10141 17133 10513 17213
tri 10513 17133 10593 17213 sw
tri 10611 17133 10691 17213 ne
rect 10691 17133 11063 17213
tri 11063 17133 11143 17213 sw
tri 11161 17133 11241 17213 ne
rect 11241 17133 11613 17213
tri 11613 17133 11693 17213 sw
tri 11711 17133 11791 17213 ne
rect 11791 17133 12163 17213
tri 12163 17133 12243 17213 sw
tri 12261 17133 12341 17213 ne
rect 12341 17133 12713 17213
tri 12713 17133 12793 17213 sw
tri 12811 17133 12891 17213 ne
rect 12891 17133 13263 17213
tri 13263 17133 13343 17213 sw
tri 13361 17133 13441 17213 ne
rect 13441 17133 13813 17213
tri 13813 17133 13893 17213 sw
tri 13911 17133 13991 17213 ne
rect 13991 17133 14363 17213
tri 14363 17133 14443 17213 sw
tri 14461 17133 14541 17213 ne
rect 14541 17133 14913 17213
tri 14913 17133 14993 17213 sw
tri 15011 17133 15091 17213 ne
rect 15091 17133 15463 17213
tri 15463 17133 15543 17213 sw
tri 15561 17133 15641 17213 ne
rect 15641 17133 16013 17213
tri 16013 17133 16093 17213 sw
tri 16111 17133 16191 17213 ne
rect 16191 17133 16563 17213
tri 16563 17133 16643 17213 sw
tri 16661 17133 16741 17213 ne
rect 16741 17133 17113 17213
tri 17113 17133 17193 17213 sw
tri 17211 17133 17291 17213 ne
rect 17291 17133 17663 17213
tri 17663 17133 17743 17213 sw
tri 17761 17133 17841 17213 ne
rect 17841 17133 18213 17213
tri 18213 17133 18293 17213 sw
tri 18311 17133 18391 17213 ne
rect 18391 17133 18763 17213
tri 18763 17133 18843 17213 sw
tri 18861 17133 18941 17213 ne
rect 18941 17133 19313 17213
tri 19313 17133 19393 17213 sw
tri 19411 17133 19491 17213 ne
rect 19491 17133 20100 17213
rect 261 17113 693 17133
rect -500 17035 163 17113
tri 163 17035 241 17113 sw
tri 261 17035 339 17113 ne
rect 339 17035 693 17113
tri 693 17035 791 17133 sw
tri 791 17035 889 17133 ne
rect 889 17035 1243 17133
tri 1243 17035 1341 17133 sw
tri 1341 17035 1439 17133 ne
rect 1439 17035 1793 17133
tri 1793 17035 1891 17133 sw
tri 1891 17035 1989 17133 ne
rect 1989 17035 2343 17133
tri 2343 17035 2441 17133 sw
tri 2441 17035 2539 17133 ne
rect 2539 17035 2893 17133
tri 2893 17035 2991 17133 sw
tri 2991 17035 3089 17133 ne
rect 3089 17035 3443 17133
tri 3443 17035 3541 17133 sw
tri 3541 17035 3639 17133 ne
rect 3639 17035 3993 17133
tri 3993 17035 4091 17133 sw
tri 4091 17035 4189 17133 ne
rect 4189 17035 4543 17133
tri 4543 17035 4641 17133 sw
tri 4641 17035 4739 17133 ne
rect 4739 17035 5093 17133
tri 5093 17035 5191 17133 sw
tri 5191 17035 5289 17133 ne
rect 5289 17035 5643 17133
tri 5643 17035 5741 17133 sw
tri 5741 17035 5839 17133 ne
rect 5839 17035 6193 17133
tri 6193 17035 6291 17133 sw
tri 6291 17035 6389 17133 ne
rect 6389 17035 6743 17133
tri 6743 17035 6841 17133 sw
tri 6841 17035 6939 17133 ne
rect 6939 17035 7293 17133
tri 7293 17035 7391 17133 sw
tri 7391 17035 7489 17133 ne
rect 7489 17035 7843 17133
tri 7843 17035 7941 17133 sw
tri 7941 17035 8039 17133 ne
rect 8039 17035 8393 17133
tri 8393 17035 8491 17133 sw
tri 8491 17035 8589 17133 ne
rect 8589 17035 8943 17133
tri 8943 17035 9041 17133 sw
tri 9041 17035 9139 17133 ne
rect 9139 17035 9493 17133
tri 9493 17035 9591 17133 sw
tri 9591 17035 9689 17133 ne
rect 9689 17035 10043 17133
tri 10043 17035 10141 17133 sw
tri 10141 17035 10239 17133 ne
rect 10239 17035 10593 17133
tri 10593 17035 10691 17133 sw
tri 10691 17035 10789 17133 ne
rect 10789 17035 11143 17133
tri 11143 17035 11241 17133 sw
tri 11241 17035 11339 17133 ne
rect 11339 17035 11693 17133
tri 11693 17035 11791 17133 sw
tri 11791 17035 11889 17133 ne
rect 11889 17035 12243 17133
tri 12243 17035 12341 17133 sw
tri 12341 17035 12439 17133 ne
rect 12439 17035 12793 17133
tri 12793 17035 12891 17133 sw
tri 12891 17035 12989 17133 ne
rect 12989 17035 13343 17133
tri 13343 17035 13441 17133 sw
tri 13441 17035 13539 17133 ne
rect 13539 17035 13893 17133
tri 13893 17035 13991 17133 sw
tri 13991 17035 14089 17133 ne
rect 14089 17035 14443 17133
tri 14443 17035 14541 17133 sw
tri 14541 17035 14639 17133 ne
rect 14639 17035 14993 17133
tri 14993 17035 15091 17133 sw
tri 15091 17035 15189 17133 ne
rect 15189 17035 15543 17133
tri 15543 17035 15641 17133 sw
tri 15641 17035 15739 17133 ne
rect 15739 17035 16093 17133
tri 16093 17035 16191 17133 sw
tri 16191 17035 16289 17133 ne
rect 16289 17035 16643 17133
tri 16643 17035 16741 17133 sw
tri 16741 17035 16839 17133 ne
rect 16839 17035 17193 17133
tri 17193 17035 17291 17133 sw
tri 17291 17035 17389 17133 ne
rect 17389 17035 17743 17133
tri 17743 17035 17841 17133 sw
tri 17841 17035 17939 17133 ne
rect 17939 17035 18293 17133
tri 18293 17035 18391 17133 sw
tri 18391 17035 18489 17133 ne
rect 18489 17035 18843 17133
tri 18843 17035 18941 17133 sw
tri 18941 17035 19039 17133 ne
rect 19039 17035 19393 17133
tri 19393 17035 19491 17133 sw
tri 19491 17035 19589 17133 ne
rect 19589 17113 20100 17133
rect 20200 17113 21800 17213
rect 19589 17035 21800 17113
rect -500 16987 241 17035
rect -500 16887 -400 16987
rect -300 16937 241 16987
tri 241 16937 339 17035 sw
tri 339 16937 437 17035 ne
rect 437 16937 791 17035
tri 791 16937 889 17035 sw
tri 889 16937 987 17035 ne
rect 987 16937 1341 17035
tri 1341 16937 1439 17035 sw
tri 1439 16937 1537 17035 ne
rect 1537 16937 1891 17035
tri 1891 16937 1989 17035 sw
tri 1989 16937 2087 17035 ne
rect 2087 16937 2441 17035
tri 2441 16937 2539 17035 sw
tri 2539 16937 2637 17035 ne
rect 2637 16937 2991 17035
tri 2991 16937 3089 17035 sw
tri 3089 16937 3187 17035 ne
rect 3187 16937 3541 17035
tri 3541 16937 3639 17035 sw
tri 3639 16937 3737 17035 ne
rect 3737 16937 4091 17035
tri 4091 16937 4189 17035 sw
tri 4189 16937 4287 17035 ne
rect 4287 16937 4641 17035
tri 4641 16937 4739 17035 sw
tri 4739 16937 4837 17035 ne
rect 4837 16937 5191 17035
tri 5191 16937 5289 17035 sw
tri 5289 16937 5387 17035 ne
rect 5387 16937 5741 17035
tri 5741 16937 5839 17035 sw
tri 5839 16937 5937 17035 ne
rect 5937 16937 6291 17035
tri 6291 16937 6389 17035 sw
tri 6389 16937 6487 17035 ne
rect 6487 16937 6841 17035
tri 6841 16937 6939 17035 sw
tri 6939 16937 7037 17035 ne
rect 7037 16937 7391 17035
tri 7391 16937 7489 17035 sw
tri 7489 16937 7587 17035 ne
rect 7587 16937 7941 17035
tri 7941 16937 8039 17035 sw
tri 8039 16937 8137 17035 ne
rect 8137 16937 8491 17035
tri 8491 16937 8589 17035 sw
tri 8589 16937 8687 17035 ne
rect 8687 16937 9041 17035
tri 9041 16937 9139 17035 sw
tri 9139 16937 9237 17035 ne
rect 9237 16937 9591 17035
tri 9591 16937 9689 17035 sw
tri 9689 16937 9787 17035 ne
rect 9787 16937 10141 17035
tri 10141 16937 10239 17035 sw
tri 10239 16937 10337 17035 ne
rect 10337 16937 10691 17035
tri 10691 16937 10789 17035 sw
tri 10789 16937 10887 17035 ne
rect 10887 16937 11241 17035
tri 11241 16937 11339 17035 sw
tri 11339 16937 11437 17035 ne
rect 11437 16937 11791 17035
tri 11791 16937 11889 17035 sw
tri 11889 16937 11987 17035 ne
rect 11987 16937 12341 17035
tri 12341 16937 12439 17035 sw
tri 12439 16937 12537 17035 ne
rect 12537 16937 12891 17035
tri 12891 16937 12989 17035 sw
tri 12989 16937 13087 17035 ne
rect 13087 16937 13441 17035
tri 13441 16937 13539 17035 sw
tri 13539 16937 13637 17035 ne
rect 13637 16937 13991 17035
tri 13991 16937 14089 17035 sw
tri 14089 16937 14187 17035 ne
rect 14187 16937 14541 17035
tri 14541 16937 14639 17035 sw
tri 14639 16937 14737 17035 ne
rect 14737 16937 15091 17035
tri 15091 16937 15189 17035 sw
tri 15189 16937 15287 17035 ne
rect 15287 16937 15641 17035
tri 15641 16937 15739 17035 sw
tri 15739 16937 15837 17035 ne
rect 15837 16937 16191 17035
tri 16191 16937 16289 17035 sw
tri 16289 16937 16387 17035 ne
rect 16387 16937 16741 17035
tri 16741 16937 16839 17035 sw
tri 16839 16937 16937 17035 ne
rect 16937 16937 17291 17035
tri 17291 16937 17389 17035 sw
tri 17389 16937 17487 17035 ne
rect 17487 16937 17841 17035
tri 17841 16937 17939 17035 sw
tri 17939 16937 18037 17035 ne
rect 18037 16937 18391 17035
tri 18391 16937 18489 17035 sw
tri 18489 16937 18587 17035 ne
rect 18587 16937 18941 17035
tri 18941 16937 19039 17035 sw
tri 19039 16937 19137 17035 ne
rect 19137 16937 19491 17035
tri 19491 16937 19589 17035 sw
tri 19589 16937 19687 17035 ne
rect 19687 16937 21800 17035
rect -300 16887 339 16937
rect -500 16839 339 16887
tri 339 16839 437 16937 sw
tri 437 16839 535 16937 ne
rect 535 16839 889 16937
tri 889 16839 987 16937 sw
tri 987 16839 1085 16937 ne
rect 1085 16839 1439 16937
tri 1439 16839 1537 16937 sw
tri 1537 16839 1635 16937 ne
rect 1635 16839 1989 16937
tri 1989 16839 2087 16937 sw
tri 2087 16839 2185 16937 ne
rect 2185 16839 2539 16937
tri 2539 16839 2637 16937 sw
tri 2637 16839 2735 16937 ne
rect 2735 16839 3089 16937
tri 3089 16839 3187 16937 sw
tri 3187 16839 3285 16937 ne
rect 3285 16839 3639 16937
tri 3639 16839 3737 16937 sw
tri 3737 16839 3835 16937 ne
rect 3835 16839 4189 16937
tri 4189 16839 4287 16937 sw
tri 4287 16839 4385 16937 ne
rect 4385 16839 4739 16937
tri 4739 16839 4837 16937 sw
tri 4837 16839 4935 16937 ne
rect 4935 16839 5289 16937
tri 5289 16839 5387 16937 sw
tri 5387 16839 5485 16937 ne
rect 5485 16839 5839 16937
tri 5839 16839 5937 16937 sw
tri 5937 16839 6035 16937 ne
rect 6035 16839 6389 16937
tri 6389 16839 6487 16937 sw
tri 6487 16839 6585 16937 ne
rect 6585 16839 6939 16937
tri 6939 16839 7037 16937 sw
tri 7037 16839 7135 16937 ne
rect 7135 16839 7489 16937
tri 7489 16839 7587 16937 sw
tri 7587 16839 7685 16937 ne
rect 7685 16839 8039 16937
tri 8039 16839 8137 16937 sw
tri 8137 16839 8235 16937 ne
rect 8235 16839 8589 16937
tri 8589 16839 8687 16937 sw
tri 8687 16839 8785 16937 ne
rect 8785 16839 9139 16937
tri 9139 16839 9237 16937 sw
tri 9237 16839 9335 16937 ne
rect 9335 16839 9689 16937
tri 9689 16839 9787 16937 sw
tri 9787 16839 9885 16937 ne
rect 9885 16839 10239 16937
tri 10239 16839 10337 16937 sw
tri 10337 16839 10435 16937 ne
rect 10435 16839 10789 16937
tri 10789 16839 10887 16937 sw
tri 10887 16839 10985 16937 ne
rect 10985 16839 11339 16937
tri 11339 16839 11437 16937 sw
tri 11437 16839 11535 16937 ne
rect 11535 16839 11889 16937
tri 11889 16839 11987 16937 sw
tri 11987 16839 12085 16937 ne
rect 12085 16839 12439 16937
tri 12439 16839 12537 16937 sw
tri 12537 16839 12635 16937 ne
rect 12635 16839 12989 16937
tri 12989 16839 13087 16937 sw
tri 13087 16839 13185 16937 ne
rect 13185 16839 13539 16937
tri 13539 16839 13637 16937 sw
tri 13637 16839 13735 16937 ne
rect 13735 16839 14089 16937
tri 14089 16839 14187 16937 sw
tri 14187 16839 14285 16937 ne
rect 14285 16839 14639 16937
tri 14639 16839 14737 16937 sw
tri 14737 16839 14835 16937 ne
rect 14835 16839 15189 16937
tri 15189 16839 15287 16937 sw
tri 15287 16839 15385 16937 ne
rect 15385 16839 15739 16937
tri 15739 16839 15837 16937 sw
tri 15837 16839 15935 16937 ne
rect 15935 16839 16289 16937
tri 16289 16839 16387 16937 sw
tri 16387 16839 16485 16937 ne
rect 16485 16839 16839 16937
tri 16839 16839 16937 16937 sw
tri 16937 16839 17035 16937 ne
rect 17035 16839 17389 16937
tri 17389 16839 17487 16937 sw
tri 17487 16839 17585 16937 ne
rect 17585 16839 17939 16937
tri 17939 16839 18037 16937 sw
tri 18037 16839 18135 16937 ne
rect 18135 16839 18489 16937
tri 18489 16839 18587 16937 sw
tri 18587 16839 18685 16937 ne
rect 18685 16839 19039 16937
tri 19039 16839 19137 16937 sw
tri 19137 16839 19235 16937 ne
rect 19235 16839 19589 16937
tri 19589 16839 19687 16937 sw
rect -500 16835 437 16839
rect -500 16715 215 16835
rect 335 16741 437 16835
tri 437 16741 535 16839 sw
tri 535 16741 633 16839 ne
rect 633 16835 987 16839
rect 633 16741 765 16835
rect 335 16715 535 16741
rect -500 16711 535 16715
tri 535 16711 565 16741 sw
tri 633 16711 663 16741 ne
rect 663 16715 765 16741
rect 885 16741 987 16835
tri 987 16741 1085 16839 sw
tri 1085 16741 1183 16839 ne
rect 1183 16835 1537 16839
rect 1183 16741 1315 16835
rect 885 16715 1085 16741
rect 663 16711 1085 16715
tri 1085 16711 1115 16741 sw
tri 1183 16711 1213 16741 ne
rect 1213 16715 1315 16741
rect 1435 16741 1537 16835
tri 1537 16741 1635 16839 sw
tri 1635 16741 1733 16839 ne
rect 1733 16835 2087 16839
rect 1733 16741 1865 16835
rect 1435 16715 1635 16741
rect 1213 16711 1635 16715
tri 1635 16711 1665 16741 sw
tri 1733 16711 1763 16741 ne
rect 1763 16715 1865 16741
rect 1985 16741 2087 16835
tri 2087 16741 2185 16839 sw
tri 2185 16741 2283 16839 ne
rect 2283 16835 2637 16839
rect 2283 16741 2415 16835
rect 1985 16715 2185 16741
rect 1763 16711 2185 16715
tri 2185 16711 2215 16741 sw
tri 2283 16711 2313 16741 ne
rect 2313 16715 2415 16741
rect 2535 16741 2637 16835
tri 2637 16741 2735 16839 sw
tri 2735 16741 2833 16839 ne
rect 2833 16835 3187 16839
rect 2833 16741 2965 16835
rect 2535 16715 2735 16741
rect 2313 16711 2735 16715
tri 2735 16711 2765 16741 sw
tri 2833 16711 2863 16741 ne
rect 2863 16715 2965 16741
rect 3085 16741 3187 16835
tri 3187 16741 3285 16839 sw
tri 3285 16741 3383 16839 ne
rect 3383 16835 3737 16839
rect 3383 16741 3515 16835
rect 3085 16715 3285 16741
rect 2863 16711 3285 16715
tri 3285 16711 3315 16741 sw
tri 3383 16711 3413 16741 ne
rect 3413 16715 3515 16741
rect 3635 16741 3737 16835
tri 3737 16741 3835 16839 sw
tri 3835 16741 3933 16839 ne
rect 3933 16835 4287 16839
rect 3933 16741 4065 16835
rect 3635 16715 3835 16741
rect 3413 16711 3835 16715
tri 3835 16711 3865 16741 sw
tri 3933 16711 3963 16741 ne
rect 3963 16715 4065 16741
rect 4185 16741 4287 16835
tri 4287 16741 4385 16839 sw
tri 4385 16741 4483 16839 ne
rect 4483 16835 4837 16839
rect 4483 16741 4615 16835
rect 4185 16715 4385 16741
rect 3963 16711 4385 16715
tri 4385 16711 4415 16741 sw
tri 4483 16711 4513 16741 ne
rect 4513 16715 4615 16741
rect 4735 16741 4837 16835
tri 4837 16741 4935 16839 sw
tri 4935 16741 5033 16839 ne
rect 5033 16835 5387 16839
rect 5033 16741 5165 16835
rect 4735 16715 4935 16741
rect 4513 16711 4935 16715
tri 4935 16711 4965 16741 sw
tri 5033 16711 5063 16741 ne
rect 5063 16715 5165 16741
rect 5285 16741 5387 16835
tri 5387 16741 5485 16839 sw
tri 5485 16741 5583 16839 ne
rect 5583 16835 5937 16839
rect 5583 16741 5715 16835
rect 5285 16715 5485 16741
rect 5063 16711 5485 16715
tri 5485 16711 5515 16741 sw
tri 5583 16711 5613 16741 ne
rect 5613 16715 5715 16741
rect 5835 16741 5937 16835
tri 5937 16741 6035 16839 sw
tri 6035 16741 6133 16839 ne
rect 6133 16835 6487 16839
rect 6133 16741 6265 16835
rect 5835 16715 6035 16741
rect 5613 16711 6035 16715
tri 6035 16711 6065 16741 sw
tri 6133 16711 6163 16741 ne
rect 6163 16715 6265 16741
rect 6385 16741 6487 16835
tri 6487 16741 6585 16839 sw
tri 6585 16741 6683 16839 ne
rect 6683 16835 7037 16839
rect 6683 16741 6815 16835
rect 6385 16715 6585 16741
rect 6163 16711 6585 16715
tri 6585 16711 6615 16741 sw
tri 6683 16711 6713 16741 ne
rect 6713 16715 6815 16741
rect 6935 16741 7037 16835
tri 7037 16741 7135 16839 sw
tri 7135 16741 7233 16839 ne
rect 7233 16835 7587 16839
rect 7233 16741 7365 16835
rect 6935 16715 7135 16741
rect 6713 16711 7135 16715
tri 7135 16711 7165 16741 sw
tri 7233 16711 7263 16741 ne
rect 7263 16715 7365 16741
rect 7485 16741 7587 16835
tri 7587 16741 7685 16839 sw
tri 7685 16741 7783 16839 ne
rect 7783 16835 8137 16839
rect 7783 16741 7915 16835
rect 7485 16715 7685 16741
rect 7263 16711 7685 16715
tri 7685 16711 7715 16741 sw
tri 7783 16711 7813 16741 ne
rect 7813 16715 7915 16741
rect 8035 16741 8137 16835
tri 8137 16741 8235 16839 sw
tri 8235 16741 8333 16839 ne
rect 8333 16835 8687 16839
rect 8333 16741 8465 16835
rect 8035 16715 8235 16741
rect 7813 16711 8235 16715
tri 8235 16711 8265 16741 sw
tri 8333 16711 8363 16741 ne
rect 8363 16715 8465 16741
rect 8585 16741 8687 16835
tri 8687 16741 8785 16839 sw
tri 8785 16741 8883 16839 ne
rect 8883 16835 9237 16839
rect 8883 16741 9015 16835
rect 8585 16715 8785 16741
rect 8363 16711 8785 16715
tri 8785 16711 8815 16741 sw
tri 8883 16711 8913 16741 ne
rect 8913 16715 9015 16741
rect 9135 16741 9237 16835
tri 9237 16741 9335 16839 sw
tri 9335 16741 9433 16839 ne
rect 9433 16835 9787 16839
rect 9433 16741 9565 16835
rect 9135 16715 9335 16741
rect 8913 16711 9335 16715
tri 9335 16711 9365 16741 sw
tri 9433 16711 9463 16741 ne
rect 9463 16715 9565 16741
rect 9685 16741 9787 16835
tri 9787 16741 9885 16839 sw
tri 9885 16741 9983 16839 ne
rect 9983 16835 10337 16839
rect 9983 16741 10115 16835
rect 9685 16715 9885 16741
rect 9463 16711 9885 16715
tri 9885 16711 9915 16741 sw
tri 9983 16711 10013 16741 ne
rect 10013 16715 10115 16741
rect 10235 16741 10337 16835
tri 10337 16741 10435 16839 sw
tri 10435 16741 10533 16839 ne
rect 10533 16835 10887 16839
rect 10533 16741 10665 16835
rect 10235 16715 10435 16741
rect 10013 16711 10435 16715
tri 10435 16711 10465 16741 sw
tri 10533 16711 10563 16741 ne
rect 10563 16715 10665 16741
rect 10785 16741 10887 16835
tri 10887 16741 10985 16839 sw
tri 10985 16741 11083 16839 ne
rect 11083 16835 11437 16839
rect 11083 16741 11215 16835
rect 10785 16715 10985 16741
rect 10563 16711 10985 16715
tri 10985 16711 11015 16741 sw
tri 11083 16711 11113 16741 ne
rect 11113 16715 11215 16741
rect 11335 16741 11437 16835
tri 11437 16741 11535 16839 sw
tri 11535 16741 11633 16839 ne
rect 11633 16835 11987 16839
rect 11633 16741 11765 16835
rect 11335 16715 11535 16741
rect 11113 16711 11535 16715
tri 11535 16711 11565 16741 sw
tri 11633 16711 11663 16741 ne
rect 11663 16715 11765 16741
rect 11885 16741 11987 16835
tri 11987 16741 12085 16839 sw
tri 12085 16741 12183 16839 ne
rect 12183 16835 12537 16839
rect 12183 16741 12315 16835
rect 11885 16715 12085 16741
rect 11663 16711 12085 16715
tri 12085 16711 12115 16741 sw
tri 12183 16711 12213 16741 ne
rect 12213 16715 12315 16741
rect 12435 16741 12537 16835
tri 12537 16741 12635 16839 sw
tri 12635 16741 12733 16839 ne
rect 12733 16835 13087 16839
rect 12733 16741 12865 16835
rect 12435 16715 12635 16741
rect 12213 16711 12635 16715
tri 12635 16711 12665 16741 sw
tri 12733 16711 12763 16741 ne
rect 12763 16715 12865 16741
rect 12985 16741 13087 16835
tri 13087 16741 13185 16839 sw
tri 13185 16741 13283 16839 ne
rect 13283 16835 13637 16839
rect 13283 16741 13415 16835
rect 12985 16715 13185 16741
rect 12763 16711 13185 16715
tri 13185 16711 13215 16741 sw
tri 13283 16711 13313 16741 ne
rect 13313 16715 13415 16741
rect 13535 16741 13637 16835
tri 13637 16741 13735 16839 sw
tri 13735 16741 13833 16839 ne
rect 13833 16835 14187 16839
rect 13833 16741 13965 16835
rect 13535 16715 13735 16741
rect 13313 16711 13735 16715
tri 13735 16711 13765 16741 sw
tri 13833 16711 13863 16741 ne
rect 13863 16715 13965 16741
rect 14085 16741 14187 16835
tri 14187 16741 14285 16839 sw
tri 14285 16741 14383 16839 ne
rect 14383 16835 14737 16839
rect 14383 16741 14515 16835
rect 14085 16715 14285 16741
rect 13863 16711 14285 16715
tri 14285 16711 14315 16741 sw
tri 14383 16711 14413 16741 ne
rect 14413 16715 14515 16741
rect 14635 16741 14737 16835
tri 14737 16741 14835 16839 sw
tri 14835 16741 14933 16839 ne
rect 14933 16835 15287 16839
rect 14933 16741 15065 16835
rect 14635 16715 14835 16741
rect 14413 16711 14835 16715
tri 14835 16711 14865 16741 sw
tri 14933 16711 14963 16741 ne
rect 14963 16715 15065 16741
rect 15185 16741 15287 16835
tri 15287 16741 15385 16839 sw
tri 15385 16741 15483 16839 ne
rect 15483 16835 15837 16839
rect 15483 16741 15615 16835
rect 15185 16715 15385 16741
rect 14963 16711 15385 16715
tri 15385 16711 15415 16741 sw
tri 15483 16711 15513 16741 ne
rect 15513 16715 15615 16741
rect 15735 16741 15837 16835
tri 15837 16741 15935 16839 sw
tri 15935 16741 16033 16839 ne
rect 16033 16835 16387 16839
rect 16033 16741 16165 16835
rect 15735 16715 15935 16741
rect 15513 16711 15935 16715
tri 15935 16711 15965 16741 sw
tri 16033 16711 16063 16741 ne
rect 16063 16715 16165 16741
rect 16285 16741 16387 16835
tri 16387 16741 16485 16839 sw
tri 16485 16741 16583 16839 ne
rect 16583 16835 16937 16839
rect 16583 16741 16715 16835
rect 16285 16715 16485 16741
rect 16063 16711 16485 16715
tri 16485 16711 16515 16741 sw
tri 16583 16711 16613 16741 ne
rect 16613 16715 16715 16741
rect 16835 16741 16937 16835
tri 16937 16741 17035 16839 sw
tri 17035 16741 17133 16839 ne
rect 17133 16835 17487 16839
rect 17133 16741 17265 16835
rect 16835 16715 17035 16741
rect 16613 16711 17035 16715
tri 17035 16711 17065 16741 sw
tri 17133 16711 17163 16741 ne
rect 17163 16715 17265 16741
rect 17385 16741 17487 16835
tri 17487 16741 17585 16839 sw
tri 17585 16741 17683 16839 ne
rect 17683 16835 18037 16839
rect 17683 16741 17815 16835
rect 17385 16715 17585 16741
rect 17163 16711 17585 16715
tri 17585 16711 17615 16741 sw
tri 17683 16711 17713 16741 ne
rect 17713 16715 17815 16741
rect 17935 16741 18037 16835
tri 18037 16741 18135 16839 sw
tri 18135 16741 18233 16839 ne
rect 18233 16835 18587 16839
rect 18233 16741 18365 16835
rect 17935 16715 18135 16741
rect 17713 16711 18135 16715
tri 18135 16711 18165 16741 sw
tri 18233 16711 18263 16741 ne
rect 18263 16715 18365 16741
rect 18485 16741 18587 16835
tri 18587 16741 18685 16839 sw
tri 18685 16741 18783 16839 ne
rect 18783 16835 19137 16839
rect 18783 16741 18915 16835
rect 18485 16715 18685 16741
rect 18263 16711 18685 16715
tri 18685 16711 18715 16741 sw
tri 18783 16711 18813 16741 ne
rect 18813 16715 18915 16741
rect 19035 16741 19137 16835
tri 19137 16741 19235 16839 sw
tri 19235 16741 19333 16839 ne
rect 19333 16835 20300 16839
rect 19333 16741 19465 16835
rect 19035 16715 19235 16741
rect 18813 16711 19235 16715
tri 19235 16711 19265 16741 sw
tri 19333 16711 19363 16741 ne
rect 19363 16715 19465 16741
rect 19585 16715 20300 16835
rect 19363 16711 20300 16715
tri 113 16613 211 16711 ne
rect 211 16613 565 16711
tri 565 16613 663 16711 sw
tri 663 16613 761 16711 ne
rect 761 16613 1115 16711
tri 1115 16613 1213 16711 sw
tri 1213 16613 1311 16711 ne
rect 1311 16613 1665 16711
tri 1665 16613 1763 16711 sw
tri 1763 16613 1861 16711 ne
rect 1861 16613 2215 16711
tri 2215 16613 2313 16711 sw
tri 2313 16613 2411 16711 ne
rect 2411 16613 2765 16711
tri 2765 16613 2863 16711 sw
tri 2863 16613 2961 16711 ne
rect 2961 16613 3315 16711
tri 3315 16613 3413 16711 sw
tri 3413 16613 3511 16711 ne
rect 3511 16613 3865 16711
tri 3865 16613 3963 16711 sw
tri 3963 16613 4061 16711 ne
rect 4061 16613 4415 16711
tri 4415 16613 4513 16711 sw
tri 4513 16613 4611 16711 ne
rect 4611 16613 4965 16711
tri 4965 16613 5063 16711 sw
tri 5063 16613 5161 16711 ne
rect 5161 16613 5515 16711
tri 5515 16613 5613 16711 sw
tri 5613 16613 5711 16711 ne
rect 5711 16613 6065 16711
tri 6065 16613 6163 16711 sw
tri 6163 16613 6261 16711 ne
rect 6261 16613 6615 16711
tri 6615 16613 6713 16711 sw
tri 6713 16613 6811 16711 ne
rect 6811 16613 7165 16711
tri 7165 16613 7263 16711 sw
tri 7263 16613 7361 16711 ne
rect 7361 16613 7715 16711
tri 7715 16613 7813 16711 sw
tri 7813 16613 7911 16711 ne
rect 7911 16613 8265 16711
tri 8265 16613 8363 16711 sw
tri 8363 16613 8461 16711 ne
rect 8461 16613 8815 16711
tri 8815 16613 8913 16711 sw
tri 8913 16613 9011 16711 ne
rect 9011 16613 9365 16711
tri 9365 16613 9463 16711 sw
tri 9463 16613 9561 16711 ne
rect 9561 16613 9915 16711
tri 9915 16613 10013 16711 sw
tri 10013 16613 10111 16711 ne
rect 10111 16613 10465 16711
tri 10465 16613 10563 16711 sw
tri 10563 16613 10661 16711 ne
rect 10661 16613 11015 16711
tri 11015 16613 11113 16711 sw
tri 11113 16613 11211 16711 ne
rect 11211 16613 11565 16711
tri 11565 16613 11663 16711 sw
tri 11663 16613 11761 16711 ne
rect 11761 16613 12115 16711
tri 12115 16613 12213 16711 sw
tri 12213 16613 12311 16711 ne
rect 12311 16613 12665 16711
tri 12665 16613 12763 16711 sw
tri 12763 16613 12861 16711 ne
rect 12861 16613 13215 16711
tri 13215 16613 13313 16711 sw
tri 13313 16613 13411 16711 ne
rect 13411 16613 13765 16711
tri 13765 16613 13863 16711 sw
tri 13863 16613 13961 16711 ne
rect 13961 16613 14315 16711
tri 14315 16613 14413 16711 sw
tri 14413 16613 14511 16711 ne
rect 14511 16613 14865 16711
tri 14865 16613 14963 16711 sw
tri 14963 16613 15061 16711 ne
rect 15061 16613 15415 16711
tri 15415 16613 15513 16711 sw
tri 15513 16613 15611 16711 ne
rect 15611 16613 15965 16711
tri 15965 16613 16063 16711 sw
tri 16063 16613 16161 16711 ne
rect 16161 16613 16515 16711
tri 16515 16613 16613 16711 sw
tri 16613 16613 16711 16711 ne
rect 16711 16613 17065 16711
tri 17065 16613 17163 16711 sw
tri 17163 16613 17261 16711 ne
rect 17261 16613 17615 16711
tri 17615 16613 17713 16711 sw
tri 17713 16613 17811 16711 ne
rect 17811 16613 18165 16711
tri 18165 16613 18263 16711 sw
tri 18263 16613 18361 16711 ne
rect 18361 16613 18715 16711
tri 18715 16613 18813 16711 sw
tri 18813 16613 18911 16711 ne
rect 18911 16613 19265 16711
tri 19265 16613 19363 16711 sw
tri 19363 16613 19461 16711 ne
rect 19461 16613 20300 16711
rect -2000 16583 113 16613
tri 113 16583 143 16613 sw
tri 211 16583 241 16613 ne
rect 241 16583 663 16613
tri 663 16583 693 16613 sw
tri 761 16583 791 16613 ne
rect 791 16583 1213 16613
tri 1213 16583 1243 16613 sw
tri 1311 16583 1341 16613 ne
rect 1341 16583 1763 16613
tri 1763 16583 1793 16613 sw
tri 1861 16583 1891 16613 ne
rect 1891 16583 2313 16613
tri 2313 16583 2343 16613 sw
tri 2411 16583 2441 16613 ne
rect 2441 16583 2863 16613
tri 2863 16583 2893 16613 sw
tri 2961 16583 2991 16613 ne
rect 2991 16583 3413 16613
tri 3413 16583 3443 16613 sw
tri 3511 16583 3541 16613 ne
rect 3541 16583 3963 16613
tri 3963 16583 3993 16613 sw
tri 4061 16583 4091 16613 ne
rect 4091 16583 4513 16613
tri 4513 16583 4543 16613 sw
tri 4611 16583 4641 16613 ne
rect 4641 16583 5063 16613
tri 5063 16583 5093 16613 sw
tri 5161 16583 5191 16613 ne
rect 5191 16583 5613 16613
tri 5613 16583 5643 16613 sw
tri 5711 16583 5741 16613 ne
rect 5741 16583 6163 16613
tri 6163 16583 6193 16613 sw
tri 6261 16583 6291 16613 ne
rect 6291 16583 6713 16613
tri 6713 16583 6743 16613 sw
tri 6811 16583 6841 16613 ne
rect 6841 16583 7263 16613
tri 7263 16583 7293 16613 sw
tri 7361 16583 7391 16613 ne
rect 7391 16583 7813 16613
tri 7813 16583 7843 16613 sw
tri 7911 16583 7941 16613 ne
rect 7941 16583 8363 16613
tri 8363 16583 8393 16613 sw
tri 8461 16583 8491 16613 ne
rect 8491 16583 8913 16613
tri 8913 16583 8943 16613 sw
tri 9011 16583 9041 16613 ne
rect 9041 16583 9463 16613
tri 9463 16583 9493 16613 sw
tri 9561 16583 9591 16613 ne
rect 9591 16583 10013 16613
tri 10013 16583 10043 16613 sw
tri 10111 16583 10141 16613 ne
rect 10141 16583 10563 16613
tri 10563 16583 10593 16613 sw
tri 10661 16583 10691 16613 ne
rect 10691 16583 11113 16613
tri 11113 16583 11143 16613 sw
tri 11211 16583 11241 16613 ne
rect 11241 16583 11663 16613
tri 11663 16583 11693 16613 sw
tri 11761 16583 11791 16613 ne
rect 11791 16583 12213 16613
tri 12213 16583 12243 16613 sw
tri 12311 16583 12341 16613 ne
rect 12341 16583 12763 16613
tri 12763 16583 12793 16613 sw
tri 12861 16583 12891 16613 ne
rect 12891 16583 13313 16613
tri 13313 16583 13343 16613 sw
tri 13411 16583 13441 16613 ne
rect 13441 16583 13863 16613
tri 13863 16583 13893 16613 sw
tri 13961 16583 13991 16613 ne
rect 13991 16583 14413 16613
tri 14413 16583 14443 16613 sw
tri 14511 16583 14541 16613 ne
rect 14541 16583 14963 16613
tri 14963 16583 14993 16613 sw
tri 15061 16583 15091 16613 ne
rect 15091 16583 15513 16613
tri 15513 16583 15543 16613 sw
tri 15611 16583 15641 16613 ne
rect 15641 16583 16063 16613
tri 16063 16583 16093 16613 sw
tri 16161 16583 16191 16613 ne
rect 16191 16583 16613 16613
tri 16613 16583 16643 16613 sw
tri 16711 16583 16741 16613 ne
rect 16741 16583 17163 16613
tri 17163 16583 17193 16613 sw
tri 17261 16583 17291 16613 ne
rect 17291 16583 17713 16613
tri 17713 16583 17743 16613 sw
tri 17811 16583 17841 16613 ne
rect 17841 16583 18263 16613
tri 18263 16583 18293 16613 sw
tri 18361 16583 18391 16613 ne
rect 18391 16583 18813 16613
tri 18813 16583 18843 16613 sw
tri 18911 16583 18941 16613 ne
rect 18941 16583 19363 16613
tri 19363 16583 19393 16613 sw
tri 19461 16583 19491 16613 ne
rect 19491 16583 20300 16613
rect -2000 16485 143 16583
tri 143 16485 241 16583 sw
tri 241 16485 339 16583 ne
rect 339 16485 693 16583
tri 693 16485 791 16583 sw
tri 791 16485 889 16583 ne
rect 889 16485 1243 16583
tri 1243 16485 1341 16583 sw
tri 1341 16485 1439 16583 ne
rect 1439 16485 1793 16583
tri 1793 16485 1891 16583 sw
tri 1891 16485 1989 16583 ne
rect 1989 16485 2343 16583
tri 2343 16485 2441 16583 sw
tri 2441 16485 2539 16583 ne
rect 2539 16485 2893 16583
tri 2893 16485 2991 16583 sw
tri 2991 16485 3089 16583 ne
rect 3089 16485 3443 16583
tri 3443 16485 3541 16583 sw
tri 3541 16485 3639 16583 ne
rect 3639 16485 3993 16583
tri 3993 16485 4091 16583 sw
tri 4091 16485 4189 16583 ne
rect 4189 16485 4543 16583
tri 4543 16485 4641 16583 sw
tri 4641 16485 4739 16583 ne
rect 4739 16485 5093 16583
tri 5093 16485 5191 16583 sw
tri 5191 16485 5289 16583 ne
rect 5289 16485 5643 16583
tri 5643 16485 5741 16583 sw
tri 5741 16485 5839 16583 ne
rect 5839 16485 6193 16583
tri 6193 16485 6291 16583 sw
tri 6291 16485 6389 16583 ne
rect 6389 16485 6743 16583
tri 6743 16485 6841 16583 sw
tri 6841 16485 6939 16583 ne
rect 6939 16485 7293 16583
tri 7293 16485 7391 16583 sw
tri 7391 16485 7489 16583 ne
rect 7489 16485 7843 16583
tri 7843 16485 7941 16583 sw
tri 7941 16485 8039 16583 ne
rect 8039 16485 8393 16583
tri 8393 16485 8491 16583 sw
tri 8491 16485 8589 16583 ne
rect 8589 16485 8943 16583
tri 8943 16485 9041 16583 sw
tri 9041 16485 9139 16583 ne
rect 9139 16485 9493 16583
tri 9493 16485 9591 16583 sw
tri 9591 16485 9689 16583 ne
rect 9689 16485 10043 16583
tri 10043 16485 10141 16583 sw
tri 10141 16485 10239 16583 ne
rect 10239 16485 10593 16583
tri 10593 16485 10691 16583 sw
tri 10691 16485 10789 16583 ne
rect 10789 16485 11143 16583
tri 11143 16485 11241 16583 sw
tri 11241 16485 11339 16583 ne
rect 11339 16485 11693 16583
tri 11693 16485 11791 16583 sw
tri 11791 16485 11889 16583 ne
rect 11889 16485 12243 16583
tri 12243 16485 12341 16583 sw
tri 12341 16485 12439 16583 ne
rect 12439 16485 12793 16583
tri 12793 16485 12891 16583 sw
tri 12891 16485 12989 16583 ne
rect 12989 16485 13343 16583
tri 13343 16485 13441 16583 sw
tri 13441 16485 13539 16583 ne
rect 13539 16485 13893 16583
tri 13893 16485 13991 16583 sw
tri 13991 16485 14089 16583 ne
rect 14089 16485 14443 16583
tri 14443 16485 14541 16583 sw
tri 14541 16485 14639 16583 ne
rect 14639 16485 14993 16583
tri 14993 16485 15091 16583 sw
tri 15091 16485 15189 16583 ne
rect 15189 16485 15543 16583
tri 15543 16485 15641 16583 sw
tri 15641 16485 15739 16583 ne
rect 15739 16485 16093 16583
tri 16093 16485 16191 16583 sw
tri 16191 16485 16289 16583 ne
rect 16289 16485 16643 16583
tri 16643 16485 16741 16583 sw
tri 16741 16485 16839 16583 ne
rect 16839 16485 17193 16583
tri 17193 16485 17291 16583 sw
tri 17291 16485 17389 16583 ne
rect 17389 16485 17743 16583
tri 17743 16485 17841 16583 sw
tri 17841 16485 17939 16583 ne
rect 17939 16485 18293 16583
tri 18293 16485 18391 16583 sw
tri 18391 16485 18489 16583 ne
rect 18489 16485 18843 16583
tri 18843 16485 18941 16583 sw
tri 18941 16485 19039 16583 ne
rect 19039 16485 19393 16583
tri 19393 16485 19491 16583 sw
tri 19491 16485 19589 16583 ne
rect 19589 16485 20300 16583
rect -2000 16387 241 16485
tri 241 16387 339 16485 sw
tri 339 16387 437 16485 ne
rect 437 16387 791 16485
tri 791 16387 889 16485 sw
tri 889 16387 987 16485 ne
rect 987 16387 1341 16485
tri 1341 16387 1439 16485 sw
tri 1439 16387 1537 16485 ne
rect 1537 16387 1891 16485
tri 1891 16387 1989 16485 sw
tri 1989 16387 2087 16485 ne
rect 2087 16387 2441 16485
tri 2441 16387 2539 16485 sw
tri 2539 16387 2637 16485 ne
rect 2637 16387 2991 16485
tri 2991 16387 3089 16485 sw
tri 3089 16387 3187 16485 ne
rect 3187 16387 3541 16485
tri 3541 16387 3639 16485 sw
tri 3639 16387 3737 16485 ne
rect 3737 16387 4091 16485
tri 4091 16387 4189 16485 sw
tri 4189 16387 4287 16485 ne
rect 4287 16387 4641 16485
tri 4641 16387 4739 16485 sw
tri 4739 16387 4837 16485 ne
rect 4837 16387 5191 16485
tri 5191 16387 5289 16485 sw
tri 5289 16387 5387 16485 ne
rect 5387 16387 5741 16485
tri 5741 16387 5839 16485 sw
tri 5839 16387 5937 16485 ne
rect 5937 16387 6291 16485
tri 6291 16387 6389 16485 sw
tri 6389 16387 6487 16485 ne
rect 6487 16387 6841 16485
tri 6841 16387 6939 16485 sw
tri 6939 16387 7037 16485 ne
rect 7037 16387 7391 16485
tri 7391 16387 7489 16485 sw
tri 7489 16387 7587 16485 ne
rect 7587 16387 7941 16485
tri 7941 16387 8039 16485 sw
tri 8039 16387 8137 16485 ne
rect 8137 16387 8491 16485
tri 8491 16387 8589 16485 sw
tri 8589 16387 8687 16485 ne
rect 8687 16387 9041 16485
tri 9041 16387 9139 16485 sw
tri 9139 16387 9237 16485 ne
rect 9237 16387 9591 16485
tri 9591 16387 9689 16485 sw
tri 9689 16387 9787 16485 ne
rect 9787 16387 10141 16485
tri 10141 16387 10239 16485 sw
tri 10239 16387 10337 16485 ne
rect 10337 16387 10691 16485
tri 10691 16387 10789 16485 sw
tri 10789 16387 10887 16485 ne
rect 10887 16387 11241 16485
tri 11241 16387 11339 16485 sw
tri 11339 16387 11437 16485 ne
rect 11437 16387 11791 16485
tri 11791 16387 11889 16485 sw
tri 11889 16387 11987 16485 ne
rect 11987 16387 12341 16485
tri 12341 16387 12439 16485 sw
tri 12439 16387 12537 16485 ne
rect 12537 16387 12891 16485
tri 12891 16387 12989 16485 sw
tri 12989 16387 13087 16485 ne
rect 13087 16387 13441 16485
tri 13441 16387 13539 16485 sw
tri 13539 16387 13637 16485 ne
rect 13637 16387 13991 16485
tri 13991 16387 14089 16485 sw
tri 14089 16387 14187 16485 ne
rect 14187 16387 14541 16485
tri 14541 16387 14639 16485 sw
tri 14639 16387 14737 16485 ne
rect 14737 16387 15091 16485
tri 15091 16387 15189 16485 sw
tri 15189 16387 15287 16485 ne
rect 15287 16387 15641 16485
tri 15641 16387 15739 16485 sw
tri 15739 16387 15837 16485 ne
rect 15837 16387 16191 16485
tri 16191 16387 16289 16485 sw
tri 16289 16387 16387 16485 ne
rect 16387 16387 16741 16485
tri 16741 16387 16839 16485 sw
tri 16839 16387 16937 16485 ne
rect 16937 16387 17291 16485
tri 17291 16387 17389 16485 sw
tri 17389 16387 17487 16485 ne
rect 17487 16387 17841 16485
tri 17841 16387 17939 16485 sw
tri 17939 16387 18037 16485 ne
rect 18037 16387 18391 16485
tri 18391 16387 18489 16485 sw
tri 18489 16387 18587 16485 ne
rect 18587 16387 18941 16485
tri 18941 16387 19039 16485 sw
tri 19039 16387 19137 16485 ne
rect 19137 16387 19491 16485
tri 19491 16387 19589 16485 sw
tri 19589 16387 19687 16485 ne
rect 19687 16387 20300 16485
rect -2000 16289 339 16387
tri 339 16289 437 16387 sw
tri 437 16289 535 16387 ne
rect 535 16289 889 16387
tri 889 16289 987 16387 sw
tri 987 16289 1085 16387 ne
rect 1085 16289 1439 16387
tri 1439 16289 1537 16387 sw
tri 1537 16289 1635 16387 ne
rect 1635 16289 1989 16387
tri 1989 16289 2087 16387 sw
tri 2087 16289 2185 16387 ne
rect 2185 16289 2539 16387
tri 2539 16289 2637 16387 sw
tri 2637 16289 2735 16387 ne
rect 2735 16289 3089 16387
tri 3089 16289 3187 16387 sw
tri 3187 16289 3285 16387 ne
rect 3285 16289 3639 16387
tri 3639 16289 3737 16387 sw
tri 3737 16289 3835 16387 ne
rect 3835 16289 4189 16387
tri 4189 16289 4287 16387 sw
tri 4287 16289 4385 16387 ne
rect 4385 16289 4739 16387
tri 4739 16289 4837 16387 sw
tri 4837 16289 4935 16387 ne
rect 4935 16289 5289 16387
tri 5289 16289 5387 16387 sw
tri 5387 16289 5485 16387 ne
rect 5485 16289 5839 16387
tri 5839 16289 5937 16387 sw
tri 5937 16289 6035 16387 ne
rect 6035 16289 6389 16387
tri 6389 16289 6487 16387 sw
tri 6487 16289 6585 16387 ne
rect 6585 16289 6939 16387
tri 6939 16289 7037 16387 sw
tri 7037 16289 7135 16387 ne
rect 7135 16289 7489 16387
tri 7489 16289 7587 16387 sw
tri 7587 16289 7685 16387 ne
rect 7685 16289 8039 16387
tri 8039 16289 8137 16387 sw
tri 8137 16289 8235 16387 ne
rect 8235 16289 8589 16387
tri 8589 16289 8687 16387 sw
tri 8687 16289 8785 16387 ne
rect 8785 16289 9139 16387
tri 9139 16289 9237 16387 sw
tri 9237 16289 9335 16387 ne
rect 9335 16289 9689 16387
tri 9689 16289 9787 16387 sw
tri 9787 16289 9885 16387 ne
rect 9885 16289 10239 16387
tri 10239 16289 10337 16387 sw
tri 10337 16289 10435 16387 ne
rect 10435 16289 10789 16387
tri 10789 16289 10887 16387 sw
tri 10887 16289 10985 16387 ne
rect 10985 16289 11339 16387
tri 11339 16289 11437 16387 sw
tri 11437 16289 11535 16387 ne
rect 11535 16289 11889 16387
tri 11889 16289 11987 16387 sw
tri 11987 16289 12085 16387 ne
rect 12085 16289 12439 16387
tri 12439 16289 12537 16387 sw
tri 12537 16289 12635 16387 ne
rect 12635 16289 12989 16387
tri 12989 16289 13087 16387 sw
tri 13087 16289 13185 16387 ne
rect 13185 16289 13539 16387
tri 13539 16289 13637 16387 sw
tri 13637 16289 13735 16387 ne
rect 13735 16289 14089 16387
tri 14089 16289 14187 16387 sw
tri 14187 16289 14285 16387 ne
rect 14285 16289 14639 16387
tri 14639 16289 14737 16387 sw
tri 14737 16289 14835 16387 ne
rect 14835 16289 15189 16387
tri 15189 16289 15287 16387 sw
tri 15287 16289 15385 16387 ne
rect 15385 16289 15739 16387
tri 15739 16289 15837 16387 sw
tri 15837 16289 15935 16387 ne
rect 15935 16289 16289 16387
tri 16289 16289 16387 16387 sw
tri 16387 16289 16485 16387 ne
rect 16485 16289 16839 16387
tri 16839 16289 16937 16387 sw
tri 16937 16289 17035 16387 ne
rect 17035 16289 17389 16387
tri 17389 16289 17487 16387 sw
tri 17487 16289 17585 16387 ne
rect 17585 16289 17939 16387
tri 17939 16289 18037 16387 sw
tri 18037 16289 18135 16387 ne
rect 18135 16289 18489 16387
tri 18489 16289 18587 16387 sw
tri 18587 16289 18685 16387 ne
rect 18685 16289 19039 16387
tri 19039 16289 19137 16387 sw
tri 19137 16289 19235 16387 ne
rect 19235 16289 19589 16387
tri 19589 16289 19687 16387 sw
rect 20800 16289 21800 16937
rect -2000 16285 437 16289
rect -2000 16165 215 16285
rect 335 16191 437 16285
tri 437 16191 535 16289 sw
tri 535 16191 633 16289 ne
rect 633 16285 987 16289
rect 633 16191 765 16285
rect 335 16165 535 16191
rect -2000 16161 535 16165
rect -2000 15513 -1000 16161
tri 113 16063 211 16161 ne
rect 211 16113 535 16161
tri 535 16113 613 16191 sw
tri 633 16113 711 16191 ne
rect 711 16165 765 16191
rect 885 16191 987 16285
tri 987 16191 1085 16289 sw
tri 1085 16191 1183 16289 ne
rect 1183 16285 1537 16289
rect 1183 16191 1315 16285
rect 885 16165 1085 16191
rect 711 16113 1085 16165
tri 1085 16113 1163 16191 sw
tri 1183 16113 1261 16191 ne
rect 1261 16165 1315 16191
rect 1435 16191 1537 16285
tri 1537 16191 1635 16289 sw
tri 1635 16191 1733 16289 ne
rect 1733 16285 2087 16289
rect 1733 16191 1865 16285
rect 1435 16165 1635 16191
rect 1261 16113 1635 16165
tri 1635 16113 1713 16191 sw
tri 1733 16113 1811 16191 ne
rect 1811 16165 1865 16191
rect 1985 16191 2087 16285
tri 2087 16191 2185 16289 sw
tri 2185 16191 2283 16289 ne
rect 2283 16285 2637 16289
rect 2283 16191 2415 16285
rect 1985 16165 2185 16191
rect 1811 16113 2185 16165
tri 2185 16113 2263 16191 sw
tri 2283 16113 2361 16191 ne
rect 2361 16165 2415 16191
rect 2535 16191 2637 16285
tri 2637 16191 2735 16289 sw
tri 2735 16191 2833 16289 ne
rect 2833 16285 3187 16289
rect 2833 16191 2965 16285
rect 2535 16165 2735 16191
rect 2361 16113 2735 16165
tri 2735 16113 2813 16191 sw
tri 2833 16113 2911 16191 ne
rect 2911 16165 2965 16191
rect 3085 16191 3187 16285
tri 3187 16191 3285 16289 sw
tri 3285 16191 3383 16289 ne
rect 3383 16285 3737 16289
rect 3383 16191 3515 16285
rect 3085 16165 3285 16191
rect 2911 16113 3285 16165
tri 3285 16113 3363 16191 sw
tri 3383 16113 3461 16191 ne
rect 3461 16165 3515 16191
rect 3635 16191 3737 16285
tri 3737 16191 3835 16289 sw
tri 3835 16191 3933 16289 ne
rect 3933 16285 4287 16289
rect 3933 16191 4065 16285
rect 3635 16165 3835 16191
rect 3461 16113 3835 16165
tri 3835 16113 3913 16191 sw
tri 3933 16113 4011 16191 ne
rect 4011 16165 4065 16191
rect 4185 16191 4287 16285
tri 4287 16191 4385 16289 sw
tri 4385 16191 4483 16289 ne
rect 4483 16285 4837 16289
rect 4483 16191 4615 16285
rect 4185 16165 4385 16191
rect 4011 16113 4385 16165
tri 4385 16113 4463 16191 sw
tri 4483 16113 4561 16191 ne
rect 4561 16165 4615 16191
rect 4735 16191 4837 16285
tri 4837 16191 4935 16289 sw
tri 4935 16191 5033 16289 ne
rect 5033 16285 5387 16289
rect 5033 16191 5165 16285
rect 4735 16165 4935 16191
rect 4561 16113 4935 16165
tri 4935 16113 5013 16191 sw
tri 5033 16113 5111 16191 ne
rect 5111 16165 5165 16191
rect 5285 16191 5387 16285
tri 5387 16191 5485 16289 sw
tri 5485 16191 5583 16289 ne
rect 5583 16285 5937 16289
rect 5583 16191 5715 16285
rect 5285 16165 5485 16191
rect 5111 16113 5485 16165
tri 5485 16113 5563 16191 sw
tri 5583 16113 5661 16191 ne
rect 5661 16165 5715 16191
rect 5835 16191 5937 16285
tri 5937 16191 6035 16289 sw
tri 6035 16191 6133 16289 ne
rect 6133 16285 6487 16289
rect 6133 16191 6265 16285
rect 5835 16165 6035 16191
rect 5661 16113 6035 16165
tri 6035 16113 6113 16191 sw
tri 6133 16113 6211 16191 ne
rect 6211 16165 6265 16191
rect 6385 16191 6487 16285
tri 6487 16191 6585 16289 sw
tri 6585 16191 6683 16289 ne
rect 6683 16285 7037 16289
rect 6683 16191 6815 16285
rect 6385 16165 6585 16191
rect 6211 16113 6585 16165
tri 6585 16113 6663 16191 sw
tri 6683 16113 6761 16191 ne
rect 6761 16165 6815 16191
rect 6935 16191 7037 16285
tri 7037 16191 7135 16289 sw
tri 7135 16191 7233 16289 ne
rect 7233 16285 7587 16289
rect 7233 16191 7365 16285
rect 6935 16165 7135 16191
rect 6761 16113 7135 16165
tri 7135 16113 7213 16191 sw
tri 7233 16113 7311 16191 ne
rect 7311 16165 7365 16191
rect 7485 16191 7587 16285
tri 7587 16191 7685 16289 sw
tri 7685 16191 7783 16289 ne
rect 7783 16285 8137 16289
rect 7783 16191 7915 16285
rect 7485 16165 7685 16191
rect 7311 16113 7685 16165
tri 7685 16113 7763 16191 sw
tri 7783 16113 7861 16191 ne
rect 7861 16165 7915 16191
rect 8035 16191 8137 16285
tri 8137 16191 8235 16289 sw
tri 8235 16191 8333 16289 ne
rect 8333 16285 8687 16289
rect 8333 16191 8465 16285
rect 8035 16165 8235 16191
rect 7861 16113 8235 16165
tri 8235 16113 8313 16191 sw
tri 8333 16113 8411 16191 ne
rect 8411 16165 8465 16191
rect 8585 16191 8687 16285
tri 8687 16191 8785 16289 sw
tri 8785 16191 8883 16289 ne
rect 8883 16285 9237 16289
rect 8883 16191 9015 16285
rect 8585 16165 8785 16191
rect 8411 16113 8785 16165
tri 8785 16113 8863 16191 sw
tri 8883 16113 8961 16191 ne
rect 8961 16165 9015 16191
rect 9135 16191 9237 16285
tri 9237 16191 9335 16289 sw
tri 9335 16191 9433 16289 ne
rect 9433 16285 9787 16289
rect 9433 16191 9565 16285
rect 9135 16165 9335 16191
rect 8961 16113 9335 16165
tri 9335 16113 9413 16191 sw
tri 9433 16113 9511 16191 ne
rect 9511 16165 9565 16191
rect 9685 16191 9787 16285
tri 9787 16191 9885 16289 sw
tri 9885 16191 9983 16289 ne
rect 9983 16285 10337 16289
rect 9983 16191 10115 16285
rect 9685 16165 9885 16191
rect 9511 16113 9885 16165
tri 9885 16113 9963 16191 sw
tri 9983 16113 10061 16191 ne
rect 10061 16165 10115 16191
rect 10235 16191 10337 16285
tri 10337 16191 10435 16289 sw
tri 10435 16191 10533 16289 ne
rect 10533 16285 10887 16289
rect 10533 16191 10665 16285
rect 10235 16165 10435 16191
rect 10061 16113 10435 16165
tri 10435 16113 10513 16191 sw
tri 10533 16113 10611 16191 ne
rect 10611 16165 10665 16191
rect 10785 16191 10887 16285
tri 10887 16191 10985 16289 sw
tri 10985 16191 11083 16289 ne
rect 11083 16285 11437 16289
rect 11083 16191 11215 16285
rect 10785 16165 10985 16191
rect 10611 16113 10985 16165
tri 10985 16113 11063 16191 sw
tri 11083 16113 11161 16191 ne
rect 11161 16165 11215 16191
rect 11335 16191 11437 16285
tri 11437 16191 11535 16289 sw
tri 11535 16191 11633 16289 ne
rect 11633 16285 11987 16289
rect 11633 16191 11765 16285
rect 11335 16165 11535 16191
rect 11161 16113 11535 16165
tri 11535 16113 11613 16191 sw
tri 11633 16113 11711 16191 ne
rect 11711 16165 11765 16191
rect 11885 16191 11987 16285
tri 11987 16191 12085 16289 sw
tri 12085 16191 12183 16289 ne
rect 12183 16285 12537 16289
rect 12183 16191 12315 16285
rect 11885 16165 12085 16191
rect 11711 16113 12085 16165
tri 12085 16113 12163 16191 sw
tri 12183 16113 12261 16191 ne
rect 12261 16165 12315 16191
rect 12435 16191 12537 16285
tri 12537 16191 12635 16289 sw
tri 12635 16191 12733 16289 ne
rect 12733 16285 13087 16289
rect 12733 16191 12865 16285
rect 12435 16165 12635 16191
rect 12261 16113 12635 16165
tri 12635 16113 12713 16191 sw
tri 12733 16113 12811 16191 ne
rect 12811 16165 12865 16191
rect 12985 16191 13087 16285
tri 13087 16191 13185 16289 sw
tri 13185 16191 13283 16289 ne
rect 13283 16285 13637 16289
rect 13283 16191 13415 16285
rect 12985 16165 13185 16191
rect 12811 16113 13185 16165
tri 13185 16113 13263 16191 sw
tri 13283 16113 13361 16191 ne
rect 13361 16165 13415 16191
rect 13535 16191 13637 16285
tri 13637 16191 13735 16289 sw
tri 13735 16191 13833 16289 ne
rect 13833 16285 14187 16289
rect 13833 16191 13965 16285
rect 13535 16165 13735 16191
rect 13361 16113 13735 16165
tri 13735 16113 13813 16191 sw
tri 13833 16113 13911 16191 ne
rect 13911 16165 13965 16191
rect 14085 16191 14187 16285
tri 14187 16191 14285 16289 sw
tri 14285 16191 14383 16289 ne
rect 14383 16285 14737 16289
rect 14383 16191 14515 16285
rect 14085 16165 14285 16191
rect 13911 16113 14285 16165
tri 14285 16113 14363 16191 sw
tri 14383 16113 14461 16191 ne
rect 14461 16165 14515 16191
rect 14635 16191 14737 16285
tri 14737 16191 14835 16289 sw
tri 14835 16191 14933 16289 ne
rect 14933 16285 15287 16289
rect 14933 16191 15065 16285
rect 14635 16165 14835 16191
rect 14461 16113 14835 16165
tri 14835 16113 14913 16191 sw
tri 14933 16113 15011 16191 ne
rect 15011 16165 15065 16191
rect 15185 16191 15287 16285
tri 15287 16191 15385 16289 sw
tri 15385 16191 15483 16289 ne
rect 15483 16285 15837 16289
rect 15483 16191 15615 16285
rect 15185 16165 15385 16191
rect 15011 16113 15385 16165
tri 15385 16113 15463 16191 sw
tri 15483 16113 15561 16191 ne
rect 15561 16165 15615 16191
rect 15735 16191 15837 16285
tri 15837 16191 15935 16289 sw
tri 15935 16191 16033 16289 ne
rect 16033 16285 16387 16289
rect 16033 16191 16165 16285
rect 15735 16165 15935 16191
rect 15561 16113 15935 16165
tri 15935 16113 16013 16191 sw
tri 16033 16113 16111 16191 ne
rect 16111 16165 16165 16191
rect 16285 16191 16387 16285
tri 16387 16191 16485 16289 sw
tri 16485 16191 16583 16289 ne
rect 16583 16285 16937 16289
rect 16583 16191 16715 16285
rect 16285 16165 16485 16191
rect 16111 16113 16485 16165
tri 16485 16113 16563 16191 sw
tri 16583 16113 16661 16191 ne
rect 16661 16165 16715 16191
rect 16835 16191 16937 16285
tri 16937 16191 17035 16289 sw
tri 17035 16191 17133 16289 ne
rect 17133 16285 17487 16289
rect 17133 16191 17265 16285
rect 16835 16165 17035 16191
rect 16661 16113 17035 16165
tri 17035 16113 17113 16191 sw
tri 17133 16113 17211 16191 ne
rect 17211 16165 17265 16191
rect 17385 16191 17487 16285
tri 17487 16191 17585 16289 sw
tri 17585 16191 17683 16289 ne
rect 17683 16285 18037 16289
rect 17683 16191 17815 16285
rect 17385 16165 17585 16191
rect 17211 16113 17585 16165
tri 17585 16113 17663 16191 sw
tri 17683 16113 17761 16191 ne
rect 17761 16165 17815 16191
rect 17935 16191 18037 16285
tri 18037 16191 18135 16289 sw
tri 18135 16191 18233 16289 ne
rect 18233 16285 18587 16289
rect 18233 16191 18365 16285
rect 17935 16165 18135 16191
rect 17761 16113 18135 16165
tri 18135 16113 18213 16191 sw
tri 18233 16113 18311 16191 ne
rect 18311 16165 18365 16191
rect 18485 16191 18587 16285
tri 18587 16191 18685 16289 sw
tri 18685 16191 18783 16289 ne
rect 18783 16285 19137 16289
rect 18783 16191 18915 16285
rect 18485 16165 18685 16191
rect 18311 16113 18685 16165
tri 18685 16113 18763 16191 sw
tri 18783 16113 18861 16191 ne
rect 18861 16165 18915 16191
rect 19035 16191 19137 16285
tri 19137 16191 19235 16289 sw
tri 19235 16191 19333 16289 ne
rect 19333 16285 21800 16289
rect 19333 16191 19465 16285
rect 19035 16165 19235 16191
rect 18861 16113 19235 16165
tri 19235 16113 19313 16191 sw
tri 19333 16113 19411 16191 ne
rect 19411 16165 19465 16191
rect 19585 16165 21800 16285
rect 19411 16113 21800 16165
rect 211 16063 613 16113
rect -500 16013 113 16063
tri 113 16013 163 16063 sw
tri 211 16013 261 16063 ne
rect 261 16033 613 16063
tri 613 16033 693 16113 sw
tri 711 16033 791 16113 ne
rect 791 16033 1163 16113
tri 1163 16033 1243 16113 sw
tri 1261 16033 1341 16113 ne
rect 1341 16033 1713 16113
tri 1713 16033 1793 16113 sw
tri 1811 16033 1891 16113 ne
rect 1891 16033 2263 16113
tri 2263 16033 2343 16113 sw
tri 2361 16033 2441 16113 ne
rect 2441 16033 2813 16113
tri 2813 16033 2893 16113 sw
tri 2911 16033 2991 16113 ne
rect 2991 16033 3363 16113
tri 3363 16033 3443 16113 sw
tri 3461 16033 3541 16113 ne
rect 3541 16033 3913 16113
tri 3913 16033 3993 16113 sw
tri 4011 16033 4091 16113 ne
rect 4091 16033 4463 16113
tri 4463 16033 4543 16113 sw
tri 4561 16033 4641 16113 ne
rect 4641 16033 5013 16113
tri 5013 16033 5093 16113 sw
tri 5111 16033 5191 16113 ne
rect 5191 16033 5563 16113
tri 5563 16033 5643 16113 sw
tri 5661 16033 5741 16113 ne
rect 5741 16033 6113 16113
tri 6113 16033 6193 16113 sw
tri 6211 16033 6291 16113 ne
rect 6291 16033 6663 16113
tri 6663 16033 6743 16113 sw
tri 6761 16033 6841 16113 ne
rect 6841 16033 7213 16113
tri 7213 16033 7293 16113 sw
tri 7311 16033 7391 16113 ne
rect 7391 16033 7763 16113
tri 7763 16033 7843 16113 sw
tri 7861 16033 7941 16113 ne
rect 7941 16033 8313 16113
tri 8313 16033 8393 16113 sw
tri 8411 16033 8491 16113 ne
rect 8491 16033 8863 16113
tri 8863 16033 8943 16113 sw
tri 8961 16033 9041 16113 ne
rect 9041 16033 9413 16113
tri 9413 16033 9493 16113 sw
tri 9511 16033 9591 16113 ne
rect 9591 16033 9963 16113
tri 9963 16033 10043 16113 sw
tri 10061 16033 10141 16113 ne
rect 10141 16033 10513 16113
tri 10513 16033 10593 16113 sw
tri 10611 16033 10691 16113 ne
rect 10691 16033 11063 16113
tri 11063 16033 11143 16113 sw
tri 11161 16033 11241 16113 ne
rect 11241 16033 11613 16113
tri 11613 16033 11693 16113 sw
tri 11711 16033 11791 16113 ne
rect 11791 16033 12163 16113
tri 12163 16033 12243 16113 sw
tri 12261 16033 12341 16113 ne
rect 12341 16033 12713 16113
tri 12713 16033 12793 16113 sw
tri 12811 16033 12891 16113 ne
rect 12891 16033 13263 16113
tri 13263 16033 13343 16113 sw
tri 13361 16033 13441 16113 ne
rect 13441 16033 13813 16113
tri 13813 16033 13893 16113 sw
tri 13911 16033 13991 16113 ne
rect 13991 16033 14363 16113
tri 14363 16033 14443 16113 sw
tri 14461 16033 14541 16113 ne
rect 14541 16033 14913 16113
tri 14913 16033 14993 16113 sw
tri 15011 16033 15091 16113 ne
rect 15091 16033 15463 16113
tri 15463 16033 15543 16113 sw
tri 15561 16033 15641 16113 ne
rect 15641 16033 16013 16113
tri 16013 16033 16093 16113 sw
tri 16111 16033 16191 16113 ne
rect 16191 16033 16563 16113
tri 16563 16033 16643 16113 sw
tri 16661 16033 16741 16113 ne
rect 16741 16033 17113 16113
tri 17113 16033 17193 16113 sw
tri 17211 16033 17291 16113 ne
rect 17291 16033 17663 16113
tri 17663 16033 17743 16113 sw
tri 17761 16033 17841 16113 ne
rect 17841 16033 18213 16113
tri 18213 16033 18293 16113 sw
tri 18311 16033 18391 16113 ne
rect 18391 16033 18763 16113
tri 18763 16033 18843 16113 sw
tri 18861 16033 18941 16113 ne
rect 18941 16033 19313 16113
tri 19313 16033 19393 16113 sw
tri 19411 16033 19491 16113 ne
rect 19491 16033 20100 16113
rect 261 16013 693 16033
rect -500 15935 163 16013
tri 163 15935 241 16013 sw
tri 261 15935 339 16013 ne
rect 339 15935 693 16013
tri 693 15935 791 16033 sw
tri 791 15935 889 16033 ne
rect 889 15935 1243 16033
tri 1243 15935 1341 16033 sw
tri 1341 15935 1439 16033 ne
rect 1439 15935 1793 16033
tri 1793 15935 1891 16033 sw
tri 1891 15935 1989 16033 ne
rect 1989 15935 2343 16033
tri 2343 15935 2441 16033 sw
tri 2441 15935 2539 16033 ne
rect 2539 15935 2893 16033
tri 2893 15935 2991 16033 sw
tri 2991 15935 3089 16033 ne
rect 3089 15935 3443 16033
tri 3443 15935 3541 16033 sw
tri 3541 15935 3639 16033 ne
rect 3639 15935 3993 16033
tri 3993 15935 4091 16033 sw
tri 4091 15935 4189 16033 ne
rect 4189 15935 4543 16033
tri 4543 15935 4641 16033 sw
tri 4641 15935 4739 16033 ne
rect 4739 15935 5093 16033
tri 5093 15935 5191 16033 sw
tri 5191 15935 5289 16033 ne
rect 5289 15935 5643 16033
tri 5643 15935 5741 16033 sw
tri 5741 15935 5839 16033 ne
rect 5839 15935 6193 16033
tri 6193 15935 6291 16033 sw
tri 6291 15935 6389 16033 ne
rect 6389 15935 6743 16033
tri 6743 15935 6841 16033 sw
tri 6841 15935 6939 16033 ne
rect 6939 15935 7293 16033
tri 7293 15935 7391 16033 sw
tri 7391 15935 7489 16033 ne
rect 7489 15935 7843 16033
tri 7843 15935 7941 16033 sw
tri 7941 15935 8039 16033 ne
rect 8039 15935 8393 16033
tri 8393 15935 8491 16033 sw
tri 8491 15935 8589 16033 ne
rect 8589 15935 8943 16033
tri 8943 15935 9041 16033 sw
tri 9041 15935 9139 16033 ne
rect 9139 15935 9493 16033
tri 9493 15935 9591 16033 sw
tri 9591 15935 9689 16033 ne
rect 9689 15935 10043 16033
tri 10043 15935 10141 16033 sw
tri 10141 15935 10239 16033 ne
rect 10239 15935 10593 16033
tri 10593 15935 10691 16033 sw
tri 10691 15935 10789 16033 ne
rect 10789 15935 11143 16033
tri 11143 15935 11241 16033 sw
tri 11241 15935 11339 16033 ne
rect 11339 15935 11693 16033
tri 11693 15935 11791 16033 sw
tri 11791 15935 11889 16033 ne
rect 11889 15935 12243 16033
tri 12243 15935 12341 16033 sw
tri 12341 15935 12439 16033 ne
rect 12439 15935 12793 16033
tri 12793 15935 12891 16033 sw
tri 12891 15935 12989 16033 ne
rect 12989 15935 13343 16033
tri 13343 15935 13441 16033 sw
tri 13441 15935 13539 16033 ne
rect 13539 15935 13893 16033
tri 13893 15935 13991 16033 sw
tri 13991 15935 14089 16033 ne
rect 14089 15935 14443 16033
tri 14443 15935 14541 16033 sw
tri 14541 15935 14639 16033 ne
rect 14639 15935 14993 16033
tri 14993 15935 15091 16033 sw
tri 15091 15935 15189 16033 ne
rect 15189 15935 15543 16033
tri 15543 15935 15641 16033 sw
tri 15641 15935 15739 16033 ne
rect 15739 15935 16093 16033
tri 16093 15935 16191 16033 sw
tri 16191 15935 16289 16033 ne
rect 16289 15935 16643 16033
tri 16643 15935 16741 16033 sw
tri 16741 15935 16839 16033 ne
rect 16839 15935 17193 16033
tri 17193 15935 17291 16033 sw
tri 17291 15935 17389 16033 ne
rect 17389 15935 17743 16033
tri 17743 15935 17841 16033 sw
tri 17841 15935 17939 16033 ne
rect 17939 15935 18293 16033
tri 18293 15935 18391 16033 sw
tri 18391 15935 18489 16033 ne
rect 18489 15935 18843 16033
tri 18843 15935 18941 16033 sw
tri 18941 15935 19039 16033 ne
rect 19039 15935 19393 16033
tri 19393 15935 19491 16033 sw
tri 19491 15935 19589 16033 ne
rect 19589 16013 20100 16033
rect 20200 16013 21800 16113
rect 19589 15935 21800 16013
rect -500 15887 241 15935
rect -500 15787 -400 15887
rect -300 15837 241 15887
tri 241 15837 339 15935 sw
tri 339 15837 437 15935 ne
rect 437 15837 791 15935
tri 791 15837 889 15935 sw
tri 889 15837 987 15935 ne
rect 987 15837 1341 15935
tri 1341 15837 1439 15935 sw
tri 1439 15837 1537 15935 ne
rect 1537 15837 1891 15935
tri 1891 15837 1989 15935 sw
tri 1989 15837 2087 15935 ne
rect 2087 15837 2441 15935
tri 2441 15837 2539 15935 sw
tri 2539 15837 2637 15935 ne
rect 2637 15837 2991 15935
tri 2991 15837 3089 15935 sw
tri 3089 15837 3187 15935 ne
rect 3187 15837 3541 15935
tri 3541 15837 3639 15935 sw
tri 3639 15837 3737 15935 ne
rect 3737 15837 4091 15935
tri 4091 15837 4189 15935 sw
tri 4189 15837 4287 15935 ne
rect 4287 15837 4641 15935
tri 4641 15837 4739 15935 sw
tri 4739 15837 4837 15935 ne
rect 4837 15837 5191 15935
tri 5191 15837 5289 15935 sw
tri 5289 15837 5387 15935 ne
rect 5387 15837 5741 15935
tri 5741 15837 5839 15935 sw
tri 5839 15837 5937 15935 ne
rect 5937 15837 6291 15935
tri 6291 15837 6389 15935 sw
tri 6389 15837 6487 15935 ne
rect 6487 15837 6841 15935
tri 6841 15837 6939 15935 sw
tri 6939 15837 7037 15935 ne
rect 7037 15837 7391 15935
tri 7391 15837 7489 15935 sw
tri 7489 15837 7587 15935 ne
rect 7587 15837 7941 15935
tri 7941 15837 8039 15935 sw
tri 8039 15837 8137 15935 ne
rect 8137 15837 8491 15935
tri 8491 15837 8589 15935 sw
tri 8589 15837 8687 15935 ne
rect 8687 15837 9041 15935
tri 9041 15837 9139 15935 sw
tri 9139 15837 9237 15935 ne
rect 9237 15837 9591 15935
tri 9591 15837 9689 15935 sw
tri 9689 15837 9787 15935 ne
rect 9787 15837 10141 15935
tri 10141 15837 10239 15935 sw
tri 10239 15837 10337 15935 ne
rect 10337 15837 10691 15935
tri 10691 15837 10789 15935 sw
tri 10789 15837 10887 15935 ne
rect 10887 15837 11241 15935
tri 11241 15837 11339 15935 sw
tri 11339 15837 11437 15935 ne
rect 11437 15837 11791 15935
tri 11791 15837 11889 15935 sw
tri 11889 15837 11987 15935 ne
rect 11987 15837 12341 15935
tri 12341 15837 12439 15935 sw
tri 12439 15837 12537 15935 ne
rect 12537 15837 12891 15935
tri 12891 15837 12989 15935 sw
tri 12989 15837 13087 15935 ne
rect 13087 15837 13441 15935
tri 13441 15837 13539 15935 sw
tri 13539 15837 13637 15935 ne
rect 13637 15837 13991 15935
tri 13991 15837 14089 15935 sw
tri 14089 15837 14187 15935 ne
rect 14187 15837 14541 15935
tri 14541 15837 14639 15935 sw
tri 14639 15837 14737 15935 ne
rect 14737 15837 15091 15935
tri 15091 15837 15189 15935 sw
tri 15189 15837 15287 15935 ne
rect 15287 15837 15641 15935
tri 15641 15837 15739 15935 sw
tri 15739 15837 15837 15935 ne
rect 15837 15837 16191 15935
tri 16191 15837 16289 15935 sw
tri 16289 15837 16387 15935 ne
rect 16387 15837 16741 15935
tri 16741 15837 16839 15935 sw
tri 16839 15837 16937 15935 ne
rect 16937 15837 17291 15935
tri 17291 15837 17389 15935 sw
tri 17389 15837 17487 15935 ne
rect 17487 15837 17841 15935
tri 17841 15837 17939 15935 sw
tri 17939 15837 18037 15935 ne
rect 18037 15837 18391 15935
tri 18391 15837 18489 15935 sw
tri 18489 15837 18587 15935 ne
rect 18587 15837 18941 15935
tri 18941 15837 19039 15935 sw
tri 19039 15837 19137 15935 ne
rect 19137 15837 19491 15935
tri 19491 15837 19589 15935 sw
tri 19589 15837 19687 15935 ne
rect 19687 15837 21800 15935
rect -300 15787 339 15837
rect -500 15739 339 15787
tri 339 15739 437 15837 sw
tri 437 15739 535 15837 ne
rect 535 15739 889 15837
tri 889 15739 987 15837 sw
tri 987 15739 1085 15837 ne
rect 1085 15739 1439 15837
tri 1439 15739 1537 15837 sw
tri 1537 15739 1635 15837 ne
rect 1635 15739 1989 15837
tri 1989 15739 2087 15837 sw
tri 2087 15739 2185 15837 ne
rect 2185 15739 2539 15837
tri 2539 15739 2637 15837 sw
tri 2637 15739 2735 15837 ne
rect 2735 15739 3089 15837
tri 3089 15739 3187 15837 sw
tri 3187 15739 3285 15837 ne
rect 3285 15739 3639 15837
tri 3639 15739 3737 15837 sw
tri 3737 15739 3835 15837 ne
rect 3835 15739 4189 15837
tri 4189 15739 4287 15837 sw
tri 4287 15739 4385 15837 ne
rect 4385 15739 4739 15837
tri 4739 15739 4837 15837 sw
tri 4837 15739 4935 15837 ne
rect 4935 15739 5289 15837
tri 5289 15739 5387 15837 sw
tri 5387 15739 5485 15837 ne
rect 5485 15739 5839 15837
tri 5839 15739 5937 15837 sw
tri 5937 15739 6035 15837 ne
rect 6035 15739 6389 15837
tri 6389 15739 6487 15837 sw
tri 6487 15739 6585 15837 ne
rect 6585 15739 6939 15837
tri 6939 15739 7037 15837 sw
tri 7037 15739 7135 15837 ne
rect 7135 15739 7489 15837
tri 7489 15739 7587 15837 sw
tri 7587 15739 7685 15837 ne
rect 7685 15739 8039 15837
tri 8039 15739 8137 15837 sw
tri 8137 15739 8235 15837 ne
rect 8235 15739 8589 15837
tri 8589 15739 8687 15837 sw
tri 8687 15739 8785 15837 ne
rect 8785 15739 9139 15837
tri 9139 15739 9237 15837 sw
tri 9237 15739 9335 15837 ne
rect 9335 15739 9689 15837
tri 9689 15739 9787 15837 sw
tri 9787 15739 9885 15837 ne
rect 9885 15739 10239 15837
tri 10239 15739 10337 15837 sw
tri 10337 15739 10435 15837 ne
rect 10435 15739 10789 15837
tri 10789 15739 10887 15837 sw
tri 10887 15739 10985 15837 ne
rect 10985 15739 11339 15837
tri 11339 15739 11437 15837 sw
tri 11437 15739 11535 15837 ne
rect 11535 15739 11889 15837
tri 11889 15739 11987 15837 sw
tri 11987 15739 12085 15837 ne
rect 12085 15739 12439 15837
tri 12439 15739 12537 15837 sw
tri 12537 15739 12635 15837 ne
rect 12635 15739 12989 15837
tri 12989 15739 13087 15837 sw
tri 13087 15739 13185 15837 ne
rect 13185 15739 13539 15837
tri 13539 15739 13637 15837 sw
tri 13637 15739 13735 15837 ne
rect 13735 15739 14089 15837
tri 14089 15739 14187 15837 sw
tri 14187 15739 14285 15837 ne
rect 14285 15739 14639 15837
tri 14639 15739 14737 15837 sw
tri 14737 15739 14835 15837 ne
rect 14835 15739 15189 15837
tri 15189 15739 15287 15837 sw
tri 15287 15739 15385 15837 ne
rect 15385 15739 15739 15837
tri 15739 15739 15837 15837 sw
tri 15837 15739 15935 15837 ne
rect 15935 15739 16289 15837
tri 16289 15739 16387 15837 sw
tri 16387 15739 16485 15837 ne
rect 16485 15739 16839 15837
tri 16839 15739 16937 15837 sw
tri 16937 15739 17035 15837 ne
rect 17035 15739 17389 15837
tri 17389 15739 17487 15837 sw
tri 17487 15739 17585 15837 ne
rect 17585 15739 17939 15837
tri 17939 15739 18037 15837 sw
tri 18037 15739 18135 15837 ne
rect 18135 15739 18489 15837
tri 18489 15739 18587 15837 sw
tri 18587 15739 18685 15837 ne
rect 18685 15739 19039 15837
tri 19039 15739 19137 15837 sw
tri 19137 15739 19235 15837 ne
rect 19235 15739 19589 15837
tri 19589 15739 19687 15837 sw
rect -500 15735 437 15739
rect -500 15615 215 15735
rect 335 15641 437 15735
tri 437 15641 535 15739 sw
tri 535 15641 633 15739 ne
rect 633 15735 987 15739
rect 633 15641 765 15735
rect 335 15615 535 15641
rect -500 15611 535 15615
tri 535 15611 565 15641 sw
tri 633 15611 663 15641 ne
rect 663 15615 765 15641
rect 885 15641 987 15735
tri 987 15641 1085 15739 sw
tri 1085 15641 1183 15739 ne
rect 1183 15735 1537 15739
rect 1183 15641 1315 15735
rect 885 15615 1085 15641
rect 663 15611 1085 15615
tri 1085 15611 1115 15641 sw
tri 1183 15611 1213 15641 ne
rect 1213 15615 1315 15641
rect 1435 15641 1537 15735
tri 1537 15641 1635 15739 sw
tri 1635 15641 1733 15739 ne
rect 1733 15735 2087 15739
rect 1733 15641 1865 15735
rect 1435 15615 1635 15641
rect 1213 15611 1635 15615
tri 1635 15611 1665 15641 sw
tri 1733 15611 1763 15641 ne
rect 1763 15615 1865 15641
rect 1985 15641 2087 15735
tri 2087 15641 2185 15739 sw
tri 2185 15641 2283 15739 ne
rect 2283 15735 2637 15739
rect 2283 15641 2415 15735
rect 1985 15615 2185 15641
rect 1763 15611 2185 15615
tri 2185 15611 2215 15641 sw
tri 2283 15611 2313 15641 ne
rect 2313 15615 2415 15641
rect 2535 15641 2637 15735
tri 2637 15641 2735 15739 sw
tri 2735 15641 2833 15739 ne
rect 2833 15735 3187 15739
rect 2833 15641 2965 15735
rect 2535 15615 2735 15641
rect 2313 15611 2735 15615
tri 2735 15611 2765 15641 sw
tri 2833 15611 2863 15641 ne
rect 2863 15615 2965 15641
rect 3085 15641 3187 15735
tri 3187 15641 3285 15739 sw
tri 3285 15641 3383 15739 ne
rect 3383 15735 3737 15739
rect 3383 15641 3515 15735
rect 3085 15615 3285 15641
rect 2863 15611 3285 15615
tri 3285 15611 3315 15641 sw
tri 3383 15611 3413 15641 ne
rect 3413 15615 3515 15641
rect 3635 15641 3737 15735
tri 3737 15641 3835 15739 sw
tri 3835 15641 3933 15739 ne
rect 3933 15735 4287 15739
rect 3933 15641 4065 15735
rect 3635 15615 3835 15641
rect 3413 15611 3835 15615
tri 3835 15611 3865 15641 sw
tri 3933 15611 3963 15641 ne
rect 3963 15615 4065 15641
rect 4185 15641 4287 15735
tri 4287 15641 4385 15739 sw
tri 4385 15641 4483 15739 ne
rect 4483 15735 4837 15739
rect 4483 15641 4615 15735
rect 4185 15615 4385 15641
rect 3963 15611 4385 15615
tri 4385 15611 4415 15641 sw
tri 4483 15611 4513 15641 ne
rect 4513 15615 4615 15641
rect 4735 15641 4837 15735
tri 4837 15641 4935 15739 sw
tri 4935 15641 5033 15739 ne
rect 5033 15735 5387 15739
rect 5033 15641 5165 15735
rect 4735 15615 4935 15641
rect 4513 15611 4935 15615
tri 4935 15611 4965 15641 sw
tri 5033 15611 5063 15641 ne
rect 5063 15615 5165 15641
rect 5285 15641 5387 15735
tri 5387 15641 5485 15739 sw
tri 5485 15641 5583 15739 ne
rect 5583 15735 5937 15739
rect 5583 15641 5715 15735
rect 5285 15615 5485 15641
rect 5063 15611 5485 15615
tri 5485 15611 5515 15641 sw
tri 5583 15611 5613 15641 ne
rect 5613 15615 5715 15641
rect 5835 15641 5937 15735
tri 5937 15641 6035 15739 sw
tri 6035 15641 6133 15739 ne
rect 6133 15735 6487 15739
rect 6133 15641 6265 15735
rect 5835 15615 6035 15641
rect 5613 15611 6035 15615
tri 6035 15611 6065 15641 sw
tri 6133 15611 6163 15641 ne
rect 6163 15615 6265 15641
rect 6385 15641 6487 15735
tri 6487 15641 6585 15739 sw
tri 6585 15641 6683 15739 ne
rect 6683 15735 7037 15739
rect 6683 15641 6815 15735
rect 6385 15615 6585 15641
rect 6163 15611 6585 15615
tri 6585 15611 6615 15641 sw
tri 6683 15611 6713 15641 ne
rect 6713 15615 6815 15641
rect 6935 15641 7037 15735
tri 7037 15641 7135 15739 sw
tri 7135 15641 7233 15739 ne
rect 7233 15735 7587 15739
rect 7233 15641 7365 15735
rect 6935 15615 7135 15641
rect 6713 15611 7135 15615
tri 7135 15611 7165 15641 sw
tri 7233 15611 7263 15641 ne
rect 7263 15615 7365 15641
rect 7485 15641 7587 15735
tri 7587 15641 7685 15739 sw
tri 7685 15641 7783 15739 ne
rect 7783 15735 8137 15739
rect 7783 15641 7915 15735
rect 7485 15615 7685 15641
rect 7263 15611 7685 15615
tri 7685 15611 7715 15641 sw
tri 7783 15611 7813 15641 ne
rect 7813 15615 7915 15641
rect 8035 15641 8137 15735
tri 8137 15641 8235 15739 sw
tri 8235 15641 8333 15739 ne
rect 8333 15735 8687 15739
rect 8333 15641 8465 15735
rect 8035 15615 8235 15641
rect 7813 15611 8235 15615
tri 8235 15611 8265 15641 sw
tri 8333 15611 8363 15641 ne
rect 8363 15615 8465 15641
rect 8585 15641 8687 15735
tri 8687 15641 8785 15739 sw
tri 8785 15641 8883 15739 ne
rect 8883 15735 9237 15739
rect 8883 15641 9015 15735
rect 8585 15615 8785 15641
rect 8363 15611 8785 15615
tri 8785 15611 8815 15641 sw
tri 8883 15611 8913 15641 ne
rect 8913 15615 9015 15641
rect 9135 15641 9237 15735
tri 9237 15641 9335 15739 sw
tri 9335 15641 9433 15739 ne
rect 9433 15735 9787 15739
rect 9433 15641 9565 15735
rect 9135 15615 9335 15641
rect 8913 15611 9335 15615
tri 9335 15611 9365 15641 sw
tri 9433 15611 9463 15641 ne
rect 9463 15615 9565 15641
rect 9685 15641 9787 15735
tri 9787 15641 9885 15739 sw
tri 9885 15641 9983 15739 ne
rect 9983 15735 10337 15739
rect 9983 15641 10115 15735
rect 9685 15615 9885 15641
rect 9463 15611 9885 15615
tri 9885 15611 9915 15641 sw
tri 9983 15611 10013 15641 ne
rect 10013 15615 10115 15641
rect 10235 15641 10337 15735
tri 10337 15641 10435 15739 sw
tri 10435 15641 10533 15739 ne
rect 10533 15735 10887 15739
rect 10533 15641 10665 15735
rect 10235 15615 10435 15641
rect 10013 15611 10435 15615
tri 10435 15611 10465 15641 sw
tri 10533 15611 10563 15641 ne
rect 10563 15615 10665 15641
rect 10785 15641 10887 15735
tri 10887 15641 10985 15739 sw
tri 10985 15641 11083 15739 ne
rect 11083 15735 11437 15739
rect 11083 15641 11215 15735
rect 10785 15615 10985 15641
rect 10563 15611 10985 15615
tri 10985 15611 11015 15641 sw
tri 11083 15611 11113 15641 ne
rect 11113 15615 11215 15641
rect 11335 15641 11437 15735
tri 11437 15641 11535 15739 sw
tri 11535 15641 11633 15739 ne
rect 11633 15735 11987 15739
rect 11633 15641 11765 15735
rect 11335 15615 11535 15641
rect 11113 15611 11535 15615
tri 11535 15611 11565 15641 sw
tri 11633 15611 11663 15641 ne
rect 11663 15615 11765 15641
rect 11885 15641 11987 15735
tri 11987 15641 12085 15739 sw
tri 12085 15641 12183 15739 ne
rect 12183 15735 12537 15739
rect 12183 15641 12315 15735
rect 11885 15615 12085 15641
rect 11663 15611 12085 15615
tri 12085 15611 12115 15641 sw
tri 12183 15611 12213 15641 ne
rect 12213 15615 12315 15641
rect 12435 15641 12537 15735
tri 12537 15641 12635 15739 sw
tri 12635 15641 12733 15739 ne
rect 12733 15735 13087 15739
rect 12733 15641 12865 15735
rect 12435 15615 12635 15641
rect 12213 15611 12635 15615
tri 12635 15611 12665 15641 sw
tri 12733 15611 12763 15641 ne
rect 12763 15615 12865 15641
rect 12985 15641 13087 15735
tri 13087 15641 13185 15739 sw
tri 13185 15641 13283 15739 ne
rect 13283 15735 13637 15739
rect 13283 15641 13415 15735
rect 12985 15615 13185 15641
rect 12763 15611 13185 15615
tri 13185 15611 13215 15641 sw
tri 13283 15611 13313 15641 ne
rect 13313 15615 13415 15641
rect 13535 15641 13637 15735
tri 13637 15641 13735 15739 sw
tri 13735 15641 13833 15739 ne
rect 13833 15735 14187 15739
rect 13833 15641 13965 15735
rect 13535 15615 13735 15641
rect 13313 15611 13735 15615
tri 13735 15611 13765 15641 sw
tri 13833 15611 13863 15641 ne
rect 13863 15615 13965 15641
rect 14085 15641 14187 15735
tri 14187 15641 14285 15739 sw
tri 14285 15641 14383 15739 ne
rect 14383 15735 14737 15739
rect 14383 15641 14515 15735
rect 14085 15615 14285 15641
rect 13863 15611 14285 15615
tri 14285 15611 14315 15641 sw
tri 14383 15611 14413 15641 ne
rect 14413 15615 14515 15641
rect 14635 15641 14737 15735
tri 14737 15641 14835 15739 sw
tri 14835 15641 14933 15739 ne
rect 14933 15735 15287 15739
rect 14933 15641 15065 15735
rect 14635 15615 14835 15641
rect 14413 15611 14835 15615
tri 14835 15611 14865 15641 sw
tri 14933 15611 14963 15641 ne
rect 14963 15615 15065 15641
rect 15185 15641 15287 15735
tri 15287 15641 15385 15739 sw
tri 15385 15641 15483 15739 ne
rect 15483 15735 15837 15739
rect 15483 15641 15615 15735
rect 15185 15615 15385 15641
rect 14963 15611 15385 15615
tri 15385 15611 15415 15641 sw
tri 15483 15611 15513 15641 ne
rect 15513 15615 15615 15641
rect 15735 15641 15837 15735
tri 15837 15641 15935 15739 sw
tri 15935 15641 16033 15739 ne
rect 16033 15735 16387 15739
rect 16033 15641 16165 15735
rect 15735 15615 15935 15641
rect 15513 15611 15935 15615
tri 15935 15611 15965 15641 sw
tri 16033 15611 16063 15641 ne
rect 16063 15615 16165 15641
rect 16285 15641 16387 15735
tri 16387 15641 16485 15739 sw
tri 16485 15641 16583 15739 ne
rect 16583 15735 16937 15739
rect 16583 15641 16715 15735
rect 16285 15615 16485 15641
rect 16063 15611 16485 15615
tri 16485 15611 16515 15641 sw
tri 16583 15611 16613 15641 ne
rect 16613 15615 16715 15641
rect 16835 15641 16937 15735
tri 16937 15641 17035 15739 sw
tri 17035 15641 17133 15739 ne
rect 17133 15735 17487 15739
rect 17133 15641 17265 15735
rect 16835 15615 17035 15641
rect 16613 15611 17035 15615
tri 17035 15611 17065 15641 sw
tri 17133 15611 17163 15641 ne
rect 17163 15615 17265 15641
rect 17385 15641 17487 15735
tri 17487 15641 17585 15739 sw
tri 17585 15641 17683 15739 ne
rect 17683 15735 18037 15739
rect 17683 15641 17815 15735
rect 17385 15615 17585 15641
rect 17163 15611 17585 15615
tri 17585 15611 17615 15641 sw
tri 17683 15611 17713 15641 ne
rect 17713 15615 17815 15641
rect 17935 15641 18037 15735
tri 18037 15641 18135 15739 sw
tri 18135 15641 18233 15739 ne
rect 18233 15735 18587 15739
rect 18233 15641 18365 15735
rect 17935 15615 18135 15641
rect 17713 15611 18135 15615
tri 18135 15611 18165 15641 sw
tri 18233 15611 18263 15641 ne
rect 18263 15615 18365 15641
rect 18485 15641 18587 15735
tri 18587 15641 18685 15739 sw
tri 18685 15641 18783 15739 ne
rect 18783 15735 19137 15739
rect 18783 15641 18915 15735
rect 18485 15615 18685 15641
rect 18263 15611 18685 15615
tri 18685 15611 18715 15641 sw
tri 18783 15611 18813 15641 ne
rect 18813 15615 18915 15641
rect 19035 15641 19137 15735
tri 19137 15641 19235 15739 sw
tri 19235 15641 19333 15739 ne
rect 19333 15735 20300 15739
rect 19333 15641 19465 15735
rect 19035 15615 19235 15641
rect 18813 15611 19235 15615
tri 19235 15611 19265 15641 sw
tri 19333 15611 19363 15641 ne
rect 19363 15615 19465 15641
rect 19585 15615 20300 15735
rect 19363 15611 20300 15615
tri 113 15513 211 15611 ne
rect 211 15513 565 15611
tri 565 15513 663 15611 sw
tri 663 15513 761 15611 ne
rect 761 15513 1115 15611
tri 1115 15513 1213 15611 sw
tri 1213 15513 1311 15611 ne
rect 1311 15513 1665 15611
tri 1665 15513 1763 15611 sw
tri 1763 15513 1861 15611 ne
rect 1861 15513 2215 15611
tri 2215 15513 2313 15611 sw
tri 2313 15513 2411 15611 ne
rect 2411 15513 2765 15611
tri 2765 15513 2863 15611 sw
tri 2863 15513 2961 15611 ne
rect 2961 15513 3315 15611
tri 3315 15513 3413 15611 sw
tri 3413 15513 3511 15611 ne
rect 3511 15513 3865 15611
tri 3865 15513 3963 15611 sw
tri 3963 15513 4061 15611 ne
rect 4061 15513 4415 15611
tri 4415 15513 4513 15611 sw
tri 4513 15513 4611 15611 ne
rect 4611 15513 4965 15611
tri 4965 15513 5063 15611 sw
tri 5063 15513 5161 15611 ne
rect 5161 15513 5515 15611
tri 5515 15513 5613 15611 sw
tri 5613 15513 5711 15611 ne
rect 5711 15513 6065 15611
tri 6065 15513 6163 15611 sw
tri 6163 15513 6261 15611 ne
rect 6261 15513 6615 15611
tri 6615 15513 6713 15611 sw
tri 6713 15513 6811 15611 ne
rect 6811 15513 7165 15611
tri 7165 15513 7263 15611 sw
tri 7263 15513 7361 15611 ne
rect 7361 15513 7715 15611
tri 7715 15513 7813 15611 sw
tri 7813 15513 7911 15611 ne
rect 7911 15513 8265 15611
tri 8265 15513 8363 15611 sw
tri 8363 15513 8461 15611 ne
rect 8461 15513 8815 15611
tri 8815 15513 8913 15611 sw
tri 8913 15513 9011 15611 ne
rect 9011 15513 9365 15611
tri 9365 15513 9463 15611 sw
tri 9463 15513 9561 15611 ne
rect 9561 15513 9915 15611
tri 9915 15513 10013 15611 sw
tri 10013 15513 10111 15611 ne
rect 10111 15513 10465 15611
tri 10465 15513 10563 15611 sw
tri 10563 15513 10661 15611 ne
rect 10661 15513 11015 15611
tri 11015 15513 11113 15611 sw
tri 11113 15513 11211 15611 ne
rect 11211 15513 11565 15611
tri 11565 15513 11663 15611 sw
tri 11663 15513 11761 15611 ne
rect 11761 15513 12115 15611
tri 12115 15513 12213 15611 sw
tri 12213 15513 12311 15611 ne
rect 12311 15513 12665 15611
tri 12665 15513 12763 15611 sw
tri 12763 15513 12861 15611 ne
rect 12861 15513 13215 15611
tri 13215 15513 13313 15611 sw
tri 13313 15513 13411 15611 ne
rect 13411 15513 13765 15611
tri 13765 15513 13863 15611 sw
tri 13863 15513 13961 15611 ne
rect 13961 15513 14315 15611
tri 14315 15513 14413 15611 sw
tri 14413 15513 14511 15611 ne
rect 14511 15513 14865 15611
tri 14865 15513 14963 15611 sw
tri 14963 15513 15061 15611 ne
rect 15061 15513 15415 15611
tri 15415 15513 15513 15611 sw
tri 15513 15513 15611 15611 ne
rect 15611 15513 15965 15611
tri 15965 15513 16063 15611 sw
tri 16063 15513 16161 15611 ne
rect 16161 15513 16515 15611
tri 16515 15513 16613 15611 sw
tri 16613 15513 16711 15611 ne
rect 16711 15513 17065 15611
tri 17065 15513 17163 15611 sw
tri 17163 15513 17261 15611 ne
rect 17261 15513 17615 15611
tri 17615 15513 17713 15611 sw
tri 17713 15513 17811 15611 ne
rect 17811 15513 18165 15611
tri 18165 15513 18263 15611 sw
tri 18263 15513 18361 15611 ne
rect 18361 15513 18715 15611
tri 18715 15513 18813 15611 sw
tri 18813 15513 18911 15611 ne
rect 18911 15513 19265 15611
tri 19265 15513 19363 15611 sw
tri 19363 15513 19461 15611 ne
rect 19461 15513 20300 15611
rect -2000 15483 113 15513
tri 113 15483 143 15513 sw
tri 211 15483 241 15513 ne
rect 241 15483 663 15513
tri 663 15483 693 15513 sw
tri 761 15483 791 15513 ne
rect 791 15483 1213 15513
tri 1213 15483 1243 15513 sw
tri 1311 15483 1341 15513 ne
rect 1341 15483 1763 15513
tri 1763 15483 1793 15513 sw
tri 1861 15483 1891 15513 ne
rect 1891 15483 2313 15513
tri 2313 15483 2343 15513 sw
tri 2411 15483 2441 15513 ne
rect 2441 15483 2863 15513
tri 2863 15483 2893 15513 sw
tri 2961 15483 2991 15513 ne
rect 2991 15483 3413 15513
tri 3413 15483 3443 15513 sw
tri 3511 15483 3541 15513 ne
rect 3541 15483 3963 15513
tri 3963 15483 3993 15513 sw
tri 4061 15483 4091 15513 ne
rect 4091 15483 4513 15513
tri 4513 15483 4543 15513 sw
tri 4611 15483 4641 15513 ne
rect 4641 15483 5063 15513
tri 5063 15483 5093 15513 sw
tri 5161 15483 5191 15513 ne
rect 5191 15483 5613 15513
tri 5613 15483 5643 15513 sw
tri 5711 15483 5741 15513 ne
rect 5741 15483 6163 15513
tri 6163 15483 6193 15513 sw
tri 6261 15483 6291 15513 ne
rect 6291 15483 6713 15513
tri 6713 15483 6743 15513 sw
tri 6811 15483 6841 15513 ne
rect 6841 15483 7263 15513
tri 7263 15483 7293 15513 sw
tri 7361 15483 7391 15513 ne
rect 7391 15483 7813 15513
tri 7813 15483 7843 15513 sw
tri 7911 15483 7941 15513 ne
rect 7941 15483 8363 15513
tri 8363 15483 8393 15513 sw
tri 8461 15483 8491 15513 ne
rect 8491 15483 8913 15513
tri 8913 15483 8943 15513 sw
tri 9011 15483 9041 15513 ne
rect 9041 15483 9463 15513
tri 9463 15483 9493 15513 sw
tri 9561 15483 9591 15513 ne
rect 9591 15483 10013 15513
tri 10013 15483 10043 15513 sw
tri 10111 15483 10141 15513 ne
rect 10141 15483 10563 15513
tri 10563 15483 10593 15513 sw
tri 10661 15483 10691 15513 ne
rect 10691 15483 11113 15513
tri 11113 15483 11143 15513 sw
tri 11211 15483 11241 15513 ne
rect 11241 15483 11663 15513
tri 11663 15483 11693 15513 sw
tri 11761 15483 11791 15513 ne
rect 11791 15483 12213 15513
tri 12213 15483 12243 15513 sw
tri 12311 15483 12341 15513 ne
rect 12341 15483 12763 15513
tri 12763 15483 12793 15513 sw
tri 12861 15483 12891 15513 ne
rect 12891 15483 13313 15513
tri 13313 15483 13343 15513 sw
tri 13411 15483 13441 15513 ne
rect 13441 15483 13863 15513
tri 13863 15483 13893 15513 sw
tri 13961 15483 13991 15513 ne
rect 13991 15483 14413 15513
tri 14413 15483 14443 15513 sw
tri 14511 15483 14541 15513 ne
rect 14541 15483 14963 15513
tri 14963 15483 14993 15513 sw
tri 15061 15483 15091 15513 ne
rect 15091 15483 15513 15513
tri 15513 15483 15543 15513 sw
tri 15611 15483 15641 15513 ne
rect 15641 15483 16063 15513
tri 16063 15483 16093 15513 sw
tri 16161 15483 16191 15513 ne
rect 16191 15483 16613 15513
tri 16613 15483 16643 15513 sw
tri 16711 15483 16741 15513 ne
rect 16741 15483 17163 15513
tri 17163 15483 17193 15513 sw
tri 17261 15483 17291 15513 ne
rect 17291 15483 17713 15513
tri 17713 15483 17743 15513 sw
tri 17811 15483 17841 15513 ne
rect 17841 15483 18263 15513
tri 18263 15483 18293 15513 sw
tri 18361 15483 18391 15513 ne
rect 18391 15483 18813 15513
tri 18813 15483 18843 15513 sw
tri 18911 15483 18941 15513 ne
rect 18941 15483 19363 15513
tri 19363 15483 19393 15513 sw
tri 19461 15483 19491 15513 ne
rect 19491 15483 20300 15513
rect -2000 15385 143 15483
tri 143 15385 241 15483 sw
tri 241 15385 339 15483 ne
rect 339 15385 693 15483
tri 693 15385 791 15483 sw
tri 791 15385 889 15483 ne
rect 889 15385 1243 15483
tri 1243 15385 1341 15483 sw
tri 1341 15385 1439 15483 ne
rect 1439 15385 1793 15483
tri 1793 15385 1891 15483 sw
tri 1891 15385 1989 15483 ne
rect 1989 15385 2343 15483
tri 2343 15385 2441 15483 sw
tri 2441 15385 2539 15483 ne
rect 2539 15385 2893 15483
tri 2893 15385 2991 15483 sw
tri 2991 15385 3089 15483 ne
rect 3089 15385 3443 15483
tri 3443 15385 3541 15483 sw
tri 3541 15385 3639 15483 ne
rect 3639 15385 3993 15483
tri 3993 15385 4091 15483 sw
tri 4091 15385 4189 15483 ne
rect 4189 15385 4543 15483
tri 4543 15385 4641 15483 sw
tri 4641 15385 4739 15483 ne
rect 4739 15385 5093 15483
tri 5093 15385 5191 15483 sw
tri 5191 15385 5289 15483 ne
rect 5289 15385 5643 15483
tri 5643 15385 5741 15483 sw
tri 5741 15385 5839 15483 ne
rect 5839 15385 6193 15483
tri 6193 15385 6291 15483 sw
tri 6291 15385 6389 15483 ne
rect 6389 15385 6743 15483
tri 6743 15385 6841 15483 sw
tri 6841 15385 6939 15483 ne
rect 6939 15385 7293 15483
tri 7293 15385 7391 15483 sw
tri 7391 15385 7489 15483 ne
rect 7489 15385 7843 15483
tri 7843 15385 7941 15483 sw
tri 7941 15385 8039 15483 ne
rect 8039 15385 8393 15483
tri 8393 15385 8491 15483 sw
tri 8491 15385 8589 15483 ne
rect 8589 15385 8943 15483
tri 8943 15385 9041 15483 sw
tri 9041 15385 9139 15483 ne
rect 9139 15385 9493 15483
tri 9493 15385 9591 15483 sw
tri 9591 15385 9689 15483 ne
rect 9689 15385 10043 15483
tri 10043 15385 10141 15483 sw
tri 10141 15385 10239 15483 ne
rect 10239 15385 10593 15483
tri 10593 15385 10691 15483 sw
tri 10691 15385 10789 15483 ne
rect 10789 15385 11143 15483
tri 11143 15385 11241 15483 sw
tri 11241 15385 11339 15483 ne
rect 11339 15385 11693 15483
tri 11693 15385 11791 15483 sw
tri 11791 15385 11889 15483 ne
rect 11889 15385 12243 15483
tri 12243 15385 12341 15483 sw
tri 12341 15385 12439 15483 ne
rect 12439 15385 12793 15483
tri 12793 15385 12891 15483 sw
tri 12891 15385 12989 15483 ne
rect 12989 15385 13343 15483
tri 13343 15385 13441 15483 sw
tri 13441 15385 13539 15483 ne
rect 13539 15385 13893 15483
tri 13893 15385 13991 15483 sw
tri 13991 15385 14089 15483 ne
rect 14089 15385 14443 15483
tri 14443 15385 14541 15483 sw
tri 14541 15385 14639 15483 ne
rect 14639 15385 14993 15483
tri 14993 15385 15091 15483 sw
tri 15091 15385 15189 15483 ne
rect 15189 15385 15543 15483
tri 15543 15385 15641 15483 sw
tri 15641 15385 15739 15483 ne
rect 15739 15385 16093 15483
tri 16093 15385 16191 15483 sw
tri 16191 15385 16289 15483 ne
rect 16289 15385 16643 15483
tri 16643 15385 16741 15483 sw
tri 16741 15385 16839 15483 ne
rect 16839 15385 17193 15483
tri 17193 15385 17291 15483 sw
tri 17291 15385 17389 15483 ne
rect 17389 15385 17743 15483
tri 17743 15385 17841 15483 sw
tri 17841 15385 17939 15483 ne
rect 17939 15385 18293 15483
tri 18293 15385 18391 15483 sw
tri 18391 15385 18489 15483 ne
rect 18489 15385 18843 15483
tri 18843 15385 18941 15483 sw
tri 18941 15385 19039 15483 ne
rect 19039 15385 19393 15483
tri 19393 15385 19491 15483 sw
tri 19491 15385 19589 15483 ne
rect 19589 15385 20300 15483
rect -2000 15287 241 15385
tri 241 15287 339 15385 sw
tri 339 15287 437 15385 ne
rect 437 15287 791 15385
tri 791 15287 889 15385 sw
tri 889 15287 987 15385 ne
rect 987 15287 1341 15385
tri 1341 15287 1439 15385 sw
tri 1439 15287 1537 15385 ne
rect 1537 15287 1891 15385
tri 1891 15287 1989 15385 sw
tri 1989 15287 2087 15385 ne
rect 2087 15287 2441 15385
tri 2441 15287 2539 15385 sw
tri 2539 15287 2637 15385 ne
rect 2637 15287 2991 15385
tri 2991 15287 3089 15385 sw
tri 3089 15287 3187 15385 ne
rect 3187 15287 3541 15385
tri 3541 15287 3639 15385 sw
tri 3639 15287 3737 15385 ne
rect 3737 15287 4091 15385
tri 4091 15287 4189 15385 sw
tri 4189 15287 4287 15385 ne
rect 4287 15287 4641 15385
tri 4641 15287 4739 15385 sw
tri 4739 15287 4837 15385 ne
rect 4837 15287 5191 15385
tri 5191 15287 5289 15385 sw
tri 5289 15287 5387 15385 ne
rect 5387 15287 5741 15385
tri 5741 15287 5839 15385 sw
tri 5839 15287 5937 15385 ne
rect 5937 15287 6291 15385
tri 6291 15287 6389 15385 sw
tri 6389 15287 6487 15385 ne
rect 6487 15287 6841 15385
tri 6841 15287 6939 15385 sw
tri 6939 15287 7037 15385 ne
rect 7037 15287 7391 15385
tri 7391 15287 7489 15385 sw
tri 7489 15287 7587 15385 ne
rect 7587 15287 7941 15385
tri 7941 15287 8039 15385 sw
tri 8039 15287 8137 15385 ne
rect 8137 15287 8491 15385
tri 8491 15287 8589 15385 sw
tri 8589 15287 8687 15385 ne
rect 8687 15287 9041 15385
tri 9041 15287 9139 15385 sw
tri 9139 15287 9237 15385 ne
rect 9237 15287 9591 15385
tri 9591 15287 9689 15385 sw
tri 9689 15287 9787 15385 ne
rect 9787 15287 10141 15385
tri 10141 15287 10239 15385 sw
tri 10239 15287 10337 15385 ne
rect 10337 15287 10691 15385
tri 10691 15287 10789 15385 sw
tri 10789 15287 10887 15385 ne
rect 10887 15287 11241 15385
tri 11241 15287 11339 15385 sw
tri 11339 15287 11437 15385 ne
rect 11437 15287 11791 15385
tri 11791 15287 11889 15385 sw
tri 11889 15287 11987 15385 ne
rect 11987 15287 12341 15385
tri 12341 15287 12439 15385 sw
tri 12439 15287 12537 15385 ne
rect 12537 15287 12891 15385
tri 12891 15287 12989 15385 sw
tri 12989 15287 13087 15385 ne
rect 13087 15287 13441 15385
tri 13441 15287 13539 15385 sw
tri 13539 15287 13637 15385 ne
rect 13637 15287 13991 15385
tri 13991 15287 14089 15385 sw
tri 14089 15287 14187 15385 ne
rect 14187 15287 14541 15385
tri 14541 15287 14639 15385 sw
tri 14639 15287 14737 15385 ne
rect 14737 15287 15091 15385
tri 15091 15287 15189 15385 sw
tri 15189 15287 15287 15385 ne
rect 15287 15287 15641 15385
tri 15641 15287 15739 15385 sw
tri 15739 15287 15837 15385 ne
rect 15837 15287 16191 15385
tri 16191 15287 16289 15385 sw
tri 16289 15287 16387 15385 ne
rect 16387 15287 16741 15385
tri 16741 15287 16839 15385 sw
tri 16839 15287 16937 15385 ne
rect 16937 15287 17291 15385
tri 17291 15287 17389 15385 sw
tri 17389 15287 17487 15385 ne
rect 17487 15287 17841 15385
tri 17841 15287 17939 15385 sw
tri 17939 15287 18037 15385 ne
rect 18037 15287 18391 15385
tri 18391 15287 18489 15385 sw
tri 18489 15287 18587 15385 ne
rect 18587 15287 18941 15385
tri 18941 15287 19039 15385 sw
tri 19039 15287 19137 15385 ne
rect 19137 15287 19491 15385
tri 19491 15287 19589 15385 sw
tri 19589 15287 19687 15385 ne
rect 19687 15287 20300 15385
rect -2000 15189 339 15287
tri 339 15189 437 15287 sw
tri 437 15189 535 15287 ne
rect 535 15189 889 15287
tri 889 15189 987 15287 sw
tri 987 15189 1085 15287 ne
rect 1085 15189 1439 15287
tri 1439 15189 1537 15287 sw
tri 1537 15189 1635 15287 ne
rect 1635 15189 1989 15287
tri 1989 15189 2087 15287 sw
tri 2087 15189 2185 15287 ne
rect 2185 15189 2539 15287
tri 2539 15189 2637 15287 sw
tri 2637 15189 2735 15287 ne
rect 2735 15189 3089 15287
tri 3089 15189 3187 15287 sw
tri 3187 15189 3285 15287 ne
rect 3285 15189 3639 15287
tri 3639 15189 3737 15287 sw
tri 3737 15189 3835 15287 ne
rect 3835 15189 4189 15287
tri 4189 15189 4287 15287 sw
tri 4287 15189 4385 15287 ne
rect 4385 15189 4739 15287
tri 4739 15189 4837 15287 sw
tri 4837 15189 4935 15287 ne
rect 4935 15189 5289 15287
tri 5289 15189 5387 15287 sw
tri 5387 15189 5485 15287 ne
rect 5485 15189 5839 15287
tri 5839 15189 5937 15287 sw
tri 5937 15189 6035 15287 ne
rect 6035 15189 6389 15287
tri 6389 15189 6487 15287 sw
tri 6487 15189 6585 15287 ne
rect 6585 15189 6939 15287
tri 6939 15189 7037 15287 sw
tri 7037 15189 7135 15287 ne
rect 7135 15189 7489 15287
tri 7489 15189 7587 15287 sw
tri 7587 15189 7685 15287 ne
rect 7685 15189 8039 15287
tri 8039 15189 8137 15287 sw
tri 8137 15189 8235 15287 ne
rect 8235 15189 8589 15287
tri 8589 15189 8687 15287 sw
tri 8687 15189 8785 15287 ne
rect 8785 15189 9139 15287
tri 9139 15189 9237 15287 sw
tri 9237 15189 9335 15287 ne
rect 9335 15189 9689 15287
tri 9689 15189 9787 15287 sw
tri 9787 15189 9885 15287 ne
rect 9885 15189 10239 15287
tri 10239 15189 10337 15287 sw
tri 10337 15189 10435 15287 ne
rect 10435 15189 10789 15287
tri 10789 15189 10887 15287 sw
tri 10887 15189 10985 15287 ne
rect 10985 15189 11339 15287
tri 11339 15189 11437 15287 sw
tri 11437 15189 11535 15287 ne
rect 11535 15189 11889 15287
tri 11889 15189 11987 15287 sw
tri 11987 15189 12085 15287 ne
rect 12085 15189 12439 15287
tri 12439 15189 12537 15287 sw
tri 12537 15189 12635 15287 ne
rect 12635 15189 12989 15287
tri 12989 15189 13087 15287 sw
tri 13087 15189 13185 15287 ne
rect 13185 15189 13539 15287
tri 13539 15189 13637 15287 sw
tri 13637 15189 13735 15287 ne
rect 13735 15189 14089 15287
tri 14089 15189 14187 15287 sw
tri 14187 15189 14285 15287 ne
rect 14285 15189 14639 15287
tri 14639 15189 14737 15287 sw
tri 14737 15189 14835 15287 ne
rect 14835 15189 15189 15287
tri 15189 15189 15287 15287 sw
tri 15287 15189 15385 15287 ne
rect 15385 15189 15739 15287
tri 15739 15189 15837 15287 sw
tri 15837 15189 15935 15287 ne
rect 15935 15189 16289 15287
tri 16289 15189 16387 15287 sw
tri 16387 15189 16485 15287 ne
rect 16485 15189 16839 15287
tri 16839 15189 16937 15287 sw
tri 16937 15189 17035 15287 ne
rect 17035 15189 17389 15287
tri 17389 15189 17487 15287 sw
tri 17487 15189 17585 15287 ne
rect 17585 15189 17939 15287
tri 17939 15189 18037 15287 sw
tri 18037 15189 18135 15287 ne
rect 18135 15189 18489 15287
tri 18489 15189 18587 15287 sw
tri 18587 15189 18685 15287 ne
rect 18685 15189 19039 15287
tri 19039 15189 19137 15287 sw
tri 19137 15189 19235 15287 ne
rect 19235 15189 19589 15287
tri 19589 15189 19687 15287 sw
rect 20800 15189 21800 15837
rect -2000 15185 437 15189
rect -2000 15065 215 15185
rect 335 15091 437 15185
tri 437 15091 535 15189 sw
tri 535 15091 633 15189 ne
rect 633 15185 987 15189
rect 633 15091 765 15185
rect 335 15065 535 15091
rect -2000 15061 535 15065
rect -2000 14413 -1000 15061
tri 113 14963 211 15061 ne
rect 211 15013 535 15061
tri 535 15013 613 15091 sw
tri 633 15013 711 15091 ne
rect 711 15065 765 15091
rect 885 15091 987 15185
tri 987 15091 1085 15189 sw
tri 1085 15091 1183 15189 ne
rect 1183 15185 1537 15189
rect 1183 15091 1315 15185
rect 885 15065 1085 15091
rect 711 15013 1085 15065
tri 1085 15013 1163 15091 sw
tri 1183 15013 1261 15091 ne
rect 1261 15065 1315 15091
rect 1435 15091 1537 15185
tri 1537 15091 1635 15189 sw
tri 1635 15091 1733 15189 ne
rect 1733 15185 2087 15189
rect 1733 15091 1865 15185
rect 1435 15065 1635 15091
rect 1261 15013 1635 15065
tri 1635 15013 1713 15091 sw
tri 1733 15013 1811 15091 ne
rect 1811 15065 1865 15091
rect 1985 15091 2087 15185
tri 2087 15091 2185 15189 sw
tri 2185 15091 2283 15189 ne
rect 2283 15185 2637 15189
rect 2283 15091 2415 15185
rect 1985 15065 2185 15091
rect 1811 15013 2185 15065
tri 2185 15013 2263 15091 sw
tri 2283 15013 2361 15091 ne
rect 2361 15065 2415 15091
rect 2535 15091 2637 15185
tri 2637 15091 2735 15189 sw
tri 2735 15091 2833 15189 ne
rect 2833 15185 3187 15189
rect 2833 15091 2965 15185
rect 2535 15065 2735 15091
rect 2361 15013 2735 15065
tri 2735 15013 2813 15091 sw
tri 2833 15013 2911 15091 ne
rect 2911 15065 2965 15091
rect 3085 15091 3187 15185
tri 3187 15091 3285 15189 sw
tri 3285 15091 3383 15189 ne
rect 3383 15185 3737 15189
rect 3383 15091 3515 15185
rect 3085 15065 3285 15091
rect 2911 15013 3285 15065
tri 3285 15013 3363 15091 sw
tri 3383 15013 3461 15091 ne
rect 3461 15065 3515 15091
rect 3635 15091 3737 15185
tri 3737 15091 3835 15189 sw
tri 3835 15091 3933 15189 ne
rect 3933 15185 4287 15189
rect 3933 15091 4065 15185
rect 3635 15065 3835 15091
rect 3461 15013 3835 15065
tri 3835 15013 3913 15091 sw
tri 3933 15013 4011 15091 ne
rect 4011 15065 4065 15091
rect 4185 15091 4287 15185
tri 4287 15091 4385 15189 sw
tri 4385 15091 4483 15189 ne
rect 4483 15185 4837 15189
rect 4483 15091 4615 15185
rect 4185 15065 4385 15091
rect 4011 15013 4385 15065
tri 4385 15013 4463 15091 sw
tri 4483 15013 4561 15091 ne
rect 4561 15065 4615 15091
rect 4735 15091 4837 15185
tri 4837 15091 4935 15189 sw
tri 4935 15091 5033 15189 ne
rect 5033 15185 5387 15189
rect 5033 15091 5165 15185
rect 4735 15065 4935 15091
rect 4561 15013 4935 15065
tri 4935 15013 5013 15091 sw
tri 5033 15013 5111 15091 ne
rect 5111 15065 5165 15091
rect 5285 15091 5387 15185
tri 5387 15091 5485 15189 sw
tri 5485 15091 5583 15189 ne
rect 5583 15185 5937 15189
rect 5583 15091 5715 15185
rect 5285 15065 5485 15091
rect 5111 15013 5485 15065
tri 5485 15013 5563 15091 sw
tri 5583 15013 5661 15091 ne
rect 5661 15065 5715 15091
rect 5835 15091 5937 15185
tri 5937 15091 6035 15189 sw
tri 6035 15091 6133 15189 ne
rect 6133 15185 6487 15189
rect 6133 15091 6265 15185
rect 5835 15065 6035 15091
rect 5661 15013 6035 15065
tri 6035 15013 6113 15091 sw
tri 6133 15013 6211 15091 ne
rect 6211 15065 6265 15091
rect 6385 15091 6487 15185
tri 6487 15091 6585 15189 sw
tri 6585 15091 6683 15189 ne
rect 6683 15185 7037 15189
rect 6683 15091 6815 15185
rect 6385 15065 6585 15091
rect 6211 15013 6585 15065
tri 6585 15013 6663 15091 sw
tri 6683 15013 6761 15091 ne
rect 6761 15065 6815 15091
rect 6935 15091 7037 15185
tri 7037 15091 7135 15189 sw
tri 7135 15091 7233 15189 ne
rect 7233 15185 7587 15189
rect 7233 15091 7365 15185
rect 6935 15065 7135 15091
rect 6761 15013 7135 15065
tri 7135 15013 7213 15091 sw
tri 7233 15013 7311 15091 ne
rect 7311 15065 7365 15091
rect 7485 15091 7587 15185
tri 7587 15091 7685 15189 sw
tri 7685 15091 7783 15189 ne
rect 7783 15185 8137 15189
rect 7783 15091 7915 15185
rect 7485 15065 7685 15091
rect 7311 15013 7685 15065
tri 7685 15013 7763 15091 sw
tri 7783 15013 7861 15091 ne
rect 7861 15065 7915 15091
rect 8035 15091 8137 15185
tri 8137 15091 8235 15189 sw
tri 8235 15091 8333 15189 ne
rect 8333 15185 8687 15189
rect 8333 15091 8465 15185
rect 8035 15065 8235 15091
rect 7861 15013 8235 15065
tri 8235 15013 8313 15091 sw
tri 8333 15013 8411 15091 ne
rect 8411 15065 8465 15091
rect 8585 15091 8687 15185
tri 8687 15091 8785 15189 sw
tri 8785 15091 8883 15189 ne
rect 8883 15185 9237 15189
rect 8883 15091 9015 15185
rect 8585 15065 8785 15091
rect 8411 15013 8785 15065
tri 8785 15013 8863 15091 sw
tri 8883 15013 8961 15091 ne
rect 8961 15065 9015 15091
rect 9135 15091 9237 15185
tri 9237 15091 9335 15189 sw
tri 9335 15091 9433 15189 ne
rect 9433 15185 9787 15189
rect 9433 15091 9565 15185
rect 9135 15065 9335 15091
rect 8961 15013 9335 15065
tri 9335 15013 9413 15091 sw
tri 9433 15013 9511 15091 ne
rect 9511 15065 9565 15091
rect 9685 15091 9787 15185
tri 9787 15091 9885 15189 sw
tri 9885 15091 9983 15189 ne
rect 9983 15185 10337 15189
rect 9983 15091 10115 15185
rect 9685 15065 9885 15091
rect 9511 15013 9885 15065
tri 9885 15013 9963 15091 sw
tri 9983 15013 10061 15091 ne
rect 10061 15065 10115 15091
rect 10235 15091 10337 15185
tri 10337 15091 10435 15189 sw
tri 10435 15091 10533 15189 ne
rect 10533 15185 10887 15189
rect 10533 15091 10665 15185
rect 10235 15065 10435 15091
rect 10061 15013 10435 15065
tri 10435 15013 10513 15091 sw
tri 10533 15013 10611 15091 ne
rect 10611 15065 10665 15091
rect 10785 15091 10887 15185
tri 10887 15091 10985 15189 sw
tri 10985 15091 11083 15189 ne
rect 11083 15185 11437 15189
rect 11083 15091 11215 15185
rect 10785 15065 10985 15091
rect 10611 15013 10985 15065
tri 10985 15013 11063 15091 sw
tri 11083 15013 11161 15091 ne
rect 11161 15065 11215 15091
rect 11335 15091 11437 15185
tri 11437 15091 11535 15189 sw
tri 11535 15091 11633 15189 ne
rect 11633 15185 11987 15189
rect 11633 15091 11765 15185
rect 11335 15065 11535 15091
rect 11161 15013 11535 15065
tri 11535 15013 11613 15091 sw
tri 11633 15013 11711 15091 ne
rect 11711 15065 11765 15091
rect 11885 15091 11987 15185
tri 11987 15091 12085 15189 sw
tri 12085 15091 12183 15189 ne
rect 12183 15185 12537 15189
rect 12183 15091 12315 15185
rect 11885 15065 12085 15091
rect 11711 15013 12085 15065
tri 12085 15013 12163 15091 sw
tri 12183 15013 12261 15091 ne
rect 12261 15065 12315 15091
rect 12435 15091 12537 15185
tri 12537 15091 12635 15189 sw
tri 12635 15091 12733 15189 ne
rect 12733 15185 13087 15189
rect 12733 15091 12865 15185
rect 12435 15065 12635 15091
rect 12261 15013 12635 15065
tri 12635 15013 12713 15091 sw
tri 12733 15013 12811 15091 ne
rect 12811 15065 12865 15091
rect 12985 15091 13087 15185
tri 13087 15091 13185 15189 sw
tri 13185 15091 13283 15189 ne
rect 13283 15185 13637 15189
rect 13283 15091 13415 15185
rect 12985 15065 13185 15091
rect 12811 15013 13185 15065
tri 13185 15013 13263 15091 sw
tri 13283 15013 13361 15091 ne
rect 13361 15065 13415 15091
rect 13535 15091 13637 15185
tri 13637 15091 13735 15189 sw
tri 13735 15091 13833 15189 ne
rect 13833 15185 14187 15189
rect 13833 15091 13965 15185
rect 13535 15065 13735 15091
rect 13361 15013 13735 15065
tri 13735 15013 13813 15091 sw
tri 13833 15013 13911 15091 ne
rect 13911 15065 13965 15091
rect 14085 15091 14187 15185
tri 14187 15091 14285 15189 sw
tri 14285 15091 14383 15189 ne
rect 14383 15185 14737 15189
rect 14383 15091 14515 15185
rect 14085 15065 14285 15091
rect 13911 15013 14285 15065
tri 14285 15013 14363 15091 sw
tri 14383 15013 14461 15091 ne
rect 14461 15065 14515 15091
rect 14635 15091 14737 15185
tri 14737 15091 14835 15189 sw
tri 14835 15091 14933 15189 ne
rect 14933 15185 15287 15189
rect 14933 15091 15065 15185
rect 14635 15065 14835 15091
rect 14461 15013 14835 15065
tri 14835 15013 14913 15091 sw
tri 14933 15013 15011 15091 ne
rect 15011 15065 15065 15091
rect 15185 15091 15287 15185
tri 15287 15091 15385 15189 sw
tri 15385 15091 15483 15189 ne
rect 15483 15185 15837 15189
rect 15483 15091 15615 15185
rect 15185 15065 15385 15091
rect 15011 15013 15385 15065
tri 15385 15013 15463 15091 sw
tri 15483 15013 15561 15091 ne
rect 15561 15065 15615 15091
rect 15735 15091 15837 15185
tri 15837 15091 15935 15189 sw
tri 15935 15091 16033 15189 ne
rect 16033 15185 16387 15189
rect 16033 15091 16165 15185
rect 15735 15065 15935 15091
rect 15561 15013 15935 15065
tri 15935 15013 16013 15091 sw
tri 16033 15013 16111 15091 ne
rect 16111 15065 16165 15091
rect 16285 15091 16387 15185
tri 16387 15091 16485 15189 sw
tri 16485 15091 16583 15189 ne
rect 16583 15185 16937 15189
rect 16583 15091 16715 15185
rect 16285 15065 16485 15091
rect 16111 15013 16485 15065
tri 16485 15013 16563 15091 sw
tri 16583 15013 16661 15091 ne
rect 16661 15065 16715 15091
rect 16835 15091 16937 15185
tri 16937 15091 17035 15189 sw
tri 17035 15091 17133 15189 ne
rect 17133 15185 17487 15189
rect 17133 15091 17265 15185
rect 16835 15065 17035 15091
rect 16661 15013 17035 15065
tri 17035 15013 17113 15091 sw
tri 17133 15013 17211 15091 ne
rect 17211 15065 17265 15091
rect 17385 15091 17487 15185
tri 17487 15091 17585 15189 sw
tri 17585 15091 17683 15189 ne
rect 17683 15185 18037 15189
rect 17683 15091 17815 15185
rect 17385 15065 17585 15091
rect 17211 15013 17585 15065
tri 17585 15013 17663 15091 sw
tri 17683 15013 17761 15091 ne
rect 17761 15065 17815 15091
rect 17935 15091 18037 15185
tri 18037 15091 18135 15189 sw
tri 18135 15091 18233 15189 ne
rect 18233 15185 18587 15189
rect 18233 15091 18365 15185
rect 17935 15065 18135 15091
rect 17761 15013 18135 15065
tri 18135 15013 18213 15091 sw
tri 18233 15013 18311 15091 ne
rect 18311 15065 18365 15091
rect 18485 15091 18587 15185
tri 18587 15091 18685 15189 sw
tri 18685 15091 18783 15189 ne
rect 18783 15185 19137 15189
rect 18783 15091 18915 15185
rect 18485 15065 18685 15091
rect 18311 15013 18685 15065
tri 18685 15013 18763 15091 sw
tri 18783 15013 18861 15091 ne
rect 18861 15065 18915 15091
rect 19035 15091 19137 15185
tri 19137 15091 19235 15189 sw
tri 19235 15091 19333 15189 ne
rect 19333 15185 21800 15189
rect 19333 15091 19465 15185
rect 19035 15065 19235 15091
rect 18861 15013 19235 15065
tri 19235 15013 19313 15091 sw
tri 19333 15013 19411 15091 ne
rect 19411 15065 19465 15091
rect 19585 15065 21800 15185
rect 19411 15013 21800 15065
rect 211 14963 613 15013
rect -500 14913 113 14963
tri 113 14913 163 14963 sw
tri 211 14913 261 14963 ne
rect 261 14933 613 14963
tri 613 14933 693 15013 sw
tri 711 14933 791 15013 ne
rect 791 14933 1163 15013
tri 1163 14933 1243 15013 sw
tri 1261 14933 1341 15013 ne
rect 1341 14933 1713 15013
tri 1713 14933 1793 15013 sw
tri 1811 14933 1891 15013 ne
rect 1891 14933 2263 15013
tri 2263 14933 2343 15013 sw
tri 2361 14933 2441 15013 ne
rect 2441 14933 2813 15013
tri 2813 14933 2893 15013 sw
tri 2911 14933 2991 15013 ne
rect 2991 14933 3363 15013
tri 3363 14933 3443 15013 sw
tri 3461 14933 3541 15013 ne
rect 3541 14933 3913 15013
tri 3913 14933 3993 15013 sw
tri 4011 14933 4091 15013 ne
rect 4091 14933 4463 15013
tri 4463 14933 4543 15013 sw
tri 4561 14933 4641 15013 ne
rect 4641 14933 5013 15013
tri 5013 14933 5093 15013 sw
tri 5111 14933 5191 15013 ne
rect 5191 14933 5563 15013
tri 5563 14933 5643 15013 sw
tri 5661 14933 5741 15013 ne
rect 5741 14933 6113 15013
tri 6113 14933 6193 15013 sw
tri 6211 14933 6291 15013 ne
rect 6291 14933 6663 15013
tri 6663 14933 6743 15013 sw
tri 6761 14933 6841 15013 ne
rect 6841 14933 7213 15013
tri 7213 14933 7293 15013 sw
tri 7311 14933 7391 15013 ne
rect 7391 14933 7763 15013
tri 7763 14933 7843 15013 sw
tri 7861 14933 7941 15013 ne
rect 7941 14933 8313 15013
tri 8313 14933 8393 15013 sw
tri 8411 14933 8491 15013 ne
rect 8491 14933 8863 15013
tri 8863 14933 8943 15013 sw
tri 8961 14933 9041 15013 ne
rect 9041 14933 9413 15013
tri 9413 14933 9493 15013 sw
tri 9511 14933 9591 15013 ne
rect 9591 14933 9963 15013
tri 9963 14933 10043 15013 sw
tri 10061 14933 10141 15013 ne
rect 10141 14933 10513 15013
tri 10513 14933 10593 15013 sw
tri 10611 14933 10691 15013 ne
rect 10691 14933 11063 15013
tri 11063 14933 11143 15013 sw
tri 11161 14933 11241 15013 ne
rect 11241 14933 11613 15013
tri 11613 14933 11693 15013 sw
tri 11711 14933 11791 15013 ne
rect 11791 14933 12163 15013
tri 12163 14933 12243 15013 sw
tri 12261 14933 12341 15013 ne
rect 12341 14933 12713 15013
tri 12713 14933 12793 15013 sw
tri 12811 14933 12891 15013 ne
rect 12891 14933 13263 15013
tri 13263 14933 13343 15013 sw
tri 13361 14933 13441 15013 ne
rect 13441 14933 13813 15013
tri 13813 14933 13893 15013 sw
tri 13911 14933 13991 15013 ne
rect 13991 14933 14363 15013
tri 14363 14933 14443 15013 sw
tri 14461 14933 14541 15013 ne
rect 14541 14933 14913 15013
tri 14913 14933 14993 15013 sw
tri 15011 14933 15091 15013 ne
rect 15091 14933 15463 15013
tri 15463 14933 15543 15013 sw
tri 15561 14933 15641 15013 ne
rect 15641 14933 16013 15013
tri 16013 14933 16093 15013 sw
tri 16111 14933 16191 15013 ne
rect 16191 14933 16563 15013
tri 16563 14933 16643 15013 sw
tri 16661 14933 16741 15013 ne
rect 16741 14933 17113 15013
tri 17113 14933 17193 15013 sw
tri 17211 14933 17291 15013 ne
rect 17291 14933 17663 15013
tri 17663 14933 17743 15013 sw
tri 17761 14933 17841 15013 ne
rect 17841 14933 18213 15013
tri 18213 14933 18293 15013 sw
tri 18311 14933 18391 15013 ne
rect 18391 14933 18763 15013
tri 18763 14933 18843 15013 sw
tri 18861 14933 18941 15013 ne
rect 18941 14933 19313 15013
tri 19313 14933 19393 15013 sw
tri 19411 14933 19491 15013 ne
rect 19491 14933 20100 15013
rect 261 14913 693 14933
rect -500 14835 163 14913
tri 163 14835 241 14913 sw
tri 261 14835 339 14913 ne
rect 339 14835 693 14913
tri 693 14835 791 14933 sw
tri 791 14835 889 14933 ne
rect 889 14835 1243 14933
tri 1243 14835 1341 14933 sw
tri 1341 14835 1439 14933 ne
rect 1439 14835 1793 14933
tri 1793 14835 1891 14933 sw
tri 1891 14835 1989 14933 ne
rect 1989 14835 2343 14933
tri 2343 14835 2441 14933 sw
tri 2441 14835 2539 14933 ne
rect 2539 14835 2893 14933
tri 2893 14835 2991 14933 sw
tri 2991 14835 3089 14933 ne
rect 3089 14835 3443 14933
tri 3443 14835 3541 14933 sw
tri 3541 14835 3639 14933 ne
rect 3639 14835 3993 14933
tri 3993 14835 4091 14933 sw
tri 4091 14835 4189 14933 ne
rect 4189 14835 4543 14933
tri 4543 14835 4641 14933 sw
tri 4641 14835 4739 14933 ne
rect 4739 14835 5093 14933
tri 5093 14835 5191 14933 sw
tri 5191 14835 5289 14933 ne
rect 5289 14835 5643 14933
tri 5643 14835 5741 14933 sw
tri 5741 14835 5839 14933 ne
rect 5839 14835 6193 14933
tri 6193 14835 6291 14933 sw
tri 6291 14835 6389 14933 ne
rect 6389 14835 6743 14933
tri 6743 14835 6841 14933 sw
tri 6841 14835 6939 14933 ne
rect 6939 14835 7293 14933
tri 7293 14835 7391 14933 sw
tri 7391 14835 7489 14933 ne
rect 7489 14835 7843 14933
tri 7843 14835 7941 14933 sw
tri 7941 14835 8039 14933 ne
rect 8039 14835 8393 14933
tri 8393 14835 8491 14933 sw
tri 8491 14835 8589 14933 ne
rect 8589 14835 8943 14933
tri 8943 14835 9041 14933 sw
tri 9041 14835 9139 14933 ne
rect 9139 14835 9493 14933
tri 9493 14835 9591 14933 sw
tri 9591 14835 9689 14933 ne
rect 9689 14835 10043 14933
tri 10043 14835 10141 14933 sw
tri 10141 14835 10239 14933 ne
rect 10239 14835 10593 14933
tri 10593 14835 10691 14933 sw
tri 10691 14835 10789 14933 ne
rect 10789 14835 11143 14933
tri 11143 14835 11241 14933 sw
tri 11241 14835 11339 14933 ne
rect 11339 14835 11693 14933
tri 11693 14835 11791 14933 sw
tri 11791 14835 11889 14933 ne
rect 11889 14835 12243 14933
tri 12243 14835 12341 14933 sw
tri 12341 14835 12439 14933 ne
rect 12439 14835 12793 14933
tri 12793 14835 12891 14933 sw
tri 12891 14835 12989 14933 ne
rect 12989 14835 13343 14933
tri 13343 14835 13441 14933 sw
tri 13441 14835 13539 14933 ne
rect 13539 14835 13893 14933
tri 13893 14835 13991 14933 sw
tri 13991 14835 14089 14933 ne
rect 14089 14835 14443 14933
tri 14443 14835 14541 14933 sw
tri 14541 14835 14639 14933 ne
rect 14639 14835 14993 14933
tri 14993 14835 15091 14933 sw
tri 15091 14835 15189 14933 ne
rect 15189 14835 15543 14933
tri 15543 14835 15641 14933 sw
tri 15641 14835 15739 14933 ne
rect 15739 14835 16093 14933
tri 16093 14835 16191 14933 sw
tri 16191 14835 16289 14933 ne
rect 16289 14835 16643 14933
tri 16643 14835 16741 14933 sw
tri 16741 14835 16839 14933 ne
rect 16839 14835 17193 14933
tri 17193 14835 17291 14933 sw
tri 17291 14835 17389 14933 ne
rect 17389 14835 17743 14933
tri 17743 14835 17841 14933 sw
tri 17841 14835 17939 14933 ne
rect 17939 14835 18293 14933
tri 18293 14835 18391 14933 sw
tri 18391 14835 18489 14933 ne
rect 18489 14835 18843 14933
tri 18843 14835 18941 14933 sw
tri 18941 14835 19039 14933 ne
rect 19039 14835 19393 14933
tri 19393 14835 19491 14933 sw
tri 19491 14835 19589 14933 ne
rect 19589 14913 20100 14933
rect 20200 14913 21800 15013
rect 19589 14835 21800 14913
rect -500 14787 241 14835
rect -500 14687 -400 14787
rect -300 14737 241 14787
tri 241 14737 339 14835 sw
tri 339 14737 437 14835 ne
rect 437 14737 791 14835
tri 791 14737 889 14835 sw
tri 889 14737 987 14835 ne
rect 987 14737 1341 14835
tri 1341 14737 1439 14835 sw
tri 1439 14737 1537 14835 ne
rect 1537 14737 1891 14835
tri 1891 14737 1989 14835 sw
tri 1989 14737 2087 14835 ne
rect 2087 14737 2441 14835
tri 2441 14737 2539 14835 sw
tri 2539 14737 2637 14835 ne
rect 2637 14737 2991 14835
tri 2991 14737 3089 14835 sw
tri 3089 14737 3187 14835 ne
rect 3187 14737 3541 14835
tri 3541 14737 3639 14835 sw
tri 3639 14737 3737 14835 ne
rect 3737 14737 4091 14835
tri 4091 14737 4189 14835 sw
tri 4189 14737 4287 14835 ne
rect 4287 14737 4641 14835
tri 4641 14737 4739 14835 sw
tri 4739 14737 4837 14835 ne
rect 4837 14737 5191 14835
tri 5191 14737 5289 14835 sw
tri 5289 14737 5387 14835 ne
rect 5387 14737 5741 14835
tri 5741 14737 5839 14835 sw
tri 5839 14737 5937 14835 ne
rect 5937 14737 6291 14835
tri 6291 14737 6389 14835 sw
tri 6389 14737 6487 14835 ne
rect 6487 14737 6841 14835
tri 6841 14737 6939 14835 sw
tri 6939 14737 7037 14835 ne
rect 7037 14737 7391 14835
tri 7391 14737 7489 14835 sw
tri 7489 14737 7587 14835 ne
rect 7587 14737 7941 14835
tri 7941 14737 8039 14835 sw
tri 8039 14737 8137 14835 ne
rect 8137 14737 8491 14835
tri 8491 14737 8589 14835 sw
tri 8589 14737 8687 14835 ne
rect 8687 14737 9041 14835
tri 9041 14737 9139 14835 sw
tri 9139 14737 9237 14835 ne
rect 9237 14737 9591 14835
tri 9591 14737 9689 14835 sw
tri 9689 14737 9787 14835 ne
rect 9787 14737 10141 14835
tri 10141 14737 10239 14835 sw
tri 10239 14737 10337 14835 ne
rect 10337 14737 10691 14835
tri 10691 14737 10789 14835 sw
tri 10789 14737 10887 14835 ne
rect 10887 14737 11241 14835
tri 11241 14737 11339 14835 sw
tri 11339 14737 11437 14835 ne
rect 11437 14737 11791 14835
tri 11791 14737 11889 14835 sw
tri 11889 14737 11987 14835 ne
rect 11987 14737 12341 14835
tri 12341 14737 12439 14835 sw
tri 12439 14737 12537 14835 ne
rect 12537 14737 12891 14835
tri 12891 14737 12989 14835 sw
tri 12989 14737 13087 14835 ne
rect 13087 14737 13441 14835
tri 13441 14737 13539 14835 sw
tri 13539 14737 13637 14835 ne
rect 13637 14737 13991 14835
tri 13991 14737 14089 14835 sw
tri 14089 14737 14187 14835 ne
rect 14187 14737 14541 14835
tri 14541 14737 14639 14835 sw
tri 14639 14737 14737 14835 ne
rect 14737 14737 15091 14835
tri 15091 14737 15189 14835 sw
tri 15189 14737 15287 14835 ne
rect 15287 14737 15641 14835
tri 15641 14737 15739 14835 sw
tri 15739 14737 15837 14835 ne
rect 15837 14737 16191 14835
tri 16191 14737 16289 14835 sw
tri 16289 14737 16387 14835 ne
rect 16387 14737 16741 14835
tri 16741 14737 16839 14835 sw
tri 16839 14737 16937 14835 ne
rect 16937 14737 17291 14835
tri 17291 14737 17389 14835 sw
tri 17389 14737 17487 14835 ne
rect 17487 14737 17841 14835
tri 17841 14737 17939 14835 sw
tri 17939 14737 18037 14835 ne
rect 18037 14737 18391 14835
tri 18391 14737 18489 14835 sw
tri 18489 14737 18587 14835 ne
rect 18587 14737 18941 14835
tri 18941 14737 19039 14835 sw
tri 19039 14737 19137 14835 ne
rect 19137 14737 19491 14835
tri 19491 14737 19589 14835 sw
tri 19589 14737 19687 14835 ne
rect 19687 14737 21800 14835
rect -300 14687 339 14737
rect -500 14639 339 14687
tri 339 14639 437 14737 sw
tri 437 14639 535 14737 ne
rect 535 14639 889 14737
tri 889 14639 987 14737 sw
tri 987 14639 1085 14737 ne
rect 1085 14639 1439 14737
tri 1439 14639 1537 14737 sw
tri 1537 14639 1635 14737 ne
rect 1635 14639 1989 14737
tri 1989 14639 2087 14737 sw
tri 2087 14639 2185 14737 ne
rect 2185 14639 2539 14737
tri 2539 14639 2637 14737 sw
tri 2637 14639 2735 14737 ne
rect 2735 14639 3089 14737
tri 3089 14639 3187 14737 sw
tri 3187 14639 3285 14737 ne
rect 3285 14639 3639 14737
tri 3639 14639 3737 14737 sw
tri 3737 14639 3835 14737 ne
rect 3835 14639 4189 14737
tri 4189 14639 4287 14737 sw
tri 4287 14639 4385 14737 ne
rect 4385 14639 4739 14737
tri 4739 14639 4837 14737 sw
tri 4837 14639 4935 14737 ne
rect 4935 14639 5289 14737
tri 5289 14639 5387 14737 sw
tri 5387 14639 5485 14737 ne
rect 5485 14639 5839 14737
tri 5839 14639 5937 14737 sw
tri 5937 14639 6035 14737 ne
rect 6035 14639 6389 14737
tri 6389 14639 6487 14737 sw
tri 6487 14639 6585 14737 ne
rect 6585 14639 6939 14737
tri 6939 14639 7037 14737 sw
tri 7037 14639 7135 14737 ne
rect 7135 14639 7489 14737
tri 7489 14639 7587 14737 sw
tri 7587 14639 7685 14737 ne
rect 7685 14639 8039 14737
tri 8039 14639 8137 14737 sw
tri 8137 14639 8235 14737 ne
rect 8235 14639 8589 14737
tri 8589 14639 8687 14737 sw
tri 8687 14639 8785 14737 ne
rect 8785 14639 9139 14737
tri 9139 14639 9237 14737 sw
tri 9237 14639 9335 14737 ne
rect 9335 14639 9689 14737
tri 9689 14639 9787 14737 sw
tri 9787 14639 9885 14737 ne
rect 9885 14639 10239 14737
tri 10239 14639 10337 14737 sw
tri 10337 14639 10435 14737 ne
rect 10435 14639 10789 14737
tri 10789 14639 10887 14737 sw
tri 10887 14639 10985 14737 ne
rect 10985 14639 11339 14737
tri 11339 14639 11437 14737 sw
tri 11437 14639 11535 14737 ne
rect 11535 14639 11889 14737
tri 11889 14639 11987 14737 sw
tri 11987 14639 12085 14737 ne
rect 12085 14639 12439 14737
tri 12439 14639 12537 14737 sw
tri 12537 14639 12635 14737 ne
rect 12635 14639 12989 14737
tri 12989 14639 13087 14737 sw
tri 13087 14639 13185 14737 ne
rect 13185 14639 13539 14737
tri 13539 14639 13637 14737 sw
tri 13637 14639 13735 14737 ne
rect 13735 14639 14089 14737
tri 14089 14639 14187 14737 sw
tri 14187 14639 14285 14737 ne
rect 14285 14639 14639 14737
tri 14639 14639 14737 14737 sw
tri 14737 14639 14835 14737 ne
rect 14835 14639 15189 14737
tri 15189 14639 15287 14737 sw
tri 15287 14639 15385 14737 ne
rect 15385 14639 15739 14737
tri 15739 14639 15837 14737 sw
tri 15837 14639 15935 14737 ne
rect 15935 14639 16289 14737
tri 16289 14639 16387 14737 sw
tri 16387 14639 16485 14737 ne
rect 16485 14639 16839 14737
tri 16839 14639 16937 14737 sw
tri 16937 14639 17035 14737 ne
rect 17035 14639 17389 14737
tri 17389 14639 17487 14737 sw
tri 17487 14639 17585 14737 ne
rect 17585 14639 17939 14737
tri 17939 14639 18037 14737 sw
tri 18037 14639 18135 14737 ne
rect 18135 14639 18489 14737
tri 18489 14639 18587 14737 sw
tri 18587 14639 18685 14737 ne
rect 18685 14639 19039 14737
tri 19039 14639 19137 14737 sw
tri 19137 14639 19235 14737 ne
rect 19235 14639 19589 14737
tri 19589 14639 19687 14737 sw
rect -500 14635 437 14639
rect -500 14515 215 14635
rect 335 14541 437 14635
tri 437 14541 535 14639 sw
tri 535 14541 633 14639 ne
rect 633 14635 987 14639
rect 633 14541 765 14635
rect 335 14515 535 14541
rect -500 14511 535 14515
tri 535 14511 565 14541 sw
tri 633 14511 663 14541 ne
rect 663 14515 765 14541
rect 885 14541 987 14635
tri 987 14541 1085 14639 sw
tri 1085 14541 1183 14639 ne
rect 1183 14635 1537 14639
rect 1183 14541 1315 14635
rect 885 14515 1085 14541
rect 663 14511 1085 14515
tri 1085 14511 1115 14541 sw
tri 1183 14511 1213 14541 ne
rect 1213 14515 1315 14541
rect 1435 14541 1537 14635
tri 1537 14541 1635 14639 sw
tri 1635 14541 1733 14639 ne
rect 1733 14635 2087 14639
rect 1733 14541 1865 14635
rect 1435 14515 1635 14541
rect 1213 14511 1635 14515
tri 1635 14511 1665 14541 sw
tri 1733 14511 1763 14541 ne
rect 1763 14515 1865 14541
rect 1985 14541 2087 14635
tri 2087 14541 2185 14639 sw
tri 2185 14541 2283 14639 ne
rect 2283 14635 2637 14639
rect 2283 14541 2415 14635
rect 1985 14515 2185 14541
rect 1763 14511 2185 14515
tri 2185 14511 2215 14541 sw
tri 2283 14511 2313 14541 ne
rect 2313 14515 2415 14541
rect 2535 14541 2637 14635
tri 2637 14541 2735 14639 sw
tri 2735 14541 2833 14639 ne
rect 2833 14635 3187 14639
rect 2833 14541 2965 14635
rect 2535 14515 2735 14541
rect 2313 14511 2735 14515
tri 2735 14511 2765 14541 sw
tri 2833 14511 2863 14541 ne
rect 2863 14515 2965 14541
rect 3085 14541 3187 14635
tri 3187 14541 3285 14639 sw
tri 3285 14541 3383 14639 ne
rect 3383 14635 3737 14639
rect 3383 14541 3515 14635
rect 3085 14515 3285 14541
rect 2863 14511 3285 14515
tri 3285 14511 3315 14541 sw
tri 3383 14511 3413 14541 ne
rect 3413 14515 3515 14541
rect 3635 14541 3737 14635
tri 3737 14541 3835 14639 sw
tri 3835 14541 3933 14639 ne
rect 3933 14635 4287 14639
rect 3933 14541 4065 14635
rect 3635 14515 3835 14541
rect 3413 14511 3835 14515
tri 3835 14511 3865 14541 sw
tri 3933 14511 3963 14541 ne
rect 3963 14515 4065 14541
rect 4185 14541 4287 14635
tri 4287 14541 4385 14639 sw
tri 4385 14541 4483 14639 ne
rect 4483 14635 4837 14639
rect 4483 14541 4615 14635
rect 4185 14515 4385 14541
rect 3963 14511 4385 14515
tri 4385 14511 4415 14541 sw
tri 4483 14511 4513 14541 ne
rect 4513 14515 4615 14541
rect 4735 14541 4837 14635
tri 4837 14541 4935 14639 sw
tri 4935 14541 5033 14639 ne
rect 5033 14635 5387 14639
rect 5033 14541 5165 14635
rect 4735 14515 4935 14541
rect 4513 14511 4935 14515
tri 4935 14511 4965 14541 sw
tri 5033 14511 5063 14541 ne
rect 5063 14515 5165 14541
rect 5285 14541 5387 14635
tri 5387 14541 5485 14639 sw
tri 5485 14541 5583 14639 ne
rect 5583 14635 5937 14639
rect 5583 14541 5715 14635
rect 5285 14515 5485 14541
rect 5063 14511 5485 14515
tri 5485 14511 5515 14541 sw
tri 5583 14511 5613 14541 ne
rect 5613 14515 5715 14541
rect 5835 14541 5937 14635
tri 5937 14541 6035 14639 sw
tri 6035 14541 6133 14639 ne
rect 6133 14635 6487 14639
rect 6133 14541 6265 14635
rect 5835 14515 6035 14541
rect 5613 14511 6035 14515
tri 6035 14511 6065 14541 sw
tri 6133 14511 6163 14541 ne
rect 6163 14515 6265 14541
rect 6385 14541 6487 14635
tri 6487 14541 6585 14639 sw
tri 6585 14541 6683 14639 ne
rect 6683 14635 7037 14639
rect 6683 14541 6815 14635
rect 6385 14515 6585 14541
rect 6163 14511 6585 14515
tri 6585 14511 6615 14541 sw
tri 6683 14511 6713 14541 ne
rect 6713 14515 6815 14541
rect 6935 14541 7037 14635
tri 7037 14541 7135 14639 sw
tri 7135 14541 7233 14639 ne
rect 7233 14635 7587 14639
rect 7233 14541 7365 14635
rect 6935 14515 7135 14541
rect 6713 14511 7135 14515
tri 7135 14511 7165 14541 sw
tri 7233 14511 7263 14541 ne
rect 7263 14515 7365 14541
rect 7485 14541 7587 14635
tri 7587 14541 7685 14639 sw
tri 7685 14541 7783 14639 ne
rect 7783 14635 8137 14639
rect 7783 14541 7915 14635
rect 7485 14515 7685 14541
rect 7263 14511 7685 14515
tri 7685 14511 7715 14541 sw
tri 7783 14511 7813 14541 ne
rect 7813 14515 7915 14541
rect 8035 14541 8137 14635
tri 8137 14541 8235 14639 sw
tri 8235 14541 8333 14639 ne
rect 8333 14635 8687 14639
rect 8333 14541 8465 14635
rect 8035 14515 8235 14541
rect 7813 14511 8235 14515
tri 8235 14511 8265 14541 sw
tri 8333 14511 8363 14541 ne
rect 8363 14515 8465 14541
rect 8585 14541 8687 14635
tri 8687 14541 8785 14639 sw
tri 8785 14541 8883 14639 ne
rect 8883 14635 9237 14639
rect 8883 14541 9015 14635
rect 8585 14515 8785 14541
rect 8363 14511 8785 14515
tri 8785 14511 8815 14541 sw
tri 8883 14511 8913 14541 ne
rect 8913 14515 9015 14541
rect 9135 14541 9237 14635
tri 9237 14541 9335 14639 sw
tri 9335 14541 9433 14639 ne
rect 9433 14635 9787 14639
rect 9433 14541 9565 14635
rect 9135 14515 9335 14541
rect 8913 14511 9335 14515
tri 9335 14511 9365 14541 sw
tri 9433 14511 9463 14541 ne
rect 9463 14515 9565 14541
rect 9685 14541 9787 14635
tri 9787 14541 9885 14639 sw
tri 9885 14541 9983 14639 ne
rect 9983 14635 10337 14639
rect 9983 14541 10115 14635
rect 9685 14515 9885 14541
rect 9463 14511 9885 14515
tri 9885 14511 9915 14541 sw
tri 9983 14511 10013 14541 ne
rect 10013 14515 10115 14541
rect 10235 14541 10337 14635
tri 10337 14541 10435 14639 sw
tri 10435 14541 10533 14639 ne
rect 10533 14635 10887 14639
rect 10533 14541 10665 14635
rect 10235 14515 10435 14541
rect 10013 14511 10435 14515
tri 10435 14511 10465 14541 sw
tri 10533 14511 10563 14541 ne
rect 10563 14515 10665 14541
rect 10785 14541 10887 14635
tri 10887 14541 10985 14639 sw
tri 10985 14541 11083 14639 ne
rect 11083 14635 11437 14639
rect 11083 14541 11215 14635
rect 10785 14515 10985 14541
rect 10563 14511 10985 14515
tri 10985 14511 11015 14541 sw
tri 11083 14511 11113 14541 ne
rect 11113 14515 11215 14541
rect 11335 14541 11437 14635
tri 11437 14541 11535 14639 sw
tri 11535 14541 11633 14639 ne
rect 11633 14635 11987 14639
rect 11633 14541 11765 14635
rect 11335 14515 11535 14541
rect 11113 14511 11535 14515
tri 11535 14511 11565 14541 sw
tri 11633 14511 11663 14541 ne
rect 11663 14515 11765 14541
rect 11885 14541 11987 14635
tri 11987 14541 12085 14639 sw
tri 12085 14541 12183 14639 ne
rect 12183 14635 12537 14639
rect 12183 14541 12315 14635
rect 11885 14515 12085 14541
rect 11663 14511 12085 14515
tri 12085 14511 12115 14541 sw
tri 12183 14511 12213 14541 ne
rect 12213 14515 12315 14541
rect 12435 14541 12537 14635
tri 12537 14541 12635 14639 sw
tri 12635 14541 12733 14639 ne
rect 12733 14635 13087 14639
rect 12733 14541 12865 14635
rect 12435 14515 12635 14541
rect 12213 14511 12635 14515
tri 12635 14511 12665 14541 sw
tri 12733 14511 12763 14541 ne
rect 12763 14515 12865 14541
rect 12985 14541 13087 14635
tri 13087 14541 13185 14639 sw
tri 13185 14541 13283 14639 ne
rect 13283 14635 13637 14639
rect 13283 14541 13415 14635
rect 12985 14515 13185 14541
rect 12763 14511 13185 14515
tri 13185 14511 13215 14541 sw
tri 13283 14511 13313 14541 ne
rect 13313 14515 13415 14541
rect 13535 14541 13637 14635
tri 13637 14541 13735 14639 sw
tri 13735 14541 13833 14639 ne
rect 13833 14635 14187 14639
rect 13833 14541 13965 14635
rect 13535 14515 13735 14541
rect 13313 14511 13735 14515
tri 13735 14511 13765 14541 sw
tri 13833 14511 13863 14541 ne
rect 13863 14515 13965 14541
rect 14085 14541 14187 14635
tri 14187 14541 14285 14639 sw
tri 14285 14541 14383 14639 ne
rect 14383 14635 14737 14639
rect 14383 14541 14515 14635
rect 14085 14515 14285 14541
rect 13863 14511 14285 14515
tri 14285 14511 14315 14541 sw
tri 14383 14511 14413 14541 ne
rect 14413 14515 14515 14541
rect 14635 14541 14737 14635
tri 14737 14541 14835 14639 sw
tri 14835 14541 14933 14639 ne
rect 14933 14635 15287 14639
rect 14933 14541 15065 14635
rect 14635 14515 14835 14541
rect 14413 14511 14835 14515
tri 14835 14511 14865 14541 sw
tri 14933 14511 14963 14541 ne
rect 14963 14515 15065 14541
rect 15185 14541 15287 14635
tri 15287 14541 15385 14639 sw
tri 15385 14541 15483 14639 ne
rect 15483 14635 15837 14639
rect 15483 14541 15615 14635
rect 15185 14515 15385 14541
rect 14963 14511 15385 14515
tri 15385 14511 15415 14541 sw
tri 15483 14511 15513 14541 ne
rect 15513 14515 15615 14541
rect 15735 14541 15837 14635
tri 15837 14541 15935 14639 sw
tri 15935 14541 16033 14639 ne
rect 16033 14635 16387 14639
rect 16033 14541 16165 14635
rect 15735 14515 15935 14541
rect 15513 14511 15935 14515
tri 15935 14511 15965 14541 sw
tri 16033 14511 16063 14541 ne
rect 16063 14515 16165 14541
rect 16285 14541 16387 14635
tri 16387 14541 16485 14639 sw
tri 16485 14541 16583 14639 ne
rect 16583 14635 16937 14639
rect 16583 14541 16715 14635
rect 16285 14515 16485 14541
rect 16063 14511 16485 14515
tri 16485 14511 16515 14541 sw
tri 16583 14511 16613 14541 ne
rect 16613 14515 16715 14541
rect 16835 14541 16937 14635
tri 16937 14541 17035 14639 sw
tri 17035 14541 17133 14639 ne
rect 17133 14635 17487 14639
rect 17133 14541 17265 14635
rect 16835 14515 17035 14541
rect 16613 14511 17035 14515
tri 17035 14511 17065 14541 sw
tri 17133 14511 17163 14541 ne
rect 17163 14515 17265 14541
rect 17385 14541 17487 14635
tri 17487 14541 17585 14639 sw
tri 17585 14541 17683 14639 ne
rect 17683 14635 18037 14639
rect 17683 14541 17815 14635
rect 17385 14515 17585 14541
rect 17163 14511 17585 14515
tri 17585 14511 17615 14541 sw
tri 17683 14511 17713 14541 ne
rect 17713 14515 17815 14541
rect 17935 14541 18037 14635
tri 18037 14541 18135 14639 sw
tri 18135 14541 18233 14639 ne
rect 18233 14635 18587 14639
rect 18233 14541 18365 14635
rect 17935 14515 18135 14541
rect 17713 14511 18135 14515
tri 18135 14511 18165 14541 sw
tri 18233 14511 18263 14541 ne
rect 18263 14515 18365 14541
rect 18485 14541 18587 14635
tri 18587 14541 18685 14639 sw
tri 18685 14541 18783 14639 ne
rect 18783 14635 19137 14639
rect 18783 14541 18915 14635
rect 18485 14515 18685 14541
rect 18263 14511 18685 14515
tri 18685 14511 18715 14541 sw
tri 18783 14511 18813 14541 ne
rect 18813 14515 18915 14541
rect 19035 14541 19137 14635
tri 19137 14541 19235 14639 sw
tri 19235 14541 19333 14639 ne
rect 19333 14635 20300 14639
rect 19333 14541 19465 14635
rect 19035 14515 19235 14541
rect 18813 14511 19235 14515
tri 19235 14511 19265 14541 sw
tri 19333 14511 19363 14541 ne
rect 19363 14515 19465 14541
rect 19585 14515 20300 14635
rect 19363 14511 20300 14515
tri 113 14413 211 14511 ne
rect 211 14413 565 14511
tri 565 14413 663 14511 sw
tri 663 14413 761 14511 ne
rect 761 14413 1115 14511
tri 1115 14413 1213 14511 sw
tri 1213 14413 1311 14511 ne
rect 1311 14413 1665 14511
tri 1665 14413 1763 14511 sw
tri 1763 14413 1861 14511 ne
rect 1861 14413 2215 14511
tri 2215 14413 2313 14511 sw
tri 2313 14413 2411 14511 ne
rect 2411 14413 2765 14511
tri 2765 14413 2863 14511 sw
tri 2863 14413 2961 14511 ne
rect 2961 14413 3315 14511
tri 3315 14413 3413 14511 sw
tri 3413 14413 3511 14511 ne
rect 3511 14413 3865 14511
tri 3865 14413 3963 14511 sw
tri 3963 14413 4061 14511 ne
rect 4061 14413 4415 14511
tri 4415 14413 4513 14511 sw
tri 4513 14413 4611 14511 ne
rect 4611 14413 4965 14511
tri 4965 14413 5063 14511 sw
tri 5063 14413 5161 14511 ne
rect 5161 14413 5515 14511
tri 5515 14413 5613 14511 sw
tri 5613 14413 5711 14511 ne
rect 5711 14413 6065 14511
tri 6065 14413 6163 14511 sw
tri 6163 14413 6261 14511 ne
rect 6261 14413 6615 14511
tri 6615 14413 6713 14511 sw
tri 6713 14413 6811 14511 ne
rect 6811 14413 7165 14511
tri 7165 14413 7263 14511 sw
tri 7263 14413 7361 14511 ne
rect 7361 14413 7715 14511
tri 7715 14413 7813 14511 sw
tri 7813 14413 7911 14511 ne
rect 7911 14413 8265 14511
tri 8265 14413 8363 14511 sw
tri 8363 14413 8461 14511 ne
rect 8461 14413 8815 14511
tri 8815 14413 8913 14511 sw
tri 8913 14413 9011 14511 ne
rect 9011 14413 9365 14511
tri 9365 14413 9463 14511 sw
tri 9463 14413 9561 14511 ne
rect 9561 14413 9915 14511
tri 9915 14413 10013 14511 sw
tri 10013 14413 10111 14511 ne
rect 10111 14413 10465 14511
tri 10465 14413 10563 14511 sw
tri 10563 14413 10661 14511 ne
rect 10661 14413 11015 14511
tri 11015 14413 11113 14511 sw
tri 11113 14413 11211 14511 ne
rect 11211 14413 11565 14511
tri 11565 14413 11663 14511 sw
tri 11663 14413 11761 14511 ne
rect 11761 14413 12115 14511
tri 12115 14413 12213 14511 sw
tri 12213 14413 12311 14511 ne
rect 12311 14413 12665 14511
tri 12665 14413 12763 14511 sw
tri 12763 14413 12861 14511 ne
rect 12861 14413 13215 14511
tri 13215 14413 13313 14511 sw
tri 13313 14413 13411 14511 ne
rect 13411 14413 13765 14511
tri 13765 14413 13863 14511 sw
tri 13863 14413 13961 14511 ne
rect 13961 14413 14315 14511
tri 14315 14413 14413 14511 sw
tri 14413 14413 14511 14511 ne
rect 14511 14413 14865 14511
tri 14865 14413 14963 14511 sw
tri 14963 14413 15061 14511 ne
rect 15061 14413 15415 14511
tri 15415 14413 15513 14511 sw
tri 15513 14413 15611 14511 ne
rect 15611 14413 15965 14511
tri 15965 14413 16063 14511 sw
tri 16063 14413 16161 14511 ne
rect 16161 14413 16515 14511
tri 16515 14413 16613 14511 sw
tri 16613 14413 16711 14511 ne
rect 16711 14413 17065 14511
tri 17065 14413 17163 14511 sw
tri 17163 14413 17261 14511 ne
rect 17261 14413 17615 14511
tri 17615 14413 17713 14511 sw
tri 17713 14413 17811 14511 ne
rect 17811 14413 18165 14511
tri 18165 14413 18263 14511 sw
tri 18263 14413 18361 14511 ne
rect 18361 14413 18715 14511
tri 18715 14413 18813 14511 sw
tri 18813 14413 18911 14511 ne
rect 18911 14413 19265 14511
tri 19265 14413 19363 14511 sw
tri 19363 14413 19461 14511 ne
rect 19461 14413 20300 14511
rect -2000 14383 113 14413
tri 113 14383 143 14413 sw
tri 211 14383 241 14413 ne
rect 241 14383 663 14413
tri 663 14383 693 14413 sw
tri 761 14383 791 14413 ne
rect 791 14383 1213 14413
tri 1213 14383 1243 14413 sw
tri 1311 14383 1341 14413 ne
rect 1341 14383 1763 14413
tri 1763 14383 1793 14413 sw
tri 1861 14383 1891 14413 ne
rect 1891 14383 2313 14413
tri 2313 14383 2343 14413 sw
tri 2411 14383 2441 14413 ne
rect 2441 14383 2863 14413
tri 2863 14383 2893 14413 sw
tri 2961 14383 2991 14413 ne
rect 2991 14383 3413 14413
tri 3413 14383 3443 14413 sw
tri 3511 14383 3541 14413 ne
rect 3541 14383 3963 14413
tri 3963 14383 3993 14413 sw
tri 4061 14383 4091 14413 ne
rect 4091 14383 4513 14413
tri 4513 14383 4543 14413 sw
tri 4611 14383 4641 14413 ne
rect 4641 14383 5063 14413
tri 5063 14383 5093 14413 sw
tri 5161 14383 5191 14413 ne
rect 5191 14383 5613 14413
tri 5613 14383 5643 14413 sw
tri 5711 14383 5741 14413 ne
rect 5741 14383 6163 14413
tri 6163 14383 6193 14413 sw
tri 6261 14383 6291 14413 ne
rect 6291 14383 6713 14413
tri 6713 14383 6743 14413 sw
tri 6811 14383 6841 14413 ne
rect 6841 14383 7263 14413
tri 7263 14383 7293 14413 sw
tri 7361 14383 7391 14413 ne
rect 7391 14383 7813 14413
tri 7813 14383 7843 14413 sw
tri 7911 14383 7941 14413 ne
rect 7941 14383 8363 14413
tri 8363 14383 8393 14413 sw
tri 8461 14383 8491 14413 ne
rect 8491 14383 8913 14413
tri 8913 14383 8943 14413 sw
tri 9011 14383 9041 14413 ne
rect 9041 14383 9463 14413
tri 9463 14383 9493 14413 sw
tri 9561 14383 9591 14413 ne
rect 9591 14383 10013 14413
tri 10013 14383 10043 14413 sw
tri 10111 14383 10141 14413 ne
rect 10141 14383 10563 14413
tri 10563 14383 10593 14413 sw
tri 10661 14383 10691 14413 ne
rect 10691 14383 11113 14413
tri 11113 14383 11143 14413 sw
tri 11211 14383 11241 14413 ne
rect 11241 14383 11663 14413
tri 11663 14383 11693 14413 sw
tri 11761 14383 11791 14413 ne
rect 11791 14383 12213 14413
tri 12213 14383 12243 14413 sw
tri 12311 14383 12341 14413 ne
rect 12341 14383 12763 14413
tri 12763 14383 12793 14413 sw
tri 12861 14383 12891 14413 ne
rect 12891 14383 13313 14413
tri 13313 14383 13343 14413 sw
tri 13411 14383 13441 14413 ne
rect 13441 14383 13863 14413
tri 13863 14383 13893 14413 sw
tri 13961 14383 13991 14413 ne
rect 13991 14383 14413 14413
tri 14413 14383 14443 14413 sw
tri 14511 14383 14541 14413 ne
rect 14541 14383 14963 14413
tri 14963 14383 14993 14413 sw
tri 15061 14383 15091 14413 ne
rect 15091 14383 15513 14413
tri 15513 14383 15543 14413 sw
tri 15611 14383 15641 14413 ne
rect 15641 14383 16063 14413
tri 16063 14383 16093 14413 sw
tri 16161 14383 16191 14413 ne
rect 16191 14383 16613 14413
tri 16613 14383 16643 14413 sw
tri 16711 14383 16741 14413 ne
rect 16741 14383 17163 14413
tri 17163 14383 17193 14413 sw
tri 17261 14383 17291 14413 ne
rect 17291 14383 17713 14413
tri 17713 14383 17743 14413 sw
tri 17811 14383 17841 14413 ne
rect 17841 14383 18263 14413
tri 18263 14383 18293 14413 sw
tri 18361 14383 18391 14413 ne
rect 18391 14383 18813 14413
tri 18813 14383 18843 14413 sw
tri 18911 14383 18941 14413 ne
rect 18941 14383 19363 14413
tri 19363 14383 19393 14413 sw
tri 19461 14383 19491 14413 ne
rect 19491 14383 20300 14413
rect -2000 14285 143 14383
tri 143 14285 241 14383 sw
tri 241 14285 339 14383 ne
rect 339 14285 693 14383
tri 693 14285 791 14383 sw
tri 791 14285 889 14383 ne
rect 889 14285 1243 14383
tri 1243 14285 1341 14383 sw
tri 1341 14285 1439 14383 ne
rect 1439 14285 1793 14383
tri 1793 14285 1891 14383 sw
tri 1891 14285 1989 14383 ne
rect 1989 14285 2343 14383
tri 2343 14285 2441 14383 sw
tri 2441 14285 2539 14383 ne
rect 2539 14285 2893 14383
tri 2893 14285 2991 14383 sw
tri 2991 14285 3089 14383 ne
rect 3089 14285 3443 14383
tri 3443 14285 3541 14383 sw
tri 3541 14285 3639 14383 ne
rect 3639 14285 3993 14383
tri 3993 14285 4091 14383 sw
tri 4091 14285 4189 14383 ne
rect 4189 14285 4543 14383
tri 4543 14285 4641 14383 sw
tri 4641 14285 4739 14383 ne
rect 4739 14285 5093 14383
tri 5093 14285 5191 14383 sw
tri 5191 14285 5289 14383 ne
rect 5289 14285 5643 14383
tri 5643 14285 5741 14383 sw
tri 5741 14285 5839 14383 ne
rect 5839 14285 6193 14383
tri 6193 14285 6291 14383 sw
tri 6291 14285 6389 14383 ne
rect 6389 14285 6743 14383
tri 6743 14285 6841 14383 sw
tri 6841 14285 6939 14383 ne
rect 6939 14285 7293 14383
tri 7293 14285 7391 14383 sw
tri 7391 14285 7489 14383 ne
rect 7489 14285 7843 14383
tri 7843 14285 7941 14383 sw
tri 7941 14285 8039 14383 ne
rect 8039 14285 8393 14383
tri 8393 14285 8491 14383 sw
tri 8491 14285 8589 14383 ne
rect 8589 14285 8943 14383
tri 8943 14285 9041 14383 sw
tri 9041 14285 9139 14383 ne
rect 9139 14285 9493 14383
tri 9493 14285 9591 14383 sw
tri 9591 14285 9689 14383 ne
rect 9689 14285 10043 14383
tri 10043 14285 10141 14383 sw
tri 10141 14285 10239 14383 ne
rect 10239 14285 10593 14383
tri 10593 14285 10691 14383 sw
tri 10691 14285 10789 14383 ne
rect 10789 14285 11143 14383
tri 11143 14285 11241 14383 sw
tri 11241 14285 11339 14383 ne
rect 11339 14285 11693 14383
tri 11693 14285 11791 14383 sw
tri 11791 14285 11889 14383 ne
rect 11889 14285 12243 14383
tri 12243 14285 12341 14383 sw
tri 12341 14285 12439 14383 ne
rect 12439 14285 12793 14383
tri 12793 14285 12891 14383 sw
tri 12891 14285 12989 14383 ne
rect 12989 14285 13343 14383
tri 13343 14285 13441 14383 sw
tri 13441 14285 13539 14383 ne
rect 13539 14285 13893 14383
tri 13893 14285 13991 14383 sw
tri 13991 14285 14089 14383 ne
rect 14089 14285 14443 14383
tri 14443 14285 14541 14383 sw
tri 14541 14285 14639 14383 ne
rect 14639 14285 14993 14383
tri 14993 14285 15091 14383 sw
tri 15091 14285 15189 14383 ne
rect 15189 14285 15543 14383
tri 15543 14285 15641 14383 sw
tri 15641 14285 15739 14383 ne
rect 15739 14285 16093 14383
tri 16093 14285 16191 14383 sw
tri 16191 14285 16289 14383 ne
rect 16289 14285 16643 14383
tri 16643 14285 16741 14383 sw
tri 16741 14285 16839 14383 ne
rect 16839 14285 17193 14383
tri 17193 14285 17291 14383 sw
tri 17291 14285 17389 14383 ne
rect 17389 14285 17743 14383
tri 17743 14285 17841 14383 sw
tri 17841 14285 17939 14383 ne
rect 17939 14285 18293 14383
tri 18293 14285 18391 14383 sw
tri 18391 14285 18489 14383 ne
rect 18489 14285 18843 14383
tri 18843 14285 18941 14383 sw
tri 18941 14285 19039 14383 ne
rect 19039 14285 19393 14383
tri 19393 14285 19491 14383 sw
tri 19491 14285 19589 14383 ne
rect 19589 14285 20300 14383
rect -2000 14187 241 14285
tri 241 14187 339 14285 sw
tri 339 14187 437 14285 ne
rect 437 14187 791 14285
tri 791 14187 889 14285 sw
tri 889 14187 987 14285 ne
rect 987 14187 1341 14285
tri 1341 14187 1439 14285 sw
tri 1439 14187 1537 14285 ne
rect 1537 14187 1891 14285
tri 1891 14187 1989 14285 sw
tri 1989 14187 2087 14285 ne
rect 2087 14187 2441 14285
tri 2441 14187 2539 14285 sw
tri 2539 14187 2637 14285 ne
rect 2637 14187 2991 14285
tri 2991 14187 3089 14285 sw
tri 3089 14187 3187 14285 ne
rect 3187 14187 3541 14285
tri 3541 14187 3639 14285 sw
tri 3639 14187 3737 14285 ne
rect 3737 14187 4091 14285
tri 4091 14187 4189 14285 sw
tri 4189 14187 4287 14285 ne
rect 4287 14187 4641 14285
tri 4641 14187 4739 14285 sw
tri 4739 14187 4837 14285 ne
rect 4837 14187 5191 14285
tri 5191 14187 5289 14285 sw
tri 5289 14187 5387 14285 ne
rect 5387 14187 5741 14285
tri 5741 14187 5839 14285 sw
tri 5839 14187 5937 14285 ne
rect 5937 14187 6291 14285
tri 6291 14187 6389 14285 sw
tri 6389 14187 6487 14285 ne
rect 6487 14187 6841 14285
tri 6841 14187 6939 14285 sw
tri 6939 14187 7037 14285 ne
rect 7037 14187 7391 14285
tri 7391 14187 7489 14285 sw
tri 7489 14187 7587 14285 ne
rect 7587 14187 7941 14285
tri 7941 14187 8039 14285 sw
tri 8039 14187 8137 14285 ne
rect 8137 14187 8491 14285
tri 8491 14187 8589 14285 sw
tri 8589 14187 8687 14285 ne
rect 8687 14187 9041 14285
tri 9041 14187 9139 14285 sw
tri 9139 14187 9237 14285 ne
rect 9237 14187 9591 14285
tri 9591 14187 9689 14285 sw
tri 9689 14187 9787 14285 ne
rect 9787 14187 10141 14285
tri 10141 14187 10239 14285 sw
tri 10239 14187 10337 14285 ne
rect 10337 14187 10691 14285
tri 10691 14187 10789 14285 sw
tri 10789 14187 10887 14285 ne
rect 10887 14187 11241 14285
tri 11241 14187 11339 14285 sw
tri 11339 14187 11437 14285 ne
rect 11437 14187 11791 14285
tri 11791 14187 11889 14285 sw
tri 11889 14187 11987 14285 ne
rect 11987 14187 12341 14285
tri 12341 14187 12439 14285 sw
tri 12439 14187 12537 14285 ne
rect 12537 14187 12891 14285
tri 12891 14187 12989 14285 sw
tri 12989 14187 13087 14285 ne
rect 13087 14187 13441 14285
tri 13441 14187 13539 14285 sw
tri 13539 14187 13637 14285 ne
rect 13637 14187 13991 14285
tri 13991 14187 14089 14285 sw
tri 14089 14187 14187 14285 ne
rect 14187 14187 14541 14285
tri 14541 14187 14639 14285 sw
tri 14639 14187 14737 14285 ne
rect 14737 14187 15091 14285
tri 15091 14187 15189 14285 sw
tri 15189 14187 15287 14285 ne
rect 15287 14187 15641 14285
tri 15641 14187 15739 14285 sw
tri 15739 14187 15837 14285 ne
rect 15837 14187 16191 14285
tri 16191 14187 16289 14285 sw
tri 16289 14187 16387 14285 ne
rect 16387 14187 16741 14285
tri 16741 14187 16839 14285 sw
tri 16839 14187 16937 14285 ne
rect 16937 14187 17291 14285
tri 17291 14187 17389 14285 sw
tri 17389 14187 17487 14285 ne
rect 17487 14187 17841 14285
tri 17841 14187 17939 14285 sw
tri 17939 14187 18037 14285 ne
rect 18037 14187 18391 14285
tri 18391 14187 18489 14285 sw
tri 18489 14187 18587 14285 ne
rect 18587 14187 18941 14285
tri 18941 14187 19039 14285 sw
tri 19039 14187 19137 14285 ne
rect 19137 14187 19491 14285
tri 19491 14187 19589 14285 sw
tri 19589 14187 19687 14285 ne
rect 19687 14187 20300 14285
rect -2000 14089 339 14187
tri 339 14089 437 14187 sw
tri 437 14089 535 14187 ne
rect 535 14089 889 14187
tri 889 14089 987 14187 sw
tri 987 14089 1085 14187 ne
rect 1085 14089 1439 14187
tri 1439 14089 1537 14187 sw
tri 1537 14089 1635 14187 ne
rect 1635 14089 1989 14187
tri 1989 14089 2087 14187 sw
tri 2087 14089 2185 14187 ne
rect 2185 14089 2539 14187
tri 2539 14089 2637 14187 sw
tri 2637 14089 2735 14187 ne
rect 2735 14089 3089 14187
tri 3089 14089 3187 14187 sw
tri 3187 14089 3285 14187 ne
rect 3285 14089 3639 14187
tri 3639 14089 3737 14187 sw
tri 3737 14089 3835 14187 ne
rect 3835 14089 4189 14187
tri 4189 14089 4287 14187 sw
tri 4287 14089 4385 14187 ne
rect 4385 14089 4739 14187
tri 4739 14089 4837 14187 sw
tri 4837 14089 4935 14187 ne
rect 4935 14089 5289 14187
tri 5289 14089 5387 14187 sw
tri 5387 14089 5485 14187 ne
rect 5485 14089 5839 14187
tri 5839 14089 5937 14187 sw
tri 5937 14089 6035 14187 ne
rect 6035 14089 6389 14187
tri 6389 14089 6487 14187 sw
tri 6487 14089 6585 14187 ne
rect 6585 14089 6939 14187
tri 6939 14089 7037 14187 sw
tri 7037 14089 7135 14187 ne
rect 7135 14089 7489 14187
tri 7489 14089 7587 14187 sw
tri 7587 14089 7685 14187 ne
rect 7685 14089 8039 14187
tri 8039 14089 8137 14187 sw
tri 8137 14089 8235 14187 ne
rect 8235 14089 8589 14187
tri 8589 14089 8687 14187 sw
tri 8687 14089 8785 14187 ne
rect 8785 14089 9139 14187
tri 9139 14089 9237 14187 sw
tri 9237 14089 9335 14187 ne
rect 9335 14089 9689 14187
tri 9689 14089 9787 14187 sw
tri 9787 14089 9885 14187 ne
rect 9885 14089 10239 14187
tri 10239 14089 10337 14187 sw
tri 10337 14089 10435 14187 ne
rect 10435 14089 10789 14187
tri 10789 14089 10887 14187 sw
tri 10887 14089 10985 14187 ne
rect 10985 14089 11339 14187
tri 11339 14089 11437 14187 sw
tri 11437 14089 11535 14187 ne
rect 11535 14089 11889 14187
tri 11889 14089 11987 14187 sw
tri 11987 14089 12085 14187 ne
rect 12085 14089 12439 14187
tri 12439 14089 12537 14187 sw
tri 12537 14089 12635 14187 ne
rect 12635 14089 12989 14187
tri 12989 14089 13087 14187 sw
tri 13087 14089 13185 14187 ne
rect 13185 14089 13539 14187
tri 13539 14089 13637 14187 sw
tri 13637 14089 13735 14187 ne
rect 13735 14089 14089 14187
tri 14089 14089 14187 14187 sw
tri 14187 14089 14285 14187 ne
rect 14285 14089 14639 14187
tri 14639 14089 14737 14187 sw
tri 14737 14089 14835 14187 ne
rect 14835 14089 15189 14187
tri 15189 14089 15287 14187 sw
tri 15287 14089 15385 14187 ne
rect 15385 14089 15739 14187
tri 15739 14089 15837 14187 sw
tri 15837 14089 15935 14187 ne
rect 15935 14089 16289 14187
tri 16289 14089 16387 14187 sw
tri 16387 14089 16485 14187 ne
rect 16485 14089 16839 14187
tri 16839 14089 16937 14187 sw
tri 16937 14089 17035 14187 ne
rect 17035 14089 17389 14187
tri 17389 14089 17487 14187 sw
tri 17487 14089 17585 14187 ne
rect 17585 14089 17939 14187
tri 17939 14089 18037 14187 sw
tri 18037 14089 18135 14187 ne
rect 18135 14089 18489 14187
tri 18489 14089 18587 14187 sw
tri 18587 14089 18685 14187 ne
rect 18685 14089 19039 14187
tri 19039 14089 19137 14187 sw
tri 19137 14089 19235 14187 ne
rect 19235 14089 19589 14187
tri 19589 14089 19687 14187 sw
rect 20800 14089 21800 14737
rect -2000 14085 437 14089
rect -2000 13965 215 14085
rect 335 13991 437 14085
tri 437 13991 535 14089 sw
tri 535 13991 633 14089 ne
rect 633 14085 987 14089
rect 633 13991 765 14085
rect 335 13965 535 13991
rect -2000 13961 535 13965
rect -2000 13313 -1000 13961
tri 113 13863 211 13961 ne
rect 211 13913 535 13961
tri 535 13913 613 13991 sw
tri 633 13913 711 13991 ne
rect 711 13965 765 13991
rect 885 13991 987 14085
tri 987 13991 1085 14089 sw
tri 1085 13991 1183 14089 ne
rect 1183 14085 1537 14089
rect 1183 13991 1315 14085
rect 885 13965 1085 13991
rect 711 13913 1085 13965
tri 1085 13913 1163 13991 sw
tri 1183 13913 1261 13991 ne
rect 1261 13965 1315 13991
rect 1435 13991 1537 14085
tri 1537 13991 1635 14089 sw
tri 1635 13991 1733 14089 ne
rect 1733 14085 2087 14089
rect 1733 13991 1865 14085
rect 1435 13965 1635 13991
rect 1261 13913 1635 13965
tri 1635 13913 1713 13991 sw
tri 1733 13913 1811 13991 ne
rect 1811 13965 1865 13991
rect 1985 13991 2087 14085
tri 2087 13991 2185 14089 sw
tri 2185 13991 2283 14089 ne
rect 2283 14085 2637 14089
rect 2283 13991 2415 14085
rect 1985 13965 2185 13991
rect 1811 13913 2185 13965
tri 2185 13913 2263 13991 sw
tri 2283 13913 2361 13991 ne
rect 2361 13965 2415 13991
rect 2535 13991 2637 14085
tri 2637 13991 2735 14089 sw
tri 2735 13991 2833 14089 ne
rect 2833 14085 3187 14089
rect 2833 13991 2965 14085
rect 2535 13965 2735 13991
rect 2361 13913 2735 13965
tri 2735 13913 2813 13991 sw
tri 2833 13913 2911 13991 ne
rect 2911 13965 2965 13991
rect 3085 13991 3187 14085
tri 3187 13991 3285 14089 sw
tri 3285 13991 3383 14089 ne
rect 3383 14085 3737 14089
rect 3383 13991 3515 14085
rect 3085 13965 3285 13991
rect 2911 13913 3285 13965
tri 3285 13913 3363 13991 sw
tri 3383 13913 3461 13991 ne
rect 3461 13965 3515 13991
rect 3635 13991 3737 14085
tri 3737 13991 3835 14089 sw
tri 3835 13991 3933 14089 ne
rect 3933 14085 4287 14089
rect 3933 13991 4065 14085
rect 3635 13965 3835 13991
rect 3461 13913 3835 13965
tri 3835 13913 3913 13991 sw
tri 3933 13913 4011 13991 ne
rect 4011 13965 4065 13991
rect 4185 13991 4287 14085
tri 4287 13991 4385 14089 sw
tri 4385 13991 4483 14089 ne
rect 4483 14085 4837 14089
rect 4483 13991 4615 14085
rect 4185 13965 4385 13991
rect 4011 13913 4385 13965
tri 4385 13913 4463 13991 sw
tri 4483 13913 4561 13991 ne
rect 4561 13965 4615 13991
rect 4735 13991 4837 14085
tri 4837 13991 4935 14089 sw
tri 4935 13991 5033 14089 ne
rect 5033 14085 5387 14089
rect 5033 13991 5165 14085
rect 4735 13965 4935 13991
rect 4561 13913 4935 13965
tri 4935 13913 5013 13991 sw
tri 5033 13913 5111 13991 ne
rect 5111 13965 5165 13991
rect 5285 13991 5387 14085
tri 5387 13991 5485 14089 sw
tri 5485 13991 5583 14089 ne
rect 5583 14085 5937 14089
rect 5583 13991 5715 14085
rect 5285 13965 5485 13991
rect 5111 13913 5485 13965
tri 5485 13913 5563 13991 sw
tri 5583 13913 5661 13991 ne
rect 5661 13965 5715 13991
rect 5835 13991 5937 14085
tri 5937 13991 6035 14089 sw
tri 6035 13991 6133 14089 ne
rect 6133 14085 6487 14089
rect 6133 13991 6265 14085
rect 5835 13965 6035 13991
rect 5661 13913 6035 13965
tri 6035 13913 6113 13991 sw
tri 6133 13913 6211 13991 ne
rect 6211 13965 6265 13991
rect 6385 13991 6487 14085
tri 6487 13991 6585 14089 sw
tri 6585 13991 6683 14089 ne
rect 6683 14085 7037 14089
rect 6683 13991 6815 14085
rect 6385 13965 6585 13991
rect 6211 13913 6585 13965
tri 6585 13913 6663 13991 sw
tri 6683 13913 6761 13991 ne
rect 6761 13965 6815 13991
rect 6935 13991 7037 14085
tri 7037 13991 7135 14089 sw
tri 7135 13991 7233 14089 ne
rect 7233 14085 7587 14089
rect 7233 13991 7365 14085
rect 6935 13965 7135 13991
rect 6761 13913 7135 13965
tri 7135 13913 7213 13991 sw
tri 7233 13913 7311 13991 ne
rect 7311 13965 7365 13991
rect 7485 13991 7587 14085
tri 7587 13991 7685 14089 sw
tri 7685 13991 7783 14089 ne
rect 7783 14085 8137 14089
rect 7783 13991 7915 14085
rect 7485 13965 7685 13991
rect 7311 13913 7685 13965
tri 7685 13913 7763 13991 sw
tri 7783 13913 7861 13991 ne
rect 7861 13965 7915 13991
rect 8035 13991 8137 14085
tri 8137 13991 8235 14089 sw
tri 8235 13991 8333 14089 ne
rect 8333 14085 8687 14089
rect 8333 13991 8465 14085
rect 8035 13965 8235 13991
rect 7861 13913 8235 13965
tri 8235 13913 8313 13991 sw
tri 8333 13913 8411 13991 ne
rect 8411 13965 8465 13991
rect 8585 13991 8687 14085
tri 8687 13991 8785 14089 sw
tri 8785 13991 8883 14089 ne
rect 8883 14085 9237 14089
rect 8883 13991 9015 14085
rect 8585 13965 8785 13991
rect 8411 13913 8785 13965
tri 8785 13913 8863 13991 sw
tri 8883 13913 8961 13991 ne
rect 8961 13965 9015 13991
rect 9135 13991 9237 14085
tri 9237 13991 9335 14089 sw
tri 9335 13991 9433 14089 ne
rect 9433 14085 9787 14089
rect 9433 13991 9565 14085
rect 9135 13965 9335 13991
rect 8961 13913 9335 13965
tri 9335 13913 9413 13991 sw
tri 9433 13913 9511 13991 ne
rect 9511 13965 9565 13991
rect 9685 13991 9787 14085
tri 9787 13991 9885 14089 sw
tri 9885 13991 9983 14089 ne
rect 9983 14085 10337 14089
rect 9983 13991 10115 14085
rect 9685 13965 9885 13991
rect 9511 13913 9885 13965
tri 9885 13913 9963 13991 sw
tri 9983 13913 10061 13991 ne
rect 10061 13965 10115 13991
rect 10235 13991 10337 14085
tri 10337 13991 10435 14089 sw
tri 10435 13991 10533 14089 ne
rect 10533 14085 10887 14089
rect 10533 13991 10665 14085
rect 10235 13965 10435 13991
rect 10061 13913 10435 13965
tri 10435 13913 10513 13991 sw
tri 10533 13913 10611 13991 ne
rect 10611 13965 10665 13991
rect 10785 13991 10887 14085
tri 10887 13991 10985 14089 sw
tri 10985 13991 11083 14089 ne
rect 11083 14085 11437 14089
rect 11083 13991 11215 14085
rect 10785 13965 10985 13991
rect 10611 13913 10985 13965
tri 10985 13913 11063 13991 sw
tri 11083 13913 11161 13991 ne
rect 11161 13965 11215 13991
rect 11335 13991 11437 14085
tri 11437 13991 11535 14089 sw
tri 11535 13991 11633 14089 ne
rect 11633 14085 11987 14089
rect 11633 13991 11765 14085
rect 11335 13965 11535 13991
rect 11161 13913 11535 13965
tri 11535 13913 11613 13991 sw
tri 11633 13913 11711 13991 ne
rect 11711 13965 11765 13991
rect 11885 13991 11987 14085
tri 11987 13991 12085 14089 sw
tri 12085 13991 12183 14089 ne
rect 12183 14085 12537 14089
rect 12183 13991 12315 14085
rect 11885 13965 12085 13991
rect 11711 13913 12085 13965
tri 12085 13913 12163 13991 sw
tri 12183 13913 12261 13991 ne
rect 12261 13965 12315 13991
rect 12435 13991 12537 14085
tri 12537 13991 12635 14089 sw
tri 12635 13991 12733 14089 ne
rect 12733 14085 13087 14089
rect 12733 13991 12865 14085
rect 12435 13965 12635 13991
rect 12261 13913 12635 13965
tri 12635 13913 12713 13991 sw
tri 12733 13913 12811 13991 ne
rect 12811 13965 12865 13991
rect 12985 13991 13087 14085
tri 13087 13991 13185 14089 sw
tri 13185 13991 13283 14089 ne
rect 13283 14085 13637 14089
rect 13283 13991 13415 14085
rect 12985 13965 13185 13991
rect 12811 13913 13185 13965
tri 13185 13913 13263 13991 sw
tri 13283 13913 13361 13991 ne
rect 13361 13965 13415 13991
rect 13535 13991 13637 14085
tri 13637 13991 13735 14089 sw
tri 13735 13991 13833 14089 ne
rect 13833 14085 14187 14089
rect 13833 13991 13965 14085
rect 13535 13965 13735 13991
rect 13361 13913 13735 13965
tri 13735 13913 13813 13991 sw
tri 13833 13913 13911 13991 ne
rect 13911 13965 13965 13991
rect 14085 13991 14187 14085
tri 14187 13991 14285 14089 sw
tri 14285 13991 14383 14089 ne
rect 14383 14085 14737 14089
rect 14383 13991 14515 14085
rect 14085 13965 14285 13991
rect 13911 13913 14285 13965
tri 14285 13913 14363 13991 sw
tri 14383 13913 14461 13991 ne
rect 14461 13965 14515 13991
rect 14635 13991 14737 14085
tri 14737 13991 14835 14089 sw
tri 14835 13991 14933 14089 ne
rect 14933 14085 15287 14089
rect 14933 13991 15065 14085
rect 14635 13965 14835 13991
rect 14461 13913 14835 13965
tri 14835 13913 14913 13991 sw
tri 14933 13913 15011 13991 ne
rect 15011 13965 15065 13991
rect 15185 13991 15287 14085
tri 15287 13991 15385 14089 sw
tri 15385 13991 15483 14089 ne
rect 15483 14085 15837 14089
rect 15483 13991 15615 14085
rect 15185 13965 15385 13991
rect 15011 13913 15385 13965
tri 15385 13913 15463 13991 sw
tri 15483 13913 15561 13991 ne
rect 15561 13965 15615 13991
rect 15735 13991 15837 14085
tri 15837 13991 15935 14089 sw
tri 15935 13991 16033 14089 ne
rect 16033 14085 16387 14089
rect 16033 13991 16165 14085
rect 15735 13965 15935 13991
rect 15561 13913 15935 13965
tri 15935 13913 16013 13991 sw
tri 16033 13913 16111 13991 ne
rect 16111 13965 16165 13991
rect 16285 13991 16387 14085
tri 16387 13991 16485 14089 sw
tri 16485 13991 16583 14089 ne
rect 16583 14085 16937 14089
rect 16583 13991 16715 14085
rect 16285 13965 16485 13991
rect 16111 13913 16485 13965
tri 16485 13913 16563 13991 sw
tri 16583 13913 16661 13991 ne
rect 16661 13965 16715 13991
rect 16835 13991 16937 14085
tri 16937 13991 17035 14089 sw
tri 17035 13991 17133 14089 ne
rect 17133 14085 17487 14089
rect 17133 13991 17265 14085
rect 16835 13965 17035 13991
rect 16661 13913 17035 13965
tri 17035 13913 17113 13991 sw
tri 17133 13913 17211 13991 ne
rect 17211 13965 17265 13991
rect 17385 13991 17487 14085
tri 17487 13991 17585 14089 sw
tri 17585 13991 17683 14089 ne
rect 17683 14085 18037 14089
rect 17683 13991 17815 14085
rect 17385 13965 17585 13991
rect 17211 13913 17585 13965
tri 17585 13913 17663 13991 sw
tri 17683 13913 17761 13991 ne
rect 17761 13965 17815 13991
rect 17935 13991 18037 14085
tri 18037 13991 18135 14089 sw
tri 18135 13991 18233 14089 ne
rect 18233 14085 18587 14089
rect 18233 13991 18365 14085
rect 17935 13965 18135 13991
rect 17761 13913 18135 13965
tri 18135 13913 18213 13991 sw
tri 18233 13913 18311 13991 ne
rect 18311 13965 18365 13991
rect 18485 13991 18587 14085
tri 18587 13991 18685 14089 sw
tri 18685 13991 18783 14089 ne
rect 18783 14085 19137 14089
rect 18783 13991 18915 14085
rect 18485 13965 18685 13991
rect 18311 13913 18685 13965
tri 18685 13913 18763 13991 sw
tri 18783 13913 18861 13991 ne
rect 18861 13965 18915 13991
rect 19035 13991 19137 14085
tri 19137 13991 19235 14089 sw
tri 19235 13991 19333 14089 ne
rect 19333 14085 21800 14089
rect 19333 13991 19465 14085
rect 19035 13965 19235 13991
rect 18861 13913 19235 13965
tri 19235 13913 19313 13991 sw
tri 19333 13913 19411 13991 ne
rect 19411 13965 19465 13991
rect 19585 13965 21800 14085
rect 19411 13913 21800 13965
rect 211 13863 613 13913
rect -500 13813 113 13863
tri 113 13813 163 13863 sw
tri 211 13813 261 13863 ne
rect 261 13833 613 13863
tri 613 13833 693 13913 sw
tri 711 13833 791 13913 ne
rect 791 13833 1163 13913
tri 1163 13833 1243 13913 sw
tri 1261 13833 1341 13913 ne
rect 1341 13833 1713 13913
tri 1713 13833 1793 13913 sw
tri 1811 13833 1891 13913 ne
rect 1891 13833 2263 13913
tri 2263 13833 2343 13913 sw
tri 2361 13833 2441 13913 ne
rect 2441 13833 2813 13913
tri 2813 13833 2893 13913 sw
tri 2911 13833 2991 13913 ne
rect 2991 13833 3363 13913
tri 3363 13833 3443 13913 sw
tri 3461 13833 3541 13913 ne
rect 3541 13833 3913 13913
tri 3913 13833 3993 13913 sw
tri 4011 13833 4091 13913 ne
rect 4091 13833 4463 13913
tri 4463 13833 4543 13913 sw
tri 4561 13833 4641 13913 ne
rect 4641 13833 5013 13913
tri 5013 13833 5093 13913 sw
tri 5111 13833 5191 13913 ne
rect 5191 13833 5563 13913
tri 5563 13833 5643 13913 sw
tri 5661 13833 5741 13913 ne
rect 5741 13833 6113 13913
tri 6113 13833 6193 13913 sw
tri 6211 13833 6291 13913 ne
rect 6291 13833 6663 13913
tri 6663 13833 6743 13913 sw
tri 6761 13833 6841 13913 ne
rect 6841 13833 7213 13913
tri 7213 13833 7293 13913 sw
tri 7311 13833 7391 13913 ne
rect 7391 13833 7763 13913
tri 7763 13833 7843 13913 sw
tri 7861 13833 7941 13913 ne
rect 7941 13833 8313 13913
tri 8313 13833 8393 13913 sw
tri 8411 13833 8491 13913 ne
rect 8491 13833 8863 13913
tri 8863 13833 8943 13913 sw
tri 8961 13833 9041 13913 ne
rect 9041 13833 9413 13913
tri 9413 13833 9493 13913 sw
tri 9511 13833 9591 13913 ne
rect 9591 13833 9963 13913
tri 9963 13833 10043 13913 sw
tri 10061 13833 10141 13913 ne
rect 10141 13833 10513 13913
tri 10513 13833 10593 13913 sw
tri 10611 13833 10691 13913 ne
rect 10691 13833 11063 13913
tri 11063 13833 11143 13913 sw
tri 11161 13833 11241 13913 ne
rect 11241 13833 11613 13913
tri 11613 13833 11693 13913 sw
tri 11711 13833 11791 13913 ne
rect 11791 13833 12163 13913
tri 12163 13833 12243 13913 sw
tri 12261 13833 12341 13913 ne
rect 12341 13833 12713 13913
tri 12713 13833 12793 13913 sw
tri 12811 13833 12891 13913 ne
rect 12891 13833 13263 13913
tri 13263 13833 13343 13913 sw
tri 13361 13833 13441 13913 ne
rect 13441 13833 13813 13913
tri 13813 13833 13893 13913 sw
tri 13911 13833 13991 13913 ne
rect 13991 13833 14363 13913
tri 14363 13833 14443 13913 sw
tri 14461 13833 14541 13913 ne
rect 14541 13833 14913 13913
tri 14913 13833 14993 13913 sw
tri 15011 13833 15091 13913 ne
rect 15091 13833 15463 13913
tri 15463 13833 15543 13913 sw
tri 15561 13833 15641 13913 ne
rect 15641 13833 16013 13913
tri 16013 13833 16093 13913 sw
tri 16111 13833 16191 13913 ne
rect 16191 13833 16563 13913
tri 16563 13833 16643 13913 sw
tri 16661 13833 16741 13913 ne
rect 16741 13833 17113 13913
tri 17113 13833 17193 13913 sw
tri 17211 13833 17291 13913 ne
rect 17291 13833 17663 13913
tri 17663 13833 17743 13913 sw
tri 17761 13833 17841 13913 ne
rect 17841 13833 18213 13913
tri 18213 13833 18293 13913 sw
tri 18311 13833 18391 13913 ne
rect 18391 13833 18763 13913
tri 18763 13833 18843 13913 sw
tri 18861 13833 18941 13913 ne
rect 18941 13833 19313 13913
tri 19313 13833 19393 13913 sw
tri 19411 13833 19491 13913 ne
rect 19491 13833 20100 13913
rect 261 13813 693 13833
rect -500 13735 163 13813
tri 163 13735 241 13813 sw
tri 261 13735 339 13813 ne
rect 339 13735 693 13813
tri 693 13735 791 13833 sw
tri 791 13735 889 13833 ne
rect 889 13735 1243 13833
tri 1243 13735 1341 13833 sw
tri 1341 13735 1439 13833 ne
rect 1439 13735 1793 13833
tri 1793 13735 1891 13833 sw
tri 1891 13735 1989 13833 ne
rect 1989 13735 2343 13833
tri 2343 13735 2441 13833 sw
tri 2441 13735 2539 13833 ne
rect 2539 13735 2893 13833
tri 2893 13735 2991 13833 sw
tri 2991 13735 3089 13833 ne
rect 3089 13735 3443 13833
tri 3443 13735 3541 13833 sw
tri 3541 13735 3639 13833 ne
rect 3639 13735 3993 13833
tri 3993 13735 4091 13833 sw
tri 4091 13735 4189 13833 ne
rect 4189 13735 4543 13833
tri 4543 13735 4641 13833 sw
tri 4641 13735 4739 13833 ne
rect 4739 13735 5093 13833
tri 5093 13735 5191 13833 sw
tri 5191 13735 5289 13833 ne
rect 5289 13735 5643 13833
tri 5643 13735 5741 13833 sw
tri 5741 13735 5839 13833 ne
rect 5839 13735 6193 13833
tri 6193 13735 6291 13833 sw
tri 6291 13735 6389 13833 ne
rect 6389 13735 6743 13833
tri 6743 13735 6841 13833 sw
tri 6841 13735 6939 13833 ne
rect 6939 13735 7293 13833
tri 7293 13735 7391 13833 sw
tri 7391 13735 7489 13833 ne
rect 7489 13735 7843 13833
tri 7843 13735 7941 13833 sw
tri 7941 13735 8039 13833 ne
rect 8039 13735 8393 13833
tri 8393 13735 8491 13833 sw
tri 8491 13735 8589 13833 ne
rect 8589 13735 8943 13833
tri 8943 13735 9041 13833 sw
tri 9041 13735 9139 13833 ne
rect 9139 13735 9493 13833
tri 9493 13735 9591 13833 sw
tri 9591 13735 9689 13833 ne
rect 9689 13735 10043 13833
tri 10043 13735 10141 13833 sw
tri 10141 13735 10239 13833 ne
rect 10239 13735 10593 13833
tri 10593 13735 10691 13833 sw
tri 10691 13735 10789 13833 ne
rect 10789 13735 11143 13833
tri 11143 13735 11241 13833 sw
tri 11241 13735 11339 13833 ne
rect 11339 13735 11693 13833
tri 11693 13735 11791 13833 sw
tri 11791 13735 11889 13833 ne
rect 11889 13735 12243 13833
tri 12243 13735 12341 13833 sw
tri 12341 13735 12439 13833 ne
rect 12439 13735 12793 13833
tri 12793 13735 12891 13833 sw
tri 12891 13735 12989 13833 ne
rect 12989 13735 13343 13833
tri 13343 13735 13441 13833 sw
tri 13441 13735 13539 13833 ne
rect 13539 13735 13893 13833
tri 13893 13735 13991 13833 sw
tri 13991 13735 14089 13833 ne
rect 14089 13735 14443 13833
tri 14443 13735 14541 13833 sw
tri 14541 13735 14639 13833 ne
rect 14639 13735 14993 13833
tri 14993 13735 15091 13833 sw
tri 15091 13735 15189 13833 ne
rect 15189 13735 15543 13833
tri 15543 13735 15641 13833 sw
tri 15641 13735 15739 13833 ne
rect 15739 13735 16093 13833
tri 16093 13735 16191 13833 sw
tri 16191 13735 16289 13833 ne
rect 16289 13735 16643 13833
tri 16643 13735 16741 13833 sw
tri 16741 13735 16839 13833 ne
rect 16839 13735 17193 13833
tri 17193 13735 17291 13833 sw
tri 17291 13735 17389 13833 ne
rect 17389 13735 17743 13833
tri 17743 13735 17841 13833 sw
tri 17841 13735 17939 13833 ne
rect 17939 13735 18293 13833
tri 18293 13735 18391 13833 sw
tri 18391 13735 18489 13833 ne
rect 18489 13735 18843 13833
tri 18843 13735 18941 13833 sw
tri 18941 13735 19039 13833 ne
rect 19039 13735 19393 13833
tri 19393 13735 19491 13833 sw
tri 19491 13735 19589 13833 ne
rect 19589 13813 20100 13833
rect 20200 13813 21800 13913
rect 19589 13735 21800 13813
rect -500 13687 241 13735
rect -500 13587 -400 13687
rect -300 13637 241 13687
tri 241 13637 339 13735 sw
tri 339 13637 437 13735 ne
rect 437 13637 791 13735
tri 791 13637 889 13735 sw
tri 889 13637 987 13735 ne
rect 987 13637 1341 13735
tri 1341 13637 1439 13735 sw
tri 1439 13637 1537 13735 ne
rect 1537 13637 1891 13735
tri 1891 13637 1989 13735 sw
tri 1989 13637 2087 13735 ne
rect 2087 13637 2441 13735
tri 2441 13637 2539 13735 sw
tri 2539 13637 2637 13735 ne
rect 2637 13637 2991 13735
tri 2991 13637 3089 13735 sw
tri 3089 13637 3187 13735 ne
rect 3187 13637 3541 13735
tri 3541 13637 3639 13735 sw
tri 3639 13637 3737 13735 ne
rect 3737 13637 4091 13735
tri 4091 13637 4189 13735 sw
tri 4189 13637 4287 13735 ne
rect 4287 13637 4641 13735
tri 4641 13637 4739 13735 sw
tri 4739 13637 4837 13735 ne
rect 4837 13637 5191 13735
tri 5191 13637 5289 13735 sw
tri 5289 13637 5387 13735 ne
rect 5387 13637 5741 13735
tri 5741 13637 5839 13735 sw
tri 5839 13637 5937 13735 ne
rect 5937 13637 6291 13735
tri 6291 13637 6389 13735 sw
tri 6389 13637 6487 13735 ne
rect 6487 13637 6841 13735
tri 6841 13637 6939 13735 sw
tri 6939 13637 7037 13735 ne
rect 7037 13637 7391 13735
tri 7391 13637 7489 13735 sw
tri 7489 13637 7587 13735 ne
rect 7587 13637 7941 13735
tri 7941 13637 8039 13735 sw
tri 8039 13637 8137 13735 ne
rect 8137 13637 8491 13735
tri 8491 13637 8589 13735 sw
tri 8589 13637 8687 13735 ne
rect 8687 13637 9041 13735
tri 9041 13637 9139 13735 sw
tri 9139 13637 9237 13735 ne
rect 9237 13637 9591 13735
tri 9591 13637 9689 13735 sw
tri 9689 13637 9787 13735 ne
rect 9787 13637 10141 13735
tri 10141 13637 10239 13735 sw
tri 10239 13637 10337 13735 ne
rect 10337 13637 10691 13735
tri 10691 13637 10789 13735 sw
tri 10789 13637 10887 13735 ne
rect 10887 13637 11241 13735
tri 11241 13637 11339 13735 sw
tri 11339 13637 11437 13735 ne
rect 11437 13637 11791 13735
tri 11791 13637 11889 13735 sw
tri 11889 13637 11987 13735 ne
rect 11987 13637 12341 13735
tri 12341 13637 12439 13735 sw
tri 12439 13637 12537 13735 ne
rect 12537 13637 12891 13735
tri 12891 13637 12989 13735 sw
tri 12989 13637 13087 13735 ne
rect 13087 13637 13441 13735
tri 13441 13637 13539 13735 sw
tri 13539 13637 13637 13735 ne
rect 13637 13637 13991 13735
tri 13991 13637 14089 13735 sw
tri 14089 13637 14187 13735 ne
rect 14187 13637 14541 13735
tri 14541 13637 14639 13735 sw
tri 14639 13637 14737 13735 ne
rect 14737 13637 15091 13735
tri 15091 13637 15189 13735 sw
tri 15189 13637 15287 13735 ne
rect 15287 13637 15641 13735
tri 15641 13637 15739 13735 sw
tri 15739 13637 15837 13735 ne
rect 15837 13637 16191 13735
tri 16191 13637 16289 13735 sw
tri 16289 13637 16387 13735 ne
rect 16387 13637 16741 13735
tri 16741 13637 16839 13735 sw
tri 16839 13637 16937 13735 ne
rect 16937 13637 17291 13735
tri 17291 13637 17389 13735 sw
tri 17389 13637 17487 13735 ne
rect 17487 13637 17841 13735
tri 17841 13637 17939 13735 sw
tri 17939 13637 18037 13735 ne
rect 18037 13637 18391 13735
tri 18391 13637 18489 13735 sw
tri 18489 13637 18587 13735 ne
rect 18587 13637 18941 13735
tri 18941 13637 19039 13735 sw
tri 19039 13637 19137 13735 ne
rect 19137 13637 19491 13735
tri 19491 13637 19589 13735 sw
tri 19589 13637 19687 13735 ne
rect 19687 13637 21800 13735
rect -300 13587 339 13637
rect -500 13539 339 13587
tri 339 13539 437 13637 sw
tri 437 13539 535 13637 ne
rect 535 13539 889 13637
tri 889 13539 987 13637 sw
tri 987 13539 1085 13637 ne
rect 1085 13539 1439 13637
tri 1439 13539 1537 13637 sw
tri 1537 13539 1635 13637 ne
rect 1635 13539 1989 13637
tri 1989 13539 2087 13637 sw
tri 2087 13539 2185 13637 ne
rect 2185 13539 2539 13637
tri 2539 13539 2637 13637 sw
tri 2637 13539 2735 13637 ne
rect 2735 13539 3089 13637
tri 3089 13539 3187 13637 sw
tri 3187 13539 3285 13637 ne
rect 3285 13539 3639 13637
tri 3639 13539 3737 13637 sw
tri 3737 13539 3835 13637 ne
rect 3835 13539 4189 13637
tri 4189 13539 4287 13637 sw
tri 4287 13539 4385 13637 ne
rect 4385 13539 4739 13637
tri 4739 13539 4837 13637 sw
tri 4837 13539 4935 13637 ne
rect 4935 13539 5289 13637
tri 5289 13539 5387 13637 sw
tri 5387 13539 5485 13637 ne
rect 5485 13539 5839 13637
tri 5839 13539 5937 13637 sw
tri 5937 13539 6035 13637 ne
rect 6035 13539 6389 13637
tri 6389 13539 6487 13637 sw
tri 6487 13539 6585 13637 ne
rect 6585 13539 6939 13637
tri 6939 13539 7037 13637 sw
tri 7037 13539 7135 13637 ne
rect 7135 13539 7489 13637
tri 7489 13539 7587 13637 sw
tri 7587 13539 7685 13637 ne
rect 7685 13539 8039 13637
tri 8039 13539 8137 13637 sw
tri 8137 13539 8235 13637 ne
rect 8235 13539 8589 13637
tri 8589 13539 8687 13637 sw
tri 8687 13539 8785 13637 ne
rect 8785 13539 9139 13637
tri 9139 13539 9237 13637 sw
tri 9237 13539 9335 13637 ne
rect 9335 13539 9689 13637
tri 9689 13539 9787 13637 sw
tri 9787 13539 9885 13637 ne
rect 9885 13539 10239 13637
tri 10239 13539 10337 13637 sw
tri 10337 13539 10435 13637 ne
rect 10435 13539 10789 13637
tri 10789 13539 10887 13637 sw
tri 10887 13539 10985 13637 ne
rect 10985 13539 11339 13637
tri 11339 13539 11437 13637 sw
tri 11437 13539 11535 13637 ne
rect 11535 13539 11889 13637
tri 11889 13539 11987 13637 sw
tri 11987 13539 12085 13637 ne
rect 12085 13539 12439 13637
tri 12439 13539 12537 13637 sw
tri 12537 13539 12635 13637 ne
rect 12635 13539 12989 13637
tri 12989 13539 13087 13637 sw
tri 13087 13539 13185 13637 ne
rect 13185 13539 13539 13637
tri 13539 13539 13637 13637 sw
tri 13637 13539 13735 13637 ne
rect 13735 13539 14089 13637
tri 14089 13539 14187 13637 sw
tri 14187 13539 14285 13637 ne
rect 14285 13539 14639 13637
tri 14639 13539 14737 13637 sw
tri 14737 13539 14835 13637 ne
rect 14835 13539 15189 13637
tri 15189 13539 15287 13637 sw
tri 15287 13539 15385 13637 ne
rect 15385 13539 15739 13637
tri 15739 13539 15837 13637 sw
tri 15837 13539 15935 13637 ne
rect 15935 13539 16289 13637
tri 16289 13539 16387 13637 sw
tri 16387 13539 16485 13637 ne
rect 16485 13539 16839 13637
tri 16839 13539 16937 13637 sw
tri 16937 13539 17035 13637 ne
rect 17035 13539 17389 13637
tri 17389 13539 17487 13637 sw
tri 17487 13539 17585 13637 ne
rect 17585 13539 17939 13637
tri 17939 13539 18037 13637 sw
tri 18037 13539 18135 13637 ne
rect 18135 13539 18489 13637
tri 18489 13539 18587 13637 sw
tri 18587 13539 18685 13637 ne
rect 18685 13539 19039 13637
tri 19039 13539 19137 13637 sw
tri 19137 13539 19235 13637 ne
rect 19235 13539 19589 13637
tri 19589 13539 19687 13637 sw
rect -500 13535 437 13539
rect -500 13415 215 13535
rect 335 13441 437 13535
tri 437 13441 535 13539 sw
tri 535 13441 633 13539 ne
rect 633 13535 987 13539
rect 633 13441 765 13535
rect 335 13415 535 13441
rect -500 13411 535 13415
tri 535 13411 565 13441 sw
tri 633 13411 663 13441 ne
rect 663 13415 765 13441
rect 885 13441 987 13535
tri 987 13441 1085 13539 sw
tri 1085 13441 1183 13539 ne
rect 1183 13535 1537 13539
rect 1183 13441 1315 13535
rect 885 13415 1085 13441
rect 663 13411 1085 13415
tri 1085 13411 1115 13441 sw
tri 1183 13411 1213 13441 ne
rect 1213 13415 1315 13441
rect 1435 13441 1537 13535
tri 1537 13441 1635 13539 sw
tri 1635 13441 1733 13539 ne
rect 1733 13535 2087 13539
rect 1733 13441 1865 13535
rect 1435 13415 1635 13441
rect 1213 13411 1635 13415
tri 1635 13411 1665 13441 sw
tri 1733 13411 1763 13441 ne
rect 1763 13415 1865 13441
rect 1985 13441 2087 13535
tri 2087 13441 2185 13539 sw
tri 2185 13441 2283 13539 ne
rect 2283 13535 2637 13539
rect 2283 13441 2415 13535
rect 1985 13415 2185 13441
rect 1763 13411 2185 13415
tri 2185 13411 2215 13441 sw
tri 2283 13411 2313 13441 ne
rect 2313 13415 2415 13441
rect 2535 13441 2637 13535
tri 2637 13441 2735 13539 sw
tri 2735 13441 2833 13539 ne
rect 2833 13535 3187 13539
rect 2833 13441 2965 13535
rect 2535 13415 2735 13441
rect 2313 13411 2735 13415
tri 2735 13411 2765 13441 sw
tri 2833 13411 2863 13441 ne
rect 2863 13415 2965 13441
rect 3085 13441 3187 13535
tri 3187 13441 3285 13539 sw
tri 3285 13441 3383 13539 ne
rect 3383 13535 3737 13539
rect 3383 13441 3515 13535
rect 3085 13415 3285 13441
rect 2863 13411 3285 13415
tri 3285 13411 3315 13441 sw
tri 3383 13411 3413 13441 ne
rect 3413 13415 3515 13441
rect 3635 13441 3737 13535
tri 3737 13441 3835 13539 sw
tri 3835 13441 3933 13539 ne
rect 3933 13535 4287 13539
rect 3933 13441 4065 13535
rect 3635 13415 3835 13441
rect 3413 13411 3835 13415
tri 3835 13411 3865 13441 sw
tri 3933 13411 3963 13441 ne
rect 3963 13415 4065 13441
rect 4185 13441 4287 13535
tri 4287 13441 4385 13539 sw
tri 4385 13441 4483 13539 ne
rect 4483 13535 4837 13539
rect 4483 13441 4615 13535
rect 4185 13415 4385 13441
rect 3963 13411 4385 13415
tri 4385 13411 4415 13441 sw
tri 4483 13411 4513 13441 ne
rect 4513 13415 4615 13441
rect 4735 13441 4837 13535
tri 4837 13441 4935 13539 sw
tri 4935 13441 5033 13539 ne
rect 5033 13535 5387 13539
rect 5033 13441 5165 13535
rect 4735 13415 4935 13441
rect 4513 13411 4935 13415
tri 4935 13411 4965 13441 sw
tri 5033 13411 5063 13441 ne
rect 5063 13415 5165 13441
rect 5285 13441 5387 13535
tri 5387 13441 5485 13539 sw
tri 5485 13441 5583 13539 ne
rect 5583 13535 5937 13539
rect 5583 13441 5715 13535
rect 5285 13415 5485 13441
rect 5063 13411 5485 13415
tri 5485 13411 5515 13441 sw
tri 5583 13411 5613 13441 ne
rect 5613 13415 5715 13441
rect 5835 13441 5937 13535
tri 5937 13441 6035 13539 sw
tri 6035 13441 6133 13539 ne
rect 6133 13535 6487 13539
rect 6133 13441 6265 13535
rect 5835 13415 6035 13441
rect 5613 13411 6035 13415
tri 6035 13411 6065 13441 sw
tri 6133 13411 6163 13441 ne
rect 6163 13415 6265 13441
rect 6385 13441 6487 13535
tri 6487 13441 6585 13539 sw
tri 6585 13441 6683 13539 ne
rect 6683 13535 7037 13539
rect 6683 13441 6815 13535
rect 6385 13415 6585 13441
rect 6163 13411 6585 13415
tri 6585 13411 6615 13441 sw
tri 6683 13411 6713 13441 ne
rect 6713 13415 6815 13441
rect 6935 13441 7037 13535
tri 7037 13441 7135 13539 sw
tri 7135 13441 7233 13539 ne
rect 7233 13535 7587 13539
rect 7233 13441 7365 13535
rect 6935 13415 7135 13441
rect 6713 13411 7135 13415
tri 7135 13411 7165 13441 sw
tri 7233 13411 7263 13441 ne
rect 7263 13415 7365 13441
rect 7485 13441 7587 13535
tri 7587 13441 7685 13539 sw
tri 7685 13441 7783 13539 ne
rect 7783 13535 8137 13539
rect 7783 13441 7915 13535
rect 7485 13415 7685 13441
rect 7263 13411 7685 13415
tri 7685 13411 7715 13441 sw
tri 7783 13411 7813 13441 ne
rect 7813 13415 7915 13441
rect 8035 13441 8137 13535
tri 8137 13441 8235 13539 sw
tri 8235 13441 8333 13539 ne
rect 8333 13535 8687 13539
rect 8333 13441 8465 13535
rect 8035 13415 8235 13441
rect 7813 13411 8235 13415
tri 8235 13411 8265 13441 sw
tri 8333 13411 8363 13441 ne
rect 8363 13415 8465 13441
rect 8585 13441 8687 13535
tri 8687 13441 8785 13539 sw
tri 8785 13441 8883 13539 ne
rect 8883 13535 9237 13539
rect 8883 13441 9015 13535
rect 8585 13415 8785 13441
rect 8363 13411 8785 13415
tri 8785 13411 8815 13441 sw
tri 8883 13411 8913 13441 ne
rect 8913 13415 9015 13441
rect 9135 13441 9237 13535
tri 9237 13441 9335 13539 sw
tri 9335 13441 9433 13539 ne
rect 9433 13535 9787 13539
rect 9433 13441 9565 13535
rect 9135 13415 9335 13441
rect 8913 13411 9335 13415
tri 9335 13411 9365 13441 sw
tri 9433 13411 9463 13441 ne
rect 9463 13415 9565 13441
rect 9685 13441 9787 13535
tri 9787 13441 9885 13539 sw
tri 9885 13441 9983 13539 ne
rect 9983 13535 10337 13539
rect 9983 13441 10115 13535
rect 9685 13415 9885 13441
rect 9463 13411 9885 13415
tri 9885 13411 9915 13441 sw
tri 9983 13411 10013 13441 ne
rect 10013 13415 10115 13441
rect 10235 13441 10337 13535
tri 10337 13441 10435 13539 sw
tri 10435 13441 10533 13539 ne
rect 10533 13535 10887 13539
rect 10533 13441 10665 13535
rect 10235 13415 10435 13441
rect 10013 13411 10435 13415
tri 10435 13411 10465 13441 sw
tri 10533 13411 10563 13441 ne
rect 10563 13415 10665 13441
rect 10785 13441 10887 13535
tri 10887 13441 10985 13539 sw
tri 10985 13441 11083 13539 ne
rect 11083 13535 11437 13539
rect 11083 13441 11215 13535
rect 10785 13415 10985 13441
rect 10563 13411 10985 13415
tri 10985 13411 11015 13441 sw
tri 11083 13411 11113 13441 ne
rect 11113 13415 11215 13441
rect 11335 13441 11437 13535
tri 11437 13441 11535 13539 sw
tri 11535 13441 11633 13539 ne
rect 11633 13535 11987 13539
rect 11633 13441 11765 13535
rect 11335 13415 11535 13441
rect 11113 13411 11535 13415
tri 11535 13411 11565 13441 sw
tri 11633 13411 11663 13441 ne
rect 11663 13415 11765 13441
rect 11885 13441 11987 13535
tri 11987 13441 12085 13539 sw
tri 12085 13441 12183 13539 ne
rect 12183 13535 12537 13539
rect 12183 13441 12315 13535
rect 11885 13415 12085 13441
rect 11663 13411 12085 13415
tri 12085 13411 12115 13441 sw
tri 12183 13411 12213 13441 ne
rect 12213 13415 12315 13441
rect 12435 13441 12537 13535
tri 12537 13441 12635 13539 sw
tri 12635 13441 12733 13539 ne
rect 12733 13535 13087 13539
rect 12733 13441 12865 13535
rect 12435 13415 12635 13441
rect 12213 13411 12635 13415
tri 12635 13411 12665 13441 sw
tri 12733 13411 12763 13441 ne
rect 12763 13415 12865 13441
rect 12985 13441 13087 13535
tri 13087 13441 13185 13539 sw
tri 13185 13441 13283 13539 ne
rect 13283 13535 13637 13539
rect 13283 13441 13415 13535
rect 12985 13415 13185 13441
rect 12763 13411 13185 13415
tri 13185 13411 13215 13441 sw
tri 13283 13411 13313 13441 ne
rect 13313 13415 13415 13441
rect 13535 13441 13637 13535
tri 13637 13441 13735 13539 sw
tri 13735 13441 13833 13539 ne
rect 13833 13535 14187 13539
rect 13833 13441 13965 13535
rect 13535 13415 13735 13441
rect 13313 13411 13735 13415
tri 13735 13411 13765 13441 sw
tri 13833 13411 13863 13441 ne
rect 13863 13415 13965 13441
rect 14085 13441 14187 13535
tri 14187 13441 14285 13539 sw
tri 14285 13441 14383 13539 ne
rect 14383 13535 14737 13539
rect 14383 13441 14515 13535
rect 14085 13415 14285 13441
rect 13863 13411 14285 13415
tri 14285 13411 14315 13441 sw
tri 14383 13411 14413 13441 ne
rect 14413 13415 14515 13441
rect 14635 13441 14737 13535
tri 14737 13441 14835 13539 sw
tri 14835 13441 14933 13539 ne
rect 14933 13535 15287 13539
rect 14933 13441 15065 13535
rect 14635 13415 14835 13441
rect 14413 13411 14835 13415
tri 14835 13411 14865 13441 sw
tri 14933 13411 14963 13441 ne
rect 14963 13415 15065 13441
rect 15185 13441 15287 13535
tri 15287 13441 15385 13539 sw
tri 15385 13441 15483 13539 ne
rect 15483 13535 15837 13539
rect 15483 13441 15615 13535
rect 15185 13415 15385 13441
rect 14963 13411 15385 13415
tri 15385 13411 15415 13441 sw
tri 15483 13411 15513 13441 ne
rect 15513 13415 15615 13441
rect 15735 13441 15837 13535
tri 15837 13441 15935 13539 sw
tri 15935 13441 16033 13539 ne
rect 16033 13535 16387 13539
rect 16033 13441 16165 13535
rect 15735 13415 15935 13441
rect 15513 13411 15935 13415
tri 15935 13411 15965 13441 sw
tri 16033 13411 16063 13441 ne
rect 16063 13415 16165 13441
rect 16285 13441 16387 13535
tri 16387 13441 16485 13539 sw
tri 16485 13441 16583 13539 ne
rect 16583 13535 16937 13539
rect 16583 13441 16715 13535
rect 16285 13415 16485 13441
rect 16063 13411 16485 13415
tri 16485 13411 16515 13441 sw
tri 16583 13411 16613 13441 ne
rect 16613 13415 16715 13441
rect 16835 13441 16937 13535
tri 16937 13441 17035 13539 sw
tri 17035 13441 17133 13539 ne
rect 17133 13535 17487 13539
rect 17133 13441 17265 13535
rect 16835 13415 17035 13441
rect 16613 13411 17035 13415
tri 17035 13411 17065 13441 sw
tri 17133 13411 17163 13441 ne
rect 17163 13415 17265 13441
rect 17385 13441 17487 13535
tri 17487 13441 17585 13539 sw
tri 17585 13441 17683 13539 ne
rect 17683 13535 18037 13539
rect 17683 13441 17815 13535
rect 17385 13415 17585 13441
rect 17163 13411 17585 13415
tri 17585 13411 17615 13441 sw
tri 17683 13411 17713 13441 ne
rect 17713 13415 17815 13441
rect 17935 13441 18037 13535
tri 18037 13441 18135 13539 sw
tri 18135 13441 18233 13539 ne
rect 18233 13535 18587 13539
rect 18233 13441 18365 13535
rect 17935 13415 18135 13441
rect 17713 13411 18135 13415
tri 18135 13411 18165 13441 sw
tri 18233 13411 18263 13441 ne
rect 18263 13415 18365 13441
rect 18485 13441 18587 13535
tri 18587 13441 18685 13539 sw
tri 18685 13441 18783 13539 ne
rect 18783 13535 19137 13539
rect 18783 13441 18915 13535
rect 18485 13415 18685 13441
rect 18263 13411 18685 13415
tri 18685 13411 18715 13441 sw
tri 18783 13411 18813 13441 ne
rect 18813 13415 18915 13441
rect 19035 13441 19137 13535
tri 19137 13441 19235 13539 sw
tri 19235 13441 19333 13539 ne
rect 19333 13535 20300 13539
rect 19333 13441 19465 13535
rect 19035 13415 19235 13441
rect 18813 13411 19235 13415
tri 19235 13411 19265 13441 sw
tri 19333 13411 19363 13441 ne
rect 19363 13415 19465 13441
rect 19585 13415 20300 13535
rect 19363 13411 20300 13415
tri 113 13313 211 13411 ne
rect 211 13313 565 13411
tri 565 13313 663 13411 sw
tri 663 13313 761 13411 ne
rect 761 13313 1115 13411
tri 1115 13313 1213 13411 sw
tri 1213 13313 1311 13411 ne
rect 1311 13313 1665 13411
tri 1665 13313 1763 13411 sw
tri 1763 13313 1861 13411 ne
rect 1861 13313 2215 13411
tri 2215 13313 2313 13411 sw
tri 2313 13313 2411 13411 ne
rect 2411 13313 2765 13411
tri 2765 13313 2863 13411 sw
tri 2863 13313 2961 13411 ne
rect 2961 13313 3315 13411
tri 3315 13313 3413 13411 sw
tri 3413 13313 3511 13411 ne
rect 3511 13313 3865 13411
tri 3865 13313 3963 13411 sw
tri 3963 13313 4061 13411 ne
rect 4061 13313 4415 13411
tri 4415 13313 4513 13411 sw
tri 4513 13313 4611 13411 ne
rect 4611 13313 4965 13411
tri 4965 13313 5063 13411 sw
tri 5063 13313 5161 13411 ne
rect 5161 13313 5515 13411
tri 5515 13313 5613 13411 sw
tri 5613 13313 5711 13411 ne
rect 5711 13313 6065 13411
tri 6065 13313 6163 13411 sw
tri 6163 13313 6261 13411 ne
rect 6261 13313 6615 13411
tri 6615 13313 6713 13411 sw
tri 6713 13313 6811 13411 ne
rect 6811 13313 7165 13411
tri 7165 13313 7263 13411 sw
tri 7263 13313 7361 13411 ne
rect 7361 13313 7715 13411
tri 7715 13313 7813 13411 sw
tri 7813 13313 7911 13411 ne
rect 7911 13313 8265 13411
tri 8265 13313 8363 13411 sw
tri 8363 13313 8461 13411 ne
rect 8461 13313 8815 13411
tri 8815 13313 8913 13411 sw
tri 8913 13313 9011 13411 ne
rect 9011 13313 9365 13411
tri 9365 13313 9463 13411 sw
tri 9463 13313 9561 13411 ne
rect 9561 13313 9915 13411
tri 9915 13313 10013 13411 sw
tri 10013 13313 10111 13411 ne
rect 10111 13313 10465 13411
tri 10465 13313 10563 13411 sw
tri 10563 13313 10661 13411 ne
rect 10661 13313 11015 13411
tri 11015 13313 11113 13411 sw
tri 11113 13313 11211 13411 ne
rect 11211 13313 11565 13411
tri 11565 13313 11663 13411 sw
tri 11663 13313 11761 13411 ne
rect 11761 13313 12115 13411
tri 12115 13313 12213 13411 sw
tri 12213 13313 12311 13411 ne
rect 12311 13313 12665 13411
tri 12665 13313 12763 13411 sw
tri 12763 13313 12861 13411 ne
rect 12861 13313 13215 13411
tri 13215 13313 13313 13411 sw
tri 13313 13313 13411 13411 ne
rect 13411 13313 13765 13411
tri 13765 13313 13863 13411 sw
tri 13863 13313 13961 13411 ne
rect 13961 13313 14315 13411
tri 14315 13313 14413 13411 sw
tri 14413 13313 14511 13411 ne
rect 14511 13313 14865 13411
tri 14865 13313 14963 13411 sw
tri 14963 13313 15061 13411 ne
rect 15061 13313 15415 13411
tri 15415 13313 15513 13411 sw
tri 15513 13313 15611 13411 ne
rect 15611 13313 15965 13411
tri 15965 13313 16063 13411 sw
tri 16063 13313 16161 13411 ne
rect 16161 13313 16515 13411
tri 16515 13313 16613 13411 sw
tri 16613 13313 16711 13411 ne
rect 16711 13313 17065 13411
tri 17065 13313 17163 13411 sw
tri 17163 13313 17261 13411 ne
rect 17261 13313 17615 13411
tri 17615 13313 17713 13411 sw
tri 17713 13313 17811 13411 ne
rect 17811 13313 18165 13411
tri 18165 13313 18263 13411 sw
tri 18263 13313 18361 13411 ne
rect 18361 13313 18715 13411
tri 18715 13313 18813 13411 sw
tri 18813 13313 18911 13411 ne
rect 18911 13313 19265 13411
tri 19265 13313 19363 13411 sw
tri 19363 13313 19461 13411 ne
rect 19461 13313 20300 13411
rect -2000 13283 113 13313
tri 113 13283 143 13313 sw
tri 211 13283 241 13313 ne
rect 241 13283 663 13313
tri 663 13283 693 13313 sw
tri 761 13283 791 13313 ne
rect 791 13283 1213 13313
tri 1213 13283 1243 13313 sw
tri 1311 13283 1341 13313 ne
rect 1341 13283 1763 13313
tri 1763 13283 1793 13313 sw
tri 1861 13283 1891 13313 ne
rect 1891 13283 2313 13313
tri 2313 13283 2343 13313 sw
tri 2411 13283 2441 13313 ne
rect 2441 13283 2863 13313
tri 2863 13283 2893 13313 sw
tri 2961 13283 2991 13313 ne
rect 2991 13283 3413 13313
tri 3413 13283 3443 13313 sw
tri 3511 13283 3541 13313 ne
rect 3541 13283 3963 13313
tri 3963 13283 3993 13313 sw
tri 4061 13283 4091 13313 ne
rect 4091 13283 4513 13313
tri 4513 13283 4543 13313 sw
tri 4611 13283 4641 13313 ne
rect 4641 13283 5063 13313
tri 5063 13283 5093 13313 sw
tri 5161 13283 5191 13313 ne
rect 5191 13283 5613 13313
tri 5613 13283 5643 13313 sw
tri 5711 13283 5741 13313 ne
rect 5741 13283 6163 13313
tri 6163 13283 6193 13313 sw
tri 6261 13283 6291 13313 ne
rect 6291 13283 6713 13313
tri 6713 13283 6743 13313 sw
tri 6811 13283 6841 13313 ne
rect 6841 13283 7263 13313
tri 7263 13283 7293 13313 sw
tri 7361 13283 7391 13313 ne
rect 7391 13283 7813 13313
tri 7813 13283 7843 13313 sw
tri 7911 13283 7941 13313 ne
rect 7941 13283 8363 13313
tri 8363 13283 8393 13313 sw
tri 8461 13283 8491 13313 ne
rect 8491 13283 8913 13313
tri 8913 13283 8943 13313 sw
tri 9011 13283 9041 13313 ne
rect 9041 13283 9463 13313
tri 9463 13283 9493 13313 sw
tri 9561 13283 9591 13313 ne
rect 9591 13283 10013 13313
tri 10013 13283 10043 13313 sw
tri 10111 13283 10141 13313 ne
rect 10141 13283 10563 13313
tri 10563 13283 10593 13313 sw
tri 10661 13283 10691 13313 ne
rect 10691 13283 11113 13313
tri 11113 13283 11143 13313 sw
tri 11211 13283 11241 13313 ne
rect 11241 13283 11663 13313
tri 11663 13283 11693 13313 sw
tri 11761 13283 11791 13313 ne
rect 11791 13283 12213 13313
tri 12213 13283 12243 13313 sw
tri 12311 13283 12341 13313 ne
rect 12341 13283 12763 13313
tri 12763 13283 12793 13313 sw
tri 12861 13283 12891 13313 ne
rect 12891 13283 13313 13313
tri 13313 13283 13343 13313 sw
tri 13411 13283 13441 13313 ne
rect 13441 13283 13863 13313
tri 13863 13283 13893 13313 sw
tri 13961 13283 13991 13313 ne
rect 13991 13283 14413 13313
tri 14413 13283 14443 13313 sw
tri 14511 13283 14541 13313 ne
rect 14541 13283 14963 13313
tri 14963 13283 14993 13313 sw
tri 15061 13283 15091 13313 ne
rect 15091 13283 15513 13313
tri 15513 13283 15543 13313 sw
tri 15611 13283 15641 13313 ne
rect 15641 13283 16063 13313
tri 16063 13283 16093 13313 sw
tri 16161 13283 16191 13313 ne
rect 16191 13283 16613 13313
tri 16613 13283 16643 13313 sw
tri 16711 13283 16741 13313 ne
rect 16741 13283 17163 13313
tri 17163 13283 17193 13313 sw
tri 17261 13283 17291 13313 ne
rect 17291 13283 17713 13313
tri 17713 13283 17743 13313 sw
tri 17811 13283 17841 13313 ne
rect 17841 13283 18263 13313
tri 18263 13283 18293 13313 sw
tri 18361 13283 18391 13313 ne
rect 18391 13283 18813 13313
tri 18813 13283 18843 13313 sw
tri 18911 13283 18941 13313 ne
rect 18941 13283 19363 13313
tri 19363 13283 19393 13313 sw
tri 19461 13283 19491 13313 ne
rect 19491 13283 20300 13313
rect -2000 13185 143 13283
tri 143 13185 241 13283 sw
tri 241 13185 339 13283 ne
rect 339 13185 693 13283
tri 693 13185 791 13283 sw
tri 791 13185 889 13283 ne
rect 889 13185 1243 13283
tri 1243 13185 1341 13283 sw
tri 1341 13185 1439 13283 ne
rect 1439 13185 1793 13283
tri 1793 13185 1891 13283 sw
tri 1891 13185 1989 13283 ne
rect 1989 13185 2343 13283
tri 2343 13185 2441 13283 sw
tri 2441 13185 2539 13283 ne
rect 2539 13185 2893 13283
tri 2893 13185 2991 13283 sw
tri 2991 13185 3089 13283 ne
rect 3089 13185 3443 13283
tri 3443 13185 3541 13283 sw
tri 3541 13185 3639 13283 ne
rect 3639 13185 3993 13283
tri 3993 13185 4091 13283 sw
tri 4091 13185 4189 13283 ne
rect 4189 13185 4543 13283
tri 4543 13185 4641 13283 sw
tri 4641 13185 4739 13283 ne
rect 4739 13185 5093 13283
tri 5093 13185 5191 13283 sw
tri 5191 13185 5289 13283 ne
rect 5289 13185 5643 13283
tri 5643 13185 5741 13283 sw
tri 5741 13185 5839 13283 ne
rect 5839 13185 6193 13283
tri 6193 13185 6291 13283 sw
tri 6291 13185 6389 13283 ne
rect 6389 13185 6743 13283
tri 6743 13185 6841 13283 sw
tri 6841 13185 6939 13283 ne
rect 6939 13185 7293 13283
tri 7293 13185 7391 13283 sw
tri 7391 13185 7489 13283 ne
rect 7489 13185 7843 13283
tri 7843 13185 7941 13283 sw
tri 7941 13185 8039 13283 ne
rect 8039 13185 8393 13283
tri 8393 13185 8491 13283 sw
tri 8491 13185 8589 13283 ne
rect 8589 13185 8943 13283
tri 8943 13185 9041 13283 sw
tri 9041 13185 9139 13283 ne
rect 9139 13185 9493 13283
tri 9493 13185 9591 13283 sw
tri 9591 13185 9689 13283 ne
rect 9689 13185 10043 13283
tri 10043 13185 10141 13283 sw
tri 10141 13185 10239 13283 ne
rect 10239 13185 10593 13283
tri 10593 13185 10691 13283 sw
tri 10691 13185 10789 13283 ne
rect 10789 13185 11143 13283
tri 11143 13185 11241 13283 sw
tri 11241 13185 11339 13283 ne
rect 11339 13185 11693 13283
tri 11693 13185 11791 13283 sw
tri 11791 13185 11889 13283 ne
rect 11889 13185 12243 13283
tri 12243 13185 12341 13283 sw
tri 12341 13185 12439 13283 ne
rect 12439 13185 12793 13283
tri 12793 13185 12891 13283 sw
tri 12891 13185 12989 13283 ne
rect 12989 13185 13343 13283
tri 13343 13185 13441 13283 sw
tri 13441 13185 13539 13283 ne
rect 13539 13185 13893 13283
tri 13893 13185 13991 13283 sw
tri 13991 13185 14089 13283 ne
rect 14089 13185 14443 13283
tri 14443 13185 14541 13283 sw
tri 14541 13185 14639 13283 ne
rect 14639 13185 14993 13283
tri 14993 13185 15091 13283 sw
tri 15091 13185 15189 13283 ne
rect 15189 13185 15543 13283
tri 15543 13185 15641 13283 sw
tri 15641 13185 15739 13283 ne
rect 15739 13185 16093 13283
tri 16093 13185 16191 13283 sw
tri 16191 13185 16289 13283 ne
rect 16289 13185 16643 13283
tri 16643 13185 16741 13283 sw
tri 16741 13185 16839 13283 ne
rect 16839 13185 17193 13283
tri 17193 13185 17291 13283 sw
tri 17291 13185 17389 13283 ne
rect 17389 13185 17743 13283
tri 17743 13185 17841 13283 sw
tri 17841 13185 17939 13283 ne
rect 17939 13185 18293 13283
tri 18293 13185 18391 13283 sw
tri 18391 13185 18489 13283 ne
rect 18489 13185 18843 13283
tri 18843 13185 18941 13283 sw
tri 18941 13185 19039 13283 ne
rect 19039 13185 19393 13283
tri 19393 13185 19491 13283 sw
tri 19491 13185 19589 13283 ne
rect 19589 13185 20300 13283
rect -2000 13087 241 13185
tri 241 13087 339 13185 sw
tri 339 13087 437 13185 ne
rect 437 13087 791 13185
tri 791 13087 889 13185 sw
tri 889 13087 987 13185 ne
rect 987 13087 1341 13185
tri 1341 13087 1439 13185 sw
tri 1439 13087 1537 13185 ne
rect 1537 13087 1891 13185
tri 1891 13087 1989 13185 sw
tri 1989 13087 2087 13185 ne
rect 2087 13087 2441 13185
tri 2441 13087 2539 13185 sw
tri 2539 13087 2637 13185 ne
rect 2637 13087 2991 13185
tri 2991 13087 3089 13185 sw
tri 3089 13087 3187 13185 ne
rect 3187 13087 3541 13185
tri 3541 13087 3639 13185 sw
tri 3639 13087 3737 13185 ne
rect 3737 13087 4091 13185
tri 4091 13087 4189 13185 sw
tri 4189 13087 4287 13185 ne
rect 4287 13087 4641 13185
tri 4641 13087 4739 13185 sw
tri 4739 13087 4837 13185 ne
rect 4837 13087 5191 13185
tri 5191 13087 5289 13185 sw
tri 5289 13087 5387 13185 ne
rect 5387 13087 5741 13185
tri 5741 13087 5839 13185 sw
tri 5839 13087 5937 13185 ne
rect 5937 13087 6291 13185
tri 6291 13087 6389 13185 sw
tri 6389 13087 6487 13185 ne
rect 6487 13087 6841 13185
tri 6841 13087 6939 13185 sw
tri 6939 13087 7037 13185 ne
rect 7037 13087 7391 13185
tri 7391 13087 7489 13185 sw
tri 7489 13087 7587 13185 ne
rect 7587 13087 7941 13185
tri 7941 13087 8039 13185 sw
tri 8039 13087 8137 13185 ne
rect 8137 13087 8491 13185
tri 8491 13087 8589 13185 sw
tri 8589 13087 8687 13185 ne
rect 8687 13087 9041 13185
tri 9041 13087 9139 13185 sw
tri 9139 13087 9237 13185 ne
rect 9237 13087 9591 13185
tri 9591 13087 9689 13185 sw
tri 9689 13087 9787 13185 ne
rect 9787 13087 10141 13185
tri 10141 13087 10239 13185 sw
tri 10239 13087 10337 13185 ne
rect 10337 13087 10691 13185
tri 10691 13087 10789 13185 sw
tri 10789 13087 10887 13185 ne
rect 10887 13087 11241 13185
tri 11241 13087 11339 13185 sw
tri 11339 13087 11437 13185 ne
rect 11437 13087 11791 13185
tri 11791 13087 11889 13185 sw
tri 11889 13087 11987 13185 ne
rect 11987 13087 12341 13185
tri 12341 13087 12439 13185 sw
tri 12439 13087 12537 13185 ne
rect 12537 13087 12891 13185
tri 12891 13087 12989 13185 sw
tri 12989 13087 13087 13185 ne
rect 13087 13087 13441 13185
tri 13441 13087 13539 13185 sw
tri 13539 13087 13637 13185 ne
rect 13637 13087 13991 13185
tri 13991 13087 14089 13185 sw
tri 14089 13087 14187 13185 ne
rect 14187 13087 14541 13185
tri 14541 13087 14639 13185 sw
tri 14639 13087 14737 13185 ne
rect 14737 13087 15091 13185
tri 15091 13087 15189 13185 sw
tri 15189 13087 15287 13185 ne
rect 15287 13087 15641 13185
tri 15641 13087 15739 13185 sw
tri 15739 13087 15837 13185 ne
rect 15837 13087 16191 13185
tri 16191 13087 16289 13185 sw
tri 16289 13087 16387 13185 ne
rect 16387 13087 16741 13185
tri 16741 13087 16839 13185 sw
tri 16839 13087 16937 13185 ne
rect 16937 13087 17291 13185
tri 17291 13087 17389 13185 sw
tri 17389 13087 17487 13185 ne
rect 17487 13087 17841 13185
tri 17841 13087 17939 13185 sw
tri 17939 13087 18037 13185 ne
rect 18037 13087 18391 13185
tri 18391 13087 18489 13185 sw
tri 18489 13087 18587 13185 ne
rect 18587 13087 18941 13185
tri 18941 13087 19039 13185 sw
tri 19039 13087 19137 13185 ne
rect 19137 13087 19491 13185
tri 19491 13087 19589 13185 sw
tri 19589 13087 19687 13185 ne
rect 19687 13087 20300 13185
rect -2000 12989 339 13087
tri 339 12989 437 13087 sw
tri 437 12989 535 13087 ne
rect 535 12989 889 13087
tri 889 12989 987 13087 sw
tri 987 12989 1085 13087 ne
rect 1085 12989 1439 13087
tri 1439 12989 1537 13087 sw
tri 1537 12989 1635 13087 ne
rect 1635 12989 1989 13087
tri 1989 12989 2087 13087 sw
tri 2087 12989 2185 13087 ne
rect 2185 12989 2539 13087
tri 2539 12989 2637 13087 sw
tri 2637 12989 2735 13087 ne
rect 2735 12989 3089 13087
tri 3089 12989 3187 13087 sw
tri 3187 12989 3285 13087 ne
rect 3285 12989 3639 13087
tri 3639 12989 3737 13087 sw
tri 3737 12989 3835 13087 ne
rect 3835 12989 4189 13087
tri 4189 12989 4287 13087 sw
tri 4287 12989 4385 13087 ne
rect 4385 12989 4739 13087
tri 4739 12989 4837 13087 sw
tri 4837 12989 4935 13087 ne
rect 4935 12989 5289 13087
tri 5289 12989 5387 13087 sw
tri 5387 12989 5485 13087 ne
rect 5485 12989 5839 13087
tri 5839 12989 5937 13087 sw
tri 5937 12989 6035 13087 ne
rect 6035 12989 6389 13087
tri 6389 12989 6487 13087 sw
tri 6487 12989 6585 13087 ne
rect 6585 12989 6939 13087
tri 6939 12989 7037 13087 sw
tri 7037 12989 7135 13087 ne
rect 7135 12989 7489 13087
tri 7489 12989 7587 13087 sw
tri 7587 12989 7685 13087 ne
rect 7685 12989 8039 13087
tri 8039 12989 8137 13087 sw
tri 8137 12989 8235 13087 ne
rect 8235 12989 8589 13087
tri 8589 12989 8687 13087 sw
tri 8687 12989 8785 13087 ne
rect 8785 12989 9139 13087
tri 9139 12989 9237 13087 sw
tri 9237 12989 9335 13087 ne
rect 9335 12989 9689 13087
tri 9689 12989 9787 13087 sw
tri 9787 12989 9885 13087 ne
rect 9885 12989 10239 13087
tri 10239 12989 10337 13087 sw
tri 10337 12989 10435 13087 ne
rect 10435 12989 10789 13087
tri 10789 12989 10887 13087 sw
tri 10887 12989 10985 13087 ne
rect 10985 12989 11339 13087
tri 11339 12989 11437 13087 sw
tri 11437 12989 11535 13087 ne
rect 11535 12989 11889 13087
tri 11889 12989 11987 13087 sw
tri 11987 12989 12085 13087 ne
rect 12085 12989 12439 13087
tri 12439 12989 12537 13087 sw
tri 12537 12989 12635 13087 ne
rect 12635 12989 12989 13087
tri 12989 12989 13087 13087 sw
tri 13087 12989 13185 13087 ne
rect 13185 12989 13539 13087
tri 13539 12989 13637 13087 sw
tri 13637 12989 13735 13087 ne
rect 13735 12989 14089 13087
tri 14089 12989 14187 13087 sw
tri 14187 12989 14285 13087 ne
rect 14285 12989 14639 13087
tri 14639 12989 14737 13087 sw
tri 14737 12989 14835 13087 ne
rect 14835 12989 15189 13087
tri 15189 12989 15287 13087 sw
tri 15287 12989 15385 13087 ne
rect 15385 12989 15739 13087
tri 15739 12989 15837 13087 sw
tri 15837 12989 15935 13087 ne
rect 15935 12989 16289 13087
tri 16289 12989 16387 13087 sw
tri 16387 12989 16485 13087 ne
rect 16485 12989 16839 13087
tri 16839 12989 16937 13087 sw
tri 16937 12989 17035 13087 ne
rect 17035 12989 17389 13087
tri 17389 12989 17487 13087 sw
tri 17487 12989 17585 13087 ne
rect 17585 12989 17939 13087
tri 17939 12989 18037 13087 sw
tri 18037 12989 18135 13087 ne
rect 18135 12989 18489 13087
tri 18489 12989 18587 13087 sw
tri 18587 12989 18685 13087 ne
rect 18685 12989 19039 13087
tri 19039 12989 19137 13087 sw
tri 19137 12989 19235 13087 ne
rect 19235 12989 19589 13087
tri 19589 12989 19687 13087 sw
rect 20800 12989 21800 13637
rect -2000 12985 437 12989
rect -2000 12865 215 12985
rect 335 12891 437 12985
tri 437 12891 535 12989 sw
tri 535 12891 633 12989 ne
rect 633 12985 987 12989
rect 633 12891 765 12985
rect 335 12865 535 12891
rect -2000 12861 535 12865
rect -2000 12213 -1000 12861
tri 113 12763 211 12861 ne
rect 211 12813 535 12861
tri 535 12813 613 12891 sw
tri 633 12813 711 12891 ne
rect 711 12865 765 12891
rect 885 12891 987 12985
tri 987 12891 1085 12989 sw
tri 1085 12891 1183 12989 ne
rect 1183 12985 1537 12989
rect 1183 12891 1315 12985
rect 885 12865 1085 12891
rect 711 12813 1085 12865
tri 1085 12813 1163 12891 sw
tri 1183 12813 1261 12891 ne
rect 1261 12865 1315 12891
rect 1435 12891 1537 12985
tri 1537 12891 1635 12989 sw
tri 1635 12891 1733 12989 ne
rect 1733 12985 2087 12989
rect 1733 12891 1865 12985
rect 1435 12865 1635 12891
rect 1261 12813 1635 12865
tri 1635 12813 1713 12891 sw
tri 1733 12813 1811 12891 ne
rect 1811 12865 1865 12891
rect 1985 12891 2087 12985
tri 2087 12891 2185 12989 sw
tri 2185 12891 2283 12989 ne
rect 2283 12985 2637 12989
rect 2283 12891 2415 12985
rect 1985 12865 2185 12891
rect 1811 12813 2185 12865
tri 2185 12813 2263 12891 sw
tri 2283 12813 2361 12891 ne
rect 2361 12865 2415 12891
rect 2535 12891 2637 12985
tri 2637 12891 2735 12989 sw
tri 2735 12891 2833 12989 ne
rect 2833 12985 3187 12989
rect 2833 12891 2965 12985
rect 2535 12865 2735 12891
rect 2361 12813 2735 12865
tri 2735 12813 2813 12891 sw
tri 2833 12813 2911 12891 ne
rect 2911 12865 2965 12891
rect 3085 12891 3187 12985
tri 3187 12891 3285 12989 sw
tri 3285 12891 3383 12989 ne
rect 3383 12985 3737 12989
rect 3383 12891 3515 12985
rect 3085 12865 3285 12891
rect 2911 12813 3285 12865
tri 3285 12813 3363 12891 sw
tri 3383 12813 3461 12891 ne
rect 3461 12865 3515 12891
rect 3635 12891 3737 12985
tri 3737 12891 3835 12989 sw
tri 3835 12891 3933 12989 ne
rect 3933 12985 4287 12989
rect 3933 12891 4065 12985
rect 3635 12865 3835 12891
rect 3461 12813 3835 12865
tri 3835 12813 3913 12891 sw
tri 3933 12813 4011 12891 ne
rect 4011 12865 4065 12891
rect 4185 12891 4287 12985
tri 4287 12891 4385 12989 sw
tri 4385 12891 4483 12989 ne
rect 4483 12985 4837 12989
rect 4483 12891 4615 12985
rect 4185 12865 4385 12891
rect 4011 12813 4385 12865
tri 4385 12813 4463 12891 sw
tri 4483 12813 4561 12891 ne
rect 4561 12865 4615 12891
rect 4735 12891 4837 12985
tri 4837 12891 4935 12989 sw
tri 4935 12891 5033 12989 ne
rect 5033 12985 5387 12989
rect 5033 12891 5165 12985
rect 4735 12865 4935 12891
rect 4561 12813 4935 12865
tri 4935 12813 5013 12891 sw
tri 5033 12813 5111 12891 ne
rect 5111 12865 5165 12891
rect 5285 12891 5387 12985
tri 5387 12891 5485 12989 sw
tri 5485 12891 5583 12989 ne
rect 5583 12985 5937 12989
rect 5583 12891 5715 12985
rect 5285 12865 5485 12891
rect 5111 12813 5485 12865
tri 5485 12813 5563 12891 sw
tri 5583 12813 5661 12891 ne
rect 5661 12865 5715 12891
rect 5835 12891 5937 12985
tri 5937 12891 6035 12989 sw
tri 6035 12891 6133 12989 ne
rect 6133 12985 6487 12989
rect 6133 12891 6265 12985
rect 5835 12865 6035 12891
rect 5661 12813 6035 12865
tri 6035 12813 6113 12891 sw
tri 6133 12813 6211 12891 ne
rect 6211 12865 6265 12891
rect 6385 12891 6487 12985
tri 6487 12891 6585 12989 sw
tri 6585 12891 6683 12989 ne
rect 6683 12985 7037 12989
rect 6683 12891 6815 12985
rect 6385 12865 6585 12891
rect 6211 12813 6585 12865
tri 6585 12813 6663 12891 sw
tri 6683 12813 6761 12891 ne
rect 6761 12865 6815 12891
rect 6935 12891 7037 12985
tri 7037 12891 7135 12989 sw
tri 7135 12891 7233 12989 ne
rect 7233 12985 7587 12989
rect 7233 12891 7365 12985
rect 6935 12865 7135 12891
rect 6761 12813 7135 12865
tri 7135 12813 7213 12891 sw
tri 7233 12813 7311 12891 ne
rect 7311 12865 7365 12891
rect 7485 12891 7587 12985
tri 7587 12891 7685 12989 sw
tri 7685 12891 7783 12989 ne
rect 7783 12985 8137 12989
rect 7783 12891 7915 12985
rect 7485 12865 7685 12891
rect 7311 12813 7685 12865
tri 7685 12813 7763 12891 sw
tri 7783 12813 7861 12891 ne
rect 7861 12865 7915 12891
rect 8035 12891 8137 12985
tri 8137 12891 8235 12989 sw
tri 8235 12891 8333 12989 ne
rect 8333 12985 8687 12989
rect 8333 12891 8465 12985
rect 8035 12865 8235 12891
rect 7861 12813 8235 12865
tri 8235 12813 8313 12891 sw
tri 8333 12813 8411 12891 ne
rect 8411 12865 8465 12891
rect 8585 12891 8687 12985
tri 8687 12891 8785 12989 sw
tri 8785 12891 8883 12989 ne
rect 8883 12985 9237 12989
rect 8883 12891 9015 12985
rect 8585 12865 8785 12891
rect 8411 12813 8785 12865
tri 8785 12813 8863 12891 sw
tri 8883 12813 8961 12891 ne
rect 8961 12865 9015 12891
rect 9135 12891 9237 12985
tri 9237 12891 9335 12989 sw
tri 9335 12891 9433 12989 ne
rect 9433 12985 9787 12989
rect 9433 12891 9565 12985
rect 9135 12865 9335 12891
rect 8961 12813 9335 12865
tri 9335 12813 9413 12891 sw
tri 9433 12813 9511 12891 ne
rect 9511 12865 9565 12891
rect 9685 12891 9787 12985
tri 9787 12891 9885 12989 sw
tri 9885 12891 9983 12989 ne
rect 9983 12985 10337 12989
rect 9983 12891 10115 12985
rect 9685 12865 9885 12891
rect 9511 12813 9885 12865
tri 9885 12813 9963 12891 sw
tri 9983 12813 10061 12891 ne
rect 10061 12865 10115 12891
rect 10235 12891 10337 12985
tri 10337 12891 10435 12989 sw
tri 10435 12891 10533 12989 ne
rect 10533 12985 10887 12989
rect 10533 12891 10665 12985
rect 10235 12865 10435 12891
rect 10061 12813 10435 12865
tri 10435 12813 10513 12891 sw
tri 10533 12813 10611 12891 ne
rect 10611 12865 10665 12891
rect 10785 12891 10887 12985
tri 10887 12891 10985 12989 sw
tri 10985 12891 11083 12989 ne
rect 11083 12985 11437 12989
rect 11083 12891 11215 12985
rect 10785 12865 10985 12891
rect 10611 12813 10985 12865
tri 10985 12813 11063 12891 sw
tri 11083 12813 11161 12891 ne
rect 11161 12865 11215 12891
rect 11335 12891 11437 12985
tri 11437 12891 11535 12989 sw
tri 11535 12891 11633 12989 ne
rect 11633 12985 11987 12989
rect 11633 12891 11765 12985
rect 11335 12865 11535 12891
rect 11161 12813 11535 12865
tri 11535 12813 11613 12891 sw
tri 11633 12813 11711 12891 ne
rect 11711 12865 11765 12891
rect 11885 12891 11987 12985
tri 11987 12891 12085 12989 sw
tri 12085 12891 12183 12989 ne
rect 12183 12985 12537 12989
rect 12183 12891 12315 12985
rect 11885 12865 12085 12891
rect 11711 12813 12085 12865
tri 12085 12813 12163 12891 sw
tri 12183 12813 12261 12891 ne
rect 12261 12865 12315 12891
rect 12435 12891 12537 12985
tri 12537 12891 12635 12989 sw
tri 12635 12891 12733 12989 ne
rect 12733 12985 13087 12989
rect 12733 12891 12865 12985
rect 12435 12865 12635 12891
rect 12261 12813 12635 12865
tri 12635 12813 12713 12891 sw
tri 12733 12813 12811 12891 ne
rect 12811 12865 12865 12891
rect 12985 12891 13087 12985
tri 13087 12891 13185 12989 sw
tri 13185 12891 13283 12989 ne
rect 13283 12985 13637 12989
rect 13283 12891 13415 12985
rect 12985 12865 13185 12891
rect 12811 12813 13185 12865
tri 13185 12813 13263 12891 sw
tri 13283 12813 13361 12891 ne
rect 13361 12865 13415 12891
rect 13535 12891 13637 12985
tri 13637 12891 13735 12989 sw
tri 13735 12891 13833 12989 ne
rect 13833 12985 14187 12989
rect 13833 12891 13965 12985
rect 13535 12865 13735 12891
rect 13361 12813 13735 12865
tri 13735 12813 13813 12891 sw
tri 13833 12813 13911 12891 ne
rect 13911 12865 13965 12891
rect 14085 12891 14187 12985
tri 14187 12891 14285 12989 sw
tri 14285 12891 14383 12989 ne
rect 14383 12985 14737 12989
rect 14383 12891 14515 12985
rect 14085 12865 14285 12891
rect 13911 12813 14285 12865
tri 14285 12813 14363 12891 sw
tri 14383 12813 14461 12891 ne
rect 14461 12865 14515 12891
rect 14635 12891 14737 12985
tri 14737 12891 14835 12989 sw
tri 14835 12891 14933 12989 ne
rect 14933 12985 15287 12989
rect 14933 12891 15065 12985
rect 14635 12865 14835 12891
rect 14461 12813 14835 12865
tri 14835 12813 14913 12891 sw
tri 14933 12813 15011 12891 ne
rect 15011 12865 15065 12891
rect 15185 12891 15287 12985
tri 15287 12891 15385 12989 sw
tri 15385 12891 15483 12989 ne
rect 15483 12985 15837 12989
rect 15483 12891 15615 12985
rect 15185 12865 15385 12891
rect 15011 12813 15385 12865
tri 15385 12813 15463 12891 sw
tri 15483 12813 15561 12891 ne
rect 15561 12865 15615 12891
rect 15735 12891 15837 12985
tri 15837 12891 15935 12989 sw
tri 15935 12891 16033 12989 ne
rect 16033 12985 16387 12989
rect 16033 12891 16165 12985
rect 15735 12865 15935 12891
rect 15561 12813 15935 12865
tri 15935 12813 16013 12891 sw
tri 16033 12813 16111 12891 ne
rect 16111 12865 16165 12891
rect 16285 12891 16387 12985
tri 16387 12891 16485 12989 sw
tri 16485 12891 16583 12989 ne
rect 16583 12985 16937 12989
rect 16583 12891 16715 12985
rect 16285 12865 16485 12891
rect 16111 12813 16485 12865
tri 16485 12813 16563 12891 sw
tri 16583 12813 16661 12891 ne
rect 16661 12865 16715 12891
rect 16835 12891 16937 12985
tri 16937 12891 17035 12989 sw
tri 17035 12891 17133 12989 ne
rect 17133 12985 17487 12989
rect 17133 12891 17265 12985
rect 16835 12865 17035 12891
rect 16661 12813 17035 12865
tri 17035 12813 17113 12891 sw
tri 17133 12813 17211 12891 ne
rect 17211 12865 17265 12891
rect 17385 12891 17487 12985
tri 17487 12891 17585 12989 sw
tri 17585 12891 17683 12989 ne
rect 17683 12985 18037 12989
rect 17683 12891 17815 12985
rect 17385 12865 17585 12891
rect 17211 12813 17585 12865
tri 17585 12813 17663 12891 sw
tri 17683 12813 17761 12891 ne
rect 17761 12865 17815 12891
rect 17935 12891 18037 12985
tri 18037 12891 18135 12989 sw
tri 18135 12891 18233 12989 ne
rect 18233 12985 18587 12989
rect 18233 12891 18365 12985
rect 17935 12865 18135 12891
rect 17761 12813 18135 12865
tri 18135 12813 18213 12891 sw
tri 18233 12813 18311 12891 ne
rect 18311 12865 18365 12891
rect 18485 12891 18587 12985
tri 18587 12891 18685 12989 sw
tri 18685 12891 18783 12989 ne
rect 18783 12985 19137 12989
rect 18783 12891 18915 12985
rect 18485 12865 18685 12891
rect 18311 12813 18685 12865
tri 18685 12813 18763 12891 sw
tri 18783 12813 18861 12891 ne
rect 18861 12865 18915 12891
rect 19035 12891 19137 12985
tri 19137 12891 19235 12989 sw
tri 19235 12891 19333 12989 ne
rect 19333 12985 21800 12989
rect 19333 12891 19465 12985
rect 19035 12865 19235 12891
rect 18861 12813 19235 12865
tri 19235 12813 19313 12891 sw
tri 19333 12813 19411 12891 ne
rect 19411 12865 19465 12891
rect 19585 12865 21800 12985
rect 19411 12813 21800 12865
rect 211 12763 613 12813
rect -500 12713 113 12763
tri 113 12713 163 12763 sw
tri 211 12713 261 12763 ne
rect 261 12733 613 12763
tri 613 12733 693 12813 sw
tri 711 12733 791 12813 ne
rect 791 12733 1163 12813
tri 1163 12733 1243 12813 sw
tri 1261 12733 1341 12813 ne
rect 1341 12733 1713 12813
tri 1713 12733 1793 12813 sw
tri 1811 12733 1891 12813 ne
rect 1891 12733 2263 12813
tri 2263 12733 2343 12813 sw
tri 2361 12733 2441 12813 ne
rect 2441 12733 2813 12813
tri 2813 12733 2893 12813 sw
tri 2911 12733 2991 12813 ne
rect 2991 12733 3363 12813
tri 3363 12733 3443 12813 sw
tri 3461 12733 3541 12813 ne
rect 3541 12733 3913 12813
tri 3913 12733 3993 12813 sw
tri 4011 12733 4091 12813 ne
rect 4091 12733 4463 12813
tri 4463 12733 4543 12813 sw
tri 4561 12733 4641 12813 ne
rect 4641 12733 5013 12813
tri 5013 12733 5093 12813 sw
tri 5111 12733 5191 12813 ne
rect 5191 12733 5563 12813
tri 5563 12733 5643 12813 sw
tri 5661 12733 5741 12813 ne
rect 5741 12733 6113 12813
tri 6113 12733 6193 12813 sw
tri 6211 12733 6291 12813 ne
rect 6291 12733 6663 12813
tri 6663 12733 6743 12813 sw
tri 6761 12733 6841 12813 ne
rect 6841 12733 7213 12813
tri 7213 12733 7293 12813 sw
tri 7311 12733 7391 12813 ne
rect 7391 12733 7763 12813
tri 7763 12733 7843 12813 sw
tri 7861 12733 7941 12813 ne
rect 7941 12733 8313 12813
tri 8313 12733 8393 12813 sw
tri 8411 12733 8491 12813 ne
rect 8491 12733 8863 12813
tri 8863 12733 8943 12813 sw
tri 8961 12733 9041 12813 ne
rect 9041 12733 9413 12813
tri 9413 12733 9493 12813 sw
tri 9511 12733 9591 12813 ne
rect 9591 12733 9963 12813
tri 9963 12733 10043 12813 sw
tri 10061 12733 10141 12813 ne
rect 10141 12733 10513 12813
tri 10513 12733 10593 12813 sw
tri 10611 12733 10691 12813 ne
rect 10691 12733 11063 12813
tri 11063 12733 11143 12813 sw
tri 11161 12733 11241 12813 ne
rect 11241 12733 11613 12813
tri 11613 12733 11693 12813 sw
tri 11711 12733 11791 12813 ne
rect 11791 12733 12163 12813
tri 12163 12733 12243 12813 sw
tri 12261 12733 12341 12813 ne
rect 12341 12733 12713 12813
tri 12713 12733 12793 12813 sw
tri 12811 12733 12891 12813 ne
rect 12891 12733 13263 12813
tri 13263 12733 13343 12813 sw
tri 13361 12733 13441 12813 ne
rect 13441 12733 13813 12813
tri 13813 12733 13893 12813 sw
tri 13911 12733 13991 12813 ne
rect 13991 12733 14363 12813
tri 14363 12733 14443 12813 sw
tri 14461 12733 14541 12813 ne
rect 14541 12733 14913 12813
tri 14913 12733 14993 12813 sw
tri 15011 12733 15091 12813 ne
rect 15091 12733 15463 12813
tri 15463 12733 15543 12813 sw
tri 15561 12733 15641 12813 ne
rect 15641 12733 16013 12813
tri 16013 12733 16093 12813 sw
tri 16111 12733 16191 12813 ne
rect 16191 12733 16563 12813
tri 16563 12733 16643 12813 sw
tri 16661 12733 16741 12813 ne
rect 16741 12733 17113 12813
tri 17113 12733 17193 12813 sw
tri 17211 12733 17291 12813 ne
rect 17291 12733 17663 12813
tri 17663 12733 17743 12813 sw
tri 17761 12733 17841 12813 ne
rect 17841 12733 18213 12813
tri 18213 12733 18293 12813 sw
tri 18311 12733 18391 12813 ne
rect 18391 12733 18763 12813
tri 18763 12733 18843 12813 sw
tri 18861 12733 18941 12813 ne
rect 18941 12733 19313 12813
tri 19313 12733 19393 12813 sw
tri 19411 12733 19491 12813 ne
rect 19491 12733 20100 12813
rect 261 12713 693 12733
rect -500 12635 163 12713
tri 163 12635 241 12713 sw
tri 261 12635 339 12713 ne
rect 339 12635 693 12713
tri 693 12635 791 12733 sw
tri 791 12635 889 12733 ne
rect 889 12635 1243 12733
tri 1243 12635 1341 12733 sw
tri 1341 12635 1439 12733 ne
rect 1439 12635 1793 12733
tri 1793 12635 1891 12733 sw
tri 1891 12635 1989 12733 ne
rect 1989 12635 2343 12733
tri 2343 12635 2441 12733 sw
tri 2441 12635 2539 12733 ne
rect 2539 12635 2893 12733
tri 2893 12635 2991 12733 sw
tri 2991 12635 3089 12733 ne
rect 3089 12635 3443 12733
tri 3443 12635 3541 12733 sw
tri 3541 12635 3639 12733 ne
rect 3639 12635 3993 12733
tri 3993 12635 4091 12733 sw
tri 4091 12635 4189 12733 ne
rect 4189 12635 4543 12733
tri 4543 12635 4641 12733 sw
tri 4641 12635 4739 12733 ne
rect 4739 12635 5093 12733
tri 5093 12635 5191 12733 sw
tri 5191 12635 5289 12733 ne
rect 5289 12635 5643 12733
tri 5643 12635 5741 12733 sw
tri 5741 12635 5839 12733 ne
rect 5839 12635 6193 12733
tri 6193 12635 6291 12733 sw
tri 6291 12635 6389 12733 ne
rect 6389 12635 6743 12733
tri 6743 12635 6841 12733 sw
tri 6841 12635 6939 12733 ne
rect 6939 12635 7293 12733
tri 7293 12635 7391 12733 sw
tri 7391 12635 7489 12733 ne
rect 7489 12635 7843 12733
tri 7843 12635 7941 12733 sw
tri 7941 12635 8039 12733 ne
rect 8039 12635 8393 12733
tri 8393 12635 8491 12733 sw
tri 8491 12635 8589 12733 ne
rect 8589 12635 8943 12733
tri 8943 12635 9041 12733 sw
tri 9041 12635 9139 12733 ne
rect 9139 12635 9493 12733
tri 9493 12635 9591 12733 sw
tri 9591 12635 9689 12733 ne
rect 9689 12635 10043 12733
tri 10043 12635 10141 12733 sw
tri 10141 12635 10239 12733 ne
rect 10239 12635 10593 12733
tri 10593 12635 10691 12733 sw
tri 10691 12635 10789 12733 ne
rect 10789 12635 11143 12733
tri 11143 12635 11241 12733 sw
tri 11241 12635 11339 12733 ne
rect 11339 12635 11693 12733
tri 11693 12635 11791 12733 sw
tri 11791 12635 11889 12733 ne
rect 11889 12635 12243 12733
tri 12243 12635 12341 12733 sw
tri 12341 12635 12439 12733 ne
rect 12439 12635 12793 12733
tri 12793 12635 12891 12733 sw
tri 12891 12635 12989 12733 ne
rect 12989 12635 13343 12733
tri 13343 12635 13441 12733 sw
tri 13441 12635 13539 12733 ne
rect 13539 12635 13893 12733
tri 13893 12635 13991 12733 sw
tri 13991 12635 14089 12733 ne
rect 14089 12635 14443 12733
tri 14443 12635 14541 12733 sw
tri 14541 12635 14639 12733 ne
rect 14639 12635 14993 12733
tri 14993 12635 15091 12733 sw
tri 15091 12635 15189 12733 ne
rect 15189 12635 15543 12733
tri 15543 12635 15641 12733 sw
tri 15641 12635 15739 12733 ne
rect 15739 12635 16093 12733
tri 16093 12635 16191 12733 sw
tri 16191 12635 16289 12733 ne
rect 16289 12635 16643 12733
tri 16643 12635 16741 12733 sw
tri 16741 12635 16839 12733 ne
rect 16839 12635 17193 12733
tri 17193 12635 17291 12733 sw
tri 17291 12635 17389 12733 ne
rect 17389 12635 17743 12733
tri 17743 12635 17841 12733 sw
tri 17841 12635 17939 12733 ne
rect 17939 12635 18293 12733
tri 18293 12635 18391 12733 sw
tri 18391 12635 18489 12733 ne
rect 18489 12635 18843 12733
tri 18843 12635 18941 12733 sw
tri 18941 12635 19039 12733 ne
rect 19039 12635 19393 12733
tri 19393 12635 19491 12733 sw
tri 19491 12635 19589 12733 ne
rect 19589 12713 20100 12733
rect 20200 12713 21800 12813
rect 19589 12635 21800 12713
rect -500 12587 241 12635
rect -500 12487 -400 12587
rect -300 12537 241 12587
tri 241 12537 339 12635 sw
tri 339 12537 437 12635 ne
rect 437 12537 791 12635
tri 791 12537 889 12635 sw
tri 889 12537 987 12635 ne
rect 987 12537 1341 12635
tri 1341 12537 1439 12635 sw
tri 1439 12537 1537 12635 ne
rect 1537 12537 1891 12635
tri 1891 12537 1989 12635 sw
tri 1989 12537 2087 12635 ne
rect 2087 12537 2441 12635
tri 2441 12537 2539 12635 sw
tri 2539 12537 2637 12635 ne
rect 2637 12537 2991 12635
tri 2991 12537 3089 12635 sw
tri 3089 12537 3187 12635 ne
rect 3187 12537 3541 12635
tri 3541 12537 3639 12635 sw
tri 3639 12537 3737 12635 ne
rect 3737 12537 4091 12635
tri 4091 12537 4189 12635 sw
tri 4189 12537 4287 12635 ne
rect 4287 12537 4641 12635
tri 4641 12537 4739 12635 sw
tri 4739 12537 4837 12635 ne
rect 4837 12537 5191 12635
tri 5191 12537 5289 12635 sw
tri 5289 12537 5387 12635 ne
rect 5387 12537 5741 12635
tri 5741 12537 5839 12635 sw
tri 5839 12537 5937 12635 ne
rect 5937 12537 6291 12635
tri 6291 12537 6389 12635 sw
tri 6389 12537 6487 12635 ne
rect 6487 12537 6841 12635
tri 6841 12537 6939 12635 sw
tri 6939 12537 7037 12635 ne
rect 7037 12537 7391 12635
tri 7391 12537 7489 12635 sw
tri 7489 12537 7587 12635 ne
rect 7587 12537 7941 12635
tri 7941 12537 8039 12635 sw
tri 8039 12537 8137 12635 ne
rect 8137 12537 8491 12635
tri 8491 12537 8589 12635 sw
tri 8589 12537 8687 12635 ne
rect 8687 12537 9041 12635
tri 9041 12537 9139 12635 sw
tri 9139 12537 9237 12635 ne
rect 9237 12537 9591 12635
tri 9591 12537 9689 12635 sw
tri 9689 12537 9787 12635 ne
rect 9787 12537 10141 12635
tri 10141 12537 10239 12635 sw
tri 10239 12537 10337 12635 ne
rect 10337 12537 10691 12635
tri 10691 12537 10789 12635 sw
tri 10789 12537 10887 12635 ne
rect 10887 12537 11241 12635
tri 11241 12537 11339 12635 sw
tri 11339 12537 11437 12635 ne
rect 11437 12537 11791 12635
tri 11791 12537 11889 12635 sw
tri 11889 12537 11987 12635 ne
rect 11987 12537 12341 12635
tri 12341 12537 12439 12635 sw
tri 12439 12537 12537 12635 ne
rect 12537 12537 12891 12635
tri 12891 12537 12989 12635 sw
tri 12989 12537 13087 12635 ne
rect 13087 12537 13441 12635
tri 13441 12537 13539 12635 sw
tri 13539 12537 13637 12635 ne
rect 13637 12537 13991 12635
tri 13991 12537 14089 12635 sw
tri 14089 12537 14187 12635 ne
rect 14187 12537 14541 12635
tri 14541 12537 14639 12635 sw
tri 14639 12537 14737 12635 ne
rect 14737 12537 15091 12635
tri 15091 12537 15189 12635 sw
tri 15189 12537 15287 12635 ne
rect 15287 12537 15641 12635
tri 15641 12537 15739 12635 sw
tri 15739 12537 15837 12635 ne
rect 15837 12537 16191 12635
tri 16191 12537 16289 12635 sw
tri 16289 12537 16387 12635 ne
rect 16387 12537 16741 12635
tri 16741 12537 16839 12635 sw
tri 16839 12537 16937 12635 ne
rect 16937 12537 17291 12635
tri 17291 12537 17389 12635 sw
tri 17389 12537 17487 12635 ne
rect 17487 12537 17841 12635
tri 17841 12537 17939 12635 sw
tri 17939 12537 18037 12635 ne
rect 18037 12537 18391 12635
tri 18391 12537 18489 12635 sw
tri 18489 12537 18587 12635 ne
rect 18587 12537 18941 12635
tri 18941 12537 19039 12635 sw
tri 19039 12537 19137 12635 ne
rect 19137 12537 19491 12635
tri 19491 12537 19589 12635 sw
tri 19589 12537 19687 12635 ne
rect 19687 12537 21800 12635
rect -300 12487 339 12537
rect -500 12439 339 12487
tri 339 12439 437 12537 sw
tri 437 12439 535 12537 ne
rect 535 12439 889 12537
tri 889 12439 987 12537 sw
tri 987 12439 1085 12537 ne
rect 1085 12439 1439 12537
tri 1439 12439 1537 12537 sw
tri 1537 12439 1635 12537 ne
rect 1635 12439 1989 12537
tri 1989 12439 2087 12537 sw
tri 2087 12439 2185 12537 ne
rect 2185 12439 2539 12537
tri 2539 12439 2637 12537 sw
tri 2637 12439 2735 12537 ne
rect 2735 12439 3089 12537
tri 3089 12439 3187 12537 sw
tri 3187 12439 3285 12537 ne
rect 3285 12439 3639 12537
tri 3639 12439 3737 12537 sw
tri 3737 12439 3835 12537 ne
rect 3835 12439 4189 12537
tri 4189 12439 4287 12537 sw
tri 4287 12439 4385 12537 ne
rect 4385 12439 4739 12537
tri 4739 12439 4837 12537 sw
tri 4837 12439 4935 12537 ne
rect 4935 12439 5289 12537
tri 5289 12439 5387 12537 sw
tri 5387 12439 5485 12537 ne
rect 5485 12439 5839 12537
tri 5839 12439 5937 12537 sw
tri 5937 12439 6035 12537 ne
rect 6035 12439 6389 12537
tri 6389 12439 6487 12537 sw
tri 6487 12439 6585 12537 ne
rect 6585 12439 6939 12537
tri 6939 12439 7037 12537 sw
tri 7037 12439 7135 12537 ne
rect 7135 12439 7489 12537
tri 7489 12439 7587 12537 sw
tri 7587 12439 7685 12537 ne
rect 7685 12439 8039 12537
tri 8039 12439 8137 12537 sw
tri 8137 12439 8235 12537 ne
rect 8235 12439 8589 12537
tri 8589 12439 8687 12537 sw
tri 8687 12439 8785 12537 ne
rect 8785 12439 9139 12537
tri 9139 12439 9237 12537 sw
tri 9237 12439 9335 12537 ne
rect 9335 12439 9689 12537
tri 9689 12439 9787 12537 sw
tri 9787 12439 9885 12537 ne
rect 9885 12439 10239 12537
tri 10239 12439 10337 12537 sw
tri 10337 12439 10435 12537 ne
rect 10435 12439 10789 12537
tri 10789 12439 10887 12537 sw
tri 10887 12439 10985 12537 ne
rect 10985 12439 11339 12537
tri 11339 12439 11437 12537 sw
tri 11437 12439 11535 12537 ne
rect 11535 12439 11889 12537
tri 11889 12439 11987 12537 sw
tri 11987 12439 12085 12537 ne
rect 12085 12439 12439 12537
tri 12439 12439 12537 12537 sw
tri 12537 12439 12635 12537 ne
rect 12635 12439 12989 12537
tri 12989 12439 13087 12537 sw
tri 13087 12439 13185 12537 ne
rect 13185 12439 13539 12537
tri 13539 12439 13637 12537 sw
tri 13637 12439 13735 12537 ne
rect 13735 12439 14089 12537
tri 14089 12439 14187 12537 sw
tri 14187 12439 14285 12537 ne
rect 14285 12439 14639 12537
tri 14639 12439 14737 12537 sw
tri 14737 12439 14835 12537 ne
rect 14835 12439 15189 12537
tri 15189 12439 15287 12537 sw
tri 15287 12439 15385 12537 ne
rect 15385 12439 15739 12537
tri 15739 12439 15837 12537 sw
tri 15837 12439 15935 12537 ne
rect 15935 12439 16289 12537
tri 16289 12439 16387 12537 sw
tri 16387 12439 16485 12537 ne
rect 16485 12439 16839 12537
tri 16839 12439 16937 12537 sw
tri 16937 12439 17035 12537 ne
rect 17035 12439 17389 12537
tri 17389 12439 17487 12537 sw
tri 17487 12439 17585 12537 ne
rect 17585 12439 17939 12537
tri 17939 12439 18037 12537 sw
tri 18037 12439 18135 12537 ne
rect 18135 12439 18489 12537
tri 18489 12439 18587 12537 sw
tri 18587 12439 18685 12537 ne
rect 18685 12439 19039 12537
tri 19039 12439 19137 12537 sw
tri 19137 12439 19235 12537 ne
rect 19235 12439 19589 12537
tri 19589 12439 19687 12537 sw
rect -500 12435 437 12439
rect -500 12315 215 12435
rect 335 12341 437 12435
tri 437 12341 535 12439 sw
tri 535 12341 633 12439 ne
rect 633 12435 987 12439
rect 633 12341 765 12435
rect 335 12315 535 12341
rect -500 12311 535 12315
tri 535 12311 565 12341 sw
tri 633 12311 663 12341 ne
rect 663 12315 765 12341
rect 885 12341 987 12435
tri 987 12341 1085 12439 sw
tri 1085 12341 1183 12439 ne
rect 1183 12435 1537 12439
rect 1183 12341 1315 12435
rect 885 12315 1085 12341
rect 663 12311 1085 12315
tri 1085 12311 1115 12341 sw
tri 1183 12311 1213 12341 ne
rect 1213 12315 1315 12341
rect 1435 12341 1537 12435
tri 1537 12341 1635 12439 sw
tri 1635 12341 1733 12439 ne
rect 1733 12435 2087 12439
rect 1733 12341 1865 12435
rect 1435 12315 1635 12341
rect 1213 12311 1635 12315
tri 1635 12311 1665 12341 sw
tri 1733 12311 1763 12341 ne
rect 1763 12315 1865 12341
rect 1985 12341 2087 12435
tri 2087 12341 2185 12439 sw
tri 2185 12341 2283 12439 ne
rect 2283 12435 2637 12439
rect 2283 12341 2415 12435
rect 1985 12315 2185 12341
rect 1763 12311 2185 12315
tri 2185 12311 2215 12341 sw
tri 2283 12311 2313 12341 ne
rect 2313 12315 2415 12341
rect 2535 12341 2637 12435
tri 2637 12341 2735 12439 sw
tri 2735 12341 2833 12439 ne
rect 2833 12435 3187 12439
rect 2833 12341 2965 12435
rect 2535 12315 2735 12341
rect 2313 12311 2735 12315
tri 2735 12311 2765 12341 sw
tri 2833 12311 2863 12341 ne
rect 2863 12315 2965 12341
rect 3085 12341 3187 12435
tri 3187 12341 3285 12439 sw
tri 3285 12341 3383 12439 ne
rect 3383 12435 3737 12439
rect 3383 12341 3515 12435
rect 3085 12315 3285 12341
rect 2863 12311 3285 12315
tri 3285 12311 3315 12341 sw
tri 3383 12311 3413 12341 ne
rect 3413 12315 3515 12341
rect 3635 12341 3737 12435
tri 3737 12341 3835 12439 sw
tri 3835 12341 3933 12439 ne
rect 3933 12435 4287 12439
rect 3933 12341 4065 12435
rect 3635 12315 3835 12341
rect 3413 12311 3835 12315
tri 3835 12311 3865 12341 sw
tri 3933 12311 3963 12341 ne
rect 3963 12315 4065 12341
rect 4185 12341 4287 12435
tri 4287 12341 4385 12439 sw
tri 4385 12341 4483 12439 ne
rect 4483 12435 4837 12439
rect 4483 12341 4615 12435
rect 4185 12315 4385 12341
rect 3963 12311 4385 12315
tri 4385 12311 4415 12341 sw
tri 4483 12311 4513 12341 ne
rect 4513 12315 4615 12341
rect 4735 12341 4837 12435
tri 4837 12341 4935 12439 sw
tri 4935 12341 5033 12439 ne
rect 5033 12435 5387 12439
rect 5033 12341 5165 12435
rect 4735 12315 4935 12341
rect 4513 12311 4935 12315
tri 4935 12311 4965 12341 sw
tri 5033 12311 5063 12341 ne
rect 5063 12315 5165 12341
rect 5285 12341 5387 12435
tri 5387 12341 5485 12439 sw
tri 5485 12341 5583 12439 ne
rect 5583 12435 5937 12439
rect 5583 12341 5715 12435
rect 5285 12315 5485 12341
rect 5063 12311 5485 12315
tri 5485 12311 5515 12341 sw
tri 5583 12311 5613 12341 ne
rect 5613 12315 5715 12341
rect 5835 12341 5937 12435
tri 5937 12341 6035 12439 sw
tri 6035 12341 6133 12439 ne
rect 6133 12435 6487 12439
rect 6133 12341 6265 12435
rect 5835 12315 6035 12341
rect 5613 12311 6035 12315
tri 6035 12311 6065 12341 sw
tri 6133 12311 6163 12341 ne
rect 6163 12315 6265 12341
rect 6385 12341 6487 12435
tri 6487 12341 6585 12439 sw
tri 6585 12341 6683 12439 ne
rect 6683 12435 7037 12439
rect 6683 12341 6815 12435
rect 6385 12315 6585 12341
rect 6163 12311 6585 12315
tri 6585 12311 6615 12341 sw
tri 6683 12311 6713 12341 ne
rect 6713 12315 6815 12341
rect 6935 12341 7037 12435
tri 7037 12341 7135 12439 sw
tri 7135 12341 7233 12439 ne
rect 7233 12435 7587 12439
rect 7233 12341 7365 12435
rect 6935 12315 7135 12341
rect 6713 12311 7135 12315
tri 7135 12311 7165 12341 sw
tri 7233 12311 7263 12341 ne
rect 7263 12315 7365 12341
rect 7485 12341 7587 12435
tri 7587 12341 7685 12439 sw
tri 7685 12341 7783 12439 ne
rect 7783 12435 8137 12439
rect 7783 12341 7915 12435
rect 7485 12315 7685 12341
rect 7263 12311 7685 12315
tri 7685 12311 7715 12341 sw
tri 7783 12311 7813 12341 ne
rect 7813 12315 7915 12341
rect 8035 12341 8137 12435
tri 8137 12341 8235 12439 sw
tri 8235 12341 8333 12439 ne
rect 8333 12435 8687 12439
rect 8333 12341 8465 12435
rect 8035 12315 8235 12341
rect 7813 12311 8235 12315
tri 8235 12311 8265 12341 sw
tri 8333 12311 8363 12341 ne
rect 8363 12315 8465 12341
rect 8585 12341 8687 12435
tri 8687 12341 8785 12439 sw
tri 8785 12341 8883 12439 ne
rect 8883 12435 9237 12439
rect 8883 12341 9015 12435
rect 8585 12315 8785 12341
rect 8363 12311 8785 12315
tri 8785 12311 8815 12341 sw
tri 8883 12311 8913 12341 ne
rect 8913 12315 9015 12341
rect 9135 12341 9237 12435
tri 9237 12341 9335 12439 sw
tri 9335 12341 9433 12439 ne
rect 9433 12435 9787 12439
rect 9433 12341 9565 12435
rect 9135 12315 9335 12341
rect 8913 12311 9335 12315
tri 9335 12311 9365 12341 sw
tri 9433 12311 9463 12341 ne
rect 9463 12315 9565 12341
rect 9685 12341 9787 12435
tri 9787 12341 9885 12439 sw
tri 9885 12341 9983 12439 ne
rect 9983 12435 10337 12439
rect 9983 12341 10115 12435
rect 9685 12315 9885 12341
rect 9463 12311 9885 12315
tri 9885 12311 9915 12341 sw
tri 9983 12311 10013 12341 ne
rect 10013 12315 10115 12341
rect 10235 12341 10337 12435
tri 10337 12341 10435 12439 sw
tri 10435 12341 10533 12439 ne
rect 10533 12435 10887 12439
rect 10533 12341 10665 12435
rect 10235 12315 10435 12341
rect 10013 12311 10435 12315
tri 10435 12311 10465 12341 sw
tri 10533 12311 10563 12341 ne
rect 10563 12315 10665 12341
rect 10785 12341 10887 12435
tri 10887 12341 10985 12439 sw
tri 10985 12341 11083 12439 ne
rect 11083 12435 11437 12439
rect 11083 12341 11215 12435
rect 10785 12315 10985 12341
rect 10563 12311 10985 12315
tri 10985 12311 11015 12341 sw
tri 11083 12311 11113 12341 ne
rect 11113 12315 11215 12341
rect 11335 12341 11437 12435
tri 11437 12341 11535 12439 sw
tri 11535 12341 11633 12439 ne
rect 11633 12435 11987 12439
rect 11633 12341 11765 12435
rect 11335 12315 11535 12341
rect 11113 12311 11535 12315
tri 11535 12311 11565 12341 sw
tri 11633 12311 11663 12341 ne
rect 11663 12315 11765 12341
rect 11885 12341 11987 12435
tri 11987 12341 12085 12439 sw
tri 12085 12341 12183 12439 ne
rect 12183 12435 12537 12439
rect 12183 12341 12315 12435
rect 11885 12315 12085 12341
rect 11663 12311 12085 12315
tri 12085 12311 12115 12341 sw
tri 12183 12311 12213 12341 ne
rect 12213 12315 12315 12341
rect 12435 12341 12537 12435
tri 12537 12341 12635 12439 sw
tri 12635 12341 12733 12439 ne
rect 12733 12435 13087 12439
rect 12733 12341 12865 12435
rect 12435 12315 12635 12341
rect 12213 12311 12635 12315
tri 12635 12311 12665 12341 sw
tri 12733 12311 12763 12341 ne
rect 12763 12315 12865 12341
rect 12985 12341 13087 12435
tri 13087 12341 13185 12439 sw
tri 13185 12341 13283 12439 ne
rect 13283 12435 13637 12439
rect 13283 12341 13415 12435
rect 12985 12315 13185 12341
rect 12763 12311 13185 12315
tri 13185 12311 13215 12341 sw
tri 13283 12311 13313 12341 ne
rect 13313 12315 13415 12341
rect 13535 12341 13637 12435
tri 13637 12341 13735 12439 sw
tri 13735 12341 13833 12439 ne
rect 13833 12435 14187 12439
rect 13833 12341 13965 12435
rect 13535 12315 13735 12341
rect 13313 12311 13735 12315
tri 13735 12311 13765 12341 sw
tri 13833 12311 13863 12341 ne
rect 13863 12315 13965 12341
rect 14085 12341 14187 12435
tri 14187 12341 14285 12439 sw
tri 14285 12341 14383 12439 ne
rect 14383 12435 14737 12439
rect 14383 12341 14515 12435
rect 14085 12315 14285 12341
rect 13863 12311 14285 12315
tri 14285 12311 14315 12341 sw
tri 14383 12311 14413 12341 ne
rect 14413 12315 14515 12341
rect 14635 12341 14737 12435
tri 14737 12341 14835 12439 sw
tri 14835 12341 14933 12439 ne
rect 14933 12435 15287 12439
rect 14933 12341 15065 12435
rect 14635 12315 14835 12341
rect 14413 12311 14835 12315
tri 14835 12311 14865 12341 sw
tri 14933 12311 14963 12341 ne
rect 14963 12315 15065 12341
rect 15185 12341 15287 12435
tri 15287 12341 15385 12439 sw
tri 15385 12341 15483 12439 ne
rect 15483 12435 15837 12439
rect 15483 12341 15615 12435
rect 15185 12315 15385 12341
rect 14963 12311 15385 12315
tri 15385 12311 15415 12341 sw
tri 15483 12311 15513 12341 ne
rect 15513 12315 15615 12341
rect 15735 12341 15837 12435
tri 15837 12341 15935 12439 sw
tri 15935 12341 16033 12439 ne
rect 16033 12435 16387 12439
rect 16033 12341 16165 12435
rect 15735 12315 15935 12341
rect 15513 12311 15935 12315
tri 15935 12311 15965 12341 sw
tri 16033 12311 16063 12341 ne
rect 16063 12315 16165 12341
rect 16285 12341 16387 12435
tri 16387 12341 16485 12439 sw
tri 16485 12341 16583 12439 ne
rect 16583 12435 16937 12439
rect 16583 12341 16715 12435
rect 16285 12315 16485 12341
rect 16063 12311 16485 12315
tri 16485 12311 16515 12341 sw
tri 16583 12311 16613 12341 ne
rect 16613 12315 16715 12341
rect 16835 12341 16937 12435
tri 16937 12341 17035 12439 sw
tri 17035 12341 17133 12439 ne
rect 17133 12435 17487 12439
rect 17133 12341 17265 12435
rect 16835 12315 17035 12341
rect 16613 12311 17035 12315
tri 17035 12311 17065 12341 sw
tri 17133 12311 17163 12341 ne
rect 17163 12315 17265 12341
rect 17385 12341 17487 12435
tri 17487 12341 17585 12439 sw
tri 17585 12341 17683 12439 ne
rect 17683 12435 18037 12439
rect 17683 12341 17815 12435
rect 17385 12315 17585 12341
rect 17163 12311 17585 12315
tri 17585 12311 17615 12341 sw
tri 17683 12311 17713 12341 ne
rect 17713 12315 17815 12341
rect 17935 12341 18037 12435
tri 18037 12341 18135 12439 sw
tri 18135 12341 18233 12439 ne
rect 18233 12435 18587 12439
rect 18233 12341 18365 12435
rect 17935 12315 18135 12341
rect 17713 12311 18135 12315
tri 18135 12311 18165 12341 sw
tri 18233 12311 18263 12341 ne
rect 18263 12315 18365 12341
rect 18485 12341 18587 12435
tri 18587 12341 18685 12439 sw
tri 18685 12341 18783 12439 ne
rect 18783 12435 19137 12439
rect 18783 12341 18915 12435
rect 18485 12315 18685 12341
rect 18263 12311 18685 12315
tri 18685 12311 18715 12341 sw
tri 18783 12311 18813 12341 ne
rect 18813 12315 18915 12341
rect 19035 12341 19137 12435
tri 19137 12341 19235 12439 sw
tri 19235 12341 19333 12439 ne
rect 19333 12435 20300 12439
rect 19333 12341 19465 12435
rect 19035 12315 19235 12341
rect 18813 12311 19235 12315
tri 19235 12311 19265 12341 sw
tri 19333 12311 19363 12341 ne
rect 19363 12315 19465 12341
rect 19585 12315 20300 12435
rect 19363 12311 20300 12315
tri 113 12213 211 12311 ne
rect 211 12213 565 12311
tri 565 12213 663 12311 sw
tri 663 12213 761 12311 ne
rect 761 12213 1115 12311
tri 1115 12213 1213 12311 sw
tri 1213 12213 1311 12311 ne
rect 1311 12213 1665 12311
tri 1665 12213 1763 12311 sw
tri 1763 12213 1861 12311 ne
rect 1861 12213 2215 12311
tri 2215 12213 2313 12311 sw
tri 2313 12213 2411 12311 ne
rect 2411 12213 2765 12311
tri 2765 12213 2863 12311 sw
tri 2863 12213 2961 12311 ne
rect 2961 12213 3315 12311
tri 3315 12213 3413 12311 sw
tri 3413 12213 3511 12311 ne
rect 3511 12213 3865 12311
tri 3865 12213 3963 12311 sw
tri 3963 12213 4061 12311 ne
rect 4061 12213 4415 12311
tri 4415 12213 4513 12311 sw
tri 4513 12213 4611 12311 ne
rect 4611 12213 4965 12311
tri 4965 12213 5063 12311 sw
tri 5063 12213 5161 12311 ne
rect 5161 12213 5515 12311
tri 5515 12213 5613 12311 sw
tri 5613 12213 5711 12311 ne
rect 5711 12213 6065 12311
tri 6065 12213 6163 12311 sw
tri 6163 12213 6261 12311 ne
rect 6261 12213 6615 12311
tri 6615 12213 6713 12311 sw
tri 6713 12213 6811 12311 ne
rect 6811 12213 7165 12311
tri 7165 12213 7263 12311 sw
tri 7263 12213 7361 12311 ne
rect 7361 12213 7715 12311
tri 7715 12213 7813 12311 sw
tri 7813 12213 7911 12311 ne
rect 7911 12213 8265 12311
tri 8265 12213 8363 12311 sw
tri 8363 12213 8461 12311 ne
rect 8461 12213 8815 12311
tri 8815 12213 8913 12311 sw
tri 8913 12213 9011 12311 ne
rect 9011 12213 9365 12311
tri 9365 12213 9463 12311 sw
tri 9463 12213 9561 12311 ne
rect 9561 12213 9915 12311
tri 9915 12213 10013 12311 sw
tri 10013 12213 10111 12311 ne
rect 10111 12213 10465 12311
tri 10465 12213 10563 12311 sw
tri 10563 12213 10661 12311 ne
rect 10661 12213 11015 12311
tri 11015 12213 11113 12311 sw
tri 11113 12213 11211 12311 ne
rect 11211 12213 11565 12311
tri 11565 12213 11663 12311 sw
tri 11663 12213 11761 12311 ne
rect 11761 12213 12115 12311
tri 12115 12213 12213 12311 sw
tri 12213 12213 12311 12311 ne
rect 12311 12213 12665 12311
tri 12665 12213 12763 12311 sw
tri 12763 12213 12861 12311 ne
rect 12861 12213 13215 12311
tri 13215 12213 13313 12311 sw
tri 13313 12213 13411 12311 ne
rect 13411 12213 13765 12311
tri 13765 12213 13863 12311 sw
tri 13863 12213 13961 12311 ne
rect 13961 12213 14315 12311
tri 14315 12213 14413 12311 sw
tri 14413 12213 14511 12311 ne
rect 14511 12213 14865 12311
tri 14865 12213 14963 12311 sw
tri 14963 12213 15061 12311 ne
rect 15061 12213 15415 12311
tri 15415 12213 15513 12311 sw
tri 15513 12213 15611 12311 ne
rect 15611 12213 15965 12311
tri 15965 12213 16063 12311 sw
tri 16063 12213 16161 12311 ne
rect 16161 12213 16515 12311
tri 16515 12213 16613 12311 sw
tri 16613 12213 16711 12311 ne
rect 16711 12213 17065 12311
tri 17065 12213 17163 12311 sw
tri 17163 12213 17261 12311 ne
rect 17261 12213 17615 12311
tri 17615 12213 17713 12311 sw
tri 17713 12213 17811 12311 ne
rect 17811 12213 18165 12311
tri 18165 12213 18263 12311 sw
tri 18263 12213 18361 12311 ne
rect 18361 12213 18715 12311
tri 18715 12213 18813 12311 sw
tri 18813 12213 18911 12311 ne
rect 18911 12213 19265 12311
tri 19265 12213 19363 12311 sw
tri 19363 12213 19461 12311 ne
rect 19461 12213 20300 12311
rect -2000 12183 113 12213
tri 113 12183 143 12213 sw
tri 211 12183 241 12213 ne
rect 241 12183 663 12213
tri 663 12183 693 12213 sw
tri 761 12183 791 12213 ne
rect 791 12183 1213 12213
tri 1213 12183 1243 12213 sw
tri 1311 12183 1341 12213 ne
rect 1341 12183 1763 12213
tri 1763 12183 1793 12213 sw
tri 1861 12183 1891 12213 ne
rect 1891 12183 2313 12213
tri 2313 12183 2343 12213 sw
tri 2411 12183 2441 12213 ne
rect 2441 12183 2863 12213
tri 2863 12183 2893 12213 sw
tri 2961 12183 2991 12213 ne
rect 2991 12183 3413 12213
tri 3413 12183 3443 12213 sw
tri 3511 12183 3541 12213 ne
rect 3541 12183 3963 12213
tri 3963 12183 3993 12213 sw
tri 4061 12183 4091 12213 ne
rect 4091 12183 4513 12213
tri 4513 12183 4543 12213 sw
tri 4611 12183 4641 12213 ne
rect 4641 12183 5063 12213
tri 5063 12183 5093 12213 sw
tri 5161 12183 5191 12213 ne
rect 5191 12183 5613 12213
tri 5613 12183 5643 12213 sw
tri 5711 12183 5741 12213 ne
rect 5741 12183 6163 12213
tri 6163 12183 6193 12213 sw
tri 6261 12183 6291 12213 ne
rect 6291 12183 6713 12213
tri 6713 12183 6743 12213 sw
tri 6811 12183 6841 12213 ne
rect 6841 12183 7263 12213
tri 7263 12183 7293 12213 sw
tri 7361 12183 7391 12213 ne
rect 7391 12183 7813 12213
tri 7813 12183 7843 12213 sw
tri 7911 12183 7941 12213 ne
rect 7941 12183 8363 12213
tri 8363 12183 8393 12213 sw
tri 8461 12183 8491 12213 ne
rect 8491 12183 8913 12213
tri 8913 12183 8943 12213 sw
tri 9011 12183 9041 12213 ne
rect 9041 12183 9463 12213
tri 9463 12183 9493 12213 sw
tri 9561 12183 9591 12213 ne
rect 9591 12183 10013 12213
tri 10013 12183 10043 12213 sw
tri 10111 12183 10141 12213 ne
rect 10141 12183 10563 12213
tri 10563 12183 10593 12213 sw
tri 10661 12183 10691 12213 ne
rect 10691 12183 11113 12213
tri 11113 12183 11143 12213 sw
tri 11211 12183 11241 12213 ne
rect 11241 12183 11663 12213
tri 11663 12183 11693 12213 sw
tri 11761 12183 11791 12213 ne
rect 11791 12183 12213 12213
tri 12213 12183 12243 12213 sw
tri 12311 12183 12341 12213 ne
rect 12341 12183 12763 12213
tri 12763 12183 12793 12213 sw
tri 12861 12183 12891 12213 ne
rect 12891 12183 13313 12213
tri 13313 12183 13343 12213 sw
tri 13411 12183 13441 12213 ne
rect 13441 12183 13863 12213
tri 13863 12183 13893 12213 sw
tri 13961 12183 13991 12213 ne
rect 13991 12183 14413 12213
tri 14413 12183 14443 12213 sw
tri 14511 12183 14541 12213 ne
rect 14541 12183 14963 12213
tri 14963 12183 14993 12213 sw
tri 15061 12183 15091 12213 ne
rect 15091 12183 15513 12213
tri 15513 12183 15543 12213 sw
tri 15611 12183 15641 12213 ne
rect 15641 12183 16063 12213
tri 16063 12183 16093 12213 sw
tri 16161 12183 16191 12213 ne
rect 16191 12183 16613 12213
tri 16613 12183 16643 12213 sw
tri 16711 12183 16741 12213 ne
rect 16741 12183 17163 12213
tri 17163 12183 17193 12213 sw
tri 17261 12183 17291 12213 ne
rect 17291 12183 17713 12213
tri 17713 12183 17743 12213 sw
tri 17811 12183 17841 12213 ne
rect 17841 12183 18263 12213
tri 18263 12183 18293 12213 sw
tri 18361 12183 18391 12213 ne
rect 18391 12183 18813 12213
tri 18813 12183 18843 12213 sw
tri 18911 12183 18941 12213 ne
rect 18941 12183 19363 12213
tri 19363 12183 19393 12213 sw
tri 19461 12183 19491 12213 ne
rect 19491 12183 20300 12213
rect -2000 12085 143 12183
tri 143 12085 241 12183 sw
tri 241 12085 339 12183 ne
rect 339 12085 693 12183
tri 693 12085 791 12183 sw
tri 791 12085 889 12183 ne
rect 889 12085 1243 12183
tri 1243 12085 1341 12183 sw
tri 1341 12085 1439 12183 ne
rect 1439 12085 1793 12183
tri 1793 12085 1891 12183 sw
tri 1891 12085 1989 12183 ne
rect 1989 12085 2343 12183
tri 2343 12085 2441 12183 sw
tri 2441 12085 2539 12183 ne
rect 2539 12085 2893 12183
tri 2893 12085 2991 12183 sw
tri 2991 12085 3089 12183 ne
rect 3089 12085 3443 12183
tri 3443 12085 3541 12183 sw
tri 3541 12085 3639 12183 ne
rect 3639 12085 3993 12183
tri 3993 12085 4091 12183 sw
tri 4091 12085 4189 12183 ne
rect 4189 12085 4543 12183
tri 4543 12085 4641 12183 sw
tri 4641 12085 4739 12183 ne
rect 4739 12085 5093 12183
tri 5093 12085 5191 12183 sw
tri 5191 12085 5289 12183 ne
rect 5289 12085 5643 12183
tri 5643 12085 5741 12183 sw
tri 5741 12085 5839 12183 ne
rect 5839 12085 6193 12183
tri 6193 12085 6291 12183 sw
tri 6291 12085 6389 12183 ne
rect 6389 12085 6743 12183
tri 6743 12085 6841 12183 sw
tri 6841 12085 6939 12183 ne
rect 6939 12085 7293 12183
tri 7293 12085 7391 12183 sw
tri 7391 12085 7489 12183 ne
rect 7489 12085 7843 12183
tri 7843 12085 7941 12183 sw
tri 7941 12085 8039 12183 ne
rect 8039 12085 8393 12183
tri 8393 12085 8491 12183 sw
tri 8491 12085 8589 12183 ne
rect 8589 12085 8943 12183
tri 8943 12085 9041 12183 sw
tri 9041 12085 9139 12183 ne
rect 9139 12085 9493 12183
tri 9493 12085 9591 12183 sw
tri 9591 12085 9689 12183 ne
rect 9689 12085 10043 12183
tri 10043 12085 10141 12183 sw
tri 10141 12085 10239 12183 ne
rect 10239 12085 10593 12183
tri 10593 12085 10691 12183 sw
tri 10691 12085 10789 12183 ne
rect 10789 12085 11143 12183
tri 11143 12085 11241 12183 sw
tri 11241 12085 11339 12183 ne
rect 11339 12085 11693 12183
tri 11693 12085 11791 12183 sw
tri 11791 12085 11889 12183 ne
rect 11889 12085 12243 12183
tri 12243 12085 12341 12183 sw
tri 12341 12085 12439 12183 ne
rect 12439 12085 12793 12183
tri 12793 12085 12891 12183 sw
tri 12891 12085 12989 12183 ne
rect 12989 12085 13343 12183
tri 13343 12085 13441 12183 sw
tri 13441 12085 13539 12183 ne
rect 13539 12085 13893 12183
tri 13893 12085 13991 12183 sw
tri 13991 12085 14089 12183 ne
rect 14089 12085 14443 12183
tri 14443 12085 14541 12183 sw
tri 14541 12085 14639 12183 ne
rect 14639 12085 14993 12183
tri 14993 12085 15091 12183 sw
tri 15091 12085 15189 12183 ne
rect 15189 12085 15543 12183
tri 15543 12085 15641 12183 sw
tri 15641 12085 15739 12183 ne
rect 15739 12085 16093 12183
tri 16093 12085 16191 12183 sw
tri 16191 12085 16289 12183 ne
rect 16289 12085 16643 12183
tri 16643 12085 16741 12183 sw
tri 16741 12085 16839 12183 ne
rect 16839 12085 17193 12183
tri 17193 12085 17291 12183 sw
tri 17291 12085 17389 12183 ne
rect 17389 12085 17743 12183
tri 17743 12085 17841 12183 sw
tri 17841 12085 17939 12183 ne
rect 17939 12085 18293 12183
tri 18293 12085 18391 12183 sw
tri 18391 12085 18489 12183 ne
rect 18489 12085 18843 12183
tri 18843 12085 18941 12183 sw
tri 18941 12085 19039 12183 ne
rect 19039 12085 19393 12183
tri 19393 12085 19491 12183 sw
tri 19491 12085 19589 12183 ne
rect 19589 12085 20300 12183
rect -2000 11987 241 12085
tri 241 11987 339 12085 sw
tri 339 11987 437 12085 ne
rect 437 11987 791 12085
tri 791 11987 889 12085 sw
tri 889 11987 987 12085 ne
rect 987 11987 1341 12085
tri 1341 11987 1439 12085 sw
tri 1439 11987 1537 12085 ne
rect 1537 11987 1891 12085
tri 1891 11987 1989 12085 sw
tri 1989 11987 2087 12085 ne
rect 2087 11987 2441 12085
tri 2441 11987 2539 12085 sw
tri 2539 11987 2637 12085 ne
rect 2637 11987 2991 12085
tri 2991 11987 3089 12085 sw
tri 3089 11987 3187 12085 ne
rect 3187 11987 3541 12085
tri 3541 11987 3639 12085 sw
tri 3639 11987 3737 12085 ne
rect 3737 11987 4091 12085
tri 4091 11987 4189 12085 sw
tri 4189 11987 4287 12085 ne
rect 4287 11987 4641 12085
tri 4641 11987 4739 12085 sw
tri 4739 11987 4837 12085 ne
rect 4837 11987 5191 12085
tri 5191 11987 5289 12085 sw
tri 5289 11987 5387 12085 ne
rect 5387 11987 5741 12085
tri 5741 11987 5839 12085 sw
tri 5839 11987 5937 12085 ne
rect 5937 11987 6291 12085
tri 6291 11987 6389 12085 sw
tri 6389 11987 6487 12085 ne
rect 6487 11987 6841 12085
tri 6841 11987 6939 12085 sw
tri 6939 11987 7037 12085 ne
rect 7037 11987 7391 12085
tri 7391 11987 7489 12085 sw
tri 7489 11987 7587 12085 ne
rect 7587 11987 7941 12085
tri 7941 11987 8039 12085 sw
tri 8039 11987 8137 12085 ne
rect 8137 11987 8491 12085
tri 8491 11987 8589 12085 sw
tri 8589 11987 8687 12085 ne
rect 8687 11987 9041 12085
tri 9041 11987 9139 12085 sw
tri 9139 11987 9237 12085 ne
rect 9237 11987 9591 12085
tri 9591 11987 9689 12085 sw
tri 9689 11987 9787 12085 ne
rect 9787 11987 10141 12085
tri 10141 11987 10239 12085 sw
tri 10239 11987 10337 12085 ne
rect 10337 11987 10691 12085
tri 10691 11987 10789 12085 sw
tri 10789 11987 10887 12085 ne
rect 10887 11987 11241 12085
tri 11241 11987 11339 12085 sw
tri 11339 11987 11437 12085 ne
rect 11437 11987 11791 12085
tri 11791 11987 11889 12085 sw
tri 11889 11987 11987 12085 ne
rect 11987 11987 12341 12085
tri 12341 11987 12439 12085 sw
tri 12439 11987 12537 12085 ne
rect 12537 11987 12891 12085
tri 12891 11987 12989 12085 sw
tri 12989 11987 13087 12085 ne
rect 13087 11987 13441 12085
tri 13441 11987 13539 12085 sw
tri 13539 11987 13637 12085 ne
rect 13637 11987 13991 12085
tri 13991 11987 14089 12085 sw
tri 14089 11987 14187 12085 ne
rect 14187 11987 14541 12085
tri 14541 11987 14639 12085 sw
tri 14639 11987 14737 12085 ne
rect 14737 11987 15091 12085
tri 15091 11987 15189 12085 sw
tri 15189 11987 15287 12085 ne
rect 15287 11987 15641 12085
tri 15641 11987 15739 12085 sw
tri 15739 11987 15837 12085 ne
rect 15837 11987 16191 12085
tri 16191 11987 16289 12085 sw
tri 16289 11987 16387 12085 ne
rect 16387 11987 16741 12085
tri 16741 11987 16839 12085 sw
tri 16839 11987 16937 12085 ne
rect 16937 11987 17291 12085
tri 17291 11987 17389 12085 sw
tri 17389 11987 17487 12085 ne
rect 17487 11987 17841 12085
tri 17841 11987 17939 12085 sw
tri 17939 11987 18037 12085 ne
rect 18037 11987 18391 12085
tri 18391 11987 18489 12085 sw
tri 18489 11987 18587 12085 ne
rect 18587 11987 18941 12085
tri 18941 11987 19039 12085 sw
tri 19039 11987 19137 12085 ne
rect 19137 11987 19491 12085
tri 19491 11987 19589 12085 sw
tri 19589 11987 19687 12085 ne
rect 19687 11987 20300 12085
rect -2000 11889 339 11987
tri 339 11889 437 11987 sw
tri 437 11889 535 11987 ne
rect 535 11889 889 11987
tri 889 11889 987 11987 sw
tri 987 11889 1085 11987 ne
rect 1085 11889 1439 11987
tri 1439 11889 1537 11987 sw
tri 1537 11889 1635 11987 ne
rect 1635 11889 1989 11987
tri 1989 11889 2087 11987 sw
tri 2087 11889 2185 11987 ne
rect 2185 11889 2539 11987
tri 2539 11889 2637 11987 sw
tri 2637 11889 2735 11987 ne
rect 2735 11889 3089 11987
tri 3089 11889 3187 11987 sw
tri 3187 11889 3285 11987 ne
rect 3285 11889 3639 11987
tri 3639 11889 3737 11987 sw
tri 3737 11889 3835 11987 ne
rect 3835 11889 4189 11987
tri 4189 11889 4287 11987 sw
tri 4287 11889 4385 11987 ne
rect 4385 11889 4739 11987
tri 4739 11889 4837 11987 sw
tri 4837 11889 4935 11987 ne
rect 4935 11889 5289 11987
tri 5289 11889 5387 11987 sw
tri 5387 11889 5485 11987 ne
rect 5485 11889 5839 11987
tri 5839 11889 5937 11987 sw
tri 5937 11889 6035 11987 ne
rect 6035 11889 6389 11987
tri 6389 11889 6487 11987 sw
tri 6487 11889 6585 11987 ne
rect 6585 11889 6939 11987
tri 6939 11889 7037 11987 sw
tri 7037 11889 7135 11987 ne
rect 7135 11889 7489 11987
tri 7489 11889 7587 11987 sw
tri 7587 11889 7685 11987 ne
rect 7685 11889 8039 11987
tri 8039 11889 8137 11987 sw
tri 8137 11889 8235 11987 ne
rect 8235 11889 8589 11987
tri 8589 11889 8687 11987 sw
tri 8687 11889 8785 11987 ne
rect 8785 11889 9139 11987
tri 9139 11889 9237 11987 sw
tri 9237 11889 9335 11987 ne
rect 9335 11889 9689 11987
tri 9689 11889 9787 11987 sw
tri 9787 11889 9885 11987 ne
rect 9885 11889 10239 11987
tri 10239 11889 10337 11987 sw
tri 10337 11889 10435 11987 ne
rect 10435 11889 10789 11987
tri 10789 11889 10887 11987 sw
tri 10887 11889 10985 11987 ne
rect 10985 11889 11339 11987
tri 11339 11889 11437 11987 sw
tri 11437 11889 11535 11987 ne
rect 11535 11889 11889 11987
tri 11889 11889 11987 11987 sw
tri 11987 11889 12085 11987 ne
rect 12085 11889 12439 11987
tri 12439 11889 12537 11987 sw
tri 12537 11889 12635 11987 ne
rect 12635 11889 12989 11987
tri 12989 11889 13087 11987 sw
tri 13087 11889 13185 11987 ne
rect 13185 11889 13539 11987
tri 13539 11889 13637 11987 sw
tri 13637 11889 13735 11987 ne
rect 13735 11889 14089 11987
tri 14089 11889 14187 11987 sw
tri 14187 11889 14285 11987 ne
rect 14285 11889 14639 11987
tri 14639 11889 14737 11987 sw
tri 14737 11889 14835 11987 ne
rect 14835 11889 15189 11987
tri 15189 11889 15287 11987 sw
tri 15287 11889 15385 11987 ne
rect 15385 11889 15739 11987
tri 15739 11889 15837 11987 sw
tri 15837 11889 15935 11987 ne
rect 15935 11889 16289 11987
tri 16289 11889 16387 11987 sw
tri 16387 11889 16485 11987 ne
rect 16485 11889 16839 11987
tri 16839 11889 16937 11987 sw
tri 16937 11889 17035 11987 ne
rect 17035 11889 17389 11987
tri 17389 11889 17487 11987 sw
tri 17487 11889 17585 11987 ne
rect 17585 11889 17939 11987
tri 17939 11889 18037 11987 sw
tri 18037 11889 18135 11987 ne
rect 18135 11889 18489 11987
tri 18489 11889 18587 11987 sw
tri 18587 11889 18685 11987 ne
rect 18685 11889 19039 11987
tri 19039 11889 19137 11987 sw
tri 19137 11889 19235 11987 ne
rect 19235 11889 19589 11987
tri 19589 11889 19687 11987 sw
rect 20800 11889 21800 12537
rect -2000 11885 437 11889
rect -2000 11765 215 11885
rect 335 11791 437 11885
tri 437 11791 535 11889 sw
tri 535 11791 633 11889 ne
rect 633 11885 987 11889
rect 633 11791 765 11885
rect 335 11765 535 11791
rect -2000 11761 535 11765
rect -2000 11113 -1000 11761
tri 113 11663 211 11761 ne
rect 211 11713 535 11761
tri 535 11713 613 11791 sw
tri 633 11713 711 11791 ne
rect 711 11765 765 11791
rect 885 11791 987 11885
tri 987 11791 1085 11889 sw
tri 1085 11791 1183 11889 ne
rect 1183 11885 1537 11889
rect 1183 11791 1315 11885
rect 885 11765 1085 11791
rect 711 11713 1085 11765
tri 1085 11713 1163 11791 sw
tri 1183 11713 1261 11791 ne
rect 1261 11765 1315 11791
rect 1435 11791 1537 11885
tri 1537 11791 1635 11889 sw
tri 1635 11791 1733 11889 ne
rect 1733 11885 2087 11889
rect 1733 11791 1865 11885
rect 1435 11765 1635 11791
rect 1261 11713 1635 11765
tri 1635 11713 1713 11791 sw
tri 1733 11713 1811 11791 ne
rect 1811 11765 1865 11791
rect 1985 11791 2087 11885
tri 2087 11791 2185 11889 sw
tri 2185 11791 2283 11889 ne
rect 2283 11885 2637 11889
rect 2283 11791 2415 11885
rect 1985 11765 2185 11791
rect 1811 11713 2185 11765
tri 2185 11713 2263 11791 sw
tri 2283 11713 2361 11791 ne
rect 2361 11765 2415 11791
rect 2535 11791 2637 11885
tri 2637 11791 2735 11889 sw
tri 2735 11791 2833 11889 ne
rect 2833 11885 3187 11889
rect 2833 11791 2965 11885
rect 2535 11765 2735 11791
rect 2361 11713 2735 11765
tri 2735 11713 2813 11791 sw
tri 2833 11713 2911 11791 ne
rect 2911 11765 2965 11791
rect 3085 11791 3187 11885
tri 3187 11791 3285 11889 sw
tri 3285 11791 3383 11889 ne
rect 3383 11885 3737 11889
rect 3383 11791 3515 11885
rect 3085 11765 3285 11791
rect 2911 11713 3285 11765
tri 3285 11713 3363 11791 sw
tri 3383 11713 3461 11791 ne
rect 3461 11765 3515 11791
rect 3635 11791 3737 11885
tri 3737 11791 3835 11889 sw
tri 3835 11791 3933 11889 ne
rect 3933 11885 4287 11889
rect 3933 11791 4065 11885
rect 3635 11765 3835 11791
rect 3461 11713 3835 11765
tri 3835 11713 3913 11791 sw
tri 3933 11713 4011 11791 ne
rect 4011 11765 4065 11791
rect 4185 11791 4287 11885
tri 4287 11791 4385 11889 sw
tri 4385 11791 4483 11889 ne
rect 4483 11885 4837 11889
rect 4483 11791 4615 11885
rect 4185 11765 4385 11791
rect 4011 11713 4385 11765
tri 4385 11713 4463 11791 sw
tri 4483 11713 4561 11791 ne
rect 4561 11765 4615 11791
rect 4735 11791 4837 11885
tri 4837 11791 4935 11889 sw
tri 4935 11791 5033 11889 ne
rect 5033 11885 5387 11889
rect 5033 11791 5165 11885
rect 4735 11765 4935 11791
rect 4561 11713 4935 11765
tri 4935 11713 5013 11791 sw
tri 5033 11713 5111 11791 ne
rect 5111 11765 5165 11791
rect 5285 11791 5387 11885
tri 5387 11791 5485 11889 sw
tri 5485 11791 5583 11889 ne
rect 5583 11885 5937 11889
rect 5583 11791 5715 11885
rect 5285 11765 5485 11791
rect 5111 11713 5485 11765
tri 5485 11713 5563 11791 sw
tri 5583 11713 5661 11791 ne
rect 5661 11765 5715 11791
rect 5835 11791 5937 11885
tri 5937 11791 6035 11889 sw
tri 6035 11791 6133 11889 ne
rect 6133 11885 6487 11889
rect 6133 11791 6265 11885
rect 5835 11765 6035 11791
rect 5661 11713 6035 11765
tri 6035 11713 6113 11791 sw
tri 6133 11713 6211 11791 ne
rect 6211 11765 6265 11791
rect 6385 11791 6487 11885
tri 6487 11791 6585 11889 sw
tri 6585 11791 6683 11889 ne
rect 6683 11885 7037 11889
rect 6683 11791 6815 11885
rect 6385 11765 6585 11791
rect 6211 11713 6585 11765
tri 6585 11713 6663 11791 sw
tri 6683 11713 6761 11791 ne
rect 6761 11765 6815 11791
rect 6935 11791 7037 11885
tri 7037 11791 7135 11889 sw
tri 7135 11791 7233 11889 ne
rect 7233 11885 7587 11889
rect 7233 11791 7365 11885
rect 6935 11765 7135 11791
rect 6761 11713 7135 11765
tri 7135 11713 7213 11791 sw
tri 7233 11713 7311 11791 ne
rect 7311 11765 7365 11791
rect 7485 11791 7587 11885
tri 7587 11791 7685 11889 sw
tri 7685 11791 7783 11889 ne
rect 7783 11885 8137 11889
rect 7783 11791 7915 11885
rect 7485 11765 7685 11791
rect 7311 11713 7685 11765
tri 7685 11713 7763 11791 sw
tri 7783 11713 7861 11791 ne
rect 7861 11765 7915 11791
rect 8035 11791 8137 11885
tri 8137 11791 8235 11889 sw
tri 8235 11791 8333 11889 ne
rect 8333 11885 8687 11889
rect 8333 11791 8465 11885
rect 8035 11765 8235 11791
rect 7861 11713 8235 11765
tri 8235 11713 8313 11791 sw
tri 8333 11713 8411 11791 ne
rect 8411 11765 8465 11791
rect 8585 11791 8687 11885
tri 8687 11791 8785 11889 sw
tri 8785 11791 8883 11889 ne
rect 8883 11885 9237 11889
rect 8883 11791 9015 11885
rect 8585 11765 8785 11791
rect 8411 11713 8785 11765
tri 8785 11713 8863 11791 sw
tri 8883 11713 8961 11791 ne
rect 8961 11765 9015 11791
rect 9135 11791 9237 11885
tri 9237 11791 9335 11889 sw
tri 9335 11791 9433 11889 ne
rect 9433 11885 9787 11889
rect 9433 11791 9565 11885
rect 9135 11765 9335 11791
rect 8961 11713 9335 11765
tri 9335 11713 9413 11791 sw
tri 9433 11713 9511 11791 ne
rect 9511 11765 9565 11791
rect 9685 11791 9787 11885
tri 9787 11791 9885 11889 sw
tri 9885 11791 9983 11889 ne
rect 9983 11885 10337 11889
rect 9983 11791 10115 11885
rect 9685 11765 9885 11791
rect 9511 11713 9885 11765
tri 9885 11713 9963 11791 sw
tri 9983 11713 10061 11791 ne
rect 10061 11765 10115 11791
rect 10235 11791 10337 11885
tri 10337 11791 10435 11889 sw
tri 10435 11791 10533 11889 ne
rect 10533 11885 10887 11889
rect 10533 11791 10665 11885
rect 10235 11765 10435 11791
rect 10061 11713 10435 11765
tri 10435 11713 10513 11791 sw
tri 10533 11713 10611 11791 ne
rect 10611 11765 10665 11791
rect 10785 11791 10887 11885
tri 10887 11791 10985 11889 sw
tri 10985 11791 11083 11889 ne
rect 11083 11885 11437 11889
rect 11083 11791 11215 11885
rect 10785 11765 10985 11791
rect 10611 11713 10985 11765
tri 10985 11713 11063 11791 sw
tri 11083 11713 11161 11791 ne
rect 11161 11765 11215 11791
rect 11335 11791 11437 11885
tri 11437 11791 11535 11889 sw
tri 11535 11791 11633 11889 ne
rect 11633 11885 11987 11889
rect 11633 11791 11765 11885
rect 11335 11765 11535 11791
rect 11161 11713 11535 11765
tri 11535 11713 11613 11791 sw
tri 11633 11713 11711 11791 ne
rect 11711 11765 11765 11791
rect 11885 11791 11987 11885
tri 11987 11791 12085 11889 sw
tri 12085 11791 12183 11889 ne
rect 12183 11885 12537 11889
rect 12183 11791 12315 11885
rect 11885 11765 12085 11791
rect 11711 11713 12085 11765
tri 12085 11713 12163 11791 sw
tri 12183 11713 12261 11791 ne
rect 12261 11765 12315 11791
rect 12435 11791 12537 11885
tri 12537 11791 12635 11889 sw
tri 12635 11791 12733 11889 ne
rect 12733 11885 13087 11889
rect 12733 11791 12865 11885
rect 12435 11765 12635 11791
rect 12261 11713 12635 11765
tri 12635 11713 12713 11791 sw
tri 12733 11713 12811 11791 ne
rect 12811 11765 12865 11791
rect 12985 11791 13087 11885
tri 13087 11791 13185 11889 sw
tri 13185 11791 13283 11889 ne
rect 13283 11885 13637 11889
rect 13283 11791 13415 11885
rect 12985 11765 13185 11791
rect 12811 11713 13185 11765
tri 13185 11713 13263 11791 sw
tri 13283 11713 13361 11791 ne
rect 13361 11765 13415 11791
rect 13535 11791 13637 11885
tri 13637 11791 13735 11889 sw
tri 13735 11791 13833 11889 ne
rect 13833 11885 14187 11889
rect 13833 11791 13965 11885
rect 13535 11765 13735 11791
rect 13361 11713 13735 11765
tri 13735 11713 13813 11791 sw
tri 13833 11713 13911 11791 ne
rect 13911 11765 13965 11791
rect 14085 11791 14187 11885
tri 14187 11791 14285 11889 sw
tri 14285 11791 14383 11889 ne
rect 14383 11885 14737 11889
rect 14383 11791 14515 11885
rect 14085 11765 14285 11791
rect 13911 11713 14285 11765
tri 14285 11713 14363 11791 sw
tri 14383 11713 14461 11791 ne
rect 14461 11765 14515 11791
rect 14635 11791 14737 11885
tri 14737 11791 14835 11889 sw
tri 14835 11791 14933 11889 ne
rect 14933 11885 15287 11889
rect 14933 11791 15065 11885
rect 14635 11765 14835 11791
rect 14461 11713 14835 11765
tri 14835 11713 14913 11791 sw
tri 14933 11713 15011 11791 ne
rect 15011 11765 15065 11791
rect 15185 11791 15287 11885
tri 15287 11791 15385 11889 sw
tri 15385 11791 15483 11889 ne
rect 15483 11885 15837 11889
rect 15483 11791 15615 11885
rect 15185 11765 15385 11791
rect 15011 11713 15385 11765
tri 15385 11713 15463 11791 sw
tri 15483 11713 15561 11791 ne
rect 15561 11765 15615 11791
rect 15735 11791 15837 11885
tri 15837 11791 15935 11889 sw
tri 15935 11791 16033 11889 ne
rect 16033 11885 16387 11889
rect 16033 11791 16165 11885
rect 15735 11765 15935 11791
rect 15561 11713 15935 11765
tri 15935 11713 16013 11791 sw
tri 16033 11713 16111 11791 ne
rect 16111 11765 16165 11791
rect 16285 11791 16387 11885
tri 16387 11791 16485 11889 sw
tri 16485 11791 16583 11889 ne
rect 16583 11885 16937 11889
rect 16583 11791 16715 11885
rect 16285 11765 16485 11791
rect 16111 11713 16485 11765
tri 16485 11713 16563 11791 sw
tri 16583 11713 16661 11791 ne
rect 16661 11765 16715 11791
rect 16835 11791 16937 11885
tri 16937 11791 17035 11889 sw
tri 17035 11791 17133 11889 ne
rect 17133 11885 17487 11889
rect 17133 11791 17265 11885
rect 16835 11765 17035 11791
rect 16661 11713 17035 11765
tri 17035 11713 17113 11791 sw
tri 17133 11713 17211 11791 ne
rect 17211 11765 17265 11791
rect 17385 11791 17487 11885
tri 17487 11791 17585 11889 sw
tri 17585 11791 17683 11889 ne
rect 17683 11885 18037 11889
rect 17683 11791 17815 11885
rect 17385 11765 17585 11791
rect 17211 11713 17585 11765
tri 17585 11713 17663 11791 sw
tri 17683 11713 17761 11791 ne
rect 17761 11765 17815 11791
rect 17935 11791 18037 11885
tri 18037 11791 18135 11889 sw
tri 18135 11791 18233 11889 ne
rect 18233 11885 18587 11889
rect 18233 11791 18365 11885
rect 17935 11765 18135 11791
rect 17761 11713 18135 11765
tri 18135 11713 18213 11791 sw
tri 18233 11713 18311 11791 ne
rect 18311 11765 18365 11791
rect 18485 11791 18587 11885
tri 18587 11791 18685 11889 sw
tri 18685 11791 18783 11889 ne
rect 18783 11885 19137 11889
rect 18783 11791 18915 11885
rect 18485 11765 18685 11791
rect 18311 11713 18685 11765
tri 18685 11713 18763 11791 sw
tri 18783 11713 18861 11791 ne
rect 18861 11765 18915 11791
rect 19035 11791 19137 11885
tri 19137 11791 19235 11889 sw
tri 19235 11791 19333 11889 ne
rect 19333 11885 21800 11889
rect 19333 11791 19465 11885
rect 19035 11765 19235 11791
rect 18861 11713 19235 11765
tri 19235 11713 19313 11791 sw
tri 19333 11713 19411 11791 ne
rect 19411 11765 19465 11791
rect 19585 11765 21800 11885
rect 19411 11713 21800 11765
rect 211 11663 613 11713
rect -500 11613 113 11663
tri 113 11613 163 11663 sw
tri 211 11613 261 11663 ne
rect 261 11633 613 11663
tri 613 11633 693 11713 sw
tri 711 11633 791 11713 ne
rect 791 11633 1163 11713
tri 1163 11633 1243 11713 sw
tri 1261 11633 1341 11713 ne
rect 1341 11633 1713 11713
tri 1713 11633 1793 11713 sw
tri 1811 11633 1891 11713 ne
rect 1891 11633 2263 11713
tri 2263 11633 2343 11713 sw
tri 2361 11633 2441 11713 ne
rect 2441 11633 2813 11713
tri 2813 11633 2893 11713 sw
tri 2911 11633 2991 11713 ne
rect 2991 11633 3363 11713
tri 3363 11633 3443 11713 sw
tri 3461 11633 3541 11713 ne
rect 3541 11633 3913 11713
tri 3913 11633 3993 11713 sw
tri 4011 11633 4091 11713 ne
rect 4091 11633 4463 11713
tri 4463 11633 4543 11713 sw
tri 4561 11633 4641 11713 ne
rect 4641 11633 5013 11713
tri 5013 11633 5093 11713 sw
tri 5111 11633 5191 11713 ne
rect 5191 11633 5563 11713
tri 5563 11633 5643 11713 sw
tri 5661 11633 5741 11713 ne
rect 5741 11633 6113 11713
tri 6113 11633 6193 11713 sw
tri 6211 11633 6291 11713 ne
rect 6291 11633 6663 11713
tri 6663 11633 6743 11713 sw
tri 6761 11633 6841 11713 ne
rect 6841 11633 7213 11713
tri 7213 11633 7293 11713 sw
tri 7311 11633 7391 11713 ne
rect 7391 11633 7763 11713
tri 7763 11633 7843 11713 sw
tri 7861 11633 7941 11713 ne
rect 7941 11633 8313 11713
tri 8313 11633 8393 11713 sw
tri 8411 11633 8491 11713 ne
rect 8491 11633 8863 11713
tri 8863 11633 8943 11713 sw
tri 8961 11633 9041 11713 ne
rect 9041 11633 9413 11713
tri 9413 11633 9493 11713 sw
tri 9511 11633 9591 11713 ne
rect 9591 11633 9963 11713
tri 9963 11633 10043 11713 sw
tri 10061 11633 10141 11713 ne
rect 10141 11633 10513 11713
tri 10513 11633 10593 11713 sw
tri 10611 11633 10691 11713 ne
rect 10691 11633 11063 11713
tri 11063 11633 11143 11713 sw
tri 11161 11633 11241 11713 ne
rect 11241 11633 11613 11713
tri 11613 11633 11693 11713 sw
tri 11711 11633 11791 11713 ne
rect 11791 11633 12163 11713
tri 12163 11633 12243 11713 sw
tri 12261 11633 12341 11713 ne
rect 12341 11633 12713 11713
tri 12713 11633 12793 11713 sw
tri 12811 11633 12891 11713 ne
rect 12891 11633 13263 11713
tri 13263 11633 13343 11713 sw
tri 13361 11633 13441 11713 ne
rect 13441 11633 13813 11713
tri 13813 11633 13893 11713 sw
tri 13911 11633 13991 11713 ne
rect 13991 11633 14363 11713
tri 14363 11633 14443 11713 sw
tri 14461 11633 14541 11713 ne
rect 14541 11633 14913 11713
tri 14913 11633 14993 11713 sw
tri 15011 11633 15091 11713 ne
rect 15091 11633 15463 11713
tri 15463 11633 15543 11713 sw
tri 15561 11633 15641 11713 ne
rect 15641 11633 16013 11713
tri 16013 11633 16093 11713 sw
tri 16111 11633 16191 11713 ne
rect 16191 11633 16563 11713
tri 16563 11633 16643 11713 sw
tri 16661 11633 16741 11713 ne
rect 16741 11633 17113 11713
tri 17113 11633 17193 11713 sw
tri 17211 11633 17291 11713 ne
rect 17291 11633 17663 11713
tri 17663 11633 17743 11713 sw
tri 17761 11633 17841 11713 ne
rect 17841 11633 18213 11713
tri 18213 11633 18293 11713 sw
tri 18311 11633 18391 11713 ne
rect 18391 11633 18763 11713
tri 18763 11633 18843 11713 sw
tri 18861 11633 18941 11713 ne
rect 18941 11633 19313 11713
tri 19313 11633 19393 11713 sw
tri 19411 11633 19491 11713 ne
rect 19491 11633 20100 11713
rect 261 11613 693 11633
rect -500 11535 163 11613
tri 163 11535 241 11613 sw
tri 261 11535 339 11613 ne
rect 339 11535 693 11613
tri 693 11535 791 11633 sw
tri 791 11535 889 11633 ne
rect 889 11535 1243 11633
tri 1243 11535 1341 11633 sw
tri 1341 11535 1439 11633 ne
rect 1439 11535 1793 11633
tri 1793 11535 1891 11633 sw
tri 1891 11535 1989 11633 ne
rect 1989 11535 2343 11633
tri 2343 11535 2441 11633 sw
tri 2441 11535 2539 11633 ne
rect 2539 11535 2893 11633
tri 2893 11535 2991 11633 sw
tri 2991 11535 3089 11633 ne
rect 3089 11535 3443 11633
tri 3443 11535 3541 11633 sw
tri 3541 11535 3639 11633 ne
rect 3639 11535 3993 11633
tri 3993 11535 4091 11633 sw
tri 4091 11535 4189 11633 ne
rect 4189 11535 4543 11633
tri 4543 11535 4641 11633 sw
tri 4641 11535 4739 11633 ne
rect 4739 11535 5093 11633
tri 5093 11535 5191 11633 sw
tri 5191 11535 5289 11633 ne
rect 5289 11535 5643 11633
tri 5643 11535 5741 11633 sw
tri 5741 11535 5839 11633 ne
rect 5839 11535 6193 11633
tri 6193 11535 6291 11633 sw
tri 6291 11535 6389 11633 ne
rect 6389 11535 6743 11633
tri 6743 11535 6841 11633 sw
tri 6841 11535 6939 11633 ne
rect 6939 11535 7293 11633
tri 7293 11535 7391 11633 sw
tri 7391 11535 7489 11633 ne
rect 7489 11535 7843 11633
tri 7843 11535 7941 11633 sw
tri 7941 11535 8039 11633 ne
rect 8039 11535 8393 11633
tri 8393 11535 8491 11633 sw
tri 8491 11535 8589 11633 ne
rect 8589 11535 8943 11633
tri 8943 11535 9041 11633 sw
tri 9041 11535 9139 11633 ne
rect 9139 11535 9493 11633
tri 9493 11535 9591 11633 sw
tri 9591 11535 9689 11633 ne
rect 9689 11535 10043 11633
tri 10043 11535 10141 11633 sw
tri 10141 11535 10239 11633 ne
rect 10239 11535 10593 11633
tri 10593 11535 10691 11633 sw
tri 10691 11535 10789 11633 ne
rect 10789 11535 11143 11633
tri 11143 11535 11241 11633 sw
tri 11241 11535 11339 11633 ne
rect 11339 11535 11693 11633
tri 11693 11535 11791 11633 sw
tri 11791 11535 11889 11633 ne
rect 11889 11535 12243 11633
tri 12243 11535 12341 11633 sw
tri 12341 11535 12439 11633 ne
rect 12439 11535 12793 11633
tri 12793 11535 12891 11633 sw
tri 12891 11535 12989 11633 ne
rect 12989 11535 13343 11633
tri 13343 11535 13441 11633 sw
tri 13441 11535 13539 11633 ne
rect 13539 11535 13893 11633
tri 13893 11535 13991 11633 sw
tri 13991 11535 14089 11633 ne
rect 14089 11535 14443 11633
tri 14443 11535 14541 11633 sw
tri 14541 11535 14639 11633 ne
rect 14639 11535 14993 11633
tri 14993 11535 15091 11633 sw
tri 15091 11535 15189 11633 ne
rect 15189 11535 15543 11633
tri 15543 11535 15641 11633 sw
tri 15641 11535 15739 11633 ne
rect 15739 11535 16093 11633
tri 16093 11535 16191 11633 sw
tri 16191 11535 16289 11633 ne
rect 16289 11535 16643 11633
tri 16643 11535 16741 11633 sw
tri 16741 11535 16839 11633 ne
rect 16839 11535 17193 11633
tri 17193 11535 17291 11633 sw
tri 17291 11535 17389 11633 ne
rect 17389 11535 17743 11633
tri 17743 11535 17841 11633 sw
tri 17841 11535 17939 11633 ne
rect 17939 11535 18293 11633
tri 18293 11535 18391 11633 sw
tri 18391 11535 18489 11633 ne
rect 18489 11535 18843 11633
tri 18843 11535 18941 11633 sw
tri 18941 11535 19039 11633 ne
rect 19039 11535 19393 11633
tri 19393 11535 19491 11633 sw
tri 19491 11535 19589 11633 ne
rect 19589 11613 20100 11633
rect 20200 11613 21800 11713
rect 19589 11535 21800 11613
rect -500 11487 241 11535
rect -500 11387 -400 11487
rect -300 11437 241 11487
tri 241 11437 339 11535 sw
tri 339 11437 437 11535 ne
rect 437 11437 791 11535
tri 791 11437 889 11535 sw
tri 889 11437 987 11535 ne
rect 987 11437 1341 11535
tri 1341 11437 1439 11535 sw
tri 1439 11437 1537 11535 ne
rect 1537 11437 1891 11535
tri 1891 11437 1989 11535 sw
tri 1989 11437 2087 11535 ne
rect 2087 11437 2441 11535
tri 2441 11437 2539 11535 sw
tri 2539 11437 2637 11535 ne
rect 2637 11437 2991 11535
tri 2991 11437 3089 11535 sw
tri 3089 11437 3187 11535 ne
rect 3187 11437 3541 11535
tri 3541 11437 3639 11535 sw
tri 3639 11437 3737 11535 ne
rect 3737 11437 4091 11535
tri 4091 11437 4189 11535 sw
tri 4189 11437 4287 11535 ne
rect 4287 11437 4641 11535
tri 4641 11437 4739 11535 sw
tri 4739 11437 4837 11535 ne
rect 4837 11437 5191 11535
tri 5191 11437 5289 11535 sw
tri 5289 11437 5387 11535 ne
rect 5387 11437 5741 11535
tri 5741 11437 5839 11535 sw
tri 5839 11437 5937 11535 ne
rect 5937 11437 6291 11535
tri 6291 11437 6389 11535 sw
tri 6389 11437 6487 11535 ne
rect 6487 11437 6841 11535
tri 6841 11437 6939 11535 sw
tri 6939 11437 7037 11535 ne
rect 7037 11437 7391 11535
tri 7391 11437 7489 11535 sw
tri 7489 11437 7587 11535 ne
rect 7587 11437 7941 11535
tri 7941 11437 8039 11535 sw
tri 8039 11437 8137 11535 ne
rect 8137 11437 8491 11535
tri 8491 11437 8589 11535 sw
tri 8589 11437 8687 11535 ne
rect 8687 11437 9041 11535
tri 9041 11437 9139 11535 sw
tri 9139 11437 9237 11535 ne
rect 9237 11437 9591 11535
tri 9591 11437 9689 11535 sw
tri 9689 11437 9787 11535 ne
rect 9787 11437 10141 11535
tri 10141 11437 10239 11535 sw
tri 10239 11437 10337 11535 ne
rect 10337 11437 10691 11535
tri 10691 11437 10789 11535 sw
tri 10789 11437 10887 11535 ne
rect 10887 11437 11241 11535
tri 11241 11437 11339 11535 sw
tri 11339 11437 11437 11535 ne
rect 11437 11437 11791 11535
tri 11791 11437 11889 11535 sw
tri 11889 11437 11987 11535 ne
rect 11987 11437 12341 11535
tri 12341 11437 12439 11535 sw
tri 12439 11437 12537 11535 ne
rect 12537 11437 12891 11535
tri 12891 11437 12989 11535 sw
tri 12989 11437 13087 11535 ne
rect 13087 11437 13441 11535
tri 13441 11437 13539 11535 sw
tri 13539 11437 13637 11535 ne
rect 13637 11437 13991 11535
tri 13991 11437 14089 11535 sw
tri 14089 11437 14187 11535 ne
rect 14187 11437 14541 11535
tri 14541 11437 14639 11535 sw
tri 14639 11437 14737 11535 ne
rect 14737 11437 15091 11535
tri 15091 11437 15189 11535 sw
tri 15189 11437 15287 11535 ne
rect 15287 11437 15641 11535
tri 15641 11437 15739 11535 sw
tri 15739 11437 15837 11535 ne
rect 15837 11437 16191 11535
tri 16191 11437 16289 11535 sw
tri 16289 11437 16387 11535 ne
rect 16387 11437 16741 11535
tri 16741 11437 16839 11535 sw
tri 16839 11437 16937 11535 ne
rect 16937 11437 17291 11535
tri 17291 11437 17389 11535 sw
tri 17389 11437 17487 11535 ne
rect 17487 11437 17841 11535
tri 17841 11437 17939 11535 sw
tri 17939 11437 18037 11535 ne
rect 18037 11437 18391 11535
tri 18391 11437 18489 11535 sw
tri 18489 11437 18587 11535 ne
rect 18587 11437 18941 11535
tri 18941 11437 19039 11535 sw
tri 19039 11437 19137 11535 ne
rect 19137 11437 19491 11535
tri 19491 11437 19589 11535 sw
tri 19589 11437 19687 11535 ne
rect 19687 11437 21800 11535
rect -300 11387 339 11437
rect -500 11339 339 11387
tri 339 11339 437 11437 sw
tri 437 11339 535 11437 ne
rect 535 11339 889 11437
tri 889 11339 987 11437 sw
tri 987 11339 1085 11437 ne
rect 1085 11339 1439 11437
tri 1439 11339 1537 11437 sw
tri 1537 11339 1635 11437 ne
rect 1635 11339 1989 11437
tri 1989 11339 2087 11437 sw
tri 2087 11339 2185 11437 ne
rect 2185 11339 2539 11437
tri 2539 11339 2637 11437 sw
tri 2637 11339 2735 11437 ne
rect 2735 11339 3089 11437
tri 3089 11339 3187 11437 sw
tri 3187 11339 3285 11437 ne
rect 3285 11339 3639 11437
tri 3639 11339 3737 11437 sw
tri 3737 11339 3835 11437 ne
rect 3835 11339 4189 11437
tri 4189 11339 4287 11437 sw
tri 4287 11339 4385 11437 ne
rect 4385 11339 4739 11437
tri 4739 11339 4837 11437 sw
tri 4837 11339 4935 11437 ne
rect 4935 11339 5289 11437
tri 5289 11339 5387 11437 sw
tri 5387 11339 5485 11437 ne
rect 5485 11339 5839 11437
tri 5839 11339 5937 11437 sw
tri 5937 11339 6035 11437 ne
rect 6035 11339 6389 11437
tri 6389 11339 6487 11437 sw
tri 6487 11339 6585 11437 ne
rect 6585 11339 6939 11437
tri 6939 11339 7037 11437 sw
tri 7037 11339 7135 11437 ne
rect 7135 11339 7489 11437
tri 7489 11339 7587 11437 sw
tri 7587 11339 7685 11437 ne
rect 7685 11339 8039 11437
tri 8039 11339 8137 11437 sw
tri 8137 11339 8235 11437 ne
rect 8235 11339 8589 11437
tri 8589 11339 8687 11437 sw
tri 8687 11339 8785 11437 ne
rect 8785 11339 9139 11437
tri 9139 11339 9237 11437 sw
tri 9237 11339 9335 11437 ne
rect 9335 11339 9689 11437
tri 9689 11339 9787 11437 sw
tri 9787 11339 9885 11437 ne
rect 9885 11339 10239 11437
tri 10239 11339 10337 11437 sw
tri 10337 11339 10435 11437 ne
rect 10435 11339 10789 11437
tri 10789 11339 10887 11437 sw
tri 10887 11339 10985 11437 ne
rect 10985 11339 11339 11437
tri 11339 11339 11437 11437 sw
tri 11437 11339 11535 11437 ne
rect 11535 11339 11889 11437
tri 11889 11339 11987 11437 sw
tri 11987 11339 12085 11437 ne
rect 12085 11339 12439 11437
tri 12439 11339 12537 11437 sw
tri 12537 11339 12635 11437 ne
rect 12635 11339 12989 11437
tri 12989 11339 13087 11437 sw
tri 13087 11339 13185 11437 ne
rect 13185 11339 13539 11437
tri 13539 11339 13637 11437 sw
tri 13637 11339 13735 11437 ne
rect 13735 11339 14089 11437
tri 14089 11339 14187 11437 sw
tri 14187 11339 14285 11437 ne
rect 14285 11339 14639 11437
tri 14639 11339 14737 11437 sw
tri 14737 11339 14835 11437 ne
rect 14835 11339 15189 11437
tri 15189 11339 15287 11437 sw
tri 15287 11339 15385 11437 ne
rect 15385 11339 15739 11437
tri 15739 11339 15837 11437 sw
tri 15837 11339 15935 11437 ne
rect 15935 11339 16289 11437
tri 16289 11339 16387 11437 sw
tri 16387 11339 16485 11437 ne
rect 16485 11339 16839 11437
tri 16839 11339 16937 11437 sw
tri 16937 11339 17035 11437 ne
rect 17035 11339 17389 11437
tri 17389 11339 17487 11437 sw
tri 17487 11339 17585 11437 ne
rect 17585 11339 17939 11437
tri 17939 11339 18037 11437 sw
tri 18037 11339 18135 11437 ne
rect 18135 11339 18489 11437
tri 18489 11339 18587 11437 sw
tri 18587 11339 18685 11437 ne
rect 18685 11339 19039 11437
tri 19039 11339 19137 11437 sw
tri 19137 11339 19235 11437 ne
rect 19235 11339 19589 11437
tri 19589 11339 19687 11437 sw
rect -500 11335 437 11339
rect -500 11215 215 11335
rect 335 11241 437 11335
tri 437 11241 535 11339 sw
tri 535 11241 633 11339 ne
rect 633 11335 987 11339
rect 633 11241 765 11335
rect 335 11215 535 11241
rect -500 11211 535 11215
tri 535 11211 565 11241 sw
tri 633 11211 663 11241 ne
rect 663 11215 765 11241
rect 885 11241 987 11335
tri 987 11241 1085 11339 sw
tri 1085 11241 1183 11339 ne
rect 1183 11335 1537 11339
rect 1183 11241 1315 11335
rect 885 11215 1085 11241
rect 663 11211 1085 11215
tri 1085 11211 1115 11241 sw
tri 1183 11211 1213 11241 ne
rect 1213 11215 1315 11241
rect 1435 11241 1537 11335
tri 1537 11241 1635 11339 sw
tri 1635 11241 1733 11339 ne
rect 1733 11335 2087 11339
rect 1733 11241 1865 11335
rect 1435 11215 1635 11241
rect 1213 11211 1635 11215
tri 1635 11211 1665 11241 sw
tri 1733 11211 1763 11241 ne
rect 1763 11215 1865 11241
rect 1985 11241 2087 11335
tri 2087 11241 2185 11339 sw
tri 2185 11241 2283 11339 ne
rect 2283 11335 2637 11339
rect 2283 11241 2415 11335
rect 1985 11215 2185 11241
rect 1763 11211 2185 11215
tri 2185 11211 2215 11241 sw
tri 2283 11211 2313 11241 ne
rect 2313 11215 2415 11241
rect 2535 11241 2637 11335
tri 2637 11241 2735 11339 sw
tri 2735 11241 2833 11339 ne
rect 2833 11335 3187 11339
rect 2833 11241 2965 11335
rect 2535 11215 2735 11241
rect 2313 11211 2735 11215
tri 2735 11211 2765 11241 sw
tri 2833 11211 2863 11241 ne
rect 2863 11215 2965 11241
rect 3085 11241 3187 11335
tri 3187 11241 3285 11339 sw
tri 3285 11241 3383 11339 ne
rect 3383 11335 3737 11339
rect 3383 11241 3515 11335
rect 3085 11215 3285 11241
rect 2863 11211 3285 11215
tri 3285 11211 3315 11241 sw
tri 3383 11211 3413 11241 ne
rect 3413 11215 3515 11241
rect 3635 11241 3737 11335
tri 3737 11241 3835 11339 sw
tri 3835 11241 3933 11339 ne
rect 3933 11335 4287 11339
rect 3933 11241 4065 11335
rect 3635 11215 3835 11241
rect 3413 11211 3835 11215
tri 3835 11211 3865 11241 sw
tri 3933 11211 3963 11241 ne
rect 3963 11215 4065 11241
rect 4185 11241 4287 11335
tri 4287 11241 4385 11339 sw
tri 4385 11241 4483 11339 ne
rect 4483 11335 4837 11339
rect 4483 11241 4615 11335
rect 4185 11215 4385 11241
rect 3963 11211 4385 11215
tri 4385 11211 4415 11241 sw
tri 4483 11211 4513 11241 ne
rect 4513 11215 4615 11241
rect 4735 11241 4837 11335
tri 4837 11241 4935 11339 sw
tri 4935 11241 5033 11339 ne
rect 5033 11335 5387 11339
rect 5033 11241 5165 11335
rect 4735 11215 4935 11241
rect 4513 11211 4935 11215
tri 4935 11211 4965 11241 sw
tri 5033 11211 5063 11241 ne
rect 5063 11215 5165 11241
rect 5285 11241 5387 11335
tri 5387 11241 5485 11339 sw
tri 5485 11241 5583 11339 ne
rect 5583 11335 5937 11339
rect 5583 11241 5715 11335
rect 5285 11215 5485 11241
rect 5063 11211 5485 11215
tri 5485 11211 5515 11241 sw
tri 5583 11211 5613 11241 ne
rect 5613 11215 5715 11241
rect 5835 11241 5937 11335
tri 5937 11241 6035 11339 sw
tri 6035 11241 6133 11339 ne
rect 6133 11335 6487 11339
rect 6133 11241 6265 11335
rect 5835 11215 6035 11241
rect 5613 11211 6035 11215
tri 6035 11211 6065 11241 sw
tri 6133 11211 6163 11241 ne
rect 6163 11215 6265 11241
rect 6385 11241 6487 11335
tri 6487 11241 6585 11339 sw
tri 6585 11241 6683 11339 ne
rect 6683 11335 7037 11339
rect 6683 11241 6815 11335
rect 6385 11215 6585 11241
rect 6163 11211 6585 11215
tri 6585 11211 6615 11241 sw
tri 6683 11211 6713 11241 ne
rect 6713 11215 6815 11241
rect 6935 11241 7037 11335
tri 7037 11241 7135 11339 sw
tri 7135 11241 7233 11339 ne
rect 7233 11335 7587 11339
rect 7233 11241 7365 11335
rect 6935 11215 7135 11241
rect 6713 11211 7135 11215
tri 7135 11211 7165 11241 sw
tri 7233 11211 7263 11241 ne
rect 7263 11215 7365 11241
rect 7485 11241 7587 11335
tri 7587 11241 7685 11339 sw
tri 7685 11241 7783 11339 ne
rect 7783 11335 8137 11339
rect 7783 11241 7915 11335
rect 7485 11215 7685 11241
rect 7263 11211 7685 11215
tri 7685 11211 7715 11241 sw
tri 7783 11211 7813 11241 ne
rect 7813 11215 7915 11241
rect 8035 11241 8137 11335
tri 8137 11241 8235 11339 sw
tri 8235 11241 8333 11339 ne
rect 8333 11335 8687 11339
rect 8333 11241 8465 11335
rect 8035 11215 8235 11241
rect 7813 11211 8235 11215
tri 8235 11211 8265 11241 sw
tri 8333 11211 8363 11241 ne
rect 8363 11215 8465 11241
rect 8585 11241 8687 11335
tri 8687 11241 8785 11339 sw
tri 8785 11241 8883 11339 ne
rect 8883 11335 9237 11339
rect 8883 11241 9015 11335
rect 8585 11215 8785 11241
rect 8363 11211 8785 11215
tri 8785 11211 8815 11241 sw
tri 8883 11211 8913 11241 ne
rect 8913 11215 9015 11241
rect 9135 11241 9237 11335
tri 9237 11241 9335 11339 sw
tri 9335 11241 9433 11339 ne
rect 9433 11335 9787 11339
rect 9433 11241 9565 11335
rect 9135 11215 9335 11241
rect 8913 11211 9335 11215
tri 9335 11211 9365 11241 sw
tri 9433 11211 9463 11241 ne
rect 9463 11215 9565 11241
rect 9685 11241 9787 11335
tri 9787 11241 9885 11339 sw
tri 9885 11241 9983 11339 ne
rect 9983 11335 10337 11339
rect 9983 11241 10115 11335
rect 9685 11215 9885 11241
rect 9463 11211 9885 11215
tri 9885 11211 9915 11241 sw
tri 9983 11211 10013 11241 ne
rect 10013 11215 10115 11241
rect 10235 11241 10337 11335
tri 10337 11241 10435 11339 sw
tri 10435 11241 10533 11339 ne
rect 10533 11335 10887 11339
rect 10533 11241 10665 11335
rect 10235 11215 10435 11241
rect 10013 11211 10435 11215
tri 10435 11211 10465 11241 sw
tri 10533 11211 10563 11241 ne
rect 10563 11215 10665 11241
rect 10785 11241 10887 11335
tri 10887 11241 10985 11339 sw
tri 10985 11241 11083 11339 ne
rect 11083 11335 11437 11339
rect 11083 11241 11215 11335
rect 10785 11215 10985 11241
rect 10563 11211 10985 11215
tri 10985 11211 11015 11241 sw
tri 11083 11211 11113 11241 ne
rect 11113 11215 11215 11241
rect 11335 11241 11437 11335
tri 11437 11241 11535 11339 sw
tri 11535 11241 11633 11339 ne
rect 11633 11335 11987 11339
rect 11633 11241 11765 11335
rect 11335 11215 11535 11241
rect 11113 11211 11535 11215
tri 11535 11211 11565 11241 sw
tri 11633 11211 11663 11241 ne
rect 11663 11215 11765 11241
rect 11885 11241 11987 11335
tri 11987 11241 12085 11339 sw
tri 12085 11241 12183 11339 ne
rect 12183 11335 12537 11339
rect 12183 11241 12315 11335
rect 11885 11215 12085 11241
rect 11663 11211 12085 11215
tri 12085 11211 12115 11241 sw
tri 12183 11211 12213 11241 ne
rect 12213 11215 12315 11241
rect 12435 11241 12537 11335
tri 12537 11241 12635 11339 sw
tri 12635 11241 12733 11339 ne
rect 12733 11335 13087 11339
rect 12733 11241 12865 11335
rect 12435 11215 12635 11241
rect 12213 11211 12635 11215
tri 12635 11211 12665 11241 sw
tri 12733 11211 12763 11241 ne
rect 12763 11215 12865 11241
rect 12985 11241 13087 11335
tri 13087 11241 13185 11339 sw
tri 13185 11241 13283 11339 ne
rect 13283 11335 13637 11339
rect 13283 11241 13415 11335
rect 12985 11215 13185 11241
rect 12763 11211 13185 11215
tri 13185 11211 13215 11241 sw
tri 13283 11211 13313 11241 ne
rect 13313 11215 13415 11241
rect 13535 11241 13637 11335
tri 13637 11241 13735 11339 sw
tri 13735 11241 13833 11339 ne
rect 13833 11335 14187 11339
rect 13833 11241 13965 11335
rect 13535 11215 13735 11241
rect 13313 11211 13735 11215
tri 13735 11211 13765 11241 sw
tri 13833 11211 13863 11241 ne
rect 13863 11215 13965 11241
rect 14085 11241 14187 11335
tri 14187 11241 14285 11339 sw
tri 14285 11241 14383 11339 ne
rect 14383 11335 14737 11339
rect 14383 11241 14515 11335
rect 14085 11215 14285 11241
rect 13863 11211 14285 11215
tri 14285 11211 14315 11241 sw
tri 14383 11211 14413 11241 ne
rect 14413 11215 14515 11241
rect 14635 11241 14737 11335
tri 14737 11241 14835 11339 sw
tri 14835 11241 14933 11339 ne
rect 14933 11335 15287 11339
rect 14933 11241 15065 11335
rect 14635 11215 14835 11241
rect 14413 11211 14835 11215
tri 14835 11211 14865 11241 sw
tri 14933 11211 14963 11241 ne
rect 14963 11215 15065 11241
rect 15185 11241 15287 11335
tri 15287 11241 15385 11339 sw
tri 15385 11241 15483 11339 ne
rect 15483 11335 15837 11339
rect 15483 11241 15615 11335
rect 15185 11215 15385 11241
rect 14963 11211 15385 11215
tri 15385 11211 15415 11241 sw
tri 15483 11211 15513 11241 ne
rect 15513 11215 15615 11241
rect 15735 11241 15837 11335
tri 15837 11241 15935 11339 sw
tri 15935 11241 16033 11339 ne
rect 16033 11335 16387 11339
rect 16033 11241 16165 11335
rect 15735 11215 15935 11241
rect 15513 11211 15935 11215
tri 15935 11211 15965 11241 sw
tri 16033 11211 16063 11241 ne
rect 16063 11215 16165 11241
rect 16285 11241 16387 11335
tri 16387 11241 16485 11339 sw
tri 16485 11241 16583 11339 ne
rect 16583 11335 16937 11339
rect 16583 11241 16715 11335
rect 16285 11215 16485 11241
rect 16063 11211 16485 11215
tri 16485 11211 16515 11241 sw
tri 16583 11211 16613 11241 ne
rect 16613 11215 16715 11241
rect 16835 11241 16937 11335
tri 16937 11241 17035 11339 sw
tri 17035 11241 17133 11339 ne
rect 17133 11335 17487 11339
rect 17133 11241 17265 11335
rect 16835 11215 17035 11241
rect 16613 11211 17035 11215
tri 17035 11211 17065 11241 sw
tri 17133 11211 17163 11241 ne
rect 17163 11215 17265 11241
rect 17385 11241 17487 11335
tri 17487 11241 17585 11339 sw
tri 17585 11241 17683 11339 ne
rect 17683 11335 18037 11339
rect 17683 11241 17815 11335
rect 17385 11215 17585 11241
rect 17163 11211 17585 11215
tri 17585 11211 17615 11241 sw
tri 17683 11211 17713 11241 ne
rect 17713 11215 17815 11241
rect 17935 11241 18037 11335
tri 18037 11241 18135 11339 sw
tri 18135 11241 18233 11339 ne
rect 18233 11335 18587 11339
rect 18233 11241 18365 11335
rect 17935 11215 18135 11241
rect 17713 11211 18135 11215
tri 18135 11211 18165 11241 sw
tri 18233 11211 18263 11241 ne
rect 18263 11215 18365 11241
rect 18485 11241 18587 11335
tri 18587 11241 18685 11339 sw
tri 18685 11241 18783 11339 ne
rect 18783 11335 19137 11339
rect 18783 11241 18915 11335
rect 18485 11215 18685 11241
rect 18263 11211 18685 11215
tri 18685 11211 18715 11241 sw
tri 18783 11211 18813 11241 ne
rect 18813 11215 18915 11241
rect 19035 11241 19137 11335
tri 19137 11241 19235 11339 sw
tri 19235 11241 19333 11339 ne
rect 19333 11335 20300 11339
rect 19333 11241 19465 11335
rect 19035 11215 19235 11241
rect 18813 11211 19235 11215
tri 19235 11211 19265 11241 sw
tri 19333 11211 19363 11241 ne
rect 19363 11215 19465 11241
rect 19585 11215 20300 11335
rect 19363 11211 20300 11215
tri 113 11113 211 11211 ne
rect 211 11113 565 11211
tri 565 11113 663 11211 sw
tri 663 11113 761 11211 ne
rect 761 11113 1115 11211
tri 1115 11113 1213 11211 sw
tri 1213 11113 1311 11211 ne
rect 1311 11113 1665 11211
tri 1665 11113 1763 11211 sw
tri 1763 11113 1861 11211 ne
rect 1861 11113 2215 11211
tri 2215 11113 2313 11211 sw
tri 2313 11113 2411 11211 ne
rect 2411 11113 2765 11211
tri 2765 11113 2863 11211 sw
tri 2863 11113 2961 11211 ne
rect 2961 11113 3315 11211
tri 3315 11113 3413 11211 sw
tri 3413 11113 3511 11211 ne
rect 3511 11113 3865 11211
tri 3865 11113 3963 11211 sw
tri 3963 11113 4061 11211 ne
rect 4061 11113 4415 11211
tri 4415 11113 4513 11211 sw
tri 4513 11113 4611 11211 ne
rect 4611 11113 4965 11211
tri 4965 11113 5063 11211 sw
tri 5063 11113 5161 11211 ne
rect 5161 11113 5515 11211
tri 5515 11113 5613 11211 sw
tri 5613 11113 5711 11211 ne
rect 5711 11113 6065 11211
tri 6065 11113 6163 11211 sw
tri 6163 11113 6261 11211 ne
rect 6261 11113 6615 11211
tri 6615 11113 6713 11211 sw
tri 6713 11113 6811 11211 ne
rect 6811 11113 7165 11211
tri 7165 11113 7263 11211 sw
tri 7263 11113 7361 11211 ne
rect 7361 11113 7715 11211
tri 7715 11113 7813 11211 sw
tri 7813 11113 7911 11211 ne
rect 7911 11113 8265 11211
tri 8265 11113 8363 11211 sw
tri 8363 11113 8461 11211 ne
rect 8461 11113 8815 11211
tri 8815 11113 8913 11211 sw
tri 8913 11113 9011 11211 ne
rect 9011 11113 9365 11211
tri 9365 11113 9463 11211 sw
tri 9463 11113 9561 11211 ne
rect 9561 11113 9915 11211
tri 9915 11113 10013 11211 sw
tri 10013 11113 10111 11211 ne
rect 10111 11113 10465 11211
tri 10465 11113 10563 11211 sw
tri 10563 11113 10661 11211 ne
rect 10661 11113 11015 11211
tri 11015 11113 11113 11211 sw
tri 11113 11113 11211 11211 ne
rect 11211 11113 11565 11211
tri 11565 11113 11663 11211 sw
tri 11663 11113 11761 11211 ne
rect 11761 11113 12115 11211
tri 12115 11113 12213 11211 sw
tri 12213 11113 12311 11211 ne
rect 12311 11113 12665 11211
tri 12665 11113 12763 11211 sw
tri 12763 11113 12861 11211 ne
rect 12861 11113 13215 11211
tri 13215 11113 13313 11211 sw
tri 13313 11113 13411 11211 ne
rect 13411 11113 13765 11211
tri 13765 11113 13863 11211 sw
tri 13863 11113 13961 11211 ne
rect 13961 11113 14315 11211
tri 14315 11113 14413 11211 sw
tri 14413 11113 14511 11211 ne
rect 14511 11113 14865 11211
tri 14865 11113 14963 11211 sw
tri 14963 11113 15061 11211 ne
rect 15061 11113 15415 11211
tri 15415 11113 15513 11211 sw
tri 15513 11113 15611 11211 ne
rect 15611 11113 15965 11211
tri 15965 11113 16063 11211 sw
tri 16063 11113 16161 11211 ne
rect 16161 11113 16515 11211
tri 16515 11113 16613 11211 sw
tri 16613 11113 16711 11211 ne
rect 16711 11113 17065 11211
tri 17065 11113 17163 11211 sw
tri 17163 11113 17261 11211 ne
rect 17261 11113 17615 11211
tri 17615 11113 17713 11211 sw
tri 17713 11113 17811 11211 ne
rect 17811 11113 18165 11211
tri 18165 11113 18263 11211 sw
tri 18263 11113 18361 11211 ne
rect 18361 11113 18715 11211
tri 18715 11113 18813 11211 sw
tri 18813 11113 18911 11211 ne
rect 18911 11113 19265 11211
tri 19265 11113 19363 11211 sw
tri 19363 11113 19461 11211 ne
rect 19461 11113 20300 11211
rect -2000 11083 113 11113
tri 113 11083 143 11113 sw
tri 211 11083 241 11113 ne
rect 241 11083 663 11113
tri 663 11083 693 11113 sw
tri 761 11083 791 11113 ne
rect 791 11083 1213 11113
tri 1213 11083 1243 11113 sw
tri 1311 11083 1341 11113 ne
rect 1341 11083 1763 11113
tri 1763 11083 1793 11113 sw
tri 1861 11083 1891 11113 ne
rect 1891 11083 2313 11113
tri 2313 11083 2343 11113 sw
tri 2411 11083 2441 11113 ne
rect 2441 11083 2863 11113
tri 2863 11083 2893 11113 sw
tri 2961 11083 2991 11113 ne
rect 2991 11083 3413 11113
tri 3413 11083 3443 11113 sw
tri 3511 11083 3541 11113 ne
rect 3541 11083 3963 11113
tri 3963 11083 3993 11113 sw
tri 4061 11083 4091 11113 ne
rect 4091 11083 4513 11113
tri 4513 11083 4543 11113 sw
tri 4611 11083 4641 11113 ne
rect 4641 11083 5063 11113
tri 5063 11083 5093 11113 sw
tri 5161 11083 5191 11113 ne
rect 5191 11083 5613 11113
tri 5613 11083 5643 11113 sw
tri 5711 11083 5741 11113 ne
rect 5741 11083 6163 11113
tri 6163 11083 6193 11113 sw
tri 6261 11083 6291 11113 ne
rect 6291 11083 6713 11113
tri 6713 11083 6743 11113 sw
tri 6811 11083 6841 11113 ne
rect 6841 11083 7263 11113
tri 7263 11083 7293 11113 sw
tri 7361 11083 7391 11113 ne
rect 7391 11083 7813 11113
tri 7813 11083 7843 11113 sw
tri 7911 11083 7941 11113 ne
rect 7941 11083 8363 11113
tri 8363 11083 8393 11113 sw
tri 8461 11083 8491 11113 ne
rect 8491 11083 8913 11113
tri 8913 11083 8943 11113 sw
tri 9011 11083 9041 11113 ne
rect 9041 11083 9463 11113
tri 9463 11083 9493 11113 sw
tri 9561 11083 9591 11113 ne
rect 9591 11083 10013 11113
tri 10013 11083 10043 11113 sw
tri 10111 11083 10141 11113 ne
rect 10141 11083 10563 11113
tri 10563 11083 10593 11113 sw
tri 10661 11083 10691 11113 ne
rect 10691 11083 11113 11113
tri 11113 11083 11143 11113 sw
tri 11211 11083 11241 11113 ne
rect 11241 11083 11663 11113
tri 11663 11083 11693 11113 sw
tri 11761 11083 11791 11113 ne
rect 11791 11083 12213 11113
tri 12213 11083 12243 11113 sw
tri 12311 11083 12341 11113 ne
rect 12341 11083 12763 11113
tri 12763 11083 12793 11113 sw
tri 12861 11083 12891 11113 ne
rect 12891 11083 13313 11113
tri 13313 11083 13343 11113 sw
tri 13411 11083 13441 11113 ne
rect 13441 11083 13863 11113
tri 13863 11083 13893 11113 sw
tri 13961 11083 13991 11113 ne
rect 13991 11083 14413 11113
tri 14413 11083 14443 11113 sw
tri 14511 11083 14541 11113 ne
rect 14541 11083 14963 11113
tri 14963 11083 14993 11113 sw
tri 15061 11083 15091 11113 ne
rect 15091 11083 15513 11113
tri 15513 11083 15543 11113 sw
tri 15611 11083 15641 11113 ne
rect 15641 11083 16063 11113
tri 16063 11083 16093 11113 sw
tri 16161 11083 16191 11113 ne
rect 16191 11083 16613 11113
tri 16613 11083 16643 11113 sw
tri 16711 11083 16741 11113 ne
rect 16741 11083 17163 11113
tri 17163 11083 17193 11113 sw
tri 17261 11083 17291 11113 ne
rect 17291 11083 17713 11113
tri 17713 11083 17743 11113 sw
tri 17811 11083 17841 11113 ne
rect 17841 11083 18263 11113
tri 18263 11083 18293 11113 sw
tri 18361 11083 18391 11113 ne
rect 18391 11083 18813 11113
tri 18813 11083 18843 11113 sw
tri 18911 11083 18941 11113 ne
rect 18941 11083 19363 11113
tri 19363 11083 19393 11113 sw
tri 19461 11083 19491 11113 ne
rect 19491 11083 20300 11113
rect -2000 10985 143 11083
tri 143 10985 241 11083 sw
tri 241 10985 339 11083 ne
rect 339 10985 693 11083
tri 693 10985 791 11083 sw
tri 791 10985 889 11083 ne
rect 889 10985 1243 11083
tri 1243 10985 1341 11083 sw
tri 1341 10985 1439 11083 ne
rect 1439 10985 1793 11083
tri 1793 10985 1891 11083 sw
tri 1891 10985 1989 11083 ne
rect 1989 10985 2343 11083
tri 2343 10985 2441 11083 sw
tri 2441 10985 2539 11083 ne
rect 2539 10985 2893 11083
tri 2893 10985 2991 11083 sw
tri 2991 10985 3089 11083 ne
rect 3089 10985 3443 11083
tri 3443 10985 3541 11083 sw
tri 3541 10985 3639 11083 ne
rect 3639 10985 3993 11083
tri 3993 10985 4091 11083 sw
tri 4091 10985 4189 11083 ne
rect 4189 10985 4543 11083
tri 4543 10985 4641 11083 sw
tri 4641 10985 4739 11083 ne
rect 4739 10985 5093 11083
tri 5093 10985 5191 11083 sw
tri 5191 10985 5289 11083 ne
rect 5289 10985 5643 11083
tri 5643 10985 5741 11083 sw
tri 5741 10985 5839 11083 ne
rect 5839 10985 6193 11083
tri 6193 10985 6291 11083 sw
tri 6291 10985 6389 11083 ne
rect 6389 10985 6743 11083
tri 6743 10985 6841 11083 sw
tri 6841 10985 6939 11083 ne
rect 6939 10985 7293 11083
tri 7293 10985 7391 11083 sw
tri 7391 10985 7489 11083 ne
rect 7489 10985 7843 11083
tri 7843 10985 7941 11083 sw
tri 7941 10985 8039 11083 ne
rect 8039 10985 8393 11083
tri 8393 10985 8491 11083 sw
tri 8491 10985 8589 11083 ne
rect 8589 10985 8943 11083
tri 8943 10985 9041 11083 sw
tri 9041 10985 9139 11083 ne
rect 9139 10985 9493 11083
tri 9493 10985 9591 11083 sw
tri 9591 10985 9689 11083 ne
rect 9689 10985 10043 11083
tri 10043 10985 10141 11083 sw
tri 10141 10985 10239 11083 ne
rect 10239 10985 10593 11083
tri 10593 10985 10691 11083 sw
tri 10691 10985 10789 11083 ne
rect 10789 10985 11143 11083
tri 11143 10985 11241 11083 sw
tri 11241 10985 11339 11083 ne
rect 11339 10985 11693 11083
tri 11693 10985 11791 11083 sw
tri 11791 10985 11889 11083 ne
rect 11889 10985 12243 11083
tri 12243 10985 12341 11083 sw
tri 12341 10985 12439 11083 ne
rect 12439 10985 12793 11083
tri 12793 10985 12891 11083 sw
tri 12891 10985 12989 11083 ne
rect 12989 10985 13343 11083
tri 13343 10985 13441 11083 sw
tri 13441 10985 13539 11083 ne
rect 13539 10985 13893 11083
tri 13893 10985 13991 11083 sw
tri 13991 10985 14089 11083 ne
rect 14089 10985 14443 11083
tri 14443 10985 14541 11083 sw
tri 14541 10985 14639 11083 ne
rect 14639 10985 14993 11083
tri 14993 10985 15091 11083 sw
tri 15091 10985 15189 11083 ne
rect 15189 10985 15543 11083
tri 15543 10985 15641 11083 sw
tri 15641 10985 15739 11083 ne
rect 15739 10985 16093 11083
tri 16093 10985 16191 11083 sw
tri 16191 10985 16289 11083 ne
rect 16289 10985 16643 11083
tri 16643 10985 16741 11083 sw
tri 16741 10985 16839 11083 ne
rect 16839 10985 17193 11083
tri 17193 10985 17291 11083 sw
tri 17291 10985 17389 11083 ne
rect 17389 10985 17743 11083
tri 17743 10985 17841 11083 sw
tri 17841 10985 17939 11083 ne
rect 17939 10985 18293 11083
tri 18293 10985 18391 11083 sw
tri 18391 10985 18489 11083 ne
rect 18489 10985 18843 11083
tri 18843 10985 18941 11083 sw
tri 18941 10985 19039 11083 ne
rect 19039 10985 19393 11083
tri 19393 10985 19491 11083 sw
tri 19491 10985 19589 11083 ne
rect 19589 10985 20300 11083
rect -2000 10887 241 10985
tri 241 10887 339 10985 sw
tri 339 10887 437 10985 ne
rect 437 10887 791 10985
tri 791 10887 889 10985 sw
tri 889 10887 987 10985 ne
rect 987 10887 1341 10985
tri 1341 10887 1439 10985 sw
tri 1439 10887 1537 10985 ne
rect 1537 10887 1891 10985
tri 1891 10887 1989 10985 sw
tri 1989 10887 2087 10985 ne
rect 2087 10887 2441 10985
tri 2441 10887 2539 10985 sw
tri 2539 10887 2637 10985 ne
rect 2637 10887 2991 10985
tri 2991 10887 3089 10985 sw
tri 3089 10887 3187 10985 ne
rect 3187 10887 3541 10985
tri 3541 10887 3639 10985 sw
tri 3639 10887 3737 10985 ne
rect 3737 10887 4091 10985
tri 4091 10887 4189 10985 sw
tri 4189 10887 4287 10985 ne
rect 4287 10887 4641 10985
tri 4641 10887 4739 10985 sw
tri 4739 10887 4837 10985 ne
rect 4837 10887 5191 10985
tri 5191 10887 5289 10985 sw
tri 5289 10887 5387 10985 ne
rect 5387 10887 5741 10985
tri 5741 10887 5839 10985 sw
tri 5839 10887 5937 10985 ne
rect 5937 10887 6291 10985
tri 6291 10887 6389 10985 sw
tri 6389 10887 6487 10985 ne
rect 6487 10887 6841 10985
tri 6841 10887 6939 10985 sw
tri 6939 10887 7037 10985 ne
rect 7037 10887 7391 10985
tri 7391 10887 7489 10985 sw
tri 7489 10887 7587 10985 ne
rect 7587 10887 7941 10985
tri 7941 10887 8039 10985 sw
tri 8039 10887 8137 10985 ne
rect 8137 10887 8491 10985
tri 8491 10887 8589 10985 sw
tri 8589 10887 8687 10985 ne
rect 8687 10887 9041 10985
tri 9041 10887 9139 10985 sw
tri 9139 10887 9237 10985 ne
rect 9237 10887 9591 10985
tri 9591 10887 9689 10985 sw
tri 9689 10887 9787 10985 ne
rect 9787 10887 10141 10985
tri 10141 10887 10239 10985 sw
tri 10239 10887 10337 10985 ne
rect 10337 10887 10691 10985
tri 10691 10887 10789 10985 sw
tri 10789 10887 10887 10985 ne
rect 10887 10887 11241 10985
tri 11241 10887 11339 10985 sw
tri 11339 10887 11437 10985 ne
rect 11437 10887 11791 10985
tri 11791 10887 11889 10985 sw
tri 11889 10887 11987 10985 ne
rect 11987 10887 12341 10985
tri 12341 10887 12439 10985 sw
tri 12439 10887 12537 10985 ne
rect 12537 10887 12891 10985
tri 12891 10887 12989 10985 sw
tri 12989 10887 13087 10985 ne
rect 13087 10887 13441 10985
tri 13441 10887 13539 10985 sw
tri 13539 10887 13637 10985 ne
rect 13637 10887 13991 10985
tri 13991 10887 14089 10985 sw
tri 14089 10887 14187 10985 ne
rect 14187 10887 14541 10985
tri 14541 10887 14639 10985 sw
tri 14639 10887 14737 10985 ne
rect 14737 10887 15091 10985
tri 15091 10887 15189 10985 sw
tri 15189 10887 15287 10985 ne
rect 15287 10887 15641 10985
tri 15641 10887 15739 10985 sw
tri 15739 10887 15837 10985 ne
rect 15837 10887 16191 10985
tri 16191 10887 16289 10985 sw
tri 16289 10887 16387 10985 ne
rect 16387 10887 16741 10985
tri 16741 10887 16839 10985 sw
tri 16839 10887 16937 10985 ne
rect 16937 10887 17291 10985
tri 17291 10887 17389 10985 sw
tri 17389 10887 17487 10985 ne
rect 17487 10887 17841 10985
tri 17841 10887 17939 10985 sw
tri 17939 10887 18037 10985 ne
rect 18037 10887 18391 10985
tri 18391 10887 18489 10985 sw
tri 18489 10887 18587 10985 ne
rect 18587 10887 18941 10985
tri 18941 10887 19039 10985 sw
tri 19039 10887 19137 10985 ne
rect 19137 10887 19491 10985
tri 19491 10887 19589 10985 sw
tri 19589 10887 19687 10985 ne
rect 19687 10887 20300 10985
rect -2000 10789 339 10887
tri 339 10789 437 10887 sw
tri 437 10789 535 10887 ne
rect 535 10789 889 10887
tri 889 10789 987 10887 sw
tri 987 10789 1085 10887 ne
rect 1085 10789 1439 10887
tri 1439 10789 1537 10887 sw
tri 1537 10789 1635 10887 ne
rect 1635 10789 1989 10887
tri 1989 10789 2087 10887 sw
tri 2087 10789 2185 10887 ne
rect 2185 10789 2539 10887
tri 2539 10789 2637 10887 sw
tri 2637 10789 2735 10887 ne
rect 2735 10789 3089 10887
tri 3089 10789 3187 10887 sw
tri 3187 10789 3285 10887 ne
rect 3285 10789 3639 10887
tri 3639 10789 3737 10887 sw
tri 3737 10789 3835 10887 ne
rect 3835 10789 4189 10887
tri 4189 10789 4287 10887 sw
tri 4287 10789 4385 10887 ne
rect 4385 10789 4739 10887
tri 4739 10789 4837 10887 sw
tri 4837 10789 4935 10887 ne
rect 4935 10789 5289 10887
tri 5289 10789 5387 10887 sw
tri 5387 10789 5485 10887 ne
rect 5485 10789 5839 10887
tri 5839 10789 5937 10887 sw
tri 5937 10789 6035 10887 ne
rect 6035 10789 6389 10887
tri 6389 10789 6487 10887 sw
tri 6487 10789 6585 10887 ne
rect 6585 10789 6939 10887
tri 6939 10789 7037 10887 sw
tri 7037 10789 7135 10887 ne
rect 7135 10789 7489 10887
tri 7489 10789 7587 10887 sw
tri 7587 10789 7685 10887 ne
rect 7685 10789 8039 10887
tri 8039 10789 8137 10887 sw
tri 8137 10789 8235 10887 ne
rect 8235 10789 8589 10887
tri 8589 10789 8687 10887 sw
tri 8687 10789 8785 10887 ne
rect 8785 10789 9139 10887
tri 9139 10789 9237 10887 sw
tri 9237 10789 9335 10887 ne
rect 9335 10789 9689 10887
tri 9689 10789 9787 10887 sw
tri 9787 10789 9885 10887 ne
rect 9885 10789 10239 10887
tri 10239 10789 10337 10887 sw
tri 10337 10789 10435 10887 ne
rect 10435 10789 10789 10887
tri 10789 10789 10887 10887 sw
tri 10887 10789 10985 10887 ne
rect 10985 10789 11339 10887
tri 11339 10789 11437 10887 sw
tri 11437 10789 11535 10887 ne
rect 11535 10789 11889 10887
tri 11889 10789 11987 10887 sw
tri 11987 10789 12085 10887 ne
rect 12085 10789 12439 10887
tri 12439 10789 12537 10887 sw
tri 12537 10789 12635 10887 ne
rect 12635 10789 12989 10887
tri 12989 10789 13087 10887 sw
tri 13087 10789 13185 10887 ne
rect 13185 10789 13539 10887
tri 13539 10789 13637 10887 sw
tri 13637 10789 13735 10887 ne
rect 13735 10789 14089 10887
tri 14089 10789 14187 10887 sw
tri 14187 10789 14285 10887 ne
rect 14285 10789 14639 10887
tri 14639 10789 14737 10887 sw
tri 14737 10789 14835 10887 ne
rect 14835 10789 15189 10887
tri 15189 10789 15287 10887 sw
tri 15287 10789 15385 10887 ne
rect 15385 10789 15739 10887
tri 15739 10789 15837 10887 sw
tri 15837 10789 15935 10887 ne
rect 15935 10789 16289 10887
tri 16289 10789 16387 10887 sw
tri 16387 10789 16485 10887 ne
rect 16485 10789 16839 10887
tri 16839 10789 16937 10887 sw
tri 16937 10789 17035 10887 ne
rect 17035 10789 17389 10887
tri 17389 10789 17487 10887 sw
tri 17487 10789 17585 10887 ne
rect 17585 10789 17939 10887
tri 17939 10789 18037 10887 sw
tri 18037 10789 18135 10887 ne
rect 18135 10789 18489 10887
tri 18489 10789 18587 10887 sw
tri 18587 10789 18685 10887 ne
rect 18685 10789 19039 10887
tri 19039 10789 19137 10887 sw
tri 19137 10789 19235 10887 ne
rect 19235 10789 19589 10887
tri 19589 10789 19687 10887 sw
rect 20800 10789 21800 11437
rect -2000 10785 437 10789
rect -2000 10665 215 10785
rect 335 10691 437 10785
tri 437 10691 535 10789 sw
tri 535 10691 633 10789 ne
rect 633 10785 987 10789
rect 633 10691 765 10785
rect 335 10665 535 10691
rect -2000 10661 535 10665
rect -2000 10013 -1000 10661
tri 113 10563 211 10661 ne
rect 211 10613 535 10661
tri 535 10613 613 10691 sw
tri 633 10613 711 10691 ne
rect 711 10665 765 10691
rect 885 10691 987 10785
tri 987 10691 1085 10789 sw
tri 1085 10691 1183 10789 ne
rect 1183 10785 1537 10789
rect 1183 10691 1315 10785
rect 885 10665 1085 10691
rect 711 10613 1085 10665
tri 1085 10613 1163 10691 sw
tri 1183 10613 1261 10691 ne
rect 1261 10665 1315 10691
rect 1435 10691 1537 10785
tri 1537 10691 1635 10789 sw
tri 1635 10691 1733 10789 ne
rect 1733 10785 2087 10789
rect 1733 10691 1865 10785
rect 1435 10665 1635 10691
rect 1261 10613 1635 10665
tri 1635 10613 1713 10691 sw
tri 1733 10613 1811 10691 ne
rect 1811 10665 1865 10691
rect 1985 10691 2087 10785
tri 2087 10691 2185 10789 sw
tri 2185 10691 2283 10789 ne
rect 2283 10785 2637 10789
rect 2283 10691 2415 10785
rect 1985 10665 2185 10691
rect 1811 10613 2185 10665
tri 2185 10613 2263 10691 sw
tri 2283 10613 2361 10691 ne
rect 2361 10665 2415 10691
rect 2535 10691 2637 10785
tri 2637 10691 2735 10789 sw
tri 2735 10691 2833 10789 ne
rect 2833 10785 3187 10789
rect 2833 10691 2965 10785
rect 2535 10665 2735 10691
rect 2361 10613 2735 10665
tri 2735 10613 2813 10691 sw
tri 2833 10613 2911 10691 ne
rect 2911 10665 2965 10691
rect 3085 10691 3187 10785
tri 3187 10691 3285 10789 sw
tri 3285 10691 3383 10789 ne
rect 3383 10785 3737 10789
rect 3383 10691 3515 10785
rect 3085 10665 3285 10691
rect 2911 10613 3285 10665
tri 3285 10613 3363 10691 sw
tri 3383 10613 3461 10691 ne
rect 3461 10665 3515 10691
rect 3635 10691 3737 10785
tri 3737 10691 3835 10789 sw
tri 3835 10691 3933 10789 ne
rect 3933 10785 4287 10789
rect 3933 10691 4065 10785
rect 3635 10665 3835 10691
rect 3461 10613 3835 10665
tri 3835 10613 3913 10691 sw
tri 3933 10613 4011 10691 ne
rect 4011 10665 4065 10691
rect 4185 10691 4287 10785
tri 4287 10691 4385 10789 sw
tri 4385 10691 4483 10789 ne
rect 4483 10785 4837 10789
rect 4483 10691 4615 10785
rect 4185 10665 4385 10691
rect 4011 10613 4385 10665
tri 4385 10613 4463 10691 sw
tri 4483 10613 4561 10691 ne
rect 4561 10665 4615 10691
rect 4735 10691 4837 10785
tri 4837 10691 4935 10789 sw
tri 4935 10691 5033 10789 ne
rect 5033 10785 5387 10789
rect 5033 10691 5165 10785
rect 4735 10665 4935 10691
rect 4561 10613 4935 10665
tri 4935 10613 5013 10691 sw
tri 5033 10613 5111 10691 ne
rect 5111 10665 5165 10691
rect 5285 10691 5387 10785
tri 5387 10691 5485 10789 sw
tri 5485 10691 5583 10789 ne
rect 5583 10785 5937 10789
rect 5583 10691 5715 10785
rect 5285 10665 5485 10691
rect 5111 10613 5485 10665
tri 5485 10613 5563 10691 sw
tri 5583 10613 5661 10691 ne
rect 5661 10665 5715 10691
rect 5835 10691 5937 10785
tri 5937 10691 6035 10789 sw
tri 6035 10691 6133 10789 ne
rect 6133 10785 6487 10789
rect 6133 10691 6265 10785
rect 5835 10665 6035 10691
rect 5661 10613 6035 10665
tri 6035 10613 6113 10691 sw
tri 6133 10613 6211 10691 ne
rect 6211 10665 6265 10691
rect 6385 10691 6487 10785
tri 6487 10691 6585 10789 sw
tri 6585 10691 6683 10789 ne
rect 6683 10785 7037 10789
rect 6683 10691 6815 10785
rect 6385 10665 6585 10691
rect 6211 10613 6585 10665
tri 6585 10613 6663 10691 sw
tri 6683 10613 6761 10691 ne
rect 6761 10665 6815 10691
rect 6935 10691 7037 10785
tri 7037 10691 7135 10789 sw
tri 7135 10691 7233 10789 ne
rect 7233 10785 7587 10789
rect 7233 10691 7365 10785
rect 6935 10665 7135 10691
rect 6761 10613 7135 10665
tri 7135 10613 7213 10691 sw
tri 7233 10613 7311 10691 ne
rect 7311 10665 7365 10691
rect 7485 10691 7587 10785
tri 7587 10691 7685 10789 sw
tri 7685 10691 7783 10789 ne
rect 7783 10785 8137 10789
rect 7783 10691 7915 10785
rect 7485 10665 7685 10691
rect 7311 10613 7685 10665
tri 7685 10613 7763 10691 sw
tri 7783 10613 7861 10691 ne
rect 7861 10665 7915 10691
rect 8035 10691 8137 10785
tri 8137 10691 8235 10789 sw
tri 8235 10691 8333 10789 ne
rect 8333 10785 8687 10789
rect 8333 10691 8465 10785
rect 8035 10665 8235 10691
rect 7861 10613 8235 10665
tri 8235 10613 8313 10691 sw
tri 8333 10613 8411 10691 ne
rect 8411 10665 8465 10691
rect 8585 10691 8687 10785
tri 8687 10691 8785 10789 sw
tri 8785 10691 8883 10789 ne
rect 8883 10785 9237 10789
rect 8883 10691 9015 10785
rect 8585 10665 8785 10691
rect 8411 10613 8785 10665
tri 8785 10613 8863 10691 sw
tri 8883 10613 8961 10691 ne
rect 8961 10665 9015 10691
rect 9135 10691 9237 10785
tri 9237 10691 9335 10789 sw
tri 9335 10691 9433 10789 ne
rect 9433 10785 9787 10789
rect 9433 10691 9565 10785
rect 9135 10665 9335 10691
rect 8961 10613 9335 10665
tri 9335 10613 9413 10691 sw
tri 9433 10613 9511 10691 ne
rect 9511 10665 9565 10691
rect 9685 10691 9787 10785
tri 9787 10691 9885 10789 sw
tri 9885 10691 9983 10789 ne
rect 9983 10785 10337 10789
rect 9983 10691 10115 10785
rect 9685 10665 9885 10691
rect 9511 10613 9885 10665
tri 9885 10613 9963 10691 sw
tri 9983 10613 10061 10691 ne
rect 10061 10665 10115 10691
rect 10235 10691 10337 10785
tri 10337 10691 10435 10789 sw
tri 10435 10691 10533 10789 ne
rect 10533 10785 10887 10789
rect 10533 10691 10665 10785
rect 10235 10665 10435 10691
rect 10061 10613 10435 10665
tri 10435 10613 10513 10691 sw
tri 10533 10613 10611 10691 ne
rect 10611 10665 10665 10691
rect 10785 10691 10887 10785
tri 10887 10691 10985 10789 sw
tri 10985 10691 11083 10789 ne
rect 11083 10785 11437 10789
rect 11083 10691 11215 10785
rect 10785 10665 10985 10691
rect 10611 10613 10985 10665
tri 10985 10613 11063 10691 sw
tri 11083 10613 11161 10691 ne
rect 11161 10665 11215 10691
rect 11335 10691 11437 10785
tri 11437 10691 11535 10789 sw
tri 11535 10691 11633 10789 ne
rect 11633 10785 11987 10789
rect 11633 10691 11765 10785
rect 11335 10665 11535 10691
rect 11161 10613 11535 10665
tri 11535 10613 11613 10691 sw
tri 11633 10613 11711 10691 ne
rect 11711 10665 11765 10691
rect 11885 10691 11987 10785
tri 11987 10691 12085 10789 sw
tri 12085 10691 12183 10789 ne
rect 12183 10785 12537 10789
rect 12183 10691 12315 10785
rect 11885 10665 12085 10691
rect 11711 10613 12085 10665
tri 12085 10613 12163 10691 sw
tri 12183 10613 12261 10691 ne
rect 12261 10665 12315 10691
rect 12435 10691 12537 10785
tri 12537 10691 12635 10789 sw
tri 12635 10691 12733 10789 ne
rect 12733 10785 13087 10789
rect 12733 10691 12865 10785
rect 12435 10665 12635 10691
rect 12261 10613 12635 10665
tri 12635 10613 12713 10691 sw
tri 12733 10613 12811 10691 ne
rect 12811 10665 12865 10691
rect 12985 10691 13087 10785
tri 13087 10691 13185 10789 sw
tri 13185 10691 13283 10789 ne
rect 13283 10785 13637 10789
rect 13283 10691 13415 10785
rect 12985 10665 13185 10691
rect 12811 10613 13185 10665
tri 13185 10613 13263 10691 sw
tri 13283 10613 13361 10691 ne
rect 13361 10665 13415 10691
rect 13535 10691 13637 10785
tri 13637 10691 13735 10789 sw
tri 13735 10691 13833 10789 ne
rect 13833 10785 14187 10789
rect 13833 10691 13965 10785
rect 13535 10665 13735 10691
rect 13361 10613 13735 10665
tri 13735 10613 13813 10691 sw
tri 13833 10613 13911 10691 ne
rect 13911 10665 13965 10691
rect 14085 10691 14187 10785
tri 14187 10691 14285 10789 sw
tri 14285 10691 14383 10789 ne
rect 14383 10785 14737 10789
rect 14383 10691 14515 10785
rect 14085 10665 14285 10691
rect 13911 10613 14285 10665
tri 14285 10613 14363 10691 sw
tri 14383 10613 14461 10691 ne
rect 14461 10665 14515 10691
rect 14635 10691 14737 10785
tri 14737 10691 14835 10789 sw
tri 14835 10691 14933 10789 ne
rect 14933 10785 15287 10789
rect 14933 10691 15065 10785
rect 14635 10665 14835 10691
rect 14461 10613 14835 10665
tri 14835 10613 14913 10691 sw
tri 14933 10613 15011 10691 ne
rect 15011 10665 15065 10691
rect 15185 10691 15287 10785
tri 15287 10691 15385 10789 sw
tri 15385 10691 15483 10789 ne
rect 15483 10785 15837 10789
rect 15483 10691 15615 10785
rect 15185 10665 15385 10691
rect 15011 10613 15385 10665
tri 15385 10613 15463 10691 sw
tri 15483 10613 15561 10691 ne
rect 15561 10665 15615 10691
rect 15735 10691 15837 10785
tri 15837 10691 15935 10789 sw
tri 15935 10691 16033 10789 ne
rect 16033 10785 16387 10789
rect 16033 10691 16165 10785
rect 15735 10665 15935 10691
rect 15561 10613 15935 10665
tri 15935 10613 16013 10691 sw
tri 16033 10613 16111 10691 ne
rect 16111 10665 16165 10691
rect 16285 10691 16387 10785
tri 16387 10691 16485 10789 sw
tri 16485 10691 16583 10789 ne
rect 16583 10785 16937 10789
rect 16583 10691 16715 10785
rect 16285 10665 16485 10691
rect 16111 10613 16485 10665
tri 16485 10613 16563 10691 sw
tri 16583 10613 16661 10691 ne
rect 16661 10665 16715 10691
rect 16835 10691 16937 10785
tri 16937 10691 17035 10789 sw
tri 17035 10691 17133 10789 ne
rect 17133 10785 17487 10789
rect 17133 10691 17265 10785
rect 16835 10665 17035 10691
rect 16661 10613 17035 10665
tri 17035 10613 17113 10691 sw
tri 17133 10613 17211 10691 ne
rect 17211 10665 17265 10691
rect 17385 10691 17487 10785
tri 17487 10691 17585 10789 sw
tri 17585 10691 17683 10789 ne
rect 17683 10785 18037 10789
rect 17683 10691 17815 10785
rect 17385 10665 17585 10691
rect 17211 10613 17585 10665
tri 17585 10613 17663 10691 sw
tri 17683 10613 17761 10691 ne
rect 17761 10665 17815 10691
rect 17935 10691 18037 10785
tri 18037 10691 18135 10789 sw
tri 18135 10691 18233 10789 ne
rect 18233 10785 18587 10789
rect 18233 10691 18365 10785
rect 17935 10665 18135 10691
rect 17761 10613 18135 10665
tri 18135 10613 18213 10691 sw
tri 18233 10613 18311 10691 ne
rect 18311 10665 18365 10691
rect 18485 10691 18587 10785
tri 18587 10691 18685 10789 sw
tri 18685 10691 18783 10789 ne
rect 18783 10785 19137 10789
rect 18783 10691 18915 10785
rect 18485 10665 18685 10691
rect 18311 10613 18685 10665
tri 18685 10613 18763 10691 sw
tri 18783 10613 18861 10691 ne
rect 18861 10665 18915 10691
rect 19035 10691 19137 10785
tri 19137 10691 19235 10789 sw
tri 19235 10691 19333 10789 ne
rect 19333 10785 21800 10789
rect 19333 10691 19465 10785
rect 19035 10665 19235 10691
rect 18861 10613 19235 10665
tri 19235 10613 19313 10691 sw
tri 19333 10613 19411 10691 ne
rect 19411 10665 19465 10691
rect 19585 10665 21800 10785
rect 19411 10613 21800 10665
rect 211 10563 613 10613
rect -500 10513 113 10563
tri 113 10513 163 10563 sw
tri 211 10513 261 10563 ne
rect 261 10533 613 10563
tri 613 10533 693 10613 sw
tri 711 10533 791 10613 ne
rect 791 10533 1163 10613
tri 1163 10533 1243 10613 sw
tri 1261 10533 1341 10613 ne
rect 1341 10533 1713 10613
tri 1713 10533 1793 10613 sw
tri 1811 10533 1891 10613 ne
rect 1891 10533 2263 10613
tri 2263 10533 2343 10613 sw
tri 2361 10533 2441 10613 ne
rect 2441 10533 2813 10613
tri 2813 10533 2893 10613 sw
tri 2911 10533 2991 10613 ne
rect 2991 10533 3363 10613
tri 3363 10533 3443 10613 sw
tri 3461 10533 3541 10613 ne
rect 3541 10533 3913 10613
tri 3913 10533 3993 10613 sw
tri 4011 10533 4091 10613 ne
rect 4091 10533 4463 10613
tri 4463 10533 4543 10613 sw
tri 4561 10533 4641 10613 ne
rect 4641 10533 5013 10613
tri 5013 10533 5093 10613 sw
tri 5111 10533 5191 10613 ne
rect 5191 10533 5563 10613
tri 5563 10533 5643 10613 sw
tri 5661 10533 5741 10613 ne
rect 5741 10533 6113 10613
tri 6113 10533 6193 10613 sw
tri 6211 10533 6291 10613 ne
rect 6291 10533 6663 10613
tri 6663 10533 6743 10613 sw
tri 6761 10533 6841 10613 ne
rect 6841 10533 7213 10613
tri 7213 10533 7293 10613 sw
tri 7311 10533 7391 10613 ne
rect 7391 10533 7763 10613
tri 7763 10533 7843 10613 sw
tri 7861 10533 7941 10613 ne
rect 7941 10533 8313 10613
tri 8313 10533 8393 10613 sw
tri 8411 10533 8491 10613 ne
rect 8491 10533 8863 10613
tri 8863 10533 8943 10613 sw
tri 8961 10533 9041 10613 ne
rect 9041 10533 9413 10613
tri 9413 10533 9493 10613 sw
tri 9511 10533 9591 10613 ne
rect 9591 10533 9963 10613
tri 9963 10533 10043 10613 sw
tri 10061 10533 10141 10613 ne
rect 10141 10533 10513 10613
tri 10513 10533 10593 10613 sw
tri 10611 10533 10691 10613 ne
rect 10691 10533 11063 10613
tri 11063 10533 11143 10613 sw
tri 11161 10533 11241 10613 ne
rect 11241 10533 11613 10613
tri 11613 10533 11693 10613 sw
tri 11711 10533 11791 10613 ne
rect 11791 10533 12163 10613
tri 12163 10533 12243 10613 sw
tri 12261 10533 12341 10613 ne
rect 12341 10533 12713 10613
tri 12713 10533 12793 10613 sw
tri 12811 10533 12891 10613 ne
rect 12891 10533 13263 10613
tri 13263 10533 13343 10613 sw
tri 13361 10533 13441 10613 ne
rect 13441 10533 13813 10613
tri 13813 10533 13893 10613 sw
tri 13911 10533 13991 10613 ne
rect 13991 10533 14363 10613
tri 14363 10533 14443 10613 sw
tri 14461 10533 14541 10613 ne
rect 14541 10533 14913 10613
tri 14913 10533 14993 10613 sw
tri 15011 10533 15091 10613 ne
rect 15091 10533 15463 10613
tri 15463 10533 15543 10613 sw
tri 15561 10533 15641 10613 ne
rect 15641 10533 16013 10613
tri 16013 10533 16093 10613 sw
tri 16111 10533 16191 10613 ne
rect 16191 10533 16563 10613
tri 16563 10533 16643 10613 sw
tri 16661 10533 16741 10613 ne
rect 16741 10533 17113 10613
tri 17113 10533 17193 10613 sw
tri 17211 10533 17291 10613 ne
rect 17291 10533 17663 10613
tri 17663 10533 17743 10613 sw
tri 17761 10533 17841 10613 ne
rect 17841 10533 18213 10613
tri 18213 10533 18293 10613 sw
tri 18311 10533 18391 10613 ne
rect 18391 10533 18763 10613
tri 18763 10533 18843 10613 sw
tri 18861 10533 18941 10613 ne
rect 18941 10533 19313 10613
tri 19313 10533 19393 10613 sw
tri 19411 10533 19491 10613 ne
rect 19491 10533 20100 10613
rect 261 10513 693 10533
rect -500 10435 163 10513
tri 163 10435 241 10513 sw
tri 261 10435 339 10513 ne
rect 339 10435 693 10513
tri 693 10435 791 10533 sw
tri 791 10435 889 10533 ne
rect 889 10435 1243 10533
tri 1243 10435 1341 10533 sw
tri 1341 10435 1439 10533 ne
rect 1439 10435 1793 10533
tri 1793 10435 1891 10533 sw
tri 1891 10435 1989 10533 ne
rect 1989 10435 2343 10533
tri 2343 10435 2441 10533 sw
tri 2441 10435 2539 10533 ne
rect 2539 10435 2893 10533
tri 2893 10435 2991 10533 sw
tri 2991 10435 3089 10533 ne
rect 3089 10435 3443 10533
tri 3443 10435 3541 10533 sw
tri 3541 10435 3639 10533 ne
rect 3639 10435 3993 10533
tri 3993 10435 4091 10533 sw
tri 4091 10435 4189 10533 ne
rect 4189 10435 4543 10533
tri 4543 10435 4641 10533 sw
tri 4641 10435 4739 10533 ne
rect 4739 10435 5093 10533
tri 5093 10435 5191 10533 sw
tri 5191 10435 5289 10533 ne
rect 5289 10435 5643 10533
tri 5643 10435 5741 10533 sw
tri 5741 10435 5839 10533 ne
rect 5839 10435 6193 10533
tri 6193 10435 6291 10533 sw
tri 6291 10435 6389 10533 ne
rect 6389 10435 6743 10533
tri 6743 10435 6841 10533 sw
tri 6841 10435 6939 10533 ne
rect 6939 10435 7293 10533
tri 7293 10435 7391 10533 sw
tri 7391 10435 7489 10533 ne
rect 7489 10435 7843 10533
tri 7843 10435 7941 10533 sw
tri 7941 10435 8039 10533 ne
rect 8039 10435 8393 10533
tri 8393 10435 8491 10533 sw
tri 8491 10435 8589 10533 ne
rect 8589 10435 8943 10533
tri 8943 10435 9041 10533 sw
tri 9041 10435 9139 10533 ne
rect 9139 10435 9493 10533
tri 9493 10435 9591 10533 sw
tri 9591 10435 9689 10533 ne
rect 9689 10435 10043 10533
tri 10043 10435 10141 10533 sw
tri 10141 10435 10239 10533 ne
rect 10239 10435 10593 10533
tri 10593 10435 10691 10533 sw
tri 10691 10435 10789 10533 ne
rect 10789 10435 11143 10533
tri 11143 10435 11241 10533 sw
tri 11241 10435 11339 10533 ne
rect 11339 10435 11693 10533
tri 11693 10435 11791 10533 sw
tri 11791 10435 11889 10533 ne
rect 11889 10435 12243 10533
tri 12243 10435 12341 10533 sw
tri 12341 10435 12439 10533 ne
rect 12439 10435 12793 10533
tri 12793 10435 12891 10533 sw
tri 12891 10435 12989 10533 ne
rect 12989 10435 13343 10533
tri 13343 10435 13441 10533 sw
tri 13441 10435 13539 10533 ne
rect 13539 10435 13893 10533
tri 13893 10435 13991 10533 sw
tri 13991 10435 14089 10533 ne
rect 14089 10435 14443 10533
tri 14443 10435 14541 10533 sw
tri 14541 10435 14639 10533 ne
rect 14639 10435 14993 10533
tri 14993 10435 15091 10533 sw
tri 15091 10435 15189 10533 ne
rect 15189 10435 15543 10533
tri 15543 10435 15641 10533 sw
tri 15641 10435 15739 10533 ne
rect 15739 10435 16093 10533
tri 16093 10435 16191 10533 sw
tri 16191 10435 16289 10533 ne
rect 16289 10435 16643 10533
tri 16643 10435 16741 10533 sw
tri 16741 10435 16839 10533 ne
rect 16839 10435 17193 10533
tri 17193 10435 17291 10533 sw
tri 17291 10435 17389 10533 ne
rect 17389 10435 17743 10533
tri 17743 10435 17841 10533 sw
tri 17841 10435 17939 10533 ne
rect 17939 10435 18293 10533
tri 18293 10435 18391 10533 sw
tri 18391 10435 18489 10533 ne
rect 18489 10435 18843 10533
tri 18843 10435 18941 10533 sw
tri 18941 10435 19039 10533 ne
rect 19039 10435 19393 10533
tri 19393 10435 19491 10533 sw
tri 19491 10435 19589 10533 ne
rect 19589 10513 20100 10533
rect 20200 10513 21800 10613
rect 19589 10435 21800 10513
rect -500 10387 241 10435
rect -500 10287 -400 10387
rect -300 10337 241 10387
tri 241 10337 339 10435 sw
tri 339 10337 437 10435 ne
rect 437 10337 791 10435
tri 791 10337 889 10435 sw
tri 889 10337 987 10435 ne
rect 987 10337 1341 10435
tri 1341 10337 1439 10435 sw
tri 1439 10337 1537 10435 ne
rect 1537 10337 1891 10435
tri 1891 10337 1989 10435 sw
tri 1989 10337 2087 10435 ne
rect 2087 10337 2441 10435
tri 2441 10337 2539 10435 sw
tri 2539 10337 2637 10435 ne
rect 2637 10337 2991 10435
tri 2991 10337 3089 10435 sw
tri 3089 10337 3187 10435 ne
rect 3187 10337 3541 10435
tri 3541 10337 3639 10435 sw
tri 3639 10337 3737 10435 ne
rect 3737 10337 4091 10435
tri 4091 10337 4189 10435 sw
tri 4189 10337 4287 10435 ne
rect 4287 10337 4641 10435
tri 4641 10337 4739 10435 sw
tri 4739 10337 4837 10435 ne
rect 4837 10337 5191 10435
tri 5191 10337 5289 10435 sw
tri 5289 10337 5387 10435 ne
rect 5387 10337 5741 10435
tri 5741 10337 5839 10435 sw
tri 5839 10337 5937 10435 ne
rect 5937 10337 6291 10435
tri 6291 10337 6389 10435 sw
tri 6389 10337 6487 10435 ne
rect 6487 10337 6841 10435
tri 6841 10337 6939 10435 sw
tri 6939 10337 7037 10435 ne
rect 7037 10337 7391 10435
tri 7391 10337 7489 10435 sw
tri 7489 10337 7587 10435 ne
rect 7587 10337 7941 10435
tri 7941 10337 8039 10435 sw
tri 8039 10337 8137 10435 ne
rect 8137 10337 8491 10435
tri 8491 10337 8589 10435 sw
tri 8589 10337 8687 10435 ne
rect 8687 10337 9041 10435
tri 9041 10337 9139 10435 sw
tri 9139 10337 9237 10435 ne
rect 9237 10337 9591 10435
tri 9591 10337 9689 10435 sw
tri 9689 10337 9787 10435 ne
rect 9787 10337 10141 10435
tri 10141 10337 10239 10435 sw
tri 10239 10337 10337 10435 ne
rect 10337 10337 10691 10435
tri 10691 10337 10789 10435 sw
tri 10789 10337 10887 10435 ne
rect 10887 10337 11241 10435
tri 11241 10337 11339 10435 sw
tri 11339 10337 11437 10435 ne
rect 11437 10337 11791 10435
tri 11791 10337 11889 10435 sw
tri 11889 10337 11987 10435 ne
rect 11987 10337 12341 10435
tri 12341 10337 12439 10435 sw
tri 12439 10337 12537 10435 ne
rect 12537 10337 12891 10435
tri 12891 10337 12989 10435 sw
tri 12989 10337 13087 10435 ne
rect 13087 10337 13441 10435
tri 13441 10337 13539 10435 sw
tri 13539 10337 13637 10435 ne
rect 13637 10337 13991 10435
tri 13991 10337 14089 10435 sw
tri 14089 10337 14187 10435 ne
rect 14187 10337 14541 10435
tri 14541 10337 14639 10435 sw
tri 14639 10337 14737 10435 ne
rect 14737 10337 15091 10435
tri 15091 10337 15189 10435 sw
tri 15189 10337 15287 10435 ne
rect 15287 10337 15641 10435
tri 15641 10337 15739 10435 sw
tri 15739 10337 15837 10435 ne
rect 15837 10337 16191 10435
tri 16191 10337 16289 10435 sw
tri 16289 10337 16387 10435 ne
rect 16387 10337 16741 10435
tri 16741 10337 16839 10435 sw
tri 16839 10337 16937 10435 ne
rect 16937 10337 17291 10435
tri 17291 10337 17389 10435 sw
tri 17389 10337 17487 10435 ne
rect 17487 10337 17841 10435
tri 17841 10337 17939 10435 sw
tri 17939 10337 18037 10435 ne
rect 18037 10337 18391 10435
tri 18391 10337 18489 10435 sw
tri 18489 10337 18587 10435 ne
rect 18587 10337 18941 10435
tri 18941 10337 19039 10435 sw
tri 19039 10337 19137 10435 ne
rect 19137 10337 19491 10435
tri 19491 10337 19589 10435 sw
tri 19589 10337 19687 10435 ne
rect 19687 10337 21800 10435
rect -300 10287 339 10337
rect -500 10239 339 10287
tri 339 10239 437 10337 sw
tri 437 10239 535 10337 ne
rect 535 10239 889 10337
tri 889 10239 987 10337 sw
tri 987 10239 1085 10337 ne
rect 1085 10239 1439 10337
tri 1439 10239 1537 10337 sw
tri 1537 10239 1635 10337 ne
rect 1635 10239 1989 10337
tri 1989 10239 2087 10337 sw
tri 2087 10239 2185 10337 ne
rect 2185 10239 2539 10337
tri 2539 10239 2637 10337 sw
tri 2637 10239 2735 10337 ne
rect 2735 10239 3089 10337
tri 3089 10239 3187 10337 sw
tri 3187 10239 3285 10337 ne
rect 3285 10239 3639 10337
tri 3639 10239 3737 10337 sw
tri 3737 10239 3835 10337 ne
rect 3835 10239 4189 10337
tri 4189 10239 4287 10337 sw
tri 4287 10239 4385 10337 ne
rect 4385 10239 4739 10337
tri 4739 10239 4837 10337 sw
tri 4837 10239 4935 10337 ne
rect 4935 10239 5289 10337
tri 5289 10239 5387 10337 sw
tri 5387 10239 5485 10337 ne
rect 5485 10239 5839 10337
tri 5839 10239 5937 10337 sw
tri 5937 10239 6035 10337 ne
rect 6035 10239 6389 10337
tri 6389 10239 6487 10337 sw
tri 6487 10239 6585 10337 ne
rect 6585 10239 6939 10337
tri 6939 10239 7037 10337 sw
tri 7037 10239 7135 10337 ne
rect 7135 10239 7489 10337
tri 7489 10239 7587 10337 sw
tri 7587 10239 7685 10337 ne
rect 7685 10239 8039 10337
tri 8039 10239 8137 10337 sw
tri 8137 10239 8235 10337 ne
rect 8235 10239 8589 10337
tri 8589 10239 8687 10337 sw
tri 8687 10239 8785 10337 ne
rect 8785 10239 9139 10337
tri 9139 10239 9237 10337 sw
tri 9237 10239 9335 10337 ne
rect 9335 10239 9689 10337
tri 9689 10239 9787 10337 sw
tri 9787 10239 9885 10337 ne
rect 9885 10239 10239 10337
tri 10239 10239 10337 10337 sw
tri 10337 10239 10435 10337 ne
rect 10435 10239 10789 10337
tri 10789 10239 10887 10337 sw
tri 10887 10239 10985 10337 ne
rect 10985 10239 11339 10337
tri 11339 10239 11437 10337 sw
tri 11437 10239 11535 10337 ne
rect 11535 10239 11889 10337
tri 11889 10239 11987 10337 sw
tri 11987 10239 12085 10337 ne
rect 12085 10239 12439 10337
tri 12439 10239 12537 10337 sw
tri 12537 10239 12635 10337 ne
rect 12635 10239 12989 10337
tri 12989 10239 13087 10337 sw
tri 13087 10239 13185 10337 ne
rect 13185 10239 13539 10337
tri 13539 10239 13637 10337 sw
tri 13637 10239 13735 10337 ne
rect 13735 10239 14089 10337
tri 14089 10239 14187 10337 sw
tri 14187 10239 14285 10337 ne
rect 14285 10239 14639 10337
tri 14639 10239 14737 10337 sw
tri 14737 10239 14835 10337 ne
rect 14835 10239 15189 10337
tri 15189 10239 15287 10337 sw
tri 15287 10239 15385 10337 ne
rect 15385 10239 15739 10337
tri 15739 10239 15837 10337 sw
tri 15837 10239 15935 10337 ne
rect 15935 10239 16289 10337
tri 16289 10239 16387 10337 sw
tri 16387 10239 16485 10337 ne
rect 16485 10239 16839 10337
tri 16839 10239 16937 10337 sw
tri 16937 10239 17035 10337 ne
rect 17035 10239 17389 10337
tri 17389 10239 17487 10337 sw
tri 17487 10239 17585 10337 ne
rect 17585 10239 17939 10337
tri 17939 10239 18037 10337 sw
tri 18037 10239 18135 10337 ne
rect 18135 10239 18489 10337
tri 18489 10239 18587 10337 sw
tri 18587 10239 18685 10337 ne
rect 18685 10239 19039 10337
tri 19039 10239 19137 10337 sw
tri 19137 10239 19235 10337 ne
rect 19235 10239 19589 10337
tri 19589 10239 19687 10337 sw
rect -500 10235 437 10239
rect -500 10115 215 10235
rect 335 10141 437 10235
tri 437 10141 535 10239 sw
tri 535 10141 633 10239 ne
rect 633 10235 987 10239
rect 633 10141 765 10235
rect 335 10115 535 10141
rect -500 10111 535 10115
tri 535 10111 565 10141 sw
tri 633 10111 663 10141 ne
rect 663 10115 765 10141
rect 885 10141 987 10235
tri 987 10141 1085 10239 sw
tri 1085 10141 1183 10239 ne
rect 1183 10235 1537 10239
rect 1183 10141 1315 10235
rect 885 10115 1085 10141
rect 663 10111 1085 10115
tri 1085 10111 1115 10141 sw
tri 1183 10111 1213 10141 ne
rect 1213 10115 1315 10141
rect 1435 10141 1537 10235
tri 1537 10141 1635 10239 sw
tri 1635 10141 1733 10239 ne
rect 1733 10235 2087 10239
rect 1733 10141 1865 10235
rect 1435 10115 1635 10141
rect 1213 10111 1635 10115
tri 1635 10111 1665 10141 sw
tri 1733 10111 1763 10141 ne
rect 1763 10115 1865 10141
rect 1985 10141 2087 10235
tri 2087 10141 2185 10239 sw
tri 2185 10141 2283 10239 ne
rect 2283 10235 2637 10239
rect 2283 10141 2415 10235
rect 1985 10115 2185 10141
rect 1763 10111 2185 10115
tri 2185 10111 2215 10141 sw
tri 2283 10111 2313 10141 ne
rect 2313 10115 2415 10141
rect 2535 10141 2637 10235
tri 2637 10141 2735 10239 sw
tri 2735 10141 2833 10239 ne
rect 2833 10235 3187 10239
rect 2833 10141 2965 10235
rect 2535 10115 2735 10141
rect 2313 10111 2735 10115
tri 2735 10111 2765 10141 sw
tri 2833 10111 2863 10141 ne
rect 2863 10115 2965 10141
rect 3085 10141 3187 10235
tri 3187 10141 3285 10239 sw
tri 3285 10141 3383 10239 ne
rect 3383 10235 3737 10239
rect 3383 10141 3515 10235
rect 3085 10115 3285 10141
rect 2863 10111 3285 10115
tri 3285 10111 3315 10141 sw
tri 3383 10111 3413 10141 ne
rect 3413 10115 3515 10141
rect 3635 10141 3737 10235
tri 3737 10141 3835 10239 sw
tri 3835 10141 3933 10239 ne
rect 3933 10235 4287 10239
rect 3933 10141 4065 10235
rect 3635 10115 3835 10141
rect 3413 10111 3835 10115
tri 3835 10111 3865 10141 sw
tri 3933 10111 3963 10141 ne
rect 3963 10115 4065 10141
rect 4185 10141 4287 10235
tri 4287 10141 4385 10239 sw
tri 4385 10141 4483 10239 ne
rect 4483 10235 4837 10239
rect 4483 10141 4615 10235
rect 4185 10115 4385 10141
rect 3963 10111 4385 10115
tri 4385 10111 4415 10141 sw
tri 4483 10111 4513 10141 ne
rect 4513 10115 4615 10141
rect 4735 10141 4837 10235
tri 4837 10141 4935 10239 sw
tri 4935 10141 5033 10239 ne
rect 5033 10235 5387 10239
rect 5033 10141 5165 10235
rect 4735 10115 4935 10141
rect 4513 10111 4935 10115
tri 4935 10111 4965 10141 sw
tri 5033 10111 5063 10141 ne
rect 5063 10115 5165 10141
rect 5285 10141 5387 10235
tri 5387 10141 5485 10239 sw
tri 5485 10141 5583 10239 ne
rect 5583 10235 5937 10239
rect 5583 10141 5715 10235
rect 5285 10115 5485 10141
rect 5063 10111 5485 10115
tri 5485 10111 5515 10141 sw
tri 5583 10111 5613 10141 ne
rect 5613 10115 5715 10141
rect 5835 10141 5937 10235
tri 5937 10141 6035 10239 sw
tri 6035 10141 6133 10239 ne
rect 6133 10235 6487 10239
rect 6133 10141 6265 10235
rect 5835 10115 6035 10141
rect 5613 10111 6035 10115
tri 6035 10111 6065 10141 sw
tri 6133 10111 6163 10141 ne
rect 6163 10115 6265 10141
rect 6385 10141 6487 10235
tri 6487 10141 6585 10239 sw
tri 6585 10141 6683 10239 ne
rect 6683 10235 7037 10239
rect 6683 10141 6815 10235
rect 6385 10115 6585 10141
rect 6163 10111 6585 10115
tri 6585 10111 6615 10141 sw
tri 6683 10111 6713 10141 ne
rect 6713 10115 6815 10141
rect 6935 10141 7037 10235
tri 7037 10141 7135 10239 sw
tri 7135 10141 7233 10239 ne
rect 7233 10235 7587 10239
rect 7233 10141 7365 10235
rect 6935 10115 7135 10141
rect 6713 10111 7135 10115
tri 7135 10111 7165 10141 sw
tri 7233 10111 7263 10141 ne
rect 7263 10115 7365 10141
rect 7485 10141 7587 10235
tri 7587 10141 7685 10239 sw
tri 7685 10141 7783 10239 ne
rect 7783 10235 8137 10239
rect 7783 10141 7915 10235
rect 7485 10115 7685 10141
rect 7263 10111 7685 10115
tri 7685 10111 7715 10141 sw
tri 7783 10111 7813 10141 ne
rect 7813 10115 7915 10141
rect 8035 10141 8137 10235
tri 8137 10141 8235 10239 sw
tri 8235 10141 8333 10239 ne
rect 8333 10235 8687 10239
rect 8333 10141 8465 10235
rect 8035 10115 8235 10141
rect 7813 10111 8235 10115
tri 8235 10111 8265 10141 sw
tri 8333 10111 8363 10141 ne
rect 8363 10115 8465 10141
rect 8585 10141 8687 10235
tri 8687 10141 8785 10239 sw
tri 8785 10141 8883 10239 ne
rect 8883 10235 9237 10239
rect 8883 10141 9015 10235
rect 8585 10115 8785 10141
rect 8363 10111 8785 10115
tri 8785 10111 8815 10141 sw
tri 8883 10111 8913 10141 ne
rect 8913 10115 9015 10141
rect 9135 10141 9237 10235
tri 9237 10141 9335 10239 sw
tri 9335 10141 9433 10239 ne
rect 9433 10235 9787 10239
rect 9433 10141 9565 10235
rect 9135 10115 9335 10141
rect 8913 10111 9335 10115
tri 9335 10111 9365 10141 sw
tri 9433 10111 9463 10141 ne
rect 9463 10115 9565 10141
rect 9685 10141 9787 10235
tri 9787 10141 9885 10239 sw
tri 9885 10141 9983 10239 ne
rect 9983 10235 10337 10239
rect 9983 10141 10115 10235
rect 9685 10115 9885 10141
rect 9463 10111 9885 10115
tri 9885 10111 9915 10141 sw
tri 9983 10111 10013 10141 ne
rect 10013 10115 10115 10141
rect 10235 10141 10337 10235
tri 10337 10141 10435 10239 sw
tri 10435 10141 10533 10239 ne
rect 10533 10235 10887 10239
rect 10533 10141 10665 10235
rect 10235 10115 10435 10141
rect 10013 10111 10435 10115
tri 10435 10111 10465 10141 sw
tri 10533 10111 10563 10141 ne
rect 10563 10115 10665 10141
rect 10785 10141 10887 10235
tri 10887 10141 10985 10239 sw
tri 10985 10141 11083 10239 ne
rect 11083 10235 11437 10239
rect 11083 10141 11215 10235
rect 10785 10115 10985 10141
rect 10563 10111 10985 10115
tri 10985 10111 11015 10141 sw
tri 11083 10111 11113 10141 ne
rect 11113 10115 11215 10141
rect 11335 10141 11437 10235
tri 11437 10141 11535 10239 sw
tri 11535 10141 11633 10239 ne
rect 11633 10235 11987 10239
rect 11633 10141 11765 10235
rect 11335 10115 11535 10141
rect 11113 10111 11535 10115
tri 11535 10111 11565 10141 sw
tri 11633 10111 11663 10141 ne
rect 11663 10115 11765 10141
rect 11885 10141 11987 10235
tri 11987 10141 12085 10239 sw
tri 12085 10141 12183 10239 ne
rect 12183 10235 12537 10239
rect 12183 10141 12315 10235
rect 11885 10115 12085 10141
rect 11663 10111 12085 10115
tri 12085 10111 12115 10141 sw
tri 12183 10111 12213 10141 ne
rect 12213 10115 12315 10141
rect 12435 10141 12537 10235
tri 12537 10141 12635 10239 sw
tri 12635 10141 12733 10239 ne
rect 12733 10235 13087 10239
rect 12733 10141 12865 10235
rect 12435 10115 12635 10141
rect 12213 10111 12635 10115
tri 12635 10111 12665 10141 sw
tri 12733 10111 12763 10141 ne
rect 12763 10115 12865 10141
rect 12985 10141 13087 10235
tri 13087 10141 13185 10239 sw
tri 13185 10141 13283 10239 ne
rect 13283 10235 13637 10239
rect 13283 10141 13415 10235
rect 12985 10115 13185 10141
rect 12763 10111 13185 10115
tri 13185 10111 13215 10141 sw
tri 13283 10111 13313 10141 ne
rect 13313 10115 13415 10141
rect 13535 10141 13637 10235
tri 13637 10141 13735 10239 sw
tri 13735 10141 13833 10239 ne
rect 13833 10235 14187 10239
rect 13833 10141 13965 10235
rect 13535 10115 13735 10141
rect 13313 10111 13735 10115
tri 13735 10111 13765 10141 sw
tri 13833 10111 13863 10141 ne
rect 13863 10115 13965 10141
rect 14085 10141 14187 10235
tri 14187 10141 14285 10239 sw
tri 14285 10141 14383 10239 ne
rect 14383 10235 14737 10239
rect 14383 10141 14515 10235
rect 14085 10115 14285 10141
rect 13863 10111 14285 10115
tri 14285 10111 14315 10141 sw
tri 14383 10111 14413 10141 ne
rect 14413 10115 14515 10141
rect 14635 10141 14737 10235
tri 14737 10141 14835 10239 sw
tri 14835 10141 14933 10239 ne
rect 14933 10235 15287 10239
rect 14933 10141 15065 10235
rect 14635 10115 14835 10141
rect 14413 10111 14835 10115
tri 14835 10111 14865 10141 sw
tri 14933 10111 14963 10141 ne
rect 14963 10115 15065 10141
rect 15185 10141 15287 10235
tri 15287 10141 15385 10239 sw
tri 15385 10141 15483 10239 ne
rect 15483 10235 15837 10239
rect 15483 10141 15615 10235
rect 15185 10115 15385 10141
rect 14963 10111 15385 10115
tri 15385 10111 15415 10141 sw
tri 15483 10111 15513 10141 ne
rect 15513 10115 15615 10141
rect 15735 10141 15837 10235
tri 15837 10141 15935 10239 sw
tri 15935 10141 16033 10239 ne
rect 16033 10235 16387 10239
rect 16033 10141 16165 10235
rect 15735 10115 15935 10141
rect 15513 10111 15935 10115
tri 15935 10111 15965 10141 sw
tri 16033 10111 16063 10141 ne
rect 16063 10115 16165 10141
rect 16285 10141 16387 10235
tri 16387 10141 16485 10239 sw
tri 16485 10141 16583 10239 ne
rect 16583 10235 16937 10239
rect 16583 10141 16715 10235
rect 16285 10115 16485 10141
rect 16063 10111 16485 10115
tri 16485 10111 16515 10141 sw
tri 16583 10111 16613 10141 ne
rect 16613 10115 16715 10141
rect 16835 10141 16937 10235
tri 16937 10141 17035 10239 sw
tri 17035 10141 17133 10239 ne
rect 17133 10235 17487 10239
rect 17133 10141 17265 10235
rect 16835 10115 17035 10141
rect 16613 10111 17035 10115
tri 17035 10111 17065 10141 sw
tri 17133 10111 17163 10141 ne
rect 17163 10115 17265 10141
rect 17385 10141 17487 10235
tri 17487 10141 17585 10239 sw
tri 17585 10141 17683 10239 ne
rect 17683 10235 18037 10239
rect 17683 10141 17815 10235
rect 17385 10115 17585 10141
rect 17163 10111 17585 10115
tri 17585 10111 17615 10141 sw
tri 17683 10111 17713 10141 ne
rect 17713 10115 17815 10141
rect 17935 10141 18037 10235
tri 18037 10141 18135 10239 sw
tri 18135 10141 18233 10239 ne
rect 18233 10235 18587 10239
rect 18233 10141 18365 10235
rect 17935 10115 18135 10141
rect 17713 10111 18135 10115
tri 18135 10111 18165 10141 sw
tri 18233 10111 18263 10141 ne
rect 18263 10115 18365 10141
rect 18485 10141 18587 10235
tri 18587 10141 18685 10239 sw
tri 18685 10141 18783 10239 ne
rect 18783 10235 19137 10239
rect 18783 10141 18915 10235
rect 18485 10115 18685 10141
rect 18263 10111 18685 10115
tri 18685 10111 18715 10141 sw
tri 18783 10111 18813 10141 ne
rect 18813 10115 18915 10141
rect 19035 10141 19137 10235
tri 19137 10141 19235 10239 sw
tri 19235 10141 19333 10239 ne
rect 19333 10235 20300 10239
rect 19333 10141 19465 10235
rect 19035 10115 19235 10141
rect 18813 10111 19235 10115
tri 19235 10111 19265 10141 sw
tri 19333 10111 19363 10141 ne
rect 19363 10115 19465 10141
rect 19585 10115 20300 10235
rect 19363 10111 20300 10115
tri 113 10013 211 10111 ne
rect 211 10013 565 10111
tri 565 10013 663 10111 sw
tri 663 10013 761 10111 ne
rect 761 10013 1115 10111
tri 1115 10013 1213 10111 sw
tri 1213 10013 1311 10111 ne
rect 1311 10013 1665 10111
tri 1665 10013 1763 10111 sw
tri 1763 10013 1861 10111 ne
rect 1861 10013 2215 10111
tri 2215 10013 2313 10111 sw
tri 2313 10013 2411 10111 ne
rect 2411 10013 2765 10111
tri 2765 10013 2863 10111 sw
tri 2863 10013 2961 10111 ne
rect 2961 10013 3315 10111
tri 3315 10013 3413 10111 sw
tri 3413 10013 3511 10111 ne
rect 3511 10013 3865 10111
tri 3865 10013 3963 10111 sw
tri 3963 10013 4061 10111 ne
rect 4061 10013 4415 10111
tri 4415 10013 4513 10111 sw
tri 4513 10013 4611 10111 ne
rect 4611 10013 4965 10111
tri 4965 10013 5063 10111 sw
tri 5063 10013 5161 10111 ne
rect 5161 10013 5515 10111
tri 5515 10013 5613 10111 sw
tri 5613 10013 5711 10111 ne
rect 5711 10013 6065 10111
tri 6065 10013 6163 10111 sw
tri 6163 10013 6261 10111 ne
rect 6261 10013 6615 10111
tri 6615 10013 6713 10111 sw
tri 6713 10013 6811 10111 ne
rect 6811 10013 7165 10111
tri 7165 10013 7263 10111 sw
tri 7263 10013 7361 10111 ne
rect 7361 10013 7715 10111
tri 7715 10013 7813 10111 sw
tri 7813 10013 7911 10111 ne
rect 7911 10013 8265 10111
tri 8265 10013 8363 10111 sw
tri 8363 10013 8461 10111 ne
rect 8461 10013 8815 10111
tri 8815 10013 8913 10111 sw
tri 8913 10013 9011 10111 ne
rect 9011 10013 9365 10111
tri 9365 10013 9463 10111 sw
tri 9463 10013 9561 10111 ne
rect 9561 10013 9915 10111
tri 9915 10013 10013 10111 sw
tri 10013 10013 10111 10111 ne
rect 10111 10013 10465 10111
tri 10465 10013 10563 10111 sw
tri 10563 10013 10661 10111 ne
rect 10661 10013 11015 10111
tri 11015 10013 11113 10111 sw
tri 11113 10013 11211 10111 ne
rect 11211 10013 11565 10111
tri 11565 10013 11663 10111 sw
tri 11663 10013 11761 10111 ne
rect 11761 10013 12115 10111
tri 12115 10013 12213 10111 sw
tri 12213 10013 12311 10111 ne
rect 12311 10013 12665 10111
tri 12665 10013 12763 10111 sw
tri 12763 10013 12861 10111 ne
rect 12861 10013 13215 10111
tri 13215 10013 13313 10111 sw
tri 13313 10013 13411 10111 ne
rect 13411 10013 13765 10111
tri 13765 10013 13863 10111 sw
tri 13863 10013 13961 10111 ne
rect 13961 10013 14315 10111
tri 14315 10013 14413 10111 sw
tri 14413 10013 14511 10111 ne
rect 14511 10013 14865 10111
tri 14865 10013 14963 10111 sw
tri 14963 10013 15061 10111 ne
rect 15061 10013 15415 10111
tri 15415 10013 15513 10111 sw
tri 15513 10013 15611 10111 ne
rect 15611 10013 15965 10111
tri 15965 10013 16063 10111 sw
tri 16063 10013 16161 10111 ne
rect 16161 10013 16515 10111
tri 16515 10013 16613 10111 sw
tri 16613 10013 16711 10111 ne
rect 16711 10013 17065 10111
tri 17065 10013 17163 10111 sw
tri 17163 10013 17261 10111 ne
rect 17261 10013 17615 10111
tri 17615 10013 17713 10111 sw
tri 17713 10013 17811 10111 ne
rect 17811 10013 18165 10111
tri 18165 10013 18263 10111 sw
tri 18263 10013 18361 10111 ne
rect 18361 10013 18715 10111
tri 18715 10013 18813 10111 sw
tri 18813 10013 18911 10111 ne
rect 18911 10013 19265 10111
tri 19265 10013 19363 10111 sw
tri 19363 10013 19461 10111 ne
rect 19461 10013 20300 10111
rect -2000 9983 113 10013
tri 113 9983 143 10013 sw
tri 211 9983 241 10013 ne
rect 241 9983 663 10013
tri 663 9983 693 10013 sw
tri 761 9983 791 10013 ne
rect 791 9983 1213 10013
tri 1213 9983 1243 10013 sw
tri 1311 9983 1341 10013 ne
rect 1341 9983 1763 10013
tri 1763 9983 1793 10013 sw
tri 1861 9983 1891 10013 ne
rect 1891 9983 2313 10013
tri 2313 9983 2343 10013 sw
tri 2411 9983 2441 10013 ne
rect 2441 9983 2863 10013
tri 2863 9983 2893 10013 sw
tri 2961 9983 2991 10013 ne
rect 2991 9983 3413 10013
tri 3413 9983 3443 10013 sw
tri 3511 9983 3541 10013 ne
rect 3541 9983 3963 10013
tri 3963 9983 3993 10013 sw
tri 4061 9983 4091 10013 ne
rect 4091 9983 4513 10013
tri 4513 9983 4543 10013 sw
tri 4611 9983 4641 10013 ne
rect 4641 9983 5063 10013
tri 5063 9983 5093 10013 sw
tri 5161 9983 5191 10013 ne
rect 5191 9983 5613 10013
tri 5613 9983 5643 10013 sw
tri 5711 9983 5741 10013 ne
rect 5741 9983 6163 10013
tri 6163 9983 6193 10013 sw
tri 6261 9983 6291 10013 ne
rect 6291 9983 6713 10013
tri 6713 9983 6743 10013 sw
tri 6811 9983 6841 10013 ne
rect 6841 9983 7263 10013
tri 7263 9983 7293 10013 sw
tri 7361 9983 7391 10013 ne
rect 7391 9983 7813 10013
tri 7813 9983 7843 10013 sw
tri 7911 9983 7941 10013 ne
rect 7941 9983 8363 10013
tri 8363 9983 8393 10013 sw
tri 8461 9983 8491 10013 ne
rect 8491 9983 8913 10013
tri 8913 9983 8943 10013 sw
tri 9011 9983 9041 10013 ne
rect 9041 9983 9463 10013
tri 9463 9983 9493 10013 sw
tri 9561 9983 9591 10013 ne
rect 9591 9983 10013 10013
tri 10013 9983 10043 10013 sw
tri 10111 9983 10141 10013 ne
rect 10141 9983 10563 10013
tri 10563 9983 10593 10013 sw
tri 10661 9983 10691 10013 ne
rect 10691 9983 11113 10013
tri 11113 9983 11143 10013 sw
tri 11211 9983 11241 10013 ne
rect 11241 9983 11663 10013
tri 11663 9983 11693 10013 sw
tri 11761 9983 11791 10013 ne
rect 11791 9983 12213 10013
tri 12213 9983 12243 10013 sw
tri 12311 9983 12341 10013 ne
rect 12341 9983 12763 10013
tri 12763 9983 12793 10013 sw
tri 12861 9983 12891 10013 ne
rect 12891 9983 13313 10013
tri 13313 9983 13343 10013 sw
tri 13411 9983 13441 10013 ne
rect 13441 9983 13863 10013
tri 13863 9983 13893 10013 sw
tri 13961 9983 13991 10013 ne
rect 13991 9983 14413 10013
tri 14413 9983 14443 10013 sw
tri 14511 9983 14541 10013 ne
rect 14541 9983 14963 10013
tri 14963 9983 14993 10013 sw
tri 15061 9983 15091 10013 ne
rect 15091 9983 15513 10013
tri 15513 9983 15543 10013 sw
tri 15611 9983 15641 10013 ne
rect 15641 9983 16063 10013
tri 16063 9983 16093 10013 sw
tri 16161 9983 16191 10013 ne
rect 16191 9983 16613 10013
tri 16613 9983 16643 10013 sw
tri 16711 9983 16741 10013 ne
rect 16741 9983 17163 10013
tri 17163 9983 17193 10013 sw
tri 17261 9983 17291 10013 ne
rect 17291 9983 17713 10013
tri 17713 9983 17743 10013 sw
tri 17811 9983 17841 10013 ne
rect 17841 9983 18263 10013
tri 18263 9983 18293 10013 sw
tri 18361 9983 18391 10013 ne
rect 18391 9983 18813 10013
tri 18813 9983 18843 10013 sw
tri 18911 9983 18941 10013 ne
rect 18941 9983 19363 10013
tri 19363 9983 19393 10013 sw
tri 19461 9983 19491 10013 ne
rect 19491 9983 20300 10013
rect -2000 9885 143 9983
tri 143 9885 241 9983 sw
tri 241 9885 339 9983 ne
rect 339 9885 693 9983
tri 693 9885 791 9983 sw
tri 791 9885 889 9983 ne
rect 889 9885 1243 9983
tri 1243 9885 1341 9983 sw
tri 1341 9885 1439 9983 ne
rect 1439 9885 1793 9983
tri 1793 9885 1891 9983 sw
tri 1891 9885 1989 9983 ne
rect 1989 9885 2343 9983
tri 2343 9885 2441 9983 sw
tri 2441 9885 2539 9983 ne
rect 2539 9885 2893 9983
tri 2893 9885 2991 9983 sw
tri 2991 9885 3089 9983 ne
rect 3089 9885 3443 9983
tri 3443 9885 3541 9983 sw
tri 3541 9885 3639 9983 ne
rect 3639 9885 3993 9983
tri 3993 9885 4091 9983 sw
tri 4091 9885 4189 9983 ne
rect 4189 9885 4543 9983
tri 4543 9885 4641 9983 sw
tri 4641 9885 4739 9983 ne
rect 4739 9885 5093 9983
tri 5093 9885 5191 9983 sw
tri 5191 9885 5289 9983 ne
rect 5289 9885 5643 9983
tri 5643 9885 5741 9983 sw
tri 5741 9885 5839 9983 ne
rect 5839 9885 6193 9983
tri 6193 9885 6291 9983 sw
tri 6291 9885 6389 9983 ne
rect 6389 9885 6743 9983
tri 6743 9885 6841 9983 sw
tri 6841 9885 6939 9983 ne
rect 6939 9885 7293 9983
tri 7293 9885 7391 9983 sw
tri 7391 9885 7489 9983 ne
rect 7489 9885 7843 9983
tri 7843 9885 7941 9983 sw
tri 7941 9885 8039 9983 ne
rect 8039 9885 8393 9983
tri 8393 9885 8491 9983 sw
tri 8491 9885 8589 9983 ne
rect 8589 9885 8943 9983
tri 8943 9885 9041 9983 sw
tri 9041 9885 9139 9983 ne
rect 9139 9885 9493 9983
tri 9493 9885 9591 9983 sw
tri 9591 9885 9689 9983 ne
rect 9689 9885 10043 9983
tri 10043 9885 10141 9983 sw
tri 10141 9885 10239 9983 ne
rect 10239 9885 10593 9983
tri 10593 9885 10691 9983 sw
tri 10691 9885 10789 9983 ne
rect 10789 9885 11143 9983
tri 11143 9885 11241 9983 sw
tri 11241 9885 11339 9983 ne
rect 11339 9885 11693 9983
tri 11693 9885 11791 9983 sw
tri 11791 9885 11889 9983 ne
rect 11889 9885 12243 9983
tri 12243 9885 12341 9983 sw
tri 12341 9885 12439 9983 ne
rect 12439 9885 12793 9983
tri 12793 9885 12891 9983 sw
tri 12891 9885 12989 9983 ne
rect 12989 9885 13343 9983
tri 13343 9885 13441 9983 sw
tri 13441 9885 13539 9983 ne
rect 13539 9885 13893 9983
tri 13893 9885 13991 9983 sw
tri 13991 9885 14089 9983 ne
rect 14089 9885 14443 9983
tri 14443 9885 14541 9983 sw
tri 14541 9885 14639 9983 ne
rect 14639 9885 14993 9983
tri 14993 9885 15091 9983 sw
tri 15091 9885 15189 9983 ne
rect 15189 9885 15543 9983
tri 15543 9885 15641 9983 sw
tri 15641 9885 15739 9983 ne
rect 15739 9885 16093 9983
tri 16093 9885 16191 9983 sw
tri 16191 9885 16289 9983 ne
rect 16289 9885 16643 9983
tri 16643 9885 16741 9983 sw
tri 16741 9885 16839 9983 ne
rect 16839 9885 17193 9983
tri 17193 9885 17291 9983 sw
tri 17291 9885 17389 9983 ne
rect 17389 9885 17743 9983
tri 17743 9885 17841 9983 sw
tri 17841 9885 17939 9983 ne
rect 17939 9885 18293 9983
tri 18293 9885 18391 9983 sw
tri 18391 9885 18489 9983 ne
rect 18489 9885 18843 9983
tri 18843 9885 18941 9983 sw
tri 18941 9885 19039 9983 ne
rect 19039 9885 19393 9983
tri 19393 9885 19491 9983 sw
tri 19491 9885 19589 9983 ne
rect 19589 9885 20300 9983
rect -2000 9787 241 9885
tri 241 9787 339 9885 sw
tri 339 9787 437 9885 ne
rect 437 9787 791 9885
tri 791 9787 889 9885 sw
tri 889 9787 987 9885 ne
rect 987 9787 1341 9885
tri 1341 9787 1439 9885 sw
tri 1439 9787 1537 9885 ne
rect 1537 9787 1891 9885
tri 1891 9787 1989 9885 sw
tri 1989 9787 2087 9885 ne
rect 2087 9787 2441 9885
tri 2441 9787 2539 9885 sw
tri 2539 9787 2637 9885 ne
rect 2637 9787 2991 9885
tri 2991 9787 3089 9885 sw
tri 3089 9787 3187 9885 ne
rect 3187 9787 3541 9885
tri 3541 9787 3639 9885 sw
tri 3639 9787 3737 9885 ne
rect 3737 9787 4091 9885
tri 4091 9787 4189 9885 sw
tri 4189 9787 4287 9885 ne
rect 4287 9787 4641 9885
tri 4641 9787 4739 9885 sw
tri 4739 9787 4837 9885 ne
rect 4837 9787 5191 9885
tri 5191 9787 5289 9885 sw
tri 5289 9787 5387 9885 ne
rect 5387 9787 5741 9885
tri 5741 9787 5839 9885 sw
tri 5839 9787 5937 9885 ne
rect 5937 9787 6291 9885
tri 6291 9787 6389 9885 sw
tri 6389 9787 6487 9885 ne
rect 6487 9787 6841 9885
tri 6841 9787 6939 9885 sw
tri 6939 9787 7037 9885 ne
rect 7037 9787 7391 9885
tri 7391 9787 7489 9885 sw
tri 7489 9787 7587 9885 ne
rect 7587 9787 7941 9885
tri 7941 9787 8039 9885 sw
tri 8039 9787 8137 9885 ne
rect 8137 9787 8491 9885
tri 8491 9787 8589 9885 sw
tri 8589 9787 8687 9885 ne
rect 8687 9787 9041 9885
tri 9041 9787 9139 9885 sw
tri 9139 9787 9237 9885 ne
rect 9237 9787 9591 9885
tri 9591 9787 9689 9885 sw
tri 9689 9787 9787 9885 ne
rect 9787 9787 10141 9885
tri 10141 9787 10239 9885 sw
tri 10239 9787 10337 9885 ne
rect 10337 9787 10691 9885
tri 10691 9787 10789 9885 sw
tri 10789 9787 10887 9885 ne
rect 10887 9787 11241 9885
tri 11241 9787 11339 9885 sw
tri 11339 9787 11437 9885 ne
rect 11437 9787 11791 9885
tri 11791 9787 11889 9885 sw
tri 11889 9787 11987 9885 ne
rect 11987 9787 12341 9885
tri 12341 9787 12439 9885 sw
tri 12439 9787 12537 9885 ne
rect 12537 9787 12891 9885
tri 12891 9787 12989 9885 sw
tri 12989 9787 13087 9885 ne
rect 13087 9787 13441 9885
tri 13441 9787 13539 9885 sw
tri 13539 9787 13637 9885 ne
rect 13637 9787 13991 9885
tri 13991 9787 14089 9885 sw
tri 14089 9787 14187 9885 ne
rect 14187 9787 14541 9885
tri 14541 9787 14639 9885 sw
tri 14639 9787 14737 9885 ne
rect 14737 9787 15091 9885
tri 15091 9787 15189 9885 sw
tri 15189 9787 15287 9885 ne
rect 15287 9787 15641 9885
tri 15641 9787 15739 9885 sw
tri 15739 9787 15837 9885 ne
rect 15837 9787 16191 9885
tri 16191 9787 16289 9885 sw
tri 16289 9787 16387 9885 ne
rect 16387 9787 16741 9885
tri 16741 9787 16839 9885 sw
tri 16839 9787 16937 9885 ne
rect 16937 9787 17291 9885
tri 17291 9787 17389 9885 sw
tri 17389 9787 17487 9885 ne
rect 17487 9787 17841 9885
tri 17841 9787 17939 9885 sw
tri 17939 9787 18037 9885 ne
rect 18037 9787 18391 9885
tri 18391 9787 18489 9885 sw
tri 18489 9787 18587 9885 ne
rect 18587 9787 18941 9885
tri 18941 9787 19039 9885 sw
tri 19039 9787 19137 9885 ne
rect 19137 9787 19491 9885
tri 19491 9787 19589 9885 sw
tri 19589 9787 19687 9885 ne
rect 19687 9787 20300 9885
rect -2000 9689 339 9787
tri 339 9689 437 9787 sw
tri 437 9689 535 9787 ne
rect 535 9689 889 9787
tri 889 9689 987 9787 sw
tri 987 9689 1085 9787 ne
rect 1085 9689 1439 9787
tri 1439 9689 1537 9787 sw
tri 1537 9689 1635 9787 ne
rect 1635 9689 1989 9787
tri 1989 9689 2087 9787 sw
tri 2087 9689 2185 9787 ne
rect 2185 9689 2539 9787
tri 2539 9689 2637 9787 sw
tri 2637 9689 2735 9787 ne
rect 2735 9689 3089 9787
tri 3089 9689 3187 9787 sw
tri 3187 9689 3285 9787 ne
rect 3285 9689 3639 9787
tri 3639 9689 3737 9787 sw
tri 3737 9689 3835 9787 ne
rect 3835 9689 4189 9787
tri 4189 9689 4287 9787 sw
tri 4287 9689 4385 9787 ne
rect 4385 9689 4739 9787
tri 4739 9689 4837 9787 sw
tri 4837 9689 4935 9787 ne
rect 4935 9689 5289 9787
tri 5289 9689 5387 9787 sw
tri 5387 9689 5485 9787 ne
rect 5485 9689 5839 9787
tri 5839 9689 5937 9787 sw
tri 5937 9689 6035 9787 ne
rect 6035 9689 6389 9787
tri 6389 9689 6487 9787 sw
tri 6487 9689 6585 9787 ne
rect 6585 9689 6939 9787
tri 6939 9689 7037 9787 sw
tri 7037 9689 7135 9787 ne
rect 7135 9689 7489 9787
tri 7489 9689 7587 9787 sw
tri 7587 9689 7685 9787 ne
rect 7685 9689 8039 9787
tri 8039 9689 8137 9787 sw
tri 8137 9689 8235 9787 ne
rect 8235 9689 8589 9787
tri 8589 9689 8687 9787 sw
tri 8687 9689 8785 9787 ne
rect 8785 9689 9139 9787
tri 9139 9689 9237 9787 sw
tri 9237 9689 9335 9787 ne
rect 9335 9689 9689 9787
tri 9689 9689 9787 9787 sw
tri 9787 9689 9885 9787 ne
rect 9885 9689 10239 9787
tri 10239 9689 10337 9787 sw
tri 10337 9689 10435 9787 ne
rect 10435 9689 10789 9787
tri 10789 9689 10887 9787 sw
tri 10887 9689 10985 9787 ne
rect 10985 9689 11339 9787
tri 11339 9689 11437 9787 sw
tri 11437 9689 11535 9787 ne
rect 11535 9689 11889 9787
tri 11889 9689 11987 9787 sw
tri 11987 9689 12085 9787 ne
rect 12085 9689 12439 9787
tri 12439 9689 12537 9787 sw
tri 12537 9689 12635 9787 ne
rect 12635 9689 12989 9787
tri 12989 9689 13087 9787 sw
tri 13087 9689 13185 9787 ne
rect 13185 9689 13539 9787
tri 13539 9689 13637 9787 sw
tri 13637 9689 13735 9787 ne
rect 13735 9689 14089 9787
tri 14089 9689 14187 9787 sw
tri 14187 9689 14285 9787 ne
rect 14285 9689 14639 9787
tri 14639 9689 14737 9787 sw
tri 14737 9689 14835 9787 ne
rect 14835 9689 15189 9787
tri 15189 9689 15287 9787 sw
tri 15287 9689 15385 9787 ne
rect 15385 9689 15739 9787
tri 15739 9689 15837 9787 sw
tri 15837 9689 15935 9787 ne
rect 15935 9689 16289 9787
tri 16289 9689 16387 9787 sw
tri 16387 9689 16485 9787 ne
rect 16485 9689 16839 9787
tri 16839 9689 16937 9787 sw
tri 16937 9689 17035 9787 ne
rect 17035 9689 17389 9787
tri 17389 9689 17487 9787 sw
tri 17487 9689 17585 9787 ne
rect 17585 9689 17939 9787
tri 17939 9689 18037 9787 sw
tri 18037 9689 18135 9787 ne
rect 18135 9689 18489 9787
tri 18489 9689 18587 9787 sw
tri 18587 9689 18685 9787 ne
rect 18685 9689 19039 9787
tri 19039 9689 19137 9787 sw
tri 19137 9689 19235 9787 ne
rect 19235 9689 19589 9787
tri 19589 9689 19687 9787 sw
rect 20800 9689 21800 10337
rect -2000 9685 437 9689
rect -2000 9565 215 9685
rect 335 9591 437 9685
tri 437 9591 535 9689 sw
tri 535 9591 633 9689 ne
rect 633 9685 987 9689
rect 633 9591 765 9685
rect 335 9565 535 9591
rect -2000 9561 535 9565
rect -2000 8913 -1000 9561
tri 113 9463 211 9561 ne
rect 211 9513 535 9561
tri 535 9513 613 9591 sw
tri 633 9513 711 9591 ne
rect 711 9565 765 9591
rect 885 9591 987 9685
tri 987 9591 1085 9689 sw
tri 1085 9591 1183 9689 ne
rect 1183 9685 1537 9689
rect 1183 9591 1315 9685
rect 885 9565 1085 9591
rect 711 9513 1085 9565
tri 1085 9513 1163 9591 sw
tri 1183 9513 1261 9591 ne
rect 1261 9565 1315 9591
rect 1435 9591 1537 9685
tri 1537 9591 1635 9689 sw
tri 1635 9591 1733 9689 ne
rect 1733 9685 2087 9689
rect 1733 9591 1865 9685
rect 1435 9565 1635 9591
rect 1261 9513 1635 9565
tri 1635 9513 1713 9591 sw
tri 1733 9513 1811 9591 ne
rect 1811 9565 1865 9591
rect 1985 9591 2087 9685
tri 2087 9591 2185 9689 sw
tri 2185 9591 2283 9689 ne
rect 2283 9685 2637 9689
rect 2283 9591 2415 9685
rect 1985 9565 2185 9591
rect 1811 9513 2185 9565
tri 2185 9513 2263 9591 sw
tri 2283 9513 2361 9591 ne
rect 2361 9565 2415 9591
rect 2535 9591 2637 9685
tri 2637 9591 2735 9689 sw
tri 2735 9591 2833 9689 ne
rect 2833 9685 3187 9689
rect 2833 9591 2965 9685
rect 2535 9565 2735 9591
rect 2361 9513 2735 9565
tri 2735 9513 2813 9591 sw
tri 2833 9513 2911 9591 ne
rect 2911 9565 2965 9591
rect 3085 9591 3187 9685
tri 3187 9591 3285 9689 sw
tri 3285 9591 3383 9689 ne
rect 3383 9685 3737 9689
rect 3383 9591 3515 9685
rect 3085 9565 3285 9591
rect 2911 9513 3285 9565
tri 3285 9513 3363 9591 sw
tri 3383 9513 3461 9591 ne
rect 3461 9565 3515 9591
rect 3635 9591 3737 9685
tri 3737 9591 3835 9689 sw
tri 3835 9591 3933 9689 ne
rect 3933 9685 4287 9689
rect 3933 9591 4065 9685
rect 3635 9565 3835 9591
rect 3461 9513 3835 9565
tri 3835 9513 3913 9591 sw
tri 3933 9513 4011 9591 ne
rect 4011 9565 4065 9591
rect 4185 9591 4287 9685
tri 4287 9591 4385 9689 sw
tri 4385 9591 4483 9689 ne
rect 4483 9685 4837 9689
rect 4483 9591 4615 9685
rect 4185 9565 4385 9591
rect 4011 9513 4385 9565
tri 4385 9513 4463 9591 sw
tri 4483 9513 4561 9591 ne
rect 4561 9565 4615 9591
rect 4735 9591 4837 9685
tri 4837 9591 4935 9689 sw
tri 4935 9591 5033 9689 ne
rect 5033 9685 5387 9689
rect 5033 9591 5165 9685
rect 4735 9565 4935 9591
rect 4561 9513 4935 9565
tri 4935 9513 5013 9591 sw
tri 5033 9513 5111 9591 ne
rect 5111 9565 5165 9591
rect 5285 9591 5387 9685
tri 5387 9591 5485 9689 sw
tri 5485 9591 5583 9689 ne
rect 5583 9685 5937 9689
rect 5583 9591 5715 9685
rect 5285 9565 5485 9591
rect 5111 9513 5485 9565
tri 5485 9513 5563 9591 sw
tri 5583 9513 5661 9591 ne
rect 5661 9565 5715 9591
rect 5835 9591 5937 9685
tri 5937 9591 6035 9689 sw
tri 6035 9591 6133 9689 ne
rect 6133 9685 6487 9689
rect 6133 9591 6265 9685
rect 5835 9565 6035 9591
rect 5661 9513 6035 9565
tri 6035 9513 6113 9591 sw
tri 6133 9513 6211 9591 ne
rect 6211 9565 6265 9591
rect 6385 9591 6487 9685
tri 6487 9591 6585 9689 sw
tri 6585 9591 6683 9689 ne
rect 6683 9685 7037 9689
rect 6683 9591 6815 9685
rect 6385 9565 6585 9591
rect 6211 9513 6585 9565
tri 6585 9513 6663 9591 sw
tri 6683 9513 6761 9591 ne
rect 6761 9565 6815 9591
rect 6935 9591 7037 9685
tri 7037 9591 7135 9689 sw
tri 7135 9591 7233 9689 ne
rect 7233 9685 7587 9689
rect 7233 9591 7365 9685
rect 6935 9565 7135 9591
rect 6761 9513 7135 9565
tri 7135 9513 7213 9591 sw
tri 7233 9513 7311 9591 ne
rect 7311 9565 7365 9591
rect 7485 9591 7587 9685
tri 7587 9591 7685 9689 sw
tri 7685 9591 7783 9689 ne
rect 7783 9685 8137 9689
rect 7783 9591 7915 9685
rect 7485 9565 7685 9591
rect 7311 9513 7685 9565
tri 7685 9513 7763 9591 sw
tri 7783 9513 7861 9591 ne
rect 7861 9565 7915 9591
rect 8035 9591 8137 9685
tri 8137 9591 8235 9689 sw
tri 8235 9591 8333 9689 ne
rect 8333 9685 8687 9689
rect 8333 9591 8465 9685
rect 8035 9565 8235 9591
rect 7861 9513 8235 9565
tri 8235 9513 8313 9591 sw
tri 8333 9513 8411 9591 ne
rect 8411 9565 8465 9591
rect 8585 9591 8687 9685
tri 8687 9591 8785 9689 sw
tri 8785 9591 8883 9689 ne
rect 8883 9685 9237 9689
rect 8883 9591 9015 9685
rect 8585 9565 8785 9591
rect 8411 9513 8785 9565
tri 8785 9513 8863 9591 sw
tri 8883 9513 8961 9591 ne
rect 8961 9565 9015 9591
rect 9135 9591 9237 9685
tri 9237 9591 9335 9689 sw
tri 9335 9591 9433 9689 ne
rect 9433 9685 9787 9689
rect 9433 9591 9565 9685
rect 9135 9565 9335 9591
rect 8961 9513 9335 9565
tri 9335 9513 9413 9591 sw
tri 9433 9513 9511 9591 ne
rect 9511 9565 9565 9591
rect 9685 9591 9787 9685
tri 9787 9591 9885 9689 sw
tri 9885 9591 9983 9689 ne
rect 9983 9685 10337 9689
rect 9983 9591 10115 9685
rect 9685 9565 9885 9591
rect 9511 9513 9885 9565
tri 9885 9513 9963 9591 sw
tri 9983 9513 10061 9591 ne
rect 10061 9565 10115 9591
rect 10235 9591 10337 9685
tri 10337 9591 10435 9689 sw
tri 10435 9591 10533 9689 ne
rect 10533 9685 10887 9689
rect 10533 9591 10665 9685
rect 10235 9565 10435 9591
rect 10061 9513 10435 9565
tri 10435 9513 10513 9591 sw
tri 10533 9513 10611 9591 ne
rect 10611 9565 10665 9591
rect 10785 9591 10887 9685
tri 10887 9591 10985 9689 sw
tri 10985 9591 11083 9689 ne
rect 11083 9685 11437 9689
rect 11083 9591 11215 9685
rect 10785 9565 10985 9591
rect 10611 9513 10985 9565
tri 10985 9513 11063 9591 sw
tri 11083 9513 11161 9591 ne
rect 11161 9565 11215 9591
rect 11335 9591 11437 9685
tri 11437 9591 11535 9689 sw
tri 11535 9591 11633 9689 ne
rect 11633 9685 11987 9689
rect 11633 9591 11765 9685
rect 11335 9565 11535 9591
rect 11161 9513 11535 9565
tri 11535 9513 11613 9591 sw
tri 11633 9513 11711 9591 ne
rect 11711 9565 11765 9591
rect 11885 9591 11987 9685
tri 11987 9591 12085 9689 sw
tri 12085 9591 12183 9689 ne
rect 12183 9685 12537 9689
rect 12183 9591 12315 9685
rect 11885 9565 12085 9591
rect 11711 9513 12085 9565
tri 12085 9513 12163 9591 sw
tri 12183 9513 12261 9591 ne
rect 12261 9565 12315 9591
rect 12435 9591 12537 9685
tri 12537 9591 12635 9689 sw
tri 12635 9591 12733 9689 ne
rect 12733 9685 13087 9689
rect 12733 9591 12865 9685
rect 12435 9565 12635 9591
rect 12261 9513 12635 9565
tri 12635 9513 12713 9591 sw
tri 12733 9513 12811 9591 ne
rect 12811 9565 12865 9591
rect 12985 9591 13087 9685
tri 13087 9591 13185 9689 sw
tri 13185 9591 13283 9689 ne
rect 13283 9685 13637 9689
rect 13283 9591 13415 9685
rect 12985 9565 13185 9591
rect 12811 9513 13185 9565
tri 13185 9513 13263 9591 sw
tri 13283 9513 13361 9591 ne
rect 13361 9565 13415 9591
rect 13535 9591 13637 9685
tri 13637 9591 13735 9689 sw
tri 13735 9591 13833 9689 ne
rect 13833 9685 14187 9689
rect 13833 9591 13965 9685
rect 13535 9565 13735 9591
rect 13361 9513 13735 9565
tri 13735 9513 13813 9591 sw
tri 13833 9513 13911 9591 ne
rect 13911 9565 13965 9591
rect 14085 9591 14187 9685
tri 14187 9591 14285 9689 sw
tri 14285 9591 14383 9689 ne
rect 14383 9685 14737 9689
rect 14383 9591 14515 9685
rect 14085 9565 14285 9591
rect 13911 9513 14285 9565
tri 14285 9513 14363 9591 sw
tri 14383 9513 14461 9591 ne
rect 14461 9565 14515 9591
rect 14635 9591 14737 9685
tri 14737 9591 14835 9689 sw
tri 14835 9591 14933 9689 ne
rect 14933 9685 15287 9689
rect 14933 9591 15065 9685
rect 14635 9565 14835 9591
rect 14461 9513 14835 9565
tri 14835 9513 14913 9591 sw
tri 14933 9513 15011 9591 ne
rect 15011 9565 15065 9591
rect 15185 9591 15287 9685
tri 15287 9591 15385 9689 sw
tri 15385 9591 15483 9689 ne
rect 15483 9685 15837 9689
rect 15483 9591 15615 9685
rect 15185 9565 15385 9591
rect 15011 9513 15385 9565
tri 15385 9513 15463 9591 sw
tri 15483 9513 15561 9591 ne
rect 15561 9565 15615 9591
rect 15735 9591 15837 9685
tri 15837 9591 15935 9689 sw
tri 15935 9591 16033 9689 ne
rect 16033 9685 16387 9689
rect 16033 9591 16165 9685
rect 15735 9565 15935 9591
rect 15561 9513 15935 9565
tri 15935 9513 16013 9591 sw
tri 16033 9513 16111 9591 ne
rect 16111 9565 16165 9591
rect 16285 9591 16387 9685
tri 16387 9591 16485 9689 sw
tri 16485 9591 16583 9689 ne
rect 16583 9685 16937 9689
rect 16583 9591 16715 9685
rect 16285 9565 16485 9591
rect 16111 9513 16485 9565
tri 16485 9513 16563 9591 sw
tri 16583 9513 16661 9591 ne
rect 16661 9565 16715 9591
rect 16835 9591 16937 9685
tri 16937 9591 17035 9689 sw
tri 17035 9591 17133 9689 ne
rect 17133 9685 17487 9689
rect 17133 9591 17265 9685
rect 16835 9565 17035 9591
rect 16661 9513 17035 9565
tri 17035 9513 17113 9591 sw
tri 17133 9513 17211 9591 ne
rect 17211 9565 17265 9591
rect 17385 9591 17487 9685
tri 17487 9591 17585 9689 sw
tri 17585 9591 17683 9689 ne
rect 17683 9685 18037 9689
rect 17683 9591 17815 9685
rect 17385 9565 17585 9591
rect 17211 9513 17585 9565
tri 17585 9513 17663 9591 sw
tri 17683 9513 17761 9591 ne
rect 17761 9565 17815 9591
rect 17935 9591 18037 9685
tri 18037 9591 18135 9689 sw
tri 18135 9591 18233 9689 ne
rect 18233 9685 18587 9689
rect 18233 9591 18365 9685
rect 17935 9565 18135 9591
rect 17761 9513 18135 9565
tri 18135 9513 18213 9591 sw
tri 18233 9513 18311 9591 ne
rect 18311 9565 18365 9591
rect 18485 9591 18587 9685
tri 18587 9591 18685 9689 sw
tri 18685 9591 18783 9689 ne
rect 18783 9685 19137 9689
rect 18783 9591 18915 9685
rect 18485 9565 18685 9591
rect 18311 9513 18685 9565
tri 18685 9513 18763 9591 sw
tri 18783 9513 18861 9591 ne
rect 18861 9565 18915 9591
rect 19035 9591 19137 9685
tri 19137 9591 19235 9689 sw
tri 19235 9591 19333 9689 ne
rect 19333 9685 21800 9689
rect 19333 9591 19465 9685
rect 19035 9565 19235 9591
rect 18861 9513 19235 9565
tri 19235 9513 19313 9591 sw
tri 19333 9513 19411 9591 ne
rect 19411 9565 19465 9591
rect 19585 9565 21800 9685
rect 19411 9513 21800 9565
rect 211 9463 613 9513
rect -500 9413 113 9463
tri 113 9413 163 9463 sw
tri 211 9413 261 9463 ne
rect 261 9433 613 9463
tri 613 9433 693 9513 sw
tri 711 9433 791 9513 ne
rect 791 9433 1163 9513
tri 1163 9433 1243 9513 sw
tri 1261 9433 1341 9513 ne
rect 1341 9433 1713 9513
tri 1713 9433 1793 9513 sw
tri 1811 9433 1891 9513 ne
rect 1891 9433 2263 9513
tri 2263 9433 2343 9513 sw
tri 2361 9433 2441 9513 ne
rect 2441 9433 2813 9513
tri 2813 9433 2893 9513 sw
tri 2911 9433 2991 9513 ne
rect 2991 9433 3363 9513
tri 3363 9433 3443 9513 sw
tri 3461 9433 3541 9513 ne
rect 3541 9433 3913 9513
tri 3913 9433 3993 9513 sw
tri 4011 9433 4091 9513 ne
rect 4091 9433 4463 9513
tri 4463 9433 4543 9513 sw
tri 4561 9433 4641 9513 ne
rect 4641 9433 5013 9513
tri 5013 9433 5093 9513 sw
tri 5111 9433 5191 9513 ne
rect 5191 9433 5563 9513
tri 5563 9433 5643 9513 sw
tri 5661 9433 5741 9513 ne
rect 5741 9433 6113 9513
tri 6113 9433 6193 9513 sw
tri 6211 9433 6291 9513 ne
rect 6291 9433 6663 9513
tri 6663 9433 6743 9513 sw
tri 6761 9433 6841 9513 ne
rect 6841 9433 7213 9513
tri 7213 9433 7293 9513 sw
tri 7311 9433 7391 9513 ne
rect 7391 9433 7763 9513
tri 7763 9433 7843 9513 sw
tri 7861 9433 7941 9513 ne
rect 7941 9433 8313 9513
tri 8313 9433 8393 9513 sw
tri 8411 9433 8491 9513 ne
rect 8491 9433 8863 9513
tri 8863 9433 8943 9513 sw
tri 8961 9433 9041 9513 ne
rect 9041 9433 9413 9513
tri 9413 9433 9493 9513 sw
tri 9511 9433 9591 9513 ne
rect 9591 9433 9963 9513
tri 9963 9433 10043 9513 sw
tri 10061 9433 10141 9513 ne
rect 10141 9433 10513 9513
tri 10513 9433 10593 9513 sw
tri 10611 9433 10691 9513 ne
rect 10691 9433 11063 9513
tri 11063 9433 11143 9513 sw
tri 11161 9433 11241 9513 ne
rect 11241 9433 11613 9513
tri 11613 9433 11693 9513 sw
tri 11711 9433 11791 9513 ne
rect 11791 9433 12163 9513
tri 12163 9433 12243 9513 sw
tri 12261 9433 12341 9513 ne
rect 12341 9433 12713 9513
tri 12713 9433 12793 9513 sw
tri 12811 9433 12891 9513 ne
rect 12891 9433 13263 9513
tri 13263 9433 13343 9513 sw
tri 13361 9433 13441 9513 ne
rect 13441 9433 13813 9513
tri 13813 9433 13893 9513 sw
tri 13911 9433 13991 9513 ne
rect 13991 9433 14363 9513
tri 14363 9433 14443 9513 sw
tri 14461 9433 14541 9513 ne
rect 14541 9433 14913 9513
tri 14913 9433 14993 9513 sw
tri 15011 9433 15091 9513 ne
rect 15091 9433 15463 9513
tri 15463 9433 15543 9513 sw
tri 15561 9433 15641 9513 ne
rect 15641 9433 16013 9513
tri 16013 9433 16093 9513 sw
tri 16111 9433 16191 9513 ne
rect 16191 9433 16563 9513
tri 16563 9433 16643 9513 sw
tri 16661 9433 16741 9513 ne
rect 16741 9433 17113 9513
tri 17113 9433 17193 9513 sw
tri 17211 9433 17291 9513 ne
rect 17291 9433 17663 9513
tri 17663 9433 17743 9513 sw
tri 17761 9433 17841 9513 ne
rect 17841 9433 18213 9513
tri 18213 9433 18293 9513 sw
tri 18311 9433 18391 9513 ne
rect 18391 9433 18763 9513
tri 18763 9433 18843 9513 sw
tri 18861 9433 18941 9513 ne
rect 18941 9433 19313 9513
tri 19313 9433 19393 9513 sw
tri 19411 9433 19491 9513 ne
rect 19491 9433 20100 9513
rect 261 9413 693 9433
rect -500 9335 163 9413
tri 163 9335 241 9413 sw
tri 261 9335 339 9413 ne
rect 339 9335 693 9413
tri 693 9335 791 9433 sw
tri 791 9335 889 9433 ne
rect 889 9335 1243 9433
tri 1243 9335 1341 9433 sw
tri 1341 9335 1439 9433 ne
rect 1439 9335 1793 9433
tri 1793 9335 1891 9433 sw
tri 1891 9335 1989 9433 ne
rect 1989 9335 2343 9433
tri 2343 9335 2441 9433 sw
tri 2441 9335 2539 9433 ne
rect 2539 9335 2893 9433
tri 2893 9335 2991 9433 sw
tri 2991 9335 3089 9433 ne
rect 3089 9335 3443 9433
tri 3443 9335 3541 9433 sw
tri 3541 9335 3639 9433 ne
rect 3639 9335 3993 9433
tri 3993 9335 4091 9433 sw
tri 4091 9335 4189 9433 ne
rect 4189 9335 4543 9433
tri 4543 9335 4641 9433 sw
tri 4641 9335 4739 9433 ne
rect 4739 9335 5093 9433
tri 5093 9335 5191 9433 sw
tri 5191 9335 5289 9433 ne
rect 5289 9335 5643 9433
tri 5643 9335 5741 9433 sw
tri 5741 9335 5839 9433 ne
rect 5839 9335 6193 9433
tri 6193 9335 6291 9433 sw
tri 6291 9335 6389 9433 ne
rect 6389 9335 6743 9433
tri 6743 9335 6841 9433 sw
tri 6841 9335 6939 9433 ne
rect 6939 9335 7293 9433
tri 7293 9335 7391 9433 sw
tri 7391 9335 7489 9433 ne
rect 7489 9335 7843 9433
tri 7843 9335 7941 9433 sw
tri 7941 9335 8039 9433 ne
rect 8039 9335 8393 9433
tri 8393 9335 8491 9433 sw
tri 8491 9335 8589 9433 ne
rect 8589 9335 8943 9433
tri 8943 9335 9041 9433 sw
tri 9041 9335 9139 9433 ne
rect 9139 9335 9493 9433
tri 9493 9335 9591 9433 sw
tri 9591 9335 9689 9433 ne
rect 9689 9335 10043 9433
tri 10043 9335 10141 9433 sw
tri 10141 9335 10239 9433 ne
rect 10239 9335 10593 9433
tri 10593 9335 10691 9433 sw
tri 10691 9335 10789 9433 ne
rect 10789 9335 11143 9433
tri 11143 9335 11241 9433 sw
tri 11241 9335 11339 9433 ne
rect 11339 9335 11693 9433
tri 11693 9335 11791 9433 sw
tri 11791 9335 11889 9433 ne
rect 11889 9335 12243 9433
tri 12243 9335 12341 9433 sw
tri 12341 9335 12439 9433 ne
rect 12439 9335 12793 9433
tri 12793 9335 12891 9433 sw
tri 12891 9335 12989 9433 ne
rect 12989 9335 13343 9433
tri 13343 9335 13441 9433 sw
tri 13441 9335 13539 9433 ne
rect 13539 9335 13893 9433
tri 13893 9335 13991 9433 sw
tri 13991 9335 14089 9433 ne
rect 14089 9335 14443 9433
tri 14443 9335 14541 9433 sw
tri 14541 9335 14639 9433 ne
rect 14639 9335 14993 9433
tri 14993 9335 15091 9433 sw
tri 15091 9335 15189 9433 ne
rect 15189 9335 15543 9433
tri 15543 9335 15641 9433 sw
tri 15641 9335 15739 9433 ne
rect 15739 9335 16093 9433
tri 16093 9335 16191 9433 sw
tri 16191 9335 16289 9433 ne
rect 16289 9335 16643 9433
tri 16643 9335 16741 9433 sw
tri 16741 9335 16839 9433 ne
rect 16839 9335 17193 9433
tri 17193 9335 17291 9433 sw
tri 17291 9335 17389 9433 ne
rect 17389 9335 17743 9433
tri 17743 9335 17841 9433 sw
tri 17841 9335 17939 9433 ne
rect 17939 9335 18293 9433
tri 18293 9335 18391 9433 sw
tri 18391 9335 18489 9433 ne
rect 18489 9335 18843 9433
tri 18843 9335 18941 9433 sw
tri 18941 9335 19039 9433 ne
rect 19039 9335 19393 9433
tri 19393 9335 19491 9433 sw
tri 19491 9335 19589 9433 ne
rect 19589 9413 20100 9433
rect 20200 9413 21800 9513
rect 19589 9335 21800 9413
rect -500 9287 241 9335
rect -500 9187 -400 9287
rect -300 9237 241 9287
tri 241 9237 339 9335 sw
tri 339 9237 437 9335 ne
rect 437 9237 791 9335
tri 791 9237 889 9335 sw
tri 889 9237 987 9335 ne
rect 987 9237 1341 9335
tri 1341 9237 1439 9335 sw
tri 1439 9237 1537 9335 ne
rect 1537 9237 1891 9335
tri 1891 9237 1989 9335 sw
tri 1989 9237 2087 9335 ne
rect 2087 9237 2441 9335
tri 2441 9237 2539 9335 sw
tri 2539 9237 2637 9335 ne
rect 2637 9237 2991 9335
tri 2991 9237 3089 9335 sw
tri 3089 9237 3187 9335 ne
rect 3187 9237 3541 9335
tri 3541 9237 3639 9335 sw
tri 3639 9237 3737 9335 ne
rect 3737 9237 4091 9335
tri 4091 9237 4189 9335 sw
tri 4189 9237 4287 9335 ne
rect 4287 9237 4641 9335
tri 4641 9237 4739 9335 sw
tri 4739 9237 4837 9335 ne
rect 4837 9237 5191 9335
tri 5191 9237 5289 9335 sw
tri 5289 9237 5387 9335 ne
rect 5387 9237 5741 9335
tri 5741 9237 5839 9335 sw
tri 5839 9237 5937 9335 ne
rect 5937 9237 6291 9335
tri 6291 9237 6389 9335 sw
tri 6389 9237 6487 9335 ne
rect 6487 9237 6841 9335
tri 6841 9237 6939 9335 sw
tri 6939 9237 7037 9335 ne
rect 7037 9237 7391 9335
tri 7391 9237 7489 9335 sw
tri 7489 9237 7587 9335 ne
rect 7587 9237 7941 9335
tri 7941 9237 8039 9335 sw
tri 8039 9237 8137 9335 ne
rect 8137 9237 8491 9335
tri 8491 9237 8589 9335 sw
tri 8589 9237 8687 9335 ne
rect 8687 9237 9041 9335
tri 9041 9237 9139 9335 sw
tri 9139 9237 9237 9335 ne
rect 9237 9237 9591 9335
tri 9591 9237 9689 9335 sw
tri 9689 9237 9787 9335 ne
rect 9787 9237 10141 9335
tri 10141 9237 10239 9335 sw
tri 10239 9237 10337 9335 ne
rect 10337 9237 10691 9335
tri 10691 9237 10789 9335 sw
tri 10789 9237 10887 9335 ne
rect 10887 9237 11241 9335
tri 11241 9237 11339 9335 sw
tri 11339 9237 11437 9335 ne
rect 11437 9237 11791 9335
tri 11791 9237 11889 9335 sw
tri 11889 9237 11987 9335 ne
rect 11987 9237 12341 9335
tri 12341 9237 12439 9335 sw
tri 12439 9237 12537 9335 ne
rect 12537 9237 12891 9335
tri 12891 9237 12989 9335 sw
tri 12989 9237 13087 9335 ne
rect 13087 9237 13441 9335
tri 13441 9237 13539 9335 sw
tri 13539 9237 13637 9335 ne
rect 13637 9237 13991 9335
tri 13991 9237 14089 9335 sw
tri 14089 9237 14187 9335 ne
rect 14187 9237 14541 9335
tri 14541 9237 14639 9335 sw
tri 14639 9237 14737 9335 ne
rect 14737 9237 15091 9335
tri 15091 9237 15189 9335 sw
tri 15189 9237 15287 9335 ne
rect 15287 9237 15641 9335
tri 15641 9237 15739 9335 sw
tri 15739 9237 15837 9335 ne
rect 15837 9237 16191 9335
tri 16191 9237 16289 9335 sw
tri 16289 9237 16387 9335 ne
rect 16387 9237 16741 9335
tri 16741 9237 16839 9335 sw
tri 16839 9237 16937 9335 ne
rect 16937 9237 17291 9335
tri 17291 9237 17389 9335 sw
tri 17389 9237 17487 9335 ne
rect 17487 9237 17841 9335
tri 17841 9237 17939 9335 sw
tri 17939 9237 18037 9335 ne
rect 18037 9237 18391 9335
tri 18391 9237 18489 9335 sw
tri 18489 9237 18587 9335 ne
rect 18587 9237 18941 9335
tri 18941 9237 19039 9335 sw
tri 19039 9237 19137 9335 ne
rect 19137 9237 19491 9335
tri 19491 9237 19589 9335 sw
tri 19589 9237 19687 9335 ne
rect 19687 9237 21800 9335
rect -300 9187 339 9237
rect -500 9139 339 9187
tri 339 9139 437 9237 sw
tri 437 9139 535 9237 ne
rect 535 9139 889 9237
tri 889 9139 987 9237 sw
tri 987 9139 1085 9237 ne
rect 1085 9139 1439 9237
tri 1439 9139 1537 9237 sw
tri 1537 9139 1635 9237 ne
rect 1635 9139 1989 9237
tri 1989 9139 2087 9237 sw
tri 2087 9139 2185 9237 ne
rect 2185 9139 2539 9237
tri 2539 9139 2637 9237 sw
tri 2637 9139 2735 9237 ne
rect 2735 9139 3089 9237
tri 3089 9139 3187 9237 sw
tri 3187 9139 3285 9237 ne
rect 3285 9139 3639 9237
tri 3639 9139 3737 9237 sw
tri 3737 9139 3835 9237 ne
rect 3835 9139 4189 9237
tri 4189 9139 4287 9237 sw
tri 4287 9139 4385 9237 ne
rect 4385 9139 4739 9237
tri 4739 9139 4837 9237 sw
tri 4837 9139 4935 9237 ne
rect 4935 9139 5289 9237
tri 5289 9139 5387 9237 sw
tri 5387 9139 5485 9237 ne
rect 5485 9139 5839 9237
tri 5839 9139 5937 9237 sw
tri 5937 9139 6035 9237 ne
rect 6035 9139 6389 9237
tri 6389 9139 6487 9237 sw
tri 6487 9139 6585 9237 ne
rect 6585 9139 6939 9237
tri 6939 9139 7037 9237 sw
tri 7037 9139 7135 9237 ne
rect 7135 9139 7489 9237
tri 7489 9139 7587 9237 sw
tri 7587 9139 7685 9237 ne
rect 7685 9139 8039 9237
tri 8039 9139 8137 9237 sw
tri 8137 9139 8235 9237 ne
rect 8235 9139 8589 9237
tri 8589 9139 8687 9237 sw
tri 8687 9139 8785 9237 ne
rect 8785 9139 9139 9237
tri 9139 9139 9237 9237 sw
tri 9237 9139 9335 9237 ne
rect 9335 9139 9689 9237
tri 9689 9139 9787 9237 sw
tri 9787 9139 9885 9237 ne
rect 9885 9139 10239 9237
tri 10239 9139 10337 9237 sw
tri 10337 9139 10435 9237 ne
rect 10435 9139 10789 9237
tri 10789 9139 10887 9237 sw
tri 10887 9139 10985 9237 ne
rect 10985 9139 11339 9237
tri 11339 9139 11437 9237 sw
tri 11437 9139 11535 9237 ne
rect 11535 9139 11889 9237
tri 11889 9139 11987 9237 sw
tri 11987 9139 12085 9237 ne
rect 12085 9139 12439 9237
tri 12439 9139 12537 9237 sw
tri 12537 9139 12635 9237 ne
rect 12635 9139 12989 9237
tri 12989 9139 13087 9237 sw
tri 13087 9139 13185 9237 ne
rect 13185 9139 13539 9237
tri 13539 9139 13637 9237 sw
tri 13637 9139 13735 9237 ne
rect 13735 9139 14089 9237
tri 14089 9139 14187 9237 sw
tri 14187 9139 14285 9237 ne
rect 14285 9139 14639 9237
tri 14639 9139 14737 9237 sw
tri 14737 9139 14835 9237 ne
rect 14835 9139 15189 9237
tri 15189 9139 15287 9237 sw
tri 15287 9139 15385 9237 ne
rect 15385 9139 15739 9237
tri 15739 9139 15837 9237 sw
tri 15837 9139 15935 9237 ne
rect 15935 9139 16289 9237
tri 16289 9139 16387 9237 sw
tri 16387 9139 16485 9237 ne
rect 16485 9139 16839 9237
tri 16839 9139 16937 9237 sw
tri 16937 9139 17035 9237 ne
rect 17035 9139 17389 9237
tri 17389 9139 17487 9237 sw
tri 17487 9139 17585 9237 ne
rect 17585 9139 17939 9237
tri 17939 9139 18037 9237 sw
tri 18037 9139 18135 9237 ne
rect 18135 9139 18489 9237
tri 18489 9139 18587 9237 sw
tri 18587 9139 18685 9237 ne
rect 18685 9139 19039 9237
tri 19039 9139 19137 9237 sw
tri 19137 9139 19235 9237 ne
rect 19235 9139 19589 9237
tri 19589 9139 19687 9237 sw
rect -500 9135 437 9139
rect -500 9015 215 9135
rect 335 9041 437 9135
tri 437 9041 535 9139 sw
tri 535 9041 633 9139 ne
rect 633 9135 987 9139
rect 633 9041 765 9135
rect 335 9015 535 9041
rect -500 9011 535 9015
tri 535 9011 565 9041 sw
tri 633 9011 663 9041 ne
rect 663 9015 765 9041
rect 885 9041 987 9135
tri 987 9041 1085 9139 sw
tri 1085 9041 1183 9139 ne
rect 1183 9135 1537 9139
rect 1183 9041 1315 9135
rect 885 9015 1085 9041
rect 663 9011 1085 9015
tri 1085 9011 1115 9041 sw
tri 1183 9011 1213 9041 ne
rect 1213 9015 1315 9041
rect 1435 9041 1537 9135
tri 1537 9041 1635 9139 sw
tri 1635 9041 1733 9139 ne
rect 1733 9135 2087 9139
rect 1733 9041 1865 9135
rect 1435 9015 1635 9041
rect 1213 9011 1635 9015
tri 1635 9011 1665 9041 sw
tri 1733 9011 1763 9041 ne
rect 1763 9015 1865 9041
rect 1985 9041 2087 9135
tri 2087 9041 2185 9139 sw
tri 2185 9041 2283 9139 ne
rect 2283 9135 2637 9139
rect 2283 9041 2415 9135
rect 1985 9015 2185 9041
rect 1763 9011 2185 9015
tri 2185 9011 2215 9041 sw
tri 2283 9011 2313 9041 ne
rect 2313 9015 2415 9041
rect 2535 9041 2637 9135
tri 2637 9041 2735 9139 sw
tri 2735 9041 2833 9139 ne
rect 2833 9135 3187 9139
rect 2833 9041 2965 9135
rect 2535 9015 2735 9041
rect 2313 9011 2735 9015
tri 2735 9011 2765 9041 sw
tri 2833 9011 2863 9041 ne
rect 2863 9015 2965 9041
rect 3085 9041 3187 9135
tri 3187 9041 3285 9139 sw
tri 3285 9041 3383 9139 ne
rect 3383 9135 3737 9139
rect 3383 9041 3515 9135
rect 3085 9015 3285 9041
rect 2863 9011 3285 9015
tri 3285 9011 3315 9041 sw
tri 3383 9011 3413 9041 ne
rect 3413 9015 3515 9041
rect 3635 9041 3737 9135
tri 3737 9041 3835 9139 sw
tri 3835 9041 3933 9139 ne
rect 3933 9135 4287 9139
rect 3933 9041 4065 9135
rect 3635 9015 3835 9041
rect 3413 9011 3835 9015
tri 3835 9011 3865 9041 sw
tri 3933 9011 3963 9041 ne
rect 3963 9015 4065 9041
rect 4185 9041 4287 9135
tri 4287 9041 4385 9139 sw
tri 4385 9041 4483 9139 ne
rect 4483 9135 4837 9139
rect 4483 9041 4615 9135
rect 4185 9015 4385 9041
rect 3963 9011 4385 9015
tri 4385 9011 4415 9041 sw
tri 4483 9011 4513 9041 ne
rect 4513 9015 4615 9041
rect 4735 9041 4837 9135
tri 4837 9041 4935 9139 sw
tri 4935 9041 5033 9139 ne
rect 5033 9135 5387 9139
rect 5033 9041 5165 9135
rect 4735 9015 4935 9041
rect 4513 9011 4935 9015
tri 4935 9011 4965 9041 sw
tri 5033 9011 5063 9041 ne
rect 5063 9015 5165 9041
rect 5285 9041 5387 9135
tri 5387 9041 5485 9139 sw
tri 5485 9041 5583 9139 ne
rect 5583 9135 5937 9139
rect 5583 9041 5715 9135
rect 5285 9015 5485 9041
rect 5063 9011 5485 9015
tri 5485 9011 5515 9041 sw
tri 5583 9011 5613 9041 ne
rect 5613 9015 5715 9041
rect 5835 9041 5937 9135
tri 5937 9041 6035 9139 sw
tri 6035 9041 6133 9139 ne
rect 6133 9135 6487 9139
rect 6133 9041 6265 9135
rect 5835 9015 6035 9041
rect 5613 9011 6035 9015
tri 6035 9011 6065 9041 sw
tri 6133 9011 6163 9041 ne
rect 6163 9015 6265 9041
rect 6385 9041 6487 9135
tri 6487 9041 6585 9139 sw
tri 6585 9041 6683 9139 ne
rect 6683 9135 7037 9139
rect 6683 9041 6815 9135
rect 6385 9015 6585 9041
rect 6163 9011 6585 9015
tri 6585 9011 6615 9041 sw
tri 6683 9011 6713 9041 ne
rect 6713 9015 6815 9041
rect 6935 9041 7037 9135
tri 7037 9041 7135 9139 sw
tri 7135 9041 7233 9139 ne
rect 7233 9135 7587 9139
rect 7233 9041 7365 9135
rect 6935 9015 7135 9041
rect 6713 9011 7135 9015
tri 7135 9011 7165 9041 sw
tri 7233 9011 7263 9041 ne
rect 7263 9015 7365 9041
rect 7485 9041 7587 9135
tri 7587 9041 7685 9139 sw
tri 7685 9041 7783 9139 ne
rect 7783 9135 8137 9139
rect 7783 9041 7915 9135
rect 7485 9015 7685 9041
rect 7263 9011 7685 9015
tri 7685 9011 7715 9041 sw
tri 7783 9011 7813 9041 ne
rect 7813 9015 7915 9041
rect 8035 9041 8137 9135
tri 8137 9041 8235 9139 sw
tri 8235 9041 8333 9139 ne
rect 8333 9135 8687 9139
rect 8333 9041 8465 9135
rect 8035 9015 8235 9041
rect 7813 9011 8235 9015
tri 8235 9011 8265 9041 sw
tri 8333 9011 8363 9041 ne
rect 8363 9015 8465 9041
rect 8585 9041 8687 9135
tri 8687 9041 8785 9139 sw
tri 8785 9041 8883 9139 ne
rect 8883 9135 9237 9139
rect 8883 9041 9015 9135
rect 8585 9015 8785 9041
rect 8363 9011 8785 9015
tri 8785 9011 8815 9041 sw
tri 8883 9011 8913 9041 ne
rect 8913 9015 9015 9041
rect 9135 9041 9237 9135
tri 9237 9041 9335 9139 sw
tri 9335 9041 9433 9139 ne
rect 9433 9135 9787 9139
rect 9433 9041 9565 9135
rect 9135 9015 9335 9041
rect 8913 9011 9335 9015
tri 9335 9011 9365 9041 sw
tri 9433 9011 9463 9041 ne
rect 9463 9015 9565 9041
rect 9685 9041 9787 9135
tri 9787 9041 9885 9139 sw
tri 9885 9041 9983 9139 ne
rect 9983 9135 10337 9139
rect 9983 9041 10115 9135
rect 9685 9015 9885 9041
rect 9463 9011 9885 9015
tri 9885 9011 9915 9041 sw
tri 9983 9011 10013 9041 ne
rect 10013 9015 10115 9041
rect 10235 9041 10337 9135
tri 10337 9041 10435 9139 sw
tri 10435 9041 10533 9139 ne
rect 10533 9135 10887 9139
rect 10533 9041 10665 9135
rect 10235 9015 10435 9041
rect 10013 9011 10435 9015
tri 10435 9011 10465 9041 sw
tri 10533 9011 10563 9041 ne
rect 10563 9015 10665 9041
rect 10785 9041 10887 9135
tri 10887 9041 10985 9139 sw
tri 10985 9041 11083 9139 ne
rect 11083 9135 11437 9139
rect 11083 9041 11215 9135
rect 10785 9015 10985 9041
rect 10563 9011 10985 9015
tri 10985 9011 11015 9041 sw
tri 11083 9011 11113 9041 ne
rect 11113 9015 11215 9041
rect 11335 9041 11437 9135
tri 11437 9041 11535 9139 sw
tri 11535 9041 11633 9139 ne
rect 11633 9135 11987 9139
rect 11633 9041 11765 9135
rect 11335 9015 11535 9041
rect 11113 9011 11535 9015
tri 11535 9011 11565 9041 sw
tri 11633 9011 11663 9041 ne
rect 11663 9015 11765 9041
rect 11885 9041 11987 9135
tri 11987 9041 12085 9139 sw
tri 12085 9041 12183 9139 ne
rect 12183 9135 12537 9139
rect 12183 9041 12315 9135
rect 11885 9015 12085 9041
rect 11663 9011 12085 9015
tri 12085 9011 12115 9041 sw
tri 12183 9011 12213 9041 ne
rect 12213 9015 12315 9041
rect 12435 9041 12537 9135
tri 12537 9041 12635 9139 sw
tri 12635 9041 12733 9139 ne
rect 12733 9135 13087 9139
rect 12733 9041 12865 9135
rect 12435 9015 12635 9041
rect 12213 9011 12635 9015
tri 12635 9011 12665 9041 sw
tri 12733 9011 12763 9041 ne
rect 12763 9015 12865 9041
rect 12985 9041 13087 9135
tri 13087 9041 13185 9139 sw
tri 13185 9041 13283 9139 ne
rect 13283 9135 13637 9139
rect 13283 9041 13415 9135
rect 12985 9015 13185 9041
rect 12763 9011 13185 9015
tri 13185 9011 13215 9041 sw
tri 13283 9011 13313 9041 ne
rect 13313 9015 13415 9041
rect 13535 9041 13637 9135
tri 13637 9041 13735 9139 sw
tri 13735 9041 13833 9139 ne
rect 13833 9135 14187 9139
rect 13833 9041 13965 9135
rect 13535 9015 13735 9041
rect 13313 9011 13735 9015
tri 13735 9011 13765 9041 sw
tri 13833 9011 13863 9041 ne
rect 13863 9015 13965 9041
rect 14085 9041 14187 9135
tri 14187 9041 14285 9139 sw
tri 14285 9041 14383 9139 ne
rect 14383 9135 14737 9139
rect 14383 9041 14515 9135
rect 14085 9015 14285 9041
rect 13863 9011 14285 9015
tri 14285 9011 14315 9041 sw
tri 14383 9011 14413 9041 ne
rect 14413 9015 14515 9041
rect 14635 9041 14737 9135
tri 14737 9041 14835 9139 sw
tri 14835 9041 14933 9139 ne
rect 14933 9135 15287 9139
rect 14933 9041 15065 9135
rect 14635 9015 14835 9041
rect 14413 9011 14835 9015
tri 14835 9011 14865 9041 sw
tri 14933 9011 14963 9041 ne
rect 14963 9015 15065 9041
rect 15185 9041 15287 9135
tri 15287 9041 15385 9139 sw
tri 15385 9041 15483 9139 ne
rect 15483 9135 15837 9139
rect 15483 9041 15615 9135
rect 15185 9015 15385 9041
rect 14963 9011 15385 9015
tri 15385 9011 15415 9041 sw
tri 15483 9011 15513 9041 ne
rect 15513 9015 15615 9041
rect 15735 9041 15837 9135
tri 15837 9041 15935 9139 sw
tri 15935 9041 16033 9139 ne
rect 16033 9135 16387 9139
rect 16033 9041 16165 9135
rect 15735 9015 15935 9041
rect 15513 9011 15935 9015
tri 15935 9011 15965 9041 sw
tri 16033 9011 16063 9041 ne
rect 16063 9015 16165 9041
rect 16285 9041 16387 9135
tri 16387 9041 16485 9139 sw
tri 16485 9041 16583 9139 ne
rect 16583 9135 16937 9139
rect 16583 9041 16715 9135
rect 16285 9015 16485 9041
rect 16063 9011 16485 9015
tri 16485 9011 16515 9041 sw
tri 16583 9011 16613 9041 ne
rect 16613 9015 16715 9041
rect 16835 9041 16937 9135
tri 16937 9041 17035 9139 sw
tri 17035 9041 17133 9139 ne
rect 17133 9135 17487 9139
rect 17133 9041 17265 9135
rect 16835 9015 17035 9041
rect 16613 9011 17035 9015
tri 17035 9011 17065 9041 sw
tri 17133 9011 17163 9041 ne
rect 17163 9015 17265 9041
rect 17385 9041 17487 9135
tri 17487 9041 17585 9139 sw
tri 17585 9041 17683 9139 ne
rect 17683 9135 18037 9139
rect 17683 9041 17815 9135
rect 17385 9015 17585 9041
rect 17163 9011 17585 9015
tri 17585 9011 17615 9041 sw
tri 17683 9011 17713 9041 ne
rect 17713 9015 17815 9041
rect 17935 9041 18037 9135
tri 18037 9041 18135 9139 sw
tri 18135 9041 18233 9139 ne
rect 18233 9135 18587 9139
rect 18233 9041 18365 9135
rect 17935 9015 18135 9041
rect 17713 9011 18135 9015
tri 18135 9011 18165 9041 sw
tri 18233 9011 18263 9041 ne
rect 18263 9015 18365 9041
rect 18485 9041 18587 9135
tri 18587 9041 18685 9139 sw
tri 18685 9041 18783 9139 ne
rect 18783 9135 19137 9139
rect 18783 9041 18915 9135
rect 18485 9015 18685 9041
rect 18263 9011 18685 9015
tri 18685 9011 18715 9041 sw
tri 18783 9011 18813 9041 ne
rect 18813 9015 18915 9041
rect 19035 9041 19137 9135
tri 19137 9041 19235 9139 sw
tri 19235 9041 19333 9139 ne
rect 19333 9135 20300 9139
rect 19333 9041 19465 9135
rect 19035 9015 19235 9041
rect 18813 9011 19235 9015
tri 19235 9011 19265 9041 sw
tri 19333 9011 19363 9041 ne
rect 19363 9015 19465 9041
rect 19585 9015 20300 9135
rect 19363 9011 20300 9015
tri 113 8913 211 9011 ne
rect 211 8913 565 9011
tri 565 8913 663 9011 sw
tri 663 8913 761 9011 ne
rect 761 8913 1115 9011
tri 1115 8913 1213 9011 sw
tri 1213 8913 1311 9011 ne
rect 1311 8913 1665 9011
tri 1665 8913 1763 9011 sw
tri 1763 8913 1861 9011 ne
rect 1861 8913 2215 9011
tri 2215 8913 2313 9011 sw
tri 2313 8913 2411 9011 ne
rect 2411 8913 2765 9011
tri 2765 8913 2863 9011 sw
tri 2863 8913 2961 9011 ne
rect 2961 8913 3315 9011
tri 3315 8913 3413 9011 sw
tri 3413 8913 3511 9011 ne
rect 3511 8913 3865 9011
tri 3865 8913 3963 9011 sw
tri 3963 8913 4061 9011 ne
rect 4061 8913 4415 9011
tri 4415 8913 4513 9011 sw
tri 4513 8913 4611 9011 ne
rect 4611 8913 4965 9011
tri 4965 8913 5063 9011 sw
tri 5063 8913 5161 9011 ne
rect 5161 8913 5515 9011
tri 5515 8913 5613 9011 sw
tri 5613 8913 5711 9011 ne
rect 5711 8913 6065 9011
tri 6065 8913 6163 9011 sw
tri 6163 8913 6261 9011 ne
rect 6261 8913 6615 9011
tri 6615 8913 6713 9011 sw
tri 6713 8913 6811 9011 ne
rect 6811 8913 7165 9011
tri 7165 8913 7263 9011 sw
tri 7263 8913 7361 9011 ne
rect 7361 8913 7715 9011
tri 7715 8913 7813 9011 sw
tri 7813 8913 7911 9011 ne
rect 7911 8913 8265 9011
tri 8265 8913 8363 9011 sw
tri 8363 8913 8461 9011 ne
rect 8461 8913 8815 9011
tri 8815 8913 8913 9011 sw
tri 8913 8913 9011 9011 ne
rect 9011 8913 9365 9011
tri 9365 8913 9463 9011 sw
tri 9463 8913 9561 9011 ne
rect 9561 8913 9915 9011
tri 9915 8913 10013 9011 sw
tri 10013 8913 10111 9011 ne
rect 10111 8913 10465 9011
tri 10465 8913 10563 9011 sw
tri 10563 8913 10661 9011 ne
rect 10661 8913 11015 9011
tri 11015 8913 11113 9011 sw
tri 11113 8913 11211 9011 ne
rect 11211 8913 11565 9011
tri 11565 8913 11663 9011 sw
tri 11663 8913 11761 9011 ne
rect 11761 8913 12115 9011
tri 12115 8913 12213 9011 sw
tri 12213 8913 12311 9011 ne
rect 12311 8913 12665 9011
tri 12665 8913 12763 9011 sw
tri 12763 8913 12861 9011 ne
rect 12861 8913 13215 9011
tri 13215 8913 13313 9011 sw
tri 13313 8913 13411 9011 ne
rect 13411 8913 13765 9011
tri 13765 8913 13863 9011 sw
tri 13863 8913 13961 9011 ne
rect 13961 8913 14315 9011
tri 14315 8913 14413 9011 sw
tri 14413 8913 14511 9011 ne
rect 14511 8913 14865 9011
tri 14865 8913 14963 9011 sw
tri 14963 8913 15061 9011 ne
rect 15061 8913 15415 9011
tri 15415 8913 15513 9011 sw
tri 15513 8913 15611 9011 ne
rect 15611 8913 15965 9011
tri 15965 8913 16063 9011 sw
tri 16063 8913 16161 9011 ne
rect 16161 8913 16515 9011
tri 16515 8913 16613 9011 sw
tri 16613 8913 16711 9011 ne
rect 16711 8913 17065 9011
tri 17065 8913 17163 9011 sw
tri 17163 8913 17261 9011 ne
rect 17261 8913 17615 9011
tri 17615 8913 17713 9011 sw
tri 17713 8913 17811 9011 ne
rect 17811 8913 18165 9011
tri 18165 8913 18263 9011 sw
tri 18263 8913 18361 9011 ne
rect 18361 8913 18715 9011
tri 18715 8913 18813 9011 sw
tri 18813 8913 18911 9011 ne
rect 18911 8913 19265 9011
tri 19265 8913 19363 9011 sw
tri 19363 8913 19461 9011 ne
rect 19461 8913 20300 9011
rect -2000 8883 113 8913
tri 113 8883 143 8913 sw
tri 211 8883 241 8913 ne
rect 241 8883 663 8913
tri 663 8883 693 8913 sw
tri 761 8883 791 8913 ne
rect 791 8883 1213 8913
tri 1213 8883 1243 8913 sw
tri 1311 8883 1341 8913 ne
rect 1341 8883 1763 8913
tri 1763 8883 1793 8913 sw
tri 1861 8883 1891 8913 ne
rect 1891 8883 2313 8913
tri 2313 8883 2343 8913 sw
tri 2411 8883 2441 8913 ne
rect 2441 8883 2863 8913
tri 2863 8883 2893 8913 sw
tri 2961 8883 2991 8913 ne
rect 2991 8883 3413 8913
tri 3413 8883 3443 8913 sw
tri 3511 8883 3541 8913 ne
rect 3541 8883 3963 8913
tri 3963 8883 3993 8913 sw
tri 4061 8883 4091 8913 ne
rect 4091 8883 4513 8913
tri 4513 8883 4543 8913 sw
tri 4611 8883 4641 8913 ne
rect 4641 8883 5063 8913
tri 5063 8883 5093 8913 sw
tri 5161 8883 5191 8913 ne
rect 5191 8883 5613 8913
tri 5613 8883 5643 8913 sw
tri 5711 8883 5741 8913 ne
rect 5741 8883 6163 8913
tri 6163 8883 6193 8913 sw
tri 6261 8883 6291 8913 ne
rect 6291 8883 6713 8913
tri 6713 8883 6743 8913 sw
tri 6811 8883 6841 8913 ne
rect 6841 8883 7263 8913
tri 7263 8883 7293 8913 sw
tri 7361 8883 7391 8913 ne
rect 7391 8883 7813 8913
tri 7813 8883 7843 8913 sw
tri 7911 8883 7941 8913 ne
rect 7941 8883 8363 8913
tri 8363 8883 8393 8913 sw
tri 8461 8883 8491 8913 ne
rect 8491 8883 8913 8913
tri 8913 8883 8943 8913 sw
tri 9011 8883 9041 8913 ne
rect 9041 8883 9463 8913
tri 9463 8883 9493 8913 sw
tri 9561 8883 9591 8913 ne
rect 9591 8883 10013 8913
tri 10013 8883 10043 8913 sw
tri 10111 8883 10141 8913 ne
rect 10141 8883 10563 8913
tri 10563 8883 10593 8913 sw
tri 10661 8883 10691 8913 ne
rect 10691 8883 11113 8913
tri 11113 8883 11143 8913 sw
tri 11211 8883 11241 8913 ne
rect 11241 8883 11663 8913
tri 11663 8883 11693 8913 sw
tri 11761 8883 11791 8913 ne
rect 11791 8883 12213 8913
tri 12213 8883 12243 8913 sw
tri 12311 8883 12341 8913 ne
rect 12341 8883 12763 8913
tri 12763 8883 12793 8913 sw
tri 12861 8883 12891 8913 ne
rect 12891 8883 13313 8913
tri 13313 8883 13343 8913 sw
tri 13411 8883 13441 8913 ne
rect 13441 8883 13863 8913
tri 13863 8883 13893 8913 sw
tri 13961 8883 13991 8913 ne
rect 13991 8883 14413 8913
tri 14413 8883 14443 8913 sw
tri 14511 8883 14541 8913 ne
rect 14541 8883 14963 8913
tri 14963 8883 14993 8913 sw
tri 15061 8883 15091 8913 ne
rect 15091 8883 15513 8913
tri 15513 8883 15543 8913 sw
tri 15611 8883 15641 8913 ne
rect 15641 8883 16063 8913
tri 16063 8883 16093 8913 sw
tri 16161 8883 16191 8913 ne
rect 16191 8883 16613 8913
tri 16613 8883 16643 8913 sw
tri 16711 8883 16741 8913 ne
rect 16741 8883 17163 8913
tri 17163 8883 17193 8913 sw
tri 17261 8883 17291 8913 ne
rect 17291 8883 17713 8913
tri 17713 8883 17743 8913 sw
tri 17811 8883 17841 8913 ne
rect 17841 8883 18263 8913
tri 18263 8883 18293 8913 sw
tri 18361 8883 18391 8913 ne
rect 18391 8883 18813 8913
tri 18813 8883 18843 8913 sw
tri 18911 8883 18941 8913 ne
rect 18941 8883 19363 8913
tri 19363 8883 19393 8913 sw
tri 19461 8883 19491 8913 ne
rect 19491 8883 20300 8913
rect -2000 8785 143 8883
tri 143 8785 241 8883 sw
tri 241 8785 339 8883 ne
rect 339 8785 693 8883
tri 693 8785 791 8883 sw
tri 791 8785 889 8883 ne
rect 889 8785 1243 8883
tri 1243 8785 1341 8883 sw
tri 1341 8785 1439 8883 ne
rect 1439 8785 1793 8883
tri 1793 8785 1891 8883 sw
tri 1891 8785 1989 8883 ne
rect 1989 8785 2343 8883
tri 2343 8785 2441 8883 sw
tri 2441 8785 2539 8883 ne
rect 2539 8785 2893 8883
tri 2893 8785 2991 8883 sw
tri 2991 8785 3089 8883 ne
rect 3089 8785 3443 8883
tri 3443 8785 3541 8883 sw
tri 3541 8785 3639 8883 ne
rect 3639 8785 3993 8883
tri 3993 8785 4091 8883 sw
tri 4091 8785 4189 8883 ne
rect 4189 8785 4543 8883
tri 4543 8785 4641 8883 sw
tri 4641 8785 4739 8883 ne
rect 4739 8785 5093 8883
tri 5093 8785 5191 8883 sw
tri 5191 8785 5289 8883 ne
rect 5289 8785 5643 8883
tri 5643 8785 5741 8883 sw
tri 5741 8785 5839 8883 ne
rect 5839 8785 6193 8883
tri 6193 8785 6291 8883 sw
tri 6291 8785 6389 8883 ne
rect 6389 8785 6743 8883
tri 6743 8785 6841 8883 sw
tri 6841 8785 6939 8883 ne
rect 6939 8785 7293 8883
tri 7293 8785 7391 8883 sw
tri 7391 8785 7489 8883 ne
rect 7489 8785 7843 8883
tri 7843 8785 7941 8883 sw
tri 7941 8785 8039 8883 ne
rect 8039 8785 8393 8883
tri 8393 8785 8491 8883 sw
tri 8491 8785 8589 8883 ne
rect 8589 8785 8943 8883
tri 8943 8785 9041 8883 sw
tri 9041 8785 9139 8883 ne
rect 9139 8785 9493 8883
tri 9493 8785 9591 8883 sw
tri 9591 8785 9689 8883 ne
rect 9689 8785 10043 8883
tri 10043 8785 10141 8883 sw
tri 10141 8785 10239 8883 ne
rect 10239 8785 10593 8883
tri 10593 8785 10691 8883 sw
tri 10691 8785 10789 8883 ne
rect 10789 8785 11143 8883
tri 11143 8785 11241 8883 sw
tri 11241 8785 11339 8883 ne
rect 11339 8785 11693 8883
tri 11693 8785 11791 8883 sw
tri 11791 8785 11889 8883 ne
rect 11889 8785 12243 8883
tri 12243 8785 12341 8883 sw
tri 12341 8785 12439 8883 ne
rect 12439 8785 12793 8883
tri 12793 8785 12891 8883 sw
tri 12891 8785 12989 8883 ne
rect 12989 8785 13343 8883
tri 13343 8785 13441 8883 sw
tri 13441 8785 13539 8883 ne
rect 13539 8785 13893 8883
tri 13893 8785 13991 8883 sw
tri 13991 8785 14089 8883 ne
rect 14089 8785 14443 8883
tri 14443 8785 14541 8883 sw
tri 14541 8785 14639 8883 ne
rect 14639 8785 14993 8883
tri 14993 8785 15091 8883 sw
tri 15091 8785 15189 8883 ne
rect 15189 8785 15543 8883
tri 15543 8785 15641 8883 sw
tri 15641 8785 15739 8883 ne
rect 15739 8785 16093 8883
tri 16093 8785 16191 8883 sw
tri 16191 8785 16289 8883 ne
rect 16289 8785 16643 8883
tri 16643 8785 16741 8883 sw
tri 16741 8785 16839 8883 ne
rect 16839 8785 17193 8883
tri 17193 8785 17291 8883 sw
tri 17291 8785 17389 8883 ne
rect 17389 8785 17743 8883
tri 17743 8785 17841 8883 sw
tri 17841 8785 17939 8883 ne
rect 17939 8785 18293 8883
tri 18293 8785 18391 8883 sw
tri 18391 8785 18489 8883 ne
rect 18489 8785 18843 8883
tri 18843 8785 18941 8883 sw
tri 18941 8785 19039 8883 ne
rect 19039 8785 19393 8883
tri 19393 8785 19491 8883 sw
tri 19491 8785 19589 8883 ne
rect 19589 8785 20300 8883
rect -2000 8687 241 8785
tri 241 8687 339 8785 sw
tri 339 8687 437 8785 ne
rect 437 8687 791 8785
tri 791 8687 889 8785 sw
tri 889 8687 987 8785 ne
rect 987 8687 1341 8785
tri 1341 8687 1439 8785 sw
tri 1439 8687 1537 8785 ne
rect 1537 8687 1891 8785
tri 1891 8687 1989 8785 sw
tri 1989 8687 2087 8785 ne
rect 2087 8687 2441 8785
tri 2441 8687 2539 8785 sw
tri 2539 8687 2637 8785 ne
rect 2637 8687 2991 8785
tri 2991 8687 3089 8785 sw
tri 3089 8687 3187 8785 ne
rect 3187 8687 3541 8785
tri 3541 8687 3639 8785 sw
tri 3639 8687 3737 8785 ne
rect 3737 8687 4091 8785
tri 4091 8687 4189 8785 sw
tri 4189 8687 4287 8785 ne
rect 4287 8687 4641 8785
tri 4641 8687 4739 8785 sw
tri 4739 8687 4837 8785 ne
rect 4837 8687 5191 8785
tri 5191 8687 5289 8785 sw
tri 5289 8687 5387 8785 ne
rect 5387 8687 5741 8785
tri 5741 8687 5839 8785 sw
tri 5839 8687 5937 8785 ne
rect 5937 8687 6291 8785
tri 6291 8687 6389 8785 sw
tri 6389 8687 6487 8785 ne
rect 6487 8687 6841 8785
tri 6841 8687 6939 8785 sw
tri 6939 8687 7037 8785 ne
rect 7037 8687 7391 8785
tri 7391 8687 7489 8785 sw
tri 7489 8687 7587 8785 ne
rect 7587 8687 7941 8785
tri 7941 8687 8039 8785 sw
tri 8039 8687 8137 8785 ne
rect 8137 8687 8491 8785
tri 8491 8687 8589 8785 sw
tri 8589 8687 8687 8785 ne
rect 8687 8687 9041 8785
tri 9041 8687 9139 8785 sw
tri 9139 8687 9237 8785 ne
rect 9237 8687 9591 8785
tri 9591 8687 9689 8785 sw
tri 9689 8687 9787 8785 ne
rect 9787 8687 10141 8785
tri 10141 8687 10239 8785 sw
tri 10239 8687 10337 8785 ne
rect 10337 8687 10691 8785
tri 10691 8687 10789 8785 sw
tri 10789 8687 10887 8785 ne
rect 10887 8687 11241 8785
tri 11241 8687 11339 8785 sw
tri 11339 8687 11437 8785 ne
rect 11437 8687 11791 8785
tri 11791 8687 11889 8785 sw
tri 11889 8687 11987 8785 ne
rect 11987 8687 12341 8785
tri 12341 8687 12439 8785 sw
tri 12439 8687 12537 8785 ne
rect 12537 8687 12891 8785
tri 12891 8687 12989 8785 sw
tri 12989 8687 13087 8785 ne
rect 13087 8687 13441 8785
tri 13441 8687 13539 8785 sw
tri 13539 8687 13637 8785 ne
rect 13637 8687 13991 8785
tri 13991 8687 14089 8785 sw
tri 14089 8687 14187 8785 ne
rect 14187 8687 14541 8785
tri 14541 8687 14639 8785 sw
tri 14639 8687 14737 8785 ne
rect 14737 8687 15091 8785
tri 15091 8687 15189 8785 sw
tri 15189 8687 15287 8785 ne
rect 15287 8687 15641 8785
tri 15641 8687 15739 8785 sw
tri 15739 8687 15837 8785 ne
rect 15837 8687 16191 8785
tri 16191 8687 16289 8785 sw
tri 16289 8687 16387 8785 ne
rect 16387 8687 16741 8785
tri 16741 8687 16839 8785 sw
tri 16839 8687 16937 8785 ne
rect 16937 8687 17291 8785
tri 17291 8687 17389 8785 sw
tri 17389 8687 17487 8785 ne
rect 17487 8687 17841 8785
tri 17841 8687 17939 8785 sw
tri 17939 8687 18037 8785 ne
rect 18037 8687 18391 8785
tri 18391 8687 18489 8785 sw
tri 18489 8687 18587 8785 ne
rect 18587 8687 18941 8785
tri 18941 8687 19039 8785 sw
tri 19039 8687 19137 8785 ne
rect 19137 8687 19491 8785
tri 19491 8687 19589 8785 sw
tri 19589 8687 19687 8785 ne
rect 19687 8687 20300 8785
rect -2000 8589 339 8687
tri 339 8589 437 8687 sw
tri 437 8589 535 8687 ne
rect 535 8589 889 8687
tri 889 8589 987 8687 sw
tri 987 8589 1085 8687 ne
rect 1085 8589 1439 8687
tri 1439 8589 1537 8687 sw
tri 1537 8589 1635 8687 ne
rect 1635 8589 1989 8687
tri 1989 8589 2087 8687 sw
tri 2087 8589 2185 8687 ne
rect 2185 8589 2539 8687
tri 2539 8589 2637 8687 sw
tri 2637 8589 2735 8687 ne
rect 2735 8589 3089 8687
tri 3089 8589 3187 8687 sw
tri 3187 8589 3285 8687 ne
rect 3285 8589 3639 8687
tri 3639 8589 3737 8687 sw
tri 3737 8589 3835 8687 ne
rect 3835 8589 4189 8687
tri 4189 8589 4287 8687 sw
tri 4287 8589 4385 8687 ne
rect 4385 8589 4739 8687
tri 4739 8589 4837 8687 sw
tri 4837 8589 4935 8687 ne
rect 4935 8589 5289 8687
tri 5289 8589 5387 8687 sw
tri 5387 8589 5485 8687 ne
rect 5485 8589 5839 8687
tri 5839 8589 5937 8687 sw
tri 5937 8589 6035 8687 ne
rect 6035 8589 6389 8687
tri 6389 8589 6487 8687 sw
tri 6487 8589 6585 8687 ne
rect 6585 8589 6939 8687
tri 6939 8589 7037 8687 sw
tri 7037 8589 7135 8687 ne
rect 7135 8589 7489 8687
tri 7489 8589 7587 8687 sw
tri 7587 8589 7685 8687 ne
rect 7685 8589 8039 8687
tri 8039 8589 8137 8687 sw
tri 8137 8589 8235 8687 ne
rect 8235 8589 8589 8687
tri 8589 8589 8687 8687 sw
tri 8687 8589 8785 8687 ne
rect 8785 8589 9139 8687
tri 9139 8589 9237 8687 sw
tri 9237 8589 9335 8687 ne
rect 9335 8589 9689 8687
tri 9689 8589 9787 8687 sw
tri 9787 8589 9885 8687 ne
rect 9885 8589 10239 8687
tri 10239 8589 10337 8687 sw
tri 10337 8589 10435 8687 ne
rect 10435 8589 10789 8687
tri 10789 8589 10887 8687 sw
tri 10887 8589 10985 8687 ne
rect 10985 8589 11339 8687
tri 11339 8589 11437 8687 sw
tri 11437 8589 11535 8687 ne
rect 11535 8589 11889 8687
tri 11889 8589 11987 8687 sw
tri 11987 8589 12085 8687 ne
rect 12085 8589 12439 8687
tri 12439 8589 12537 8687 sw
tri 12537 8589 12635 8687 ne
rect 12635 8589 12989 8687
tri 12989 8589 13087 8687 sw
tri 13087 8589 13185 8687 ne
rect 13185 8589 13539 8687
tri 13539 8589 13637 8687 sw
tri 13637 8589 13735 8687 ne
rect 13735 8589 14089 8687
tri 14089 8589 14187 8687 sw
tri 14187 8589 14285 8687 ne
rect 14285 8589 14639 8687
tri 14639 8589 14737 8687 sw
tri 14737 8589 14835 8687 ne
rect 14835 8589 15189 8687
tri 15189 8589 15287 8687 sw
tri 15287 8589 15385 8687 ne
rect 15385 8589 15739 8687
tri 15739 8589 15837 8687 sw
tri 15837 8589 15935 8687 ne
rect 15935 8589 16289 8687
tri 16289 8589 16387 8687 sw
tri 16387 8589 16485 8687 ne
rect 16485 8589 16839 8687
tri 16839 8589 16937 8687 sw
tri 16937 8589 17035 8687 ne
rect 17035 8589 17389 8687
tri 17389 8589 17487 8687 sw
tri 17487 8589 17585 8687 ne
rect 17585 8589 17939 8687
tri 17939 8589 18037 8687 sw
tri 18037 8589 18135 8687 ne
rect 18135 8589 18489 8687
tri 18489 8589 18587 8687 sw
tri 18587 8589 18685 8687 ne
rect 18685 8589 19039 8687
tri 19039 8589 19137 8687 sw
tri 19137 8589 19235 8687 ne
rect 19235 8589 19589 8687
tri 19589 8589 19687 8687 sw
rect 20800 8589 21800 9237
rect -2000 8585 437 8589
rect -2000 8465 215 8585
rect 335 8491 437 8585
tri 437 8491 535 8589 sw
tri 535 8491 633 8589 ne
rect 633 8585 987 8589
rect 633 8491 765 8585
rect 335 8465 535 8491
rect -2000 8461 535 8465
rect -2000 7813 -1000 8461
tri 113 8363 211 8461 ne
rect 211 8413 535 8461
tri 535 8413 613 8491 sw
tri 633 8413 711 8491 ne
rect 711 8465 765 8491
rect 885 8491 987 8585
tri 987 8491 1085 8589 sw
tri 1085 8491 1183 8589 ne
rect 1183 8585 1537 8589
rect 1183 8491 1315 8585
rect 885 8465 1085 8491
rect 711 8413 1085 8465
tri 1085 8413 1163 8491 sw
tri 1183 8413 1261 8491 ne
rect 1261 8465 1315 8491
rect 1435 8491 1537 8585
tri 1537 8491 1635 8589 sw
tri 1635 8491 1733 8589 ne
rect 1733 8585 2087 8589
rect 1733 8491 1865 8585
rect 1435 8465 1635 8491
rect 1261 8413 1635 8465
tri 1635 8413 1713 8491 sw
tri 1733 8413 1811 8491 ne
rect 1811 8465 1865 8491
rect 1985 8491 2087 8585
tri 2087 8491 2185 8589 sw
tri 2185 8491 2283 8589 ne
rect 2283 8585 2637 8589
rect 2283 8491 2415 8585
rect 1985 8465 2185 8491
rect 1811 8413 2185 8465
tri 2185 8413 2263 8491 sw
tri 2283 8413 2361 8491 ne
rect 2361 8465 2415 8491
rect 2535 8491 2637 8585
tri 2637 8491 2735 8589 sw
tri 2735 8491 2833 8589 ne
rect 2833 8585 3187 8589
rect 2833 8491 2965 8585
rect 2535 8465 2735 8491
rect 2361 8413 2735 8465
tri 2735 8413 2813 8491 sw
tri 2833 8413 2911 8491 ne
rect 2911 8465 2965 8491
rect 3085 8491 3187 8585
tri 3187 8491 3285 8589 sw
tri 3285 8491 3383 8589 ne
rect 3383 8585 3737 8589
rect 3383 8491 3515 8585
rect 3085 8465 3285 8491
rect 2911 8413 3285 8465
tri 3285 8413 3363 8491 sw
tri 3383 8413 3461 8491 ne
rect 3461 8465 3515 8491
rect 3635 8491 3737 8585
tri 3737 8491 3835 8589 sw
tri 3835 8491 3933 8589 ne
rect 3933 8585 4287 8589
rect 3933 8491 4065 8585
rect 3635 8465 3835 8491
rect 3461 8413 3835 8465
tri 3835 8413 3913 8491 sw
tri 3933 8413 4011 8491 ne
rect 4011 8465 4065 8491
rect 4185 8491 4287 8585
tri 4287 8491 4385 8589 sw
tri 4385 8491 4483 8589 ne
rect 4483 8585 4837 8589
rect 4483 8491 4615 8585
rect 4185 8465 4385 8491
rect 4011 8413 4385 8465
tri 4385 8413 4463 8491 sw
tri 4483 8413 4561 8491 ne
rect 4561 8465 4615 8491
rect 4735 8491 4837 8585
tri 4837 8491 4935 8589 sw
tri 4935 8491 5033 8589 ne
rect 5033 8585 5387 8589
rect 5033 8491 5165 8585
rect 4735 8465 4935 8491
rect 4561 8413 4935 8465
tri 4935 8413 5013 8491 sw
tri 5033 8413 5111 8491 ne
rect 5111 8465 5165 8491
rect 5285 8491 5387 8585
tri 5387 8491 5485 8589 sw
tri 5485 8491 5583 8589 ne
rect 5583 8585 5937 8589
rect 5583 8491 5715 8585
rect 5285 8465 5485 8491
rect 5111 8413 5485 8465
tri 5485 8413 5563 8491 sw
tri 5583 8413 5661 8491 ne
rect 5661 8465 5715 8491
rect 5835 8491 5937 8585
tri 5937 8491 6035 8589 sw
tri 6035 8491 6133 8589 ne
rect 6133 8585 6487 8589
rect 6133 8491 6265 8585
rect 5835 8465 6035 8491
rect 5661 8413 6035 8465
tri 6035 8413 6113 8491 sw
tri 6133 8413 6211 8491 ne
rect 6211 8465 6265 8491
rect 6385 8491 6487 8585
tri 6487 8491 6585 8589 sw
tri 6585 8491 6683 8589 ne
rect 6683 8585 7037 8589
rect 6683 8491 6815 8585
rect 6385 8465 6585 8491
rect 6211 8413 6585 8465
tri 6585 8413 6663 8491 sw
tri 6683 8413 6761 8491 ne
rect 6761 8465 6815 8491
rect 6935 8491 7037 8585
tri 7037 8491 7135 8589 sw
tri 7135 8491 7233 8589 ne
rect 7233 8585 7587 8589
rect 7233 8491 7365 8585
rect 6935 8465 7135 8491
rect 6761 8413 7135 8465
tri 7135 8413 7213 8491 sw
tri 7233 8413 7311 8491 ne
rect 7311 8465 7365 8491
rect 7485 8491 7587 8585
tri 7587 8491 7685 8589 sw
tri 7685 8491 7783 8589 ne
rect 7783 8585 8137 8589
rect 7783 8491 7915 8585
rect 7485 8465 7685 8491
rect 7311 8413 7685 8465
tri 7685 8413 7763 8491 sw
tri 7783 8413 7861 8491 ne
rect 7861 8465 7915 8491
rect 8035 8491 8137 8585
tri 8137 8491 8235 8589 sw
tri 8235 8491 8333 8589 ne
rect 8333 8585 8687 8589
rect 8333 8491 8465 8585
rect 8035 8465 8235 8491
rect 7861 8413 8235 8465
tri 8235 8413 8313 8491 sw
tri 8333 8413 8411 8491 ne
rect 8411 8465 8465 8491
rect 8585 8491 8687 8585
tri 8687 8491 8785 8589 sw
tri 8785 8491 8883 8589 ne
rect 8883 8585 9237 8589
rect 8883 8491 9015 8585
rect 8585 8465 8785 8491
rect 8411 8413 8785 8465
tri 8785 8413 8863 8491 sw
tri 8883 8413 8961 8491 ne
rect 8961 8465 9015 8491
rect 9135 8491 9237 8585
tri 9237 8491 9335 8589 sw
tri 9335 8491 9433 8589 ne
rect 9433 8585 9787 8589
rect 9433 8491 9565 8585
rect 9135 8465 9335 8491
rect 8961 8413 9335 8465
tri 9335 8413 9413 8491 sw
tri 9433 8413 9511 8491 ne
rect 9511 8465 9565 8491
rect 9685 8491 9787 8585
tri 9787 8491 9885 8589 sw
tri 9885 8491 9983 8589 ne
rect 9983 8585 10337 8589
rect 9983 8491 10115 8585
rect 9685 8465 9885 8491
rect 9511 8413 9885 8465
tri 9885 8413 9963 8491 sw
tri 9983 8413 10061 8491 ne
rect 10061 8465 10115 8491
rect 10235 8491 10337 8585
tri 10337 8491 10435 8589 sw
tri 10435 8491 10533 8589 ne
rect 10533 8585 10887 8589
rect 10533 8491 10665 8585
rect 10235 8465 10435 8491
rect 10061 8413 10435 8465
tri 10435 8413 10513 8491 sw
tri 10533 8413 10611 8491 ne
rect 10611 8465 10665 8491
rect 10785 8491 10887 8585
tri 10887 8491 10985 8589 sw
tri 10985 8491 11083 8589 ne
rect 11083 8585 11437 8589
rect 11083 8491 11215 8585
rect 10785 8465 10985 8491
rect 10611 8413 10985 8465
tri 10985 8413 11063 8491 sw
tri 11083 8413 11161 8491 ne
rect 11161 8465 11215 8491
rect 11335 8491 11437 8585
tri 11437 8491 11535 8589 sw
tri 11535 8491 11633 8589 ne
rect 11633 8585 11987 8589
rect 11633 8491 11765 8585
rect 11335 8465 11535 8491
rect 11161 8413 11535 8465
tri 11535 8413 11613 8491 sw
tri 11633 8413 11711 8491 ne
rect 11711 8465 11765 8491
rect 11885 8491 11987 8585
tri 11987 8491 12085 8589 sw
tri 12085 8491 12183 8589 ne
rect 12183 8585 12537 8589
rect 12183 8491 12315 8585
rect 11885 8465 12085 8491
rect 11711 8413 12085 8465
tri 12085 8413 12163 8491 sw
tri 12183 8413 12261 8491 ne
rect 12261 8465 12315 8491
rect 12435 8491 12537 8585
tri 12537 8491 12635 8589 sw
tri 12635 8491 12733 8589 ne
rect 12733 8585 13087 8589
rect 12733 8491 12865 8585
rect 12435 8465 12635 8491
rect 12261 8413 12635 8465
tri 12635 8413 12713 8491 sw
tri 12733 8413 12811 8491 ne
rect 12811 8465 12865 8491
rect 12985 8491 13087 8585
tri 13087 8491 13185 8589 sw
tri 13185 8491 13283 8589 ne
rect 13283 8585 13637 8589
rect 13283 8491 13415 8585
rect 12985 8465 13185 8491
rect 12811 8413 13185 8465
tri 13185 8413 13263 8491 sw
tri 13283 8413 13361 8491 ne
rect 13361 8465 13415 8491
rect 13535 8491 13637 8585
tri 13637 8491 13735 8589 sw
tri 13735 8491 13833 8589 ne
rect 13833 8585 14187 8589
rect 13833 8491 13965 8585
rect 13535 8465 13735 8491
rect 13361 8413 13735 8465
tri 13735 8413 13813 8491 sw
tri 13833 8413 13911 8491 ne
rect 13911 8465 13965 8491
rect 14085 8491 14187 8585
tri 14187 8491 14285 8589 sw
tri 14285 8491 14383 8589 ne
rect 14383 8585 14737 8589
rect 14383 8491 14515 8585
rect 14085 8465 14285 8491
rect 13911 8413 14285 8465
tri 14285 8413 14363 8491 sw
tri 14383 8413 14461 8491 ne
rect 14461 8465 14515 8491
rect 14635 8491 14737 8585
tri 14737 8491 14835 8589 sw
tri 14835 8491 14933 8589 ne
rect 14933 8585 15287 8589
rect 14933 8491 15065 8585
rect 14635 8465 14835 8491
rect 14461 8413 14835 8465
tri 14835 8413 14913 8491 sw
tri 14933 8413 15011 8491 ne
rect 15011 8465 15065 8491
rect 15185 8491 15287 8585
tri 15287 8491 15385 8589 sw
tri 15385 8491 15483 8589 ne
rect 15483 8585 15837 8589
rect 15483 8491 15615 8585
rect 15185 8465 15385 8491
rect 15011 8413 15385 8465
tri 15385 8413 15463 8491 sw
tri 15483 8413 15561 8491 ne
rect 15561 8465 15615 8491
rect 15735 8491 15837 8585
tri 15837 8491 15935 8589 sw
tri 15935 8491 16033 8589 ne
rect 16033 8585 16387 8589
rect 16033 8491 16165 8585
rect 15735 8465 15935 8491
rect 15561 8413 15935 8465
tri 15935 8413 16013 8491 sw
tri 16033 8413 16111 8491 ne
rect 16111 8465 16165 8491
rect 16285 8491 16387 8585
tri 16387 8491 16485 8589 sw
tri 16485 8491 16583 8589 ne
rect 16583 8585 16937 8589
rect 16583 8491 16715 8585
rect 16285 8465 16485 8491
rect 16111 8413 16485 8465
tri 16485 8413 16563 8491 sw
tri 16583 8413 16661 8491 ne
rect 16661 8465 16715 8491
rect 16835 8491 16937 8585
tri 16937 8491 17035 8589 sw
tri 17035 8491 17133 8589 ne
rect 17133 8585 17487 8589
rect 17133 8491 17265 8585
rect 16835 8465 17035 8491
rect 16661 8413 17035 8465
tri 17035 8413 17113 8491 sw
tri 17133 8413 17211 8491 ne
rect 17211 8465 17265 8491
rect 17385 8491 17487 8585
tri 17487 8491 17585 8589 sw
tri 17585 8491 17683 8589 ne
rect 17683 8585 18037 8589
rect 17683 8491 17815 8585
rect 17385 8465 17585 8491
rect 17211 8413 17585 8465
tri 17585 8413 17663 8491 sw
tri 17683 8413 17761 8491 ne
rect 17761 8465 17815 8491
rect 17935 8491 18037 8585
tri 18037 8491 18135 8589 sw
tri 18135 8491 18233 8589 ne
rect 18233 8585 18587 8589
rect 18233 8491 18365 8585
rect 17935 8465 18135 8491
rect 17761 8413 18135 8465
tri 18135 8413 18213 8491 sw
tri 18233 8413 18311 8491 ne
rect 18311 8465 18365 8491
rect 18485 8491 18587 8585
tri 18587 8491 18685 8589 sw
tri 18685 8491 18783 8589 ne
rect 18783 8585 19137 8589
rect 18783 8491 18915 8585
rect 18485 8465 18685 8491
rect 18311 8413 18685 8465
tri 18685 8413 18763 8491 sw
tri 18783 8413 18861 8491 ne
rect 18861 8465 18915 8491
rect 19035 8491 19137 8585
tri 19137 8491 19235 8589 sw
tri 19235 8491 19333 8589 ne
rect 19333 8585 21800 8589
rect 19333 8491 19465 8585
rect 19035 8465 19235 8491
rect 18861 8413 19235 8465
tri 19235 8413 19313 8491 sw
tri 19333 8413 19411 8491 ne
rect 19411 8465 19465 8491
rect 19585 8465 21800 8585
rect 19411 8413 21800 8465
rect 211 8363 613 8413
rect -500 8313 113 8363
tri 113 8313 163 8363 sw
tri 211 8313 261 8363 ne
rect 261 8333 613 8363
tri 613 8333 693 8413 sw
tri 711 8333 791 8413 ne
rect 791 8333 1163 8413
tri 1163 8333 1243 8413 sw
tri 1261 8333 1341 8413 ne
rect 1341 8333 1713 8413
tri 1713 8333 1793 8413 sw
tri 1811 8333 1891 8413 ne
rect 1891 8333 2263 8413
tri 2263 8333 2343 8413 sw
tri 2361 8333 2441 8413 ne
rect 2441 8333 2813 8413
tri 2813 8333 2893 8413 sw
tri 2911 8333 2991 8413 ne
rect 2991 8333 3363 8413
tri 3363 8333 3443 8413 sw
tri 3461 8333 3541 8413 ne
rect 3541 8333 3913 8413
tri 3913 8333 3993 8413 sw
tri 4011 8333 4091 8413 ne
rect 4091 8333 4463 8413
tri 4463 8333 4543 8413 sw
tri 4561 8333 4641 8413 ne
rect 4641 8333 5013 8413
tri 5013 8333 5093 8413 sw
tri 5111 8333 5191 8413 ne
rect 5191 8333 5563 8413
tri 5563 8333 5643 8413 sw
tri 5661 8333 5741 8413 ne
rect 5741 8333 6113 8413
tri 6113 8333 6193 8413 sw
tri 6211 8333 6291 8413 ne
rect 6291 8333 6663 8413
tri 6663 8333 6743 8413 sw
tri 6761 8333 6841 8413 ne
rect 6841 8333 7213 8413
tri 7213 8333 7293 8413 sw
tri 7311 8333 7391 8413 ne
rect 7391 8333 7763 8413
tri 7763 8333 7843 8413 sw
tri 7861 8333 7941 8413 ne
rect 7941 8333 8313 8413
tri 8313 8333 8393 8413 sw
tri 8411 8333 8491 8413 ne
rect 8491 8333 8863 8413
tri 8863 8333 8943 8413 sw
tri 8961 8333 9041 8413 ne
rect 9041 8333 9413 8413
tri 9413 8333 9493 8413 sw
tri 9511 8333 9591 8413 ne
rect 9591 8333 9963 8413
tri 9963 8333 10043 8413 sw
tri 10061 8333 10141 8413 ne
rect 10141 8333 10513 8413
tri 10513 8333 10593 8413 sw
tri 10611 8333 10691 8413 ne
rect 10691 8333 11063 8413
tri 11063 8333 11143 8413 sw
tri 11161 8333 11241 8413 ne
rect 11241 8333 11613 8413
tri 11613 8333 11693 8413 sw
tri 11711 8333 11791 8413 ne
rect 11791 8333 12163 8413
tri 12163 8333 12243 8413 sw
tri 12261 8333 12341 8413 ne
rect 12341 8333 12713 8413
tri 12713 8333 12793 8413 sw
tri 12811 8333 12891 8413 ne
rect 12891 8333 13263 8413
tri 13263 8333 13343 8413 sw
tri 13361 8333 13441 8413 ne
rect 13441 8333 13813 8413
tri 13813 8333 13893 8413 sw
tri 13911 8333 13991 8413 ne
rect 13991 8333 14363 8413
tri 14363 8333 14443 8413 sw
tri 14461 8333 14541 8413 ne
rect 14541 8333 14913 8413
tri 14913 8333 14993 8413 sw
tri 15011 8333 15091 8413 ne
rect 15091 8333 15463 8413
tri 15463 8333 15543 8413 sw
tri 15561 8333 15641 8413 ne
rect 15641 8333 16013 8413
tri 16013 8333 16093 8413 sw
tri 16111 8333 16191 8413 ne
rect 16191 8333 16563 8413
tri 16563 8333 16643 8413 sw
tri 16661 8333 16741 8413 ne
rect 16741 8333 17113 8413
tri 17113 8333 17193 8413 sw
tri 17211 8333 17291 8413 ne
rect 17291 8333 17663 8413
tri 17663 8333 17743 8413 sw
tri 17761 8333 17841 8413 ne
rect 17841 8333 18213 8413
tri 18213 8333 18293 8413 sw
tri 18311 8333 18391 8413 ne
rect 18391 8333 18763 8413
tri 18763 8333 18843 8413 sw
tri 18861 8333 18941 8413 ne
rect 18941 8333 19313 8413
tri 19313 8333 19393 8413 sw
tri 19411 8333 19491 8413 ne
rect 19491 8333 20100 8413
rect 261 8313 693 8333
rect -500 8235 163 8313
tri 163 8235 241 8313 sw
tri 261 8235 339 8313 ne
rect 339 8235 693 8313
tri 693 8235 791 8333 sw
tri 791 8235 889 8333 ne
rect 889 8235 1243 8333
tri 1243 8235 1341 8333 sw
tri 1341 8235 1439 8333 ne
rect 1439 8235 1793 8333
tri 1793 8235 1891 8333 sw
tri 1891 8235 1989 8333 ne
rect 1989 8235 2343 8333
tri 2343 8235 2441 8333 sw
tri 2441 8235 2539 8333 ne
rect 2539 8235 2893 8333
tri 2893 8235 2991 8333 sw
tri 2991 8235 3089 8333 ne
rect 3089 8235 3443 8333
tri 3443 8235 3541 8333 sw
tri 3541 8235 3639 8333 ne
rect 3639 8235 3993 8333
tri 3993 8235 4091 8333 sw
tri 4091 8235 4189 8333 ne
rect 4189 8235 4543 8333
tri 4543 8235 4641 8333 sw
tri 4641 8235 4739 8333 ne
rect 4739 8235 5093 8333
tri 5093 8235 5191 8333 sw
tri 5191 8235 5289 8333 ne
rect 5289 8235 5643 8333
tri 5643 8235 5741 8333 sw
tri 5741 8235 5839 8333 ne
rect 5839 8235 6193 8333
tri 6193 8235 6291 8333 sw
tri 6291 8235 6389 8333 ne
rect 6389 8235 6743 8333
tri 6743 8235 6841 8333 sw
tri 6841 8235 6939 8333 ne
rect 6939 8235 7293 8333
tri 7293 8235 7391 8333 sw
tri 7391 8235 7489 8333 ne
rect 7489 8235 7843 8333
tri 7843 8235 7941 8333 sw
tri 7941 8235 8039 8333 ne
rect 8039 8235 8393 8333
tri 8393 8235 8491 8333 sw
tri 8491 8235 8589 8333 ne
rect 8589 8235 8943 8333
tri 8943 8235 9041 8333 sw
tri 9041 8235 9139 8333 ne
rect 9139 8235 9493 8333
tri 9493 8235 9591 8333 sw
tri 9591 8235 9689 8333 ne
rect 9689 8235 10043 8333
tri 10043 8235 10141 8333 sw
tri 10141 8235 10239 8333 ne
rect 10239 8235 10593 8333
tri 10593 8235 10691 8333 sw
tri 10691 8235 10789 8333 ne
rect 10789 8235 11143 8333
tri 11143 8235 11241 8333 sw
tri 11241 8235 11339 8333 ne
rect 11339 8235 11693 8333
tri 11693 8235 11791 8333 sw
tri 11791 8235 11889 8333 ne
rect 11889 8235 12243 8333
tri 12243 8235 12341 8333 sw
tri 12341 8235 12439 8333 ne
rect 12439 8235 12793 8333
tri 12793 8235 12891 8333 sw
tri 12891 8235 12989 8333 ne
rect 12989 8235 13343 8333
tri 13343 8235 13441 8333 sw
tri 13441 8235 13539 8333 ne
rect 13539 8235 13893 8333
tri 13893 8235 13991 8333 sw
tri 13991 8235 14089 8333 ne
rect 14089 8235 14443 8333
tri 14443 8235 14541 8333 sw
tri 14541 8235 14639 8333 ne
rect 14639 8235 14993 8333
tri 14993 8235 15091 8333 sw
tri 15091 8235 15189 8333 ne
rect 15189 8235 15543 8333
tri 15543 8235 15641 8333 sw
tri 15641 8235 15739 8333 ne
rect 15739 8235 16093 8333
tri 16093 8235 16191 8333 sw
tri 16191 8235 16289 8333 ne
rect 16289 8235 16643 8333
tri 16643 8235 16741 8333 sw
tri 16741 8235 16839 8333 ne
rect 16839 8235 17193 8333
tri 17193 8235 17291 8333 sw
tri 17291 8235 17389 8333 ne
rect 17389 8235 17743 8333
tri 17743 8235 17841 8333 sw
tri 17841 8235 17939 8333 ne
rect 17939 8235 18293 8333
tri 18293 8235 18391 8333 sw
tri 18391 8235 18489 8333 ne
rect 18489 8235 18843 8333
tri 18843 8235 18941 8333 sw
tri 18941 8235 19039 8333 ne
rect 19039 8235 19393 8333
tri 19393 8235 19491 8333 sw
tri 19491 8235 19589 8333 ne
rect 19589 8313 20100 8333
rect 20200 8313 21800 8413
rect 19589 8235 21800 8313
rect -500 8187 241 8235
rect -500 8087 -400 8187
rect -300 8137 241 8187
tri 241 8137 339 8235 sw
tri 339 8137 437 8235 ne
rect 437 8137 791 8235
tri 791 8137 889 8235 sw
tri 889 8137 987 8235 ne
rect 987 8137 1341 8235
tri 1341 8137 1439 8235 sw
tri 1439 8137 1537 8235 ne
rect 1537 8137 1891 8235
tri 1891 8137 1989 8235 sw
tri 1989 8137 2087 8235 ne
rect 2087 8137 2441 8235
tri 2441 8137 2539 8235 sw
tri 2539 8137 2637 8235 ne
rect 2637 8137 2991 8235
tri 2991 8137 3089 8235 sw
tri 3089 8137 3187 8235 ne
rect 3187 8137 3541 8235
tri 3541 8137 3639 8235 sw
tri 3639 8137 3737 8235 ne
rect 3737 8137 4091 8235
tri 4091 8137 4189 8235 sw
tri 4189 8137 4287 8235 ne
rect 4287 8137 4641 8235
tri 4641 8137 4739 8235 sw
tri 4739 8137 4837 8235 ne
rect 4837 8137 5191 8235
tri 5191 8137 5289 8235 sw
tri 5289 8137 5387 8235 ne
rect 5387 8137 5741 8235
tri 5741 8137 5839 8235 sw
tri 5839 8137 5937 8235 ne
rect 5937 8137 6291 8235
tri 6291 8137 6389 8235 sw
tri 6389 8137 6487 8235 ne
rect 6487 8137 6841 8235
tri 6841 8137 6939 8235 sw
tri 6939 8137 7037 8235 ne
rect 7037 8137 7391 8235
tri 7391 8137 7489 8235 sw
tri 7489 8137 7587 8235 ne
rect 7587 8137 7941 8235
tri 7941 8137 8039 8235 sw
tri 8039 8137 8137 8235 ne
rect 8137 8137 8491 8235
tri 8491 8137 8589 8235 sw
tri 8589 8137 8687 8235 ne
rect 8687 8137 9041 8235
tri 9041 8137 9139 8235 sw
tri 9139 8137 9237 8235 ne
rect 9237 8137 9591 8235
tri 9591 8137 9689 8235 sw
tri 9689 8137 9787 8235 ne
rect 9787 8137 10141 8235
tri 10141 8137 10239 8235 sw
tri 10239 8137 10337 8235 ne
rect 10337 8137 10691 8235
tri 10691 8137 10789 8235 sw
tri 10789 8137 10887 8235 ne
rect 10887 8137 11241 8235
tri 11241 8137 11339 8235 sw
tri 11339 8137 11437 8235 ne
rect 11437 8137 11791 8235
tri 11791 8137 11889 8235 sw
tri 11889 8137 11987 8235 ne
rect 11987 8137 12341 8235
tri 12341 8137 12439 8235 sw
tri 12439 8137 12537 8235 ne
rect 12537 8137 12891 8235
tri 12891 8137 12989 8235 sw
tri 12989 8137 13087 8235 ne
rect 13087 8137 13441 8235
tri 13441 8137 13539 8235 sw
tri 13539 8137 13637 8235 ne
rect 13637 8137 13991 8235
tri 13991 8137 14089 8235 sw
tri 14089 8137 14187 8235 ne
rect 14187 8137 14541 8235
tri 14541 8137 14639 8235 sw
tri 14639 8137 14737 8235 ne
rect 14737 8137 15091 8235
tri 15091 8137 15189 8235 sw
tri 15189 8137 15287 8235 ne
rect 15287 8137 15641 8235
tri 15641 8137 15739 8235 sw
tri 15739 8137 15837 8235 ne
rect 15837 8137 16191 8235
tri 16191 8137 16289 8235 sw
tri 16289 8137 16387 8235 ne
rect 16387 8137 16741 8235
tri 16741 8137 16839 8235 sw
tri 16839 8137 16937 8235 ne
rect 16937 8137 17291 8235
tri 17291 8137 17389 8235 sw
tri 17389 8137 17487 8235 ne
rect 17487 8137 17841 8235
tri 17841 8137 17939 8235 sw
tri 17939 8137 18037 8235 ne
rect 18037 8137 18391 8235
tri 18391 8137 18489 8235 sw
tri 18489 8137 18587 8235 ne
rect 18587 8137 18941 8235
tri 18941 8137 19039 8235 sw
tri 19039 8137 19137 8235 ne
rect 19137 8137 19491 8235
tri 19491 8137 19589 8235 sw
tri 19589 8137 19687 8235 ne
rect 19687 8137 21800 8235
rect -300 8087 339 8137
rect -500 8039 339 8087
tri 339 8039 437 8137 sw
tri 437 8039 535 8137 ne
rect 535 8039 889 8137
tri 889 8039 987 8137 sw
tri 987 8039 1085 8137 ne
rect 1085 8039 1439 8137
tri 1439 8039 1537 8137 sw
tri 1537 8039 1635 8137 ne
rect 1635 8039 1989 8137
tri 1989 8039 2087 8137 sw
tri 2087 8039 2185 8137 ne
rect 2185 8039 2539 8137
tri 2539 8039 2637 8137 sw
tri 2637 8039 2735 8137 ne
rect 2735 8039 3089 8137
tri 3089 8039 3187 8137 sw
tri 3187 8039 3285 8137 ne
rect 3285 8039 3639 8137
tri 3639 8039 3737 8137 sw
tri 3737 8039 3835 8137 ne
rect 3835 8039 4189 8137
tri 4189 8039 4287 8137 sw
tri 4287 8039 4385 8137 ne
rect 4385 8039 4739 8137
tri 4739 8039 4837 8137 sw
tri 4837 8039 4935 8137 ne
rect 4935 8039 5289 8137
tri 5289 8039 5387 8137 sw
tri 5387 8039 5485 8137 ne
rect 5485 8039 5839 8137
tri 5839 8039 5937 8137 sw
tri 5937 8039 6035 8137 ne
rect 6035 8039 6389 8137
tri 6389 8039 6487 8137 sw
tri 6487 8039 6585 8137 ne
rect 6585 8039 6939 8137
tri 6939 8039 7037 8137 sw
tri 7037 8039 7135 8137 ne
rect 7135 8039 7489 8137
tri 7489 8039 7587 8137 sw
tri 7587 8039 7685 8137 ne
rect 7685 8039 8039 8137
tri 8039 8039 8137 8137 sw
tri 8137 8039 8235 8137 ne
rect 8235 8039 8589 8137
tri 8589 8039 8687 8137 sw
tri 8687 8039 8785 8137 ne
rect 8785 8039 9139 8137
tri 9139 8039 9237 8137 sw
tri 9237 8039 9335 8137 ne
rect 9335 8039 9689 8137
tri 9689 8039 9787 8137 sw
tri 9787 8039 9885 8137 ne
rect 9885 8039 10239 8137
tri 10239 8039 10337 8137 sw
tri 10337 8039 10435 8137 ne
rect 10435 8039 10789 8137
tri 10789 8039 10887 8137 sw
tri 10887 8039 10985 8137 ne
rect 10985 8039 11339 8137
tri 11339 8039 11437 8137 sw
tri 11437 8039 11535 8137 ne
rect 11535 8039 11889 8137
tri 11889 8039 11987 8137 sw
tri 11987 8039 12085 8137 ne
rect 12085 8039 12439 8137
tri 12439 8039 12537 8137 sw
tri 12537 8039 12635 8137 ne
rect 12635 8039 12989 8137
tri 12989 8039 13087 8137 sw
tri 13087 8039 13185 8137 ne
rect 13185 8039 13539 8137
tri 13539 8039 13637 8137 sw
tri 13637 8039 13735 8137 ne
rect 13735 8039 14089 8137
tri 14089 8039 14187 8137 sw
tri 14187 8039 14285 8137 ne
rect 14285 8039 14639 8137
tri 14639 8039 14737 8137 sw
tri 14737 8039 14835 8137 ne
rect 14835 8039 15189 8137
tri 15189 8039 15287 8137 sw
tri 15287 8039 15385 8137 ne
rect 15385 8039 15739 8137
tri 15739 8039 15837 8137 sw
tri 15837 8039 15935 8137 ne
rect 15935 8039 16289 8137
tri 16289 8039 16387 8137 sw
tri 16387 8039 16485 8137 ne
rect 16485 8039 16839 8137
tri 16839 8039 16937 8137 sw
tri 16937 8039 17035 8137 ne
rect 17035 8039 17389 8137
tri 17389 8039 17487 8137 sw
tri 17487 8039 17585 8137 ne
rect 17585 8039 17939 8137
tri 17939 8039 18037 8137 sw
tri 18037 8039 18135 8137 ne
rect 18135 8039 18489 8137
tri 18489 8039 18587 8137 sw
tri 18587 8039 18685 8137 ne
rect 18685 8039 19039 8137
tri 19039 8039 19137 8137 sw
tri 19137 8039 19235 8137 ne
rect 19235 8039 19589 8137
tri 19589 8039 19687 8137 sw
rect -500 8035 437 8039
rect -500 7915 215 8035
rect 335 7941 437 8035
tri 437 7941 535 8039 sw
tri 535 7941 633 8039 ne
rect 633 8035 987 8039
rect 633 7941 765 8035
rect 335 7915 535 7941
rect -500 7911 535 7915
tri 535 7911 565 7941 sw
tri 633 7911 663 7941 ne
rect 663 7915 765 7941
rect 885 7941 987 8035
tri 987 7941 1085 8039 sw
tri 1085 7941 1183 8039 ne
rect 1183 8035 1537 8039
rect 1183 7941 1315 8035
rect 885 7915 1085 7941
rect 663 7911 1085 7915
tri 1085 7911 1115 7941 sw
tri 1183 7911 1213 7941 ne
rect 1213 7915 1315 7941
rect 1435 7941 1537 8035
tri 1537 7941 1635 8039 sw
tri 1635 7941 1733 8039 ne
rect 1733 8035 2087 8039
rect 1733 7941 1865 8035
rect 1435 7915 1635 7941
rect 1213 7911 1635 7915
tri 1635 7911 1665 7941 sw
tri 1733 7911 1763 7941 ne
rect 1763 7915 1865 7941
rect 1985 7941 2087 8035
tri 2087 7941 2185 8039 sw
tri 2185 7941 2283 8039 ne
rect 2283 8035 2637 8039
rect 2283 7941 2415 8035
rect 1985 7915 2185 7941
rect 1763 7911 2185 7915
tri 2185 7911 2215 7941 sw
tri 2283 7911 2313 7941 ne
rect 2313 7915 2415 7941
rect 2535 7941 2637 8035
tri 2637 7941 2735 8039 sw
tri 2735 7941 2833 8039 ne
rect 2833 8035 3187 8039
rect 2833 7941 2965 8035
rect 2535 7915 2735 7941
rect 2313 7911 2735 7915
tri 2735 7911 2765 7941 sw
tri 2833 7911 2863 7941 ne
rect 2863 7915 2965 7941
rect 3085 7941 3187 8035
tri 3187 7941 3285 8039 sw
tri 3285 7941 3383 8039 ne
rect 3383 8035 3737 8039
rect 3383 7941 3515 8035
rect 3085 7915 3285 7941
rect 2863 7911 3285 7915
tri 3285 7911 3315 7941 sw
tri 3383 7911 3413 7941 ne
rect 3413 7915 3515 7941
rect 3635 7941 3737 8035
tri 3737 7941 3835 8039 sw
tri 3835 7941 3933 8039 ne
rect 3933 8035 4287 8039
rect 3933 7941 4065 8035
rect 3635 7915 3835 7941
rect 3413 7911 3835 7915
tri 3835 7911 3865 7941 sw
tri 3933 7911 3963 7941 ne
rect 3963 7915 4065 7941
rect 4185 7941 4287 8035
tri 4287 7941 4385 8039 sw
tri 4385 7941 4483 8039 ne
rect 4483 8035 4837 8039
rect 4483 7941 4615 8035
rect 4185 7915 4385 7941
rect 3963 7911 4385 7915
tri 4385 7911 4415 7941 sw
tri 4483 7911 4513 7941 ne
rect 4513 7915 4615 7941
rect 4735 7941 4837 8035
tri 4837 7941 4935 8039 sw
tri 4935 7941 5033 8039 ne
rect 5033 8035 5387 8039
rect 5033 7941 5165 8035
rect 4735 7915 4935 7941
rect 4513 7911 4935 7915
tri 4935 7911 4965 7941 sw
tri 5033 7911 5063 7941 ne
rect 5063 7915 5165 7941
rect 5285 7941 5387 8035
tri 5387 7941 5485 8039 sw
tri 5485 7941 5583 8039 ne
rect 5583 8035 5937 8039
rect 5583 7941 5715 8035
rect 5285 7915 5485 7941
rect 5063 7911 5485 7915
tri 5485 7911 5515 7941 sw
tri 5583 7911 5613 7941 ne
rect 5613 7915 5715 7941
rect 5835 7941 5937 8035
tri 5937 7941 6035 8039 sw
tri 6035 7941 6133 8039 ne
rect 6133 8035 6487 8039
rect 6133 7941 6265 8035
rect 5835 7915 6035 7941
rect 5613 7911 6035 7915
tri 6035 7911 6065 7941 sw
tri 6133 7911 6163 7941 ne
rect 6163 7915 6265 7941
rect 6385 7941 6487 8035
tri 6487 7941 6585 8039 sw
tri 6585 7941 6683 8039 ne
rect 6683 8035 7037 8039
rect 6683 7941 6815 8035
rect 6385 7915 6585 7941
rect 6163 7911 6585 7915
tri 6585 7911 6615 7941 sw
tri 6683 7911 6713 7941 ne
rect 6713 7915 6815 7941
rect 6935 7941 7037 8035
tri 7037 7941 7135 8039 sw
tri 7135 7941 7233 8039 ne
rect 7233 8035 7587 8039
rect 7233 7941 7365 8035
rect 6935 7915 7135 7941
rect 6713 7911 7135 7915
tri 7135 7911 7165 7941 sw
tri 7233 7911 7263 7941 ne
rect 7263 7915 7365 7941
rect 7485 7941 7587 8035
tri 7587 7941 7685 8039 sw
tri 7685 7941 7783 8039 ne
rect 7783 8035 8137 8039
rect 7783 7941 7915 8035
rect 7485 7915 7685 7941
rect 7263 7911 7685 7915
tri 7685 7911 7715 7941 sw
tri 7783 7911 7813 7941 ne
rect 7813 7915 7915 7941
rect 8035 7941 8137 8035
tri 8137 7941 8235 8039 sw
tri 8235 7941 8333 8039 ne
rect 8333 8035 8687 8039
rect 8333 7941 8465 8035
rect 8035 7915 8235 7941
rect 7813 7911 8235 7915
tri 8235 7911 8265 7941 sw
tri 8333 7911 8363 7941 ne
rect 8363 7915 8465 7941
rect 8585 7941 8687 8035
tri 8687 7941 8785 8039 sw
tri 8785 7941 8883 8039 ne
rect 8883 8035 9237 8039
rect 8883 7941 9015 8035
rect 8585 7915 8785 7941
rect 8363 7911 8785 7915
tri 8785 7911 8815 7941 sw
tri 8883 7911 8913 7941 ne
rect 8913 7915 9015 7941
rect 9135 7941 9237 8035
tri 9237 7941 9335 8039 sw
tri 9335 7941 9433 8039 ne
rect 9433 8035 9787 8039
rect 9433 7941 9565 8035
rect 9135 7915 9335 7941
rect 8913 7911 9335 7915
tri 9335 7911 9365 7941 sw
tri 9433 7911 9463 7941 ne
rect 9463 7915 9565 7941
rect 9685 7941 9787 8035
tri 9787 7941 9885 8039 sw
tri 9885 7941 9983 8039 ne
rect 9983 8035 10337 8039
rect 9983 7941 10115 8035
rect 9685 7915 9885 7941
rect 9463 7911 9885 7915
tri 9885 7911 9915 7941 sw
tri 9983 7911 10013 7941 ne
rect 10013 7915 10115 7941
rect 10235 7941 10337 8035
tri 10337 7941 10435 8039 sw
tri 10435 7941 10533 8039 ne
rect 10533 8035 10887 8039
rect 10533 7941 10665 8035
rect 10235 7915 10435 7941
rect 10013 7911 10435 7915
tri 10435 7911 10465 7941 sw
tri 10533 7911 10563 7941 ne
rect 10563 7915 10665 7941
rect 10785 7941 10887 8035
tri 10887 7941 10985 8039 sw
tri 10985 7941 11083 8039 ne
rect 11083 8035 11437 8039
rect 11083 7941 11215 8035
rect 10785 7915 10985 7941
rect 10563 7911 10985 7915
tri 10985 7911 11015 7941 sw
tri 11083 7911 11113 7941 ne
rect 11113 7915 11215 7941
rect 11335 7941 11437 8035
tri 11437 7941 11535 8039 sw
tri 11535 7941 11633 8039 ne
rect 11633 8035 11987 8039
rect 11633 7941 11765 8035
rect 11335 7915 11535 7941
rect 11113 7911 11535 7915
tri 11535 7911 11565 7941 sw
tri 11633 7911 11663 7941 ne
rect 11663 7915 11765 7941
rect 11885 7941 11987 8035
tri 11987 7941 12085 8039 sw
tri 12085 7941 12183 8039 ne
rect 12183 8035 12537 8039
rect 12183 7941 12315 8035
rect 11885 7915 12085 7941
rect 11663 7911 12085 7915
tri 12085 7911 12115 7941 sw
tri 12183 7911 12213 7941 ne
rect 12213 7915 12315 7941
rect 12435 7941 12537 8035
tri 12537 7941 12635 8039 sw
tri 12635 7941 12733 8039 ne
rect 12733 8035 13087 8039
rect 12733 7941 12865 8035
rect 12435 7915 12635 7941
rect 12213 7911 12635 7915
tri 12635 7911 12665 7941 sw
tri 12733 7911 12763 7941 ne
rect 12763 7915 12865 7941
rect 12985 7941 13087 8035
tri 13087 7941 13185 8039 sw
tri 13185 7941 13283 8039 ne
rect 13283 8035 13637 8039
rect 13283 7941 13415 8035
rect 12985 7915 13185 7941
rect 12763 7911 13185 7915
tri 13185 7911 13215 7941 sw
tri 13283 7911 13313 7941 ne
rect 13313 7915 13415 7941
rect 13535 7941 13637 8035
tri 13637 7941 13735 8039 sw
tri 13735 7941 13833 8039 ne
rect 13833 8035 14187 8039
rect 13833 7941 13965 8035
rect 13535 7915 13735 7941
rect 13313 7911 13735 7915
tri 13735 7911 13765 7941 sw
tri 13833 7911 13863 7941 ne
rect 13863 7915 13965 7941
rect 14085 7941 14187 8035
tri 14187 7941 14285 8039 sw
tri 14285 7941 14383 8039 ne
rect 14383 8035 14737 8039
rect 14383 7941 14515 8035
rect 14085 7915 14285 7941
rect 13863 7911 14285 7915
tri 14285 7911 14315 7941 sw
tri 14383 7911 14413 7941 ne
rect 14413 7915 14515 7941
rect 14635 7941 14737 8035
tri 14737 7941 14835 8039 sw
tri 14835 7941 14933 8039 ne
rect 14933 8035 15287 8039
rect 14933 7941 15065 8035
rect 14635 7915 14835 7941
rect 14413 7911 14835 7915
tri 14835 7911 14865 7941 sw
tri 14933 7911 14963 7941 ne
rect 14963 7915 15065 7941
rect 15185 7941 15287 8035
tri 15287 7941 15385 8039 sw
tri 15385 7941 15483 8039 ne
rect 15483 8035 15837 8039
rect 15483 7941 15615 8035
rect 15185 7915 15385 7941
rect 14963 7911 15385 7915
tri 15385 7911 15415 7941 sw
tri 15483 7911 15513 7941 ne
rect 15513 7915 15615 7941
rect 15735 7941 15837 8035
tri 15837 7941 15935 8039 sw
tri 15935 7941 16033 8039 ne
rect 16033 8035 16387 8039
rect 16033 7941 16165 8035
rect 15735 7915 15935 7941
rect 15513 7911 15935 7915
tri 15935 7911 15965 7941 sw
tri 16033 7911 16063 7941 ne
rect 16063 7915 16165 7941
rect 16285 7941 16387 8035
tri 16387 7941 16485 8039 sw
tri 16485 7941 16583 8039 ne
rect 16583 8035 16937 8039
rect 16583 7941 16715 8035
rect 16285 7915 16485 7941
rect 16063 7911 16485 7915
tri 16485 7911 16515 7941 sw
tri 16583 7911 16613 7941 ne
rect 16613 7915 16715 7941
rect 16835 7941 16937 8035
tri 16937 7941 17035 8039 sw
tri 17035 7941 17133 8039 ne
rect 17133 8035 17487 8039
rect 17133 7941 17265 8035
rect 16835 7915 17035 7941
rect 16613 7911 17035 7915
tri 17035 7911 17065 7941 sw
tri 17133 7911 17163 7941 ne
rect 17163 7915 17265 7941
rect 17385 7941 17487 8035
tri 17487 7941 17585 8039 sw
tri 17585 7941 17683 8039 ne
rect 17683 8035 18037 8039
rect 17683 7941 17815 8035
rect 17385 7915 17585 7941
rect 17163 7911 17585 7915
tri 17585 7911 17615 7941 sw
tri 17683 7911 17713 7941 ne
rect 17713 7915 17815 7941
rect 17935 7941 18037 8035
tri 18037 7941 18135 8039 sw
tri 18135 7941 18233 8039 ne
rect 18233 8035 18587 8039
rect 18233 7941 18365 8035
rect 17935 7915 18135 7941
rect 17713 7911 18135 7915
tri 18135 7911 18165 7941 sw
tri 18233 7911 18263 7941 ne
rect 18263 7915 18365 7941
rect 18485 7941 18587 8035
tri 18587 7941 18685 8039 sw
tri 18685 7941 18783 8039 ne
rect 18783 8035 19137 8039
rect 18783 7941 18915 8035
rect 18485 7915 18685 7941
rect 18263 7911 18685 7915
tri 18685 7911 18715 7941 sw
tri 18783 7911 18813 7941 ne
rect 18813 7915 18915 7941
rect 19035 7941 19137 8035
tri 19137 7941 19235 8039 sw
tri 19235 7941 19333 8039 ne
rect 19333 8035 20300 8039
rect 19333 7941 19465 8035
rect 19035 7915 19235 7941
rect 18813 7911 19235 7915
tri 19235 7911 19265 7941 sw
tri 19333 7911 19363 7941 ne
rect 19363 7915 19465 7941
rect 19585 7915 20300 8035
rect 19363 7911 20300 7915
tri 113 7813 211 7911 ne
rect 211 7813 565 7911
tri 565 7813 663 7911 sw
tri 663 7813 761 7911 ne
rect 761 7813 1115 7911
tri 1115 7813 1213 7911 sw
tri 1213 7813 1311 7911 ne
rect 1311 7813 1665 7911
tri 1665 7813 1763 7911 sw
tri 1763 7813 1861 7911 ne
rect 1861 7813 2215 7911
tri 2215 7813 2313 7911 sw
tri 2313 7813 2411 7911 ne
rect 2411 7813 2765 7911
tri 2765 7813 2863 7911 sw
tri 2863 7813 2961 7911 ne
rect 2961 7813 3315 7911
tri 3315 7813 3413 7911 sw
tri 3413 7813 3511 7911 ne
rect 3511 7813 3865 7911
tri 3865 7813 3963 7911 sw
tri 3963 7813 4061 7911 ne
rect 4061 7813 4415 7911
tri 4415 7813 4513 7911 sw
tri 4513 7813 4611 7911 ne
rect 4611 7813 4965 7911
tri 4965 7813 5063 7911 sw
tri 5063 7813 5161 7911 ne
rect 5161 7813 5515 7911
tri 5515 7813 5613 7911 sw
tri 5613 7813 5711 7911 ne
rect 5711 7813 6065 7911
tri 6065 7813 6163 7911 sw
tri 6163 7813 6261 7911 ne
rect 6261 7813 6615 7911
tri 6615 7813 6713 7911 sw
tri 6713 7813 6811 7911 ne
rect 6811 7813 7165 7911
tri 7165 7813 7263 7911 sw
tri 7263 7813 7361 7911 ne
rect 7361 7813 7715 7911
tri 7715 7813 7813 7911 sw
tri 7813 7813 7911 7911 ne
rect 7911 7813 8265 7911
tri 8265 7813 8363 7911 sw
tri 8363 7813 8461 7911 ne
rect 8461 7813 8815 7911
tri 8815 7813 8913 7911 sw
tri 8913 7813 9011 7911 ne
rect 9011 7813 9365 7911
tri 9365 7813 9463 7911 sw
tri 9463 7813 9561 7911 ne
rect 9561 7813 9915 7911
tri 9915 7813 10013 7911 sw
tri 10013 7813 10111 7911 ne
rect 10111 7813 10465 7911
tri 10465 7813 10563 7911 sw
tri 10563 7813 10661 7911 ne
rect 10661 7813 11015 7911
tri 11015 7813 11113 7911 sw
tri 11113 7813 11211 7911 ne
rect 11211 7813 11565 7911
tri 11565 7813 11663 7911 sw
tri 11663 7813 11761 7911 ne
rect 11761 7813 12115 7911
tri 12115 7813 12213 7911 sw
tri 12213 7813 12311 7911 ne
rect 12311 7813 12665 7911
tri 12665 7813 12763 7911 sw
tri 12763 7813 12861 7911 ne
rect 12861 7813 13215 7911
tri 13215 7813 13313 7911 sw
tri 13313 7813 13411 7911 ne
rect 13411 7813 13765 7911
tri 13765 7813 13863 7911 sw
tri 13863 7813 13961 7911 ne
rect 13961 7813 14315 7911
tri 14315 7813 14413 7911 sw
tri 14413 7813 14511 7911 ne
rect 14511 7813 14865 7911
tri 14865 7813 14963 7911 sw
tri 14963 7813 15061 7911 ne
rect 15061 7813 15415 7911
tri 15415 7813 15513 7911 sw
tri 15513 7813 15611 7911 ne
rect 15611 7813 15965 7911
tri 15965 7813 16063 7911 sw
tri 16063 7813 16161 7911 ne
rect 16161 7813 16515 7911
tri 16515 7813 16613 7911 sw
tri 16613 7813 16711 7911 ne
rect 16711 7813 17065 7911
tri 17065 7813 17163 7911 sw
tri 17163 7813 17261 7911 ne
rect 17261 7813 17615 7911
tri 17615 7813 17713 7911 sw
tri 17713 7813 17811 7911 ne
rect 17811 7813 18165 7911
tri 18165 7813 18263 7911 sw
tri 18263 7813 18361 7911 ne
rect 18361 7813 18715 7911
tri 18715 7813 18813 7911 sw
tri 18813 7813 18911 7911 ne
rect 18911 7813 19265 7911
tri 19265 7813 19363 7911 sw
tri 19363 7813 19461 7911 ne
rect 19461 7813 20300 7911
rect -2000 7783 113 7813
tri 113 7783 143 7813 sw
tri 211 7783 241 7813 ne
rect 241 7783 663 7813
tri 663 7783 693 7813 sw
tri 761 7783 791 7813 ne
rect 791 7783 1213 7813
tri 1213 7783 1243 7813 sw
tri 1311 7783 1341 7813 ne
rect 1341 7783 1763 7813
tri 1763 7783 1793 7813 sw
tri 1861 7783 1891 7813 ne
rect 1891 7783 2313 7813
tri 2313 7783 2343 7813 sw
tri 2411 7783 2441 7813 ne
rect 2441 7783 2863 7813
tri 2863 7783 2893 7813 sw
tri 2961 7783 2991 7813 ne
rect 2991 7783 3413 7813
tri 3413 7783 3443 7813 sw
tri 3511 7783 3541 7813 ne
rect 3541 7783 3963 7813
tri 3963 7783 3993 7813 sw
tri 4061 7783 4091 7813 ne
rect 4091 7783 4513 7813
tri 4513 7783 4543 7813 sw
tri 4611 7783 4641 7813 ne
rect 4641 7783 5063 7813
tri 5063 7783 5093 7813 sw
tri 5161 7783 5191 7813 ne
rect 5191 7783 5613 7813
tri 5613 7783 5643 7813 sw
tri 5711 7783 5741 7813 ne
rect 5741 7783 6163 7813
tri 6163 7783 6193 7813 sw
tri 6261 7783 6291 7813 ne
rect 6291 7783 6713 7813
tri 6713 7783 6743 7813 sw
tri 6811 7783 6841 7813 ne
rect 6841 7783 7263 7813
tri 7263 7783 7293 7813 sw
tri 7361 7783 7391 7813 ne
rect 7391 7783 7813 7813
tri 7813 7783 7843 7813 sw
tri 7911 7783 7941 7813 ne
rect 7941 7783 8363 7813
tri 8363 7783 8393 7813 sw
tri 8461 7783 8491 7813 ne
rect 8491 7783 8913 7813
tri 8913 7783 8943 7813 sw
tri 9011 7783 9041 7813 ne
rect 9041 7783 9463 7813
tri 9463 7783 9493 7813 sw
tri 9561 7783 9591 7813 ne
rect 9591 7783 10013 7813
tri 10013 7783 10043 7813 sw
tri 10111 7783 10141 7813 ne
rect 10141 7783 10563 7813
tri 10563 7783 10593 7813 sw
tri 10661 7783 10691 7813 ne
rect 10691 7783 11113 7813
tri 11113 7783 11143 7813 sw
tri 11211 7783 11241 7813 ne
rect 11241 7783 11663 7813
tri 11663 7783 11693 7813 sw
tri 11761 7783 11791 7813 ne
rect 11791 7783 12213 7813
tri 12213 7783 12243 7813 sw
tri 12311 7783 12341 7813 ne
rect 12341 7783 12763 7813
tri 12763 7783 12793 7813 sw
tri 12861 7783 12891 7813 ne
rect 12891 7783 13313 7813
tri 13313 7783 13343 7813 sw
tri 13411 7783 13441 7813 ne
rect 13441 7783 13863 7813
tri 13863 7783 13893 7813 sw
tri 13961 7783 13991 7813 ne
rect 13991 7783 14413 7813
tri 14413 7783 14443 7813 sw
tri 14511 7783 14541 7813 ne
rect 14541 7783 14963 7813
tri 14963 7783 14993 7813 sw
tri 15061 7783 15091 7813 ne
rect 15091 7783 15513 7813
tri 15513 7783 15543 7813 sw
tri 15611 7783 15641 7813 ne
rect 15641 7783 16063 7813
tri 16063 7783 16093 7813 sw
tri 16161 7783 16191 7813 ne
rect 16191 7783 16613 7813
tri 16613 7783 16643 7813 sw
tri 16711 7783 16741 7813 ne
rect 16741 7783 17163 7813
tri 17163 7783 17193 7813 sw
tri 17261 7783 17291 7813 ne
rect 17291 7783 17713 7813
tri 17713 7783 17743 7813 sw
tri 17811 7783 17841 7813 ne
rect 17841 7783 18263 7813
tri 18263 7783 18293 7813 sw
tri 18361 7783 18391 7813 ne
rect 18391 7783 18813 7813
tri 18813 7783 18843 7813 sw
tri 18911 7783 18941 7813 ne
rect 18941 7783 19363 7813
tri 19363 7783 19393 7813 sw
tri 19461 7783 19491 7813 ne
rect 19491 7783 20300 7813
rect -2000 7685 143 7783
tri 143 7685 241 7783 sw
tri 241 7685 339 7783 ne
rect 339 7685 693 7783
tri 693 7685 791 7783 sw
tri 791 7685 889 7783 ne
rect 889 7685 1243 7783
tri 1243 7685 1341 7783 sw
tri 1341 7685 1439 7783 ne
rect 1439 7685 1793 7783
tri 1793 7685 1891 7783 sw
tri 1891 7685 1989 7783 ne
rect 1989 7685 2343 7783
tri 2343 7685 2441 7783 sw
tri 2441 7685 2539 7783 ne
rect 2539 7685 2893 7783
tri 2893 7685 2991 7783 sw
tri 2991 7685 3089 7783 ne
rect 3089 7685 3443 7783
tri 3443 7685 3541 7783 sw
tri 3541 7685 3639 7783 ne
rect 3639 7685 3993 7783
tri 3993 7685 4091 7783 sw
tri 4091 7685 4189 7783 ne
rect 4189 7685 4543 7783
tri 4543 7685 4641 7783 sw
tri 4641 7685 4739 7783 ne
rect 4739 7685 5093 7783
tri 5093 7685 5191 7783 sw
tri 5191 7685 5289 7783 ne
rect 5289 7685 5643 7783
tri 5643 7685 5741 7783 sw
tri 5741 7685 5839 7783 ne
rect 5839 7685 6193 7783
tri 6193 7685 6291 7783 sw
tri 6291 7685 6389 7783 ne
rect 6389 7685 6743 7783
tri 6743 7685 6841 7783 sw
tri 6841 7685 6939 7783 ne
rect 6939 7685 7293 7783
tri 7293 7685 7391 7783 sw
tri 7391 7685 7489 7783 ne
rect 7489 7685 7843 7783
tri 7843 7685 7941 7783 sw
tri 7941 7685 8039 7783 ne
rect 8039 7685 8393 7783
tri 8393 7685 8491 7783 sw
tri 8491 7685 8589 7783 ne
rect 8589 7685 8943 7783
tri 8943 7685 9041 7783 sw
tri 9041 7685 9139 7783 ne
rect 9139 7685 9493 7783
tri 9493 7685 9591 7783 sw
tri 9591 7685 9689 7783 ne
rect 9689 7685 10043 7783
tri 10043 7685 10141 7783 sw
tri 10141 7685 10239 7783 ne
rect 10239 7685 10593 7783
tri 10593 7685 10691 7783 sw
tri 10691 7685 10789 7783 ne
rect 10789 7685 11143 7783
tri 11143 7685 11241 7783 sw
tri 11241 7685 11339 7783 ne
rect 11339 7685 11693 7783
tri 11693 7685 11791 7783 sw
tri 11791 7685 11889 7783 ne
rect 11889 7685 12243 7783
tri 12243 7685 12341 7783 sw
tri 12341 7685 12439 7783 ne
rect 12439 7685 12793 7783
tri 12793 7685 12891 7783 sw
tri 12891 7685 12989 7783 ne
rect 12989 7685 13343 7783
tri 13343 7685 13441 7783 sw
tri 13441 7685 13539 7783 ne
rect 13539 7685 13893 7783
tri 13893 7685 13991 7783 sw
tri 13991 7685 14089 7783 ne
rect 14089 7685 14443 7783
tri 14443 7685 14541 7783 sw
tri 14541 7685 14639 7783 ne
rect 14639 7685 14993 7783
tri 14993 7685 15091 7783 sw
tri 15091 7685 15189 7783 ne
rect 15189 7685 15543 7783
tri 15543 7685 15641 7783 sw
tri 15641 7685 15739 7783 ne
rect 15739 7685 16093 7783
tri 16093 7685 16191 7783 sw
tri 16191 7685 16289 7783 ne
rect 16289 7685 16643 7783
tri 16643 7685 16741 7783 sw
tri 16741 7685 16839 7783 ne
rect 16839 7685 17193 7783
tri 17193 7685 17291 7783 sw
tri 17291 7685 17389 7783 ne
rect 17389 7685 17743 7783
tri 17743 7685 17841 7783 sw
tri 17841 7685 17939 7783 ne
rect 17939 7685 18293 7783
tri 18293 7685 18391 7783 sw
tri 18391 7685 18489 7783 ne
rect 18489 7685 18843 7783
tri 18843 7685 18941 7783 sw
tri 18941 7685 19039 7783 ne
rect 19039 7685 19393 7783
tri 19393 7685 19491 7783 sw
tri 19491 7685 19589 7783 ne
rect 19589 7685 20300 7783
rect -2000 7587 241 7685
tri 241 7587 339 7685 sw
tri 339 7587 437 7685 ne
rect 437 7587 791 7685
tri 791 7587 889 7685 sw
tri 889 7587 987 7685 ne
rect 987 7587 1341 7685
tri 1341 7587 1439 7685 sw
tri 1439 7587 1537 7685 ne
rect 1537 7587 1891 7685
tri 1891 7587 1989 7685 sw
tri 1989 7587 2087 7685 ne
rect 2087 7587 2441 7685
tri 2441 7587 2539 7685 sw
tri 2539 7587 2637 7685 ne
rect 2637 7587 2991 7685
tri 2991 7587 3089 7685 sw
tri 3089 7587 3187 7685 ne
rect 3187 7587 3541 7685
tri 3541 7587 3639 7685 sw
tri 3639 7587 3737 7685 ne
rect 3737 7587 4091 7685
tri 4091 7587 4189 7685 sw
tri 4189 7587 4287 7685 ne
rect 4287 7587 4641 7685
tri 4641 7587 4739 7685 sw
tri 4739 7587 4837 7685 ne
rect 4837 7587 5191 7685
tri 5191 7587 5289 7685 sw
tri 5289 7587 5387 7685 ne
rect 5387 7587 5741 7685
tri 5741 7587 5839 7685 sw
tri 5839 7587 5937 7685 ne
rect 5937 7587 6291 7685
tri 6291 7587 6389 7685 sw
tri 6389 7587 6487 7685 ne
rect 6487 7587 6841 7685
tri 6841 7587 6939 7685 sw
tri 6939 7587 7037 7685 ne
rect 7037 7587 7391 7685
tri 7391 7587 7489 7685 sw
tri 7489 7587 7587 7685 ne
rect 7587 7587 7941 7685
tri 7941 7587 8039 7685 sw
tri 8039 7587 8137 7685 ne
rect 8137 7587 8491 7685
tri 8491 7587 8589 7685 sw
tri 8589 7587 8687 7685 ne
rect 8687 7587 9041 7685
tri 9041 7587 9139 7685 sw
tri 9139 7587 9237 7685 ne
rect 9237 7587 9591 7685
tri 9591 7587 9689 7685 sw
tri 9689 7587 9787 7685 ne
rect 9787 7587 10141 7685
tri 10141 7587 10239 7685 sw
tri 10239 7587 10337 7685 ne
rect 10337 7587 10691 7685
tri 10691 7587 10789 7685 sw
tri 10789 7587 10887 7685 ne
rect 10887 7587 11241 7685
tri 11241 7587 11339 7685 sw
tri 11339 7587 11437 7685 ne
rect 11437 7587 11791 7685
tri 11791 7587 11889 7685 sw
tri 11889 7587 11987 7685 ne
rect 11987 7587 12341 7685
tri 12341 7587 12439 7685 sw
tri 12439 7587 12537 7685 ne
rect 12537 7587 12891 7685
tri 12891 7587 12989 7685 sw
tri 12989 7587 13087 7685 ne
rect 13087 7587 13441 7685
tri 13441 7587 13539 7685 sw
tri 13539 7587 13637 7685 ne
rect 13637 7587 13991 7685
tri 13991 7587 14089 7685 sw
tri 14089 7587 14187 7685 ne
rect 14187 7587 14541 7685
tri 14541 7587 14639 7685 sw
tri 14639 7587 14737 7685 ne
rect 14737 7587 15091 7685
tri 15091 7587 15189 7685 sw
tri 15189 7587 15287 7685 ne
rect 15287 7587 15641 7685
tri 15641 7587 15739 7685 sw
tri 15739 7587 15837 7685 ne
rect 15837 7587 16191 7685
tri 16191 7587 16289 7685 sw
tri 16289 7587 16387 7685 ne
rect 16387 7587 16741 7685
tri 16741 7587 16839 7685 sw
tri 16839 7587 16937 7685 ne
rect 16937 7587 17291 7685
tri 17291 7587 17389 7685 sw
tri 17389 7587 17487 7685 ne
rect 17487 7587 17841 7685
tri 17841 7587 17939 7685 sw
tri 17939 7587 18037 7685 ne
rect 18037 7587 18391 7685
tri 18391 7587 18489 7685 sw
tri 18489 7587 18587 7685 ne
rect 18587 7587 18941 7685
tri 18941 7587 19039 7685 sw
tri 19039 7587 19137 7685 ne
rect 19137 7587 19491 7685
tri 19491 7587 19589 7685 sw
tri 19589 7587 19687 7685 ne
rect 19687 7587 20300 7685
rect -2000 7489 339 7587
tri 339 7489 437 7587 sw
tri 437 7489 535 7587 ne
rect 535 7489 889 7587
tri 889 7489 987 7587 sw
tri 987 7489 1085 7587 ne
rect 1085 7489 1439 7587
tri 1439 7489 1537 7587 sw
tri 1537 7489 1635 7587 ne
rect 1635 7489 1989 7587
tri 1989 7489 2087 7587 sw
tri 2087 7489 2185 7587 ne
rect 2185 7489 2539 7587
tri 2539 7489 2637 7587 sw
tri 2637 7489 2735 7587 ne
rect 2735 7489 3089 7587
tri 3089 7489 3187 7587 sw
tri 3187 7489 3285 7587 ne
rect 3285 7489 3639 7587
tri 3639 7489 3737 7587 sw
tri 3737 7489 3835 7587 ne
rect 3835 7489 4189 7587
tri 4189 7489 4287 7587 sw
tri 4287 7489 4385 7587 ne
rect 4385 7489 4739 7587
tri 4739 7489 4837 7587 sw
tri 4837 7489 4935 7587 ne
rect 4935 7489 5289 7587
tri 5289 7489 5387 7587 sw
tri 5387 7489 5485 7587 ne
rect 5485 7489 5839 7587
tri 5839 7489 5937 7587 sw
tri 5937 7489 6035 7587 ne
rect 6035 7489 6389 7587
tri 6389 7489 6487 7587 sw
tri 6487 7489 6585 7587 ne
rect 6585 7489 6939 7587
tri 6939 7489 7037 7587 sw
tri 7037 7489 7135 7587 ne
rect 7135 7489 7489 7587
tri 7489 7489 7587 7587 sw
tri 7587 7489 7685 7587 ne
rect 7685 7489 8039 7587
tri 8039 7489 8137 7587 sw
tri 8137 7489 8235 7587 ne
rect 8235 7489 8589 7587
tri 8589 7489 8687 7587 sw
tri 8687 7489 8785 7587 ne
rect 8785 7489 9139 7587
tri 9139 7489 9237 7587 sw
tri 9237 7489 9335 7587 ne
rect 9335 7489 9689 7587
tri 9689 7489 9787 7587 sw
tri 9787 7489 9885 7587 ne
rect 9885 7489 10239 7587
tri 10239 7489 10337 7587 sw
tri 10337 7489 10435 7587 ne
rect 10435 7489 10789 7587
tri 10789 7489 10887 7587 sw
tri 10887 7489 10985 7587 ne
rect 10985 7489 11339 7587
tri 11339 7489 11437 7587 sw
tri 11437 7489 11535 7587 ne
rect 11535 7489 11889 7587
tri 11889 7489 11987 7587 sw
tri 11987 7489 12085 7587 ne
rect 12085 7489 12439 7587
tri 12439 7489 12537 7587 sw
tri 12537 7489 12635 7587 ne
rect 12635 7489 12989 7587
tri 12989 7489 13087 7587 sw
tri 13087 7489 13185 7587 ne
rect 13185 7489 13539 7587
tri 13539 7489 13637 7587 sw
tri 13637 7489 13735 7587 ne
rect 13735 7489 14089 7587
tri 14089 7489 14187 7587 sw
tri 14187 7489 14285 7587 ne
rect 14285 7489 14639 7587
tri 14639 7489 14737 7587 sw
tri 14737 7489 14835 7587 ne
rect 14835 7489 15189 7587
tri 15189 7489 15287 7587 sw
tri 15287 7489 15385 7587 ne
rect 15385 7489 15739 7587
tri 15739 7489 15837 7587 sw
tri 15837 7489 15935 7587 ne
rect 15935 7489 16289 7587
tri 16289 7489 16387 7587 sw
tri 16387 7489 16485 7587 ne
rect 16485 7489 16839 7587
tri 16839 7489 16937 7587 sw
tri 16937 7489 17035 7587 ne
rect 17035 7489 17389 7587
tri 17389 7489 17487 7587 sw
tri 17487 7489 17585 7587 ne
rect 17585 7489 17939 7587
tri 17939 7489 18037 7587 sw
tri 18037 7489 18135 7587 ne
rect 18135 7489 18489 7587
tri 18489 7489 18587 7587 sw
tri 18587 7489 18685 7587 ne
rect 18685 7489 19039 7587
tri 19039 7489 19137 7587 sw
tri 19137 7489 19235 7587 ne
rect 19235 7489 19589 7587
tri 19589 7489 19687 7587 sw
rect 20800 7489 21800 8137
rect -2000 7485 437 7489
rect -2000 7365 215 7485
rect 335 7391 437 7485
tri 437 7391 535 7489 sw
tri 535 7391 633 7489 ne
rect 633 7485 987 7489
rect 633 7391 765 7485
rect 335 7365 535 7391
rect -2000 7361 535 7365
rect -2000 6713 -1000 7361
tri 113 7263 211 7361 ne
rect 211 7313 535 7361
tri 535 7313 613 7391 sw
tri 633 7313 711 7391 ne
rect 711 7365 765 7391
rect 885 7391 987 7485
tri 987 7391 1085 7489 sw
tri 1085 7391 1183 7489 ne
rect 1183 7485 1537 7489
rect 1183 7391 1315 7485
rect 885 7365 1085 7391
rect 711 7313 1085 7365
tri 1085 7313 1163 7391 sw
tri 1183 7313 1261 7391 ne
rect 1261 7365 1315 7391
rect 1435 7391 1537 7485
tri 1537 7391 1635 7489 sw
tri 1635 7391 1733 7489 ne
rect 1733 7485 2087 7489
rect 1733 7391 1865 7485
rect 1435 7365 1635 7391
rect 1261 7313 1635 7365
tri 1635 7313 1713 7391 sw
tri 1733 7313 1811 7391 ne
rect 1811 7365 1865 7391
rect 1985 7391 2087 7485
tri 2087 7391 2185 7489 sw
tri 2185 7391 2283 7489 ne
rect 2283 7485 2637 7489
rect 2283 7391 2415 7485
rect 1985 7365 2185 7391
rect 1811 7313 2185 7365
tri 2185 7313 2263 7391 sw
tri 2283 7313 2361 7391 ne
rect 2361 7365 2415 7391
rect 2535 7391 2637 7485
tri 2637 7391 2735 7489 sw
tri 2735 7391 2833 7489 ne
rect 2833 7485 3187 7489
rect 2833 7391 2965 7485
rect 2535 7365 2735 7391
rect 2361 7313 2735 7365
tri 2735 7313 2813 7391 sw
tri 2833 7313 2911 7391 ne
rect 2911 7365 2965 7391
rect 3085 7391 3187 7485
tri 3187 7391 3285 7489 sw
tri 3285 7391 3383 7489 ne
rect 3383 7485 3737 7489
rect 3383 7391 3515 7485
rect 3085 7365 3285 7391
rect 2911 7313 3285 7365
tri 3285 7313 3363 7391 sw
tri 3383 7313 3461 7391 ne
rect 3461 7365 3515 7391
rect 3635 7391 3737 7485
tri 3737 7391 3835 7489 sw
tri 3835 7391 3933 7489 ne
rect 3933 7485 4287 7489
rect 3933 7391 4065 7485
rect 3635 7365 3835 7391
rect 3461 7313 3835 7365
tri 3835 7313 3913 7391 sw
tri 3933 7313 4011 7391 ne
rect 4011 7365 4065 7391
rect 4185 7391 4287 7485
tri 4287 7391 4385 7489 sw
tri 4385 7391 4483 7489 ne
rect 4483 7485 4837 7489
rect 4483 7391 4615 7485
rect 4185 7365 4385 7391
rect 4011 7313 4385 7365
tri 4385 7313 4463 7391 sw
tri 4483 7313 4561 7391 ne
rect 4561 7365 4615 7391
rect 4735 7391 4837 7485
tri 4837 7391 4935 7489 sw
tri 4935 7391 5033 7489 ne
rect 5033 7485 5387 7489
rect 5033 7391 5165 7485
rect 4735 7365 4935 7391
rect 4561 7313 4935 7365
tri 4935 7313 5013 7391 sw
tri 5033 7313 5111 7391 ne
rect 5111 7365 5165 7391
rect 5285 7391 5387 7485
tri 5387 7391 5485 7489 sw
tri 5485 7391 5583 7489 ne
rect 5583 7485 5937 7489
rect 5583 7391 5715 7485
rect 5285 7365 5485 7391
rect 5111 7313 5485 7365
tri 5485 7313 5563 7391 sw
tri 5583 7313 5661 7391 ne
rect 5661 7365 5715 7391
rect 5835 7391 5937 7485
tri 5937 7391 6035 7489 sw
tri 6035 7391 6133 7489 ne
rect 6133 7485 6487 7489
rect 6133 7391 6265 7485
rect 5835 7365 6035 7391
rect 5661 7313 6035 7365
tri 6035 7313 6113 7391 sw
tri 6133 7313 6211 7391 ne
rect 6211 7365 6265 7391
rect 6385 7391 6487 7485
tri 6487 7391 6585 7489 sw
tri 6585 7391 6683 7489 ne
rect 6683 7485 7037 7489
rect 6683 7391 6815 7485
rect 6385 7365 6585 7391
rect 6211 7313 6585 7365
tri 6585 7313 6663 7391 sw
tri 6683 7313 6761 7391 ne
rect 6761 7365 6815 7391
rect 6935 7391 7037 7485
tri 7037 7391 7135 7489 sw
tri 7135 7391 7233 7489 ne
rect 7233 7485 7587 7489
rect 7233 7391 7365 7485
rect 6935 7365 7135 7391
rect 6761 7313 7135 7365
tri 7135 7313 7213 7391 sw
tri 7233 7313 7311 7391 ne
rect 7311 7365 7365 7391
rect 7485 7391 7587 7485
tri 7587 7391 7685 7489 sw
tri 7685 7391 7783 7489 ne
rect 7783 7485 8137 7489
rect 7783 7391 7915 7485
rect 7485 7365 7685 7391
rect 7311 7313 7685 7365
tri 7685 7313 7763 7391 sw
tri 7783 7313 7861 7391 ne
rect 7861 7365 7915 7391
rect 8035 7391 8137 7485
tri 8137 7391 8235 7489 sw
tri 8235 7391 8333 7489 ne
rect 8333 7485 8687 7489
rect 8333 7391 8465 7485
rect 8035 7365 8235 7391
rect 7861 7313 8235 7365
tri 8235 7313 8313 7391 sw
tri 8333 7313 8411 7391 ne
rect 8411 7365 8465 7391
rect 8585 7391 8687 7485
tri 8687 7391 8785 7489 sw
tri 8785 7391 8883 7489 ne
rect 8883 7485 9237 7489
rect 8883 7391 9015 7485
rect 8585 7365 8785 7391
rect 8411 7313 8785 7365
tri 8785 7313 8863 7391 sw
tri 8883 7313 8961 7391 ne
rect 8961 7365 9015 7391
rect 9135 7391 9237 7485
tri 9237 7391 9335 7489 sw
tri 9335 7391 9433 7489 ne
rect 9433 7485 9787 7489
rect 9433 7391 9565 7485
rect 9135 7365 9335 7391
rect 8961 7313 9335 7365
tri 9335 7313 9413 7391 sw
tri 9433 7313 9511 7391 ne
rect 9511 7365 9565 7391
rect 9685 7391 9787 7485
tri 9787 7391 9885 7489 sw
tri 9885 7391 9983 7489 ne
rect 9983 7485 10337 7489
rect 9983 7391 10115 7485
rect 9685 7365 9885 7391
rect 9511 7313 9885 7365
tri 9885 7313 9963 7391 sw
tri 9983 7313 10061 7391 ne
rect 10061 7365 10115 7391
rect 10235 7391 10337 7485
tri 10337 7391 10435 7489 sw
tri 10435 7391 10533 7489 ne
rect 10533 7485 10887 7489
rect 10533 7391 10665 7485
rect 10235 7365 10435 7391
rect 10061 7313 10435 7365
tri 10435 7313 10513 7391 sw
tri 10533 7313 10611 7391 ne
rect 10611 7365 10665 7391
rect 10785 7391 10887 7485
tri 10887 7391 10985 7489 sw
tri 10985 7391 11083 7489 ne
rect 11083 7485 11437 7489
rect 11083 7391 11215 7485
rect 10785 7365 10985 7391
rect 10611 7313 10985 7365
tri 10985 7313 11063 7391 sw
tri 11083 7313 11161 7391 ne
rect 11161 7365 11215 7391
rect 11335 7391 11437 7485
tri 11437 7391 11535 7489 sw
tri 11535 7391 11633 7489 ne
rect 11633 7485 11987 7489
rect 11633 7391 11765 7485
rect 11335 7365 11535 7391
rect 11161 7313 11535 7365
tri 11535 7313 11613 7391 sw
tri 11633 7313 11711 7391 ne
rect 11711 7365 11765 7391
rect 11885 7391 11987 7485
tri 11987 7391 12085 7489 sw
tri 12085 7391 12183 7489 ne
rect 12183 7485 12537 7489
rect 12183 7391 12315 7485
rect 11885 7365 12085 7391
rect 11711 7313 12085 7365
tri 12085 7313 12163 7391 sw
tri 12183 7313 12261 7391 ne
rect 12261 7365 12315 7391
rect 12435 7391 12537 7485
tri 12537 7391 12635 7489 sw
tri 12635 7391 12733 7489 ne
rect 12733 7485 13087 7489
rect 12733 7391 12865 7485
rect 12435 7365 12635 7391
rect 12261 7313 12635 7365
tri 12635 7313 12713 7391 sw
tri 12733 7313 12811 7391 ne
rect 12811 7365 12865 7391
rect 12985 7391 13087 7485
tri 13087 7391 13185 7489 sw
tri 13185 7391 13283 7489 ne
rect 13283 7485 13637 7489
rect 13283 7391 13415 7485
rect 12985 7365 13185 7391
rect 12811 7313 13185 7365
tri 13185 7313 13263 7391 sw
tri 13283 7313 13361 7391 ne
rect 13361 7365 13415 7391
rect 13535 7391 13637 7485
tri 13637 7391 13735 7489 sw
tri 13735 7391 13833 7489 ne
rect 13833 7485 14187 7489
rect 13833 7391 13965 7485
rect 13535 7365 13735 7391
rect 13361 7313 13735 7365
tri 13735 7313 13813 7391 sw
tri 13833 7313 13911 7391 ne
rect 13911 7365 13965 7391
rect 14085 7391 14187 7485
tri 14187 7391 14285 7489 sw
tri 14285 7391 14383 7489 ne
rect 14383 7485 14737 7489
rect 14383 7391 14515 7485
rect 14085 7365 14285 7391
rect 13911 7313 14285 7365
tri 14285 7313 14363 7391 sw
tri 14383 7313 14461 7391 ne
rect 14461 7365 14515 7391
rect 14635 7391 14737 7485
tri 14737 7391 14835 7489 sw
tri 14835 7391 14933 7489 ne
rect 14933 7485 15287 7489
rect 14933 7391 15065 7485
rect 14635 7365 14835 7391
rect 14461 7313 14835 7365
tri 14835 7313 14913 7391 sw
tri 14933 7313 15011 7391 ne
rect 15011 7365 15065 7391
rect 15185 7391 15287 7485
tri 15287 7391 15385 7489 sw
tri 15385 7391 15483 7489 ne
rect 15483 7485 15837 7489
rect 15483 7391 15615 7485
rect 15185 7365 15385 7391
rect 15011 7313 15385 7365
tri 15385 7313 15463 7391 sw
tri 15483 7313 15561 7391 ne
rect 15561 7365 15615 7391
rect 15735 7391 15837 7485
tri 15837 7391 15935 7489 sw
tri 15935 7391 16033 7489 ne
rect 16033 7485 16387 7489
rect 16033 7391 16165 7485
rect 15735 7365 15935 7391
rect 15561 7313 15935 7365
tri 15935 7313 16013 7391 sw
tri 16033 7313 16111 7391 ne
rect 16111 7365 16165 7391
rect 16285 7391 16387 7485
tri 16387 7391 16485 7489 sw
tri 16485 7391 16583 7489 ne
rect 16583 7485 16937 7489
rect 16583 7391 16715 7485
rect 16285 7365 16485 7391
rect 16111 7313 16485 7365
tri 16485 7313 16563 7391 sw
tri 16583 7313 16661 7391 ne
rect 16661 7365 16715 7391
rect 16835 7391 16937 7485
tri 16937 7391 17035 7489 sw
tri 17035 7391 17133 7489 ne
rect 17133 7485 17487 7489
rect 17133 7391 17265 7485
rect 16835 7365 17035 7391
rect 16661 7313 17035 7365
tri 17035 7313 17113 7391 sw
tri 17133 7313 17211 7391 ne
rect 17211 7365 17265 7391
rect 17385 7391 17487 7485
tri 17487 7391 17585 7489 sw
tri 17585 7391 17683 7489 ne
rect 17683 7485 18037 7489
rect 17683 7391 17815 7485
rect 17385 7365 17585 7391
rect 17211 7313 17585 7365
tri 17585 7313 17663 7391 sw
tri 17683 7313 17761 7391 ne
rect 17761 7365 17815 7391
rect 17935 7391 18037 7485
tri 18037 7391 18135 7489 sw
tri 18135 7391 18233 7489 ne
rect 18233 7485 18587 7489
rect 18233 7391 18365 7485
rect 17935 7365 18135 7391
rect 17761 7313 18135 7365
tri 18135 7313 18213 7391 sw
tri 18233 7313 18311 7391 ne
rect 18311 7365 18365 7391
rect 18485 7391 18587 7485
tri 18587 7391 18685 7489 sw
tri 18685 7391 18783 7489 ne
rect 18783 7485 19137 7489
rect 18783 7391 18915 7485
rect 18485 7365 18685 7391
rect 18311 7313 18685 7365
tri 18685 7313 18763 7391 sw
tri 18783 7313 18861 7391 ne
rect 18861 7365 18915 7391
rect 19035 7391 19137 7485
tri 19137 7391 19235 7489 sw
tri 19235 7391 19333 7489 ne
rect 19333 7485 21800 7489
rect 19333 7391 19465 7485
rect 19035 7365 19235 7391
rect 18861 7313 19235 7365
tri 19235 7313 19313 7391 sw
tri 19333 7313 19411 7391 ne
rect 19411 7365 19465 7391
rect 19585 7365 21800 7485
rect 19411 7313 21800 7365
rect 211 7263 613 7313
rect -500 7213 113 7263
tri 113 7213 163 7263 sw
tri 211 7213 261 7263 ne
rect 261 7233 613 7263
tri 613 7233 693 7313 sw
tri 711 7233 791 7313 ne
rect 791 7233 1163 7313
tri 1163 7233 1243 7313 sw
tri 1261 7233 1341 7313 ne
rect 1341 7233 1713 7313
tri 1713 7233 1793 7313 sw
tri 1811 7233 1891 7313 ne
rect 1891 7233 2263 7313
tri 2263 7233 2343 7313 sw
tri 2361 7233 2441 7313 ne
rect 2441 7233 2813 7313
tri 2813 7233 2893 7313 sw
tri 2911 7233 2991 7313 ne
rect 2991 7233 3363 7313
tri 3363 7233 3443 7313 sw
tri 3461 7233 3541 7313 ne
rect 3541 7233 3913 7313
tri 3913 7233 3993 7313 sw
tri 4011 7233 4091 7313 ne
rect 4091 7233 4463 7313
tri 4463 7233 4543 7313 sw
tri 4561 7233 4641 7313 ne
rect 4641 7233 5013 7313
tri 5013 7233 5093 7313 sw
tri 5111 7233 5191 7313 ne
rect 5191 7233 5563 7313
tri 5563 7233 5643 7313 sw
tri 5661 7233 5741 7313 ne
rect 5741 7233 6113 7313
tri 6113 7233 6193 7313 sw
tri 6211 7233 6291 7313 ne
rect 6291 7233 6663 7313
tri 6663 7233 6743 7313 sw
tri 6761 7233 6841 7313 ne
rect 6841 7233 7213 7313
tri 7213 7233 7293 7313 sw
tri 7311 7233 7391 7313 ne
rect 7391 7233 7763 7313
tri 7763 7233 7843 7313 sw
tri 7861 7233 7941 7313 ne
rect 7941 7233 8313 7313
tri 8313 7233 8393 7313 sw
tri 8411 7233 8491 7313 ne
rect 8491 7233 8863 7313
tri 8863 7233 8943 7313 sw
tri 8961 7233 9041 7313 ne
rect 9041 7233 9413 7313
tri 9413 7233 9493 7313 sw
tri 9511 7233 9591 7313 ne
rect 9591 7233 9963 7313
tri 9963 7233 10043 7313 sw
tri 10061 7233 10141 7313 ne
rect 10141 7233 10513 7313
tri 10513 7233 10593 7313 sw
tri 10611 7233 10691 7313 ne
rect 10691 7233 11063 7313
tri 11063 7233 11143 7313 sw
tri 11161 7233 11241 7313 ne
rect 11241 7233 11613 7313
tri 11613 7233 11693 7313 sw
tri 11711 7233 11791 7313 ne
rect 11791 7233 12163 7313
tri 12163 7233 12243 7313 sw
tri 12261 7233 12341 7313 ne
rect 12341 7233 12713 7313
tri 12713 7233 12793 7313 sw
tri 12811 7233 12891 7313 ne
rect 12891 7233 13263 7313
tri 13263 7233 13343 7313 sw
tri 13361 7233 13441 7313 ne
rect 13441 7233 13813 7313
tri 13813 7233 13893 7313 sw
tri 13911 7233 13991 7313 ne
rect 13991 7233 14363 7313
tri 14363 7233 14443 7313 sw
tri 14461 7233 14541 7313 ne
rect 14541 7233 14913 7313
tri 14913 7233 14993 7313 sw
tri 15011 7233 15091 7313 ne
rect 15091 7233 15463 7313
tri 15463 7233 15543 7313 sw
tri 15561 7233 15641 7313 ne
rect 15641 7233 16013 7313
tri 16013 7233 16093 7313 sw
tri 16111 7233 16191 7313 ne
rect 16191 7233 16563 7313
tri 16563 7233 16643 7313 sw
tri 16661 7233 16741 7313 ne
rect 16741 7233 17113 7313
tri 17113 7233 17193 7313 sw
tri 17211 7233 17291 7313 ne
rect 17291 7233 17663 7313
tri 17663 7233 17743 7313 sw
tri 17761 7233 17841 7313 ne
rect 17841 7233 18213 7313
tri 18213 7233 18293 7313 sw
tri 18311 7233 18391 7313 ne
rect 18391 7233 18763 7313
tri 18763 7233 18843 7313 sw
tri 18861 7233 18941 7313 ne
rect 18941 7233 19313 7313
tri 19313 7233 19393 7313 sw
tri 19411 7233 19491 7313 ne
rect 19491 7233 20100 7313
rect 261 7213 693 7233
rect -500 7135 163 7213
tri 163 7135 241 7213 sw
tri 261 7135 339 7213 ne
rect 339 7135 693 7213
tri 693 7135 791 7233 sw
tri 791 7135 889 7233 ne
rect 889 7135 1243 7233
tri 1243 7135 1341 7233 sw
tri 1341 7135 1439 7233 ne
rect 1439 7135 1793 7233
tri 1793 7135 1891 7233 sw
tri 1891 7135 1989 7233 ne
rect 1989 7135 2343 7233
tri 2343 7135 2441 7233 sw
tri 2441 7135 2539 7233 ne
rect 2539 7135 2893 7233
tri 2893 7135 2991 7233 sw
tri 2991 7135 3089 7233 ne
rect 3089 7135 3443 7233
tri 3443 7135 3541 7233 sw
tri 3541 7135 3639 7233 ne
rect 3639 7135 3993 7233
tri 3993 7135 4091 7233 sw
tri 4091 7135 4189 7233 ne
rect 4189 7135 4543 7233
tri 4543 7135 4641 7233 sw
tri 4641 7135 4739 7233 ne
rect 4739 7135 5093 7233
tri 5093 7135 5191 7233 sw
tri 5191 7135 5289 7233 ne
rect 5289 7135 5643 7233
tri 5643 7135 5741 7233 sw
tri 5741 7135 5839 7233 ne
rect 5839 7135 6193 7233
tri 6193 7135 6291 7233 sw
tri 6291 7135 6389 7233 ne
rect 6389 7135 6743 7233
tri 6743 7135 6841 7233 sw
tri 6841 7135 6939 7233 ne
rect 6939 7135 7293 7233
tri 7293 7135 7391 7233 sw
tri 7391 7135 7489 7233 ne
rect 7489 7135 7843 7233
tri 7843 7135 7941 7233 sw
tri 7941 7135 8039 7233 ne
rect 8039 7135 8393 7233
tri 8393 7135 8491 7233 sw
tri 8491 7135 8589 7233 ne
rect 8589 7135 8943 7233
tri 8943 7135 9041 7233 sw
tri 9041 7135 9139 7233 ne
rect 9139 7135 9493 7233
tri 9493 7135 9591 7233 sw
tri 9591 7135 9689 7233 ne
rect 9689 7135 10043 7233
tri 10043 7135 10141 7233 sw
tri 10141 7135 10239 7233 ne
rect 10239 7135 10593 7233
tri 10593 7135 10691 7233 sw
tri 10691 7135 10789 7233 ne
rect 10789 7135 11143 7233
tri 11143 7135 11241 7233 sw
tri 11241 7135 11339 7233 ne
rect 11339 7135 11693 7233
tri 11693 7135 11791 7233 sw
tri 11791 7135 11889 7233 ne
rect 11889 7135 12243 7233
tri 12243 7135 12341 7233 sw
tri 12341 7135 12439 7233 ne
rect 12439 7135 12793 7233
tri 12793 7135 12891 7233 sw
tri 12891 7135 12989 7233 ne
rect 12989 7135 13343 7233
tri 13343 7135 13441 7233 sw
tri 13441 7135 13539 7233 ne
rect 13539 7135 13893 7233
tri 13893 7135 13991 7233 sw
tri 13991 7135 14089 7233 ne
rect 14089 7135 14443 7233
tri 14443 7135 14541 7233 sw
tri 14541 7135 14639 7233 ne
rect 14639 7135 14993 7233
tri 14993 7135 15091 7233 sw
tri 15091 7135 15189 7233 ne
rect 15189 7135 15543 7233
tri 15543 7135 15641 7233 sw
tri 15641 7135 15739 7233 ne
rect 15739 7135 16093 7233
tri 16093 7135 16191 7233 sw
tri 16191 7135 16289 7233 ne
rect 16289 7135 16643 7233
tri 16643 7135 16741 7233 sw
tri 16741 7135 16839 7233 ne
rect 16839 7135 17193 7233
tri 17193 7135 17291 7233 sw
tri 17291 7135 17389 7233 ne
rect 17389 7135 17743 7233
tri 17743 7135 17841 7233 sw
tri 17841 7135 17939 7233 ne
rect 17939 7135 18293 7233
tri 18293 7135 18391 7233 sw
tri 18391 7135 18489 7233 ne
rect 18489 7135 18843 7233
tri 18843 7135 18941 7233 sw
tri 18941 7135 19039 7233 ne
rect 19039 7135 19393 7233
tri 19393 7135 19491 7233 sw
tri 19491 7135 19589 7233 ne
rect 19589 7213 20100 7233
rect 20200 7213 21800 7313
rect 19589 7135 21800 7213
rect -500 7087 241 7135
rect -500 6987 -400 7087
rect -300 7037 241 7087
tri 241 7037 339 7135 sw
tri 339 7037 437 7135 ne
rect 437 7037 791 7135
tri 791 7037 889 7135 sw
tri 889 7037 987 7135 ne
rect 987 7037 1341 7135
tri 1341 7037 1439 7135 sw
tri 1439 7037 1537 7135 ne
rect 1537 7037 1891 7135
tri 1891 7037 1989 7135 sw
tri 1989 7037 2087 7135 ne
rect 2087 7037 2441 7135
tri 2441 7037 2539 7135 sw
tri 2539 7037 2637 7135 ne
rect 2637 7037 2991 7135
tri 2991 7037 3089 7135 sw
tri 3089 7037 3187 7135 ne
rect 3187 7037 3541 7135
tri 3541 7037 3639 7135 sw
tri 3639 7037 3737 7135 ne
rect 3737 7037 4091 7135
tri 4091 7037 4189 7135 sw
tri 4189 7037 4287 7135 ne
rect 4287 7037 4641 7135
tri 4641 7037 4739 7135 sw
tri 4739 7037 4837 7135 ne
rect 4837 7037 5191 7135
tri 5191 7037 5289 7135 sw
tri 5289 7037 5387 7135 ne
rect 5387 7037 5741 7135
tri 5741 7037 5839 7135 sw
tri 5839 7037 5937 7135 ne
rect 5937 7037 6291 7135
tri 6291 7037 6389 7135 sw
tri 6389 7037 6487 7135 ne
rect 6487 7037 6841 7135
tri 6841 7037 6939 7135 sw
tri 6939 7037 7037 7135 ne
rect 7037 7037 7391 7135
tri 7391 7037 7489 7135 sw
tri 7489 7037 7587 7135 ne
rect 7587 7037 7941 7135
tri 7941 7037 8039 7135 sw
tri 8039 7037 8137 7135 ne
rect 8137 7037 8491 7135
tri 8491 7037 8589 7135 sw
tri 8589 7037 8687 7135 ne
rect 8687 7037 9041 7135
tri 9041 7037 9139 7135 sw
tri 9139 7037 9237 7135 ne
rect 9237 7037 9591 7135
tri 9591 7037 9689 7135 sw
tri 9689 7037 9787 7135 ne
rect 9787 7037 10141 7135
tri 10141 7037 10239 7135 sw
tri 10239 7037 10337 7135 ne
rect 10337 7037 10691 7135
tri 10691 7037 10789 7135 sw
tri 10789 7037 10887 7135 ne
rect 10887 7037 11241 7135
tri 11241 7037 11339 7135 sw
tri 11339 7037 11437 7135 ne
rect 11437 7037 11791 7135
tri 11791 7037 11889 7135 sw
tri 11889 7037 11987 7135 ne
rect 11987 7037 12341 7135
tri 12341 7037 12439 7135 sw
tri 12439 7037 12537 7135 ne
rect 12537 7037 12891 7135
tri 12891 7037 12989 7135 sw
tri 12989 7037 13087 7135 ne
rect 13087 7037 13441 7135
tri 13441 7037 13539 7135 sw
tri 13539 7037 13637 7135 ne
rect 13637 7037 13991 7135
tri 13991 7037 14089 7135 sw
tri 14089 7037 14187 7135 ne
rect 14187 7037 14541 7135
tri 14541 7037 14639 7135 sw
tri 14639 7037 14737 7135 ne
rect 14737 7037 15091 7135
tri 15091 7037 15189 7135 sw
tri 15189 7037 15287 7135 ne
rect 15287 7037 15641 7135
tri 15641 7037 15739 7135 sw
tri 15739 7037 15837 7135 ne
rect 15837 7037 16191 7135
tri 16191 7037 16289 7135 sw
tri 16289 7037 16387 7135 ne
rect 16387 7037 16741 7135
tri 16741 7037 16839 7135 sw
tri 16839 7037 16937 7135 ne
rect 16937 7037 17291 7135
tri 17291 7037 17389 7135 sw
tri 17389 7037 17487 7135 ne
rect 17487 7037 17841 7135
tri 17841 7037 17939 7135 sw
tri 17939 7037 18037 7135 ne
rect 18037 7037 18391 7135
tri 18391 7037 18489 7135 sw
tri 18489 7037 18587 7135 ne
rect 18587 7037 18941 7135
tri 18941 7037 19039 7135 sw
tri 19039 7037 19137 7135 ne
rect 19137 7037 19491 7135
tri 19491 7037 19589 7135 sw
tri 19589 7037 19687 7135 ne
rect 19687 7037 21800 7135
rect -300 6987 339 7037
rect -500 6939 339 6987
tri 339 6939 437 7037 sw
tri 437 6939 535 7037 ne
rect 535 6939 889 7037
tri 889 6939 987 7037 sw
tri 987 6939 1085 7037 ne
rect 1085 6939 1439 7037
tri 1439 6939 1537 7037 sw
tri 1537 6939 1635 7037 ne
rect 1635 6939 1989 7037
tri 1989 6939 2087 7037 sw
tri 2087 6939 2185 7037 ne
rect 2185 6939 2539 7037
tri 2539 6939 2637 7037 sw
tri 2637 6939 2735 7037 ne
rect 2735 6939 3089 7037
tri 3089 6939 3187 7037 sw
tri 3187 6939 3285 7037 ne
rect 3285 6939 3639 7037
tri 3639 6939 3737 7037 sw
tri 3737 6939 3835 7037 ne
rect 3835 6939 4189 7037
tri 4189 6939 4287 7037 sw
tri 4287 6939 4385 7037 ne
rect 4385 6939 4739 7037
tri 4739 6939 4837 7037 sw
tri 4837 6939 4935 7037 ne
rect 4935 6939 5289 7037
tri 5289 6939 5387 7037 sw
tri 5387 6939 5485 7037 ne
rect 5485 6939 5839 7037
tri 5839 6939 5937 7037 sw
tri 5937 6939 6035 7037 ne
rect 6035 6939 6389 7037
tri 6389 6939 6487 7037 sw
tri 6487 6939 6585 7037 ne
rect 6585 6939 6939 7037
tri 6939 6939 7037 7037 sw
tri 7037 6939 7135 7037 ne
rect 7135 6939 7489 7037
tri 7489 6939 7587 7037 sw
tri 7587 6939 7685 7037 ne
rect 7685 6939 8039 7037
tri 8039 6939 8137 7037 sw
tri 8137 6939 8235 7037 ne
rect 8235 6939 8589 7037
tri 8589 6939 8687 7037 sw
tri 8687 6939 8785 7037 ne
rect 8785 6939 9139 7037
tri 9139 6939 9237 7037 sw
tri 9237 6939 9335 7037 ne
rect 9335 6939 9689 7037
tri 9689 6939 9787 7037 sw
tri 9787 6939 9885 7037 ne
rect 9885 6939 10239 7037
tri 10239 6939 10337 7037 sw
tri 10337 6939 10435 7037 ne
rect 10435 6939 10789 7037
tri 10789 6939 10887 7037 sw
tri 10887 6939 10985 7037 ne
rect 10985 6939 11339 7037
tri 11339 6939 11437 7037 sw
tri 11437 6939 11535 7037 ne
rect 11535 6939 11889 7037
tri 11889 6939 11987 7037 sw
tri 11987 6939 12085 7037 ne
rect 12085 6939 12439 7037
tri 12439 6939 12537 7037 sw
tri 12537 6939 12635 7037 ne
rect 12635 6939 12989 7037
tri 12989 6939 13087 7037 sw
tri 13087 6939 13185 7037 ne
rect 13185 6939 13539 7037
tri 13539 6939 13637 7037 sw
tri 13637 6939 13735 7037 ne
rect 13735 6939 14089 7037
tri 14089 6939 14187 7037 sw
tri 14187 6939 14285 7037 ne
rect 14285 6939 14639 7037
tri 14639 6939 14737 7037 sw
tri 14737 6939 14835 7037 ne
rect 14835 6939 15189 7037
tri 15189 6939 15287 7037 sw
tri 15287 6939 15385 7037 ne
rect 15385 6939 15739 7037
tri 15739 6939 15837 7037 sw
tri 15837 6939 15935 7037 ne
rect 15935 6939 16289 7037
tri 16289 6939 16387 7037 sw
tri 16387 6939 16485 7037 ne
rect 16485 6939 16839 7037
tri 16839 6939 16937 7037 sw
tri 16937 6939 17035 7037 ne
rect 17035 6939 17389 7037
tri 17389 6939 17487 7037 sw
tri 17487 6939 17585 7037 ne
rect 17585 6939 17939 7037
tri 17939 6939 18037 7037 sw
tri 18037 6939 18135 7037 ne
rect 18135 6939 18489 7037
tri 18489 6939 18587 7037 sw
tri 18587 6939 18685 7037 ne
rect 18685 6939 19039 7037
tri 19039 6939 19137 7037 sw
tri 19137 6939 19235 7037 ne
rect 19235 6939 19589 7037
tri 19589 6939 19687 7037 sw
rect -500 6935 437 6939
rect -500 6815 215 6935
rect 335 6841 437 6935
tri 437 6841 535 6939 sw
tri 535 6841 633 6939 ne
rect 633 6935 987 6939
rect 633 6841 765 6935
rect 335 6815 535 6841
rect -500 6811 535 6815
tri 535 6811 565 6841 sw
tri 633 6811 663 6841 ne
rect 663 6815 765 6841
rect 885 6841 987 6935
tri 987 6841 1085 6939 sw
tri 1085 6841 1183 6939 ne
rect 1183 6935 1537 6939
rect 1183 6841 1315 6935
rect 885 6815 1085 6841
rect 663 6811 1085 6815
tri 1085 6811 1115 6841 sw
tri 1183 6811 1213 6841 ne
rect 1213 6815 1315 6841
rect 1435 6841 1537 6935
tri 1537 6841 1635 6939 sw
tri 1635 6841 1733 6939 ne
rect 1733 6935 2087 6939
rect 1733 6841 1865 6935
rect 1435 6815 1635 6841
rect 1213 6811 1635 6815
tri 1635 6811 1665 6841 sw
tri 1733 6811 1763 6841 ne
rect 1763 6815 1865 6841
rect 1985 6841 2087 6935
tri 2087 6841 2185 6939 sw
tri 2185 6841 2283 6939 ne
rect 2283 6935 2637 6939
rect 2283 6841 2415 6935
rect 1985 6815 2185 6841
rect 1763 6811 2185 6815
tri 2185 6811 2215 6841 sw
tri 2283 6811 2313 6841 ne
rect 2313 6815 2415 6841
rect 2535 6841 2637 6935
tri 2637 6841 2735 6939 sw
tri 2735 6841 2833 6939 ne
rect 2833 6935 3187 6939
rect 2833 6841 2965 6935
rect 2535 6815 2735 6841
rect 2313 6811 2735 6815
tri 2735 6811 2765 6841 sw
tri 2833 6811 2863 6841 ne
rect 2863 6815 2965 6841
rect 3085 6841 3187 6935
tri 3187 6841 3285 6939 sw
tri 3285 6841 3383 6939 ne
rect 3383 6935 3737 6939
rect 3383 6841 3515 6935
rect 3085 6815 3285 6841
rect 2863 6811 3285 6815
tri 3285 6811 3315 6841 sw
tri 3383 6811 3413 6841 ne
rect 3413 6815 3515 6841
rect 3635 6841 3737 6935
tri 3737 6841 3835 6939 sw
tri 3835 6841 3933 6939 ne
rect 3933 6935 4287 6939
rect 3933 6841 4065 6935
rect 3635 6815 3835 6841
rect 3413 6811 3835 6815
tri 3835 6811 3865 6841 sw
tri 3933 6811 3963 6841 ne
rect 3963 6815 4065 6841
rect 4185 6841 4287 6935
tri 4287 6841 4385 6939 sw
tri 4385 6841 4483 6939 ne
rect 4483 6935 4837 6939
rect 4483 6841 4615 6935
rect 4185 6815 4385 6841
rect 3963 6811 4385 6815
tri 4385 6811 4415 6841 sw
tri 4483 6811 4513 6841 ne
rect 4513 6815 4615 6841
rect 4735 6841 4837 6935
tri 4837 6841 4935 6939 sw
tri 4935 6841 5033 6939 ne
rect 5033 6935 5387 6939
rect 5033 6841 5165 6935
rect 4735 6815 4935 6841
rect 4513 6811 4935 6815
tri 4935 6811 4965 6841 sw
tri 5033 6811 5063 6841 ne
rect 5063 6815 5165 6841
rect 5285 6841 5387 6935
tri 5387 6841 5485 6939 sw
tri 5485 6841 5583 6939 ne
rect 5583 6935 5937 6939
rect 5583 6841 5715 6935
rect 5285 6815 5485 6841
rect 5063 6811 5485 6815
tri 5485 6811 5515 6841 sw
tri 5583 6811 5613 6841 ne
rect 5613 6815 5715 6841
rect 5835 6841 5937 6935
tri 5937 6841 6035 6939 sw
tri 6035 6841 6133 6939 ne
rect 6133 6935 6487 6939
rect 6133 6841 6265 6935
rect 5835 6815 6035 6841
rect 5613 6811 6035 6815
tri 6035 6811 6065 6841 sw
tri 6133 6811 6163 6841 ne
rect 6163 6815 6265 6841
rect 6385 6841 6487 6935
tri 6487 6841 6585 6939 sw
tri 6585 6841 6683 6939 ne
rect 6683 6935 7037 6939
rect 6683 6841 6815 6935
rect 6385 6815 6585 6841
rect 6163 6811 6585 6815
tri 6585 6811 6615 6841 sw
tri 6683 6811 6713 6841 ne
rect 6713 6815 6815 6841
rect 6935 6841 7037 6935
tri 7037 6841 7135 6939 sw
tri 7135 6841 7233 6939 ne
rect 7233 6935 7587 6939
rect 7233 6841 7365 6935
rect 6935 6815 7135 6841
rect 6713 6811 7135 6815
tri 7135 6811 7165 6841 sw
tri 7233 6811 7263 6841 ne
rect 7263 6815 7365 6841
rect 7485 6841 7587 6935
tri 7587 6841 7685 6939 sw
tri 7685 6841 7783 6939 ne
rect 7783 6935 8137 6939
rect 7783 6841 7915 6935
rect 7485 6815 7685 6841
rect 7263 6811 7685 6815
tri 7685 6811 7715 6841 sw
tri 7783 6811 7813 6841 ne
rect 7813 6815 7915 6841
rect 8035 6841 8137 6935
tri 8137 6841 8235 6939 sw
tri 8235 6841 8333 6939 ne
rect 8333 6935 8687 6939
rect 8333 6841 8465 6935
rect 8035 6815 8235 6841
rect 7813 6811 8235 6815
tri 8235 6811 8265 6841 sw
tri 8333 6811 8363 6841 ne
rect 8363 6815 8465 6841
rect 8585 6841 8687 6935
tri 8687 6841 8785 6939 sw
tri 8785 6841 8883 6939 ne
rect 8883 6935 9237 6939
rect 8883 6841 9015 6935
rect 8585 6815 8785 6841
rect 8363 6811 8785 6815
tri 8785 6811 8815 6841 sw
tri 8883 6811 8913 6841 ne
rect 8913 6815 9015 6841
rect 9135 6841 9237 6935
tri 9237 6841 9335 6939 sw
tri 9335 6841 9433 6939 ne
rect 9433 6935 9787 6939
rect 9433 6841 9565 6935
rect 9135 6815 9335 6841
rect 8913 6811 9335 6815
tri 9335 6811 9365 6841 sw
tri 9433 6811 9463 6841 ne
rect 9463 6815 9565 6841
rect 9685 6841 9787 6935
tri 9787 6841 9885 6939 sw
tri 9885 6841 9983 6939 ne
rect 9983 6935 10337 6939
rect 9983 6841 10115 6935
rect 9685 6815 9885 6841
rect 9463 6811 9885 6815
tri 9885 6811 9915 6841 sw
tri 9983 6811 10013 6841 ne
rect 10013 6815 10115 6841
rect 10235 6841 10337 6935
tri 10337 6841 10435 6939 sw
tri 10435 6841 10533 6939 ne
rect 10533 6935 10887 6939
rect 10533 6841 10665 6935
rect 10235 6815 10435 6841
rect 10013 6811 10435 6815
tri 10435 6811 10465 6841 sw
tri 10533 6811 10563 6841 ne
rect 10563 6815 10665 6841
rect 10785 6841 10887 6935
tri 10887 6841 10985 6939 sw
tri 10985 6841 11083 6939 ne
rect 11083 6935 11437 6939
rect 11083 6841 11215 6935
rect 10785 6815 10985 6841
rect 10563 6811 10985 6815
tri 10985 6811 11015 6841 sw
tri 11083 6811 11113 6841 ne
rect 11113 6815 11215 6841
rect 11335 6841 11437 6935
tri 11437 6841 11535 6939 sw
tri 11535 6841 11633 6939 ne
rect 11633 6935 11987 6939
rect 11633 6841 11765 6935
rect 11335 6815 11535 6841
rect 11113 6811 11535 6815
tri 11535 6811 11565 6841 sw
tri 11633 6811 11663 6841 ne
rect 11663 6815 11765 6841
rect 11885 6841 11987 6935
tri 11987 6841 12085 6939 sw
tri 12085 6841 12183 6939 ne
rect 12183 6935 12537 6939
rect 12183 6841 12315 6935
rect 11885 6815 12085 6841
rect 11663 6811 12085 6815
tri 12085 6811 12115 6841 sw
tri 12183 6811 12213 6841 ne
rect 12213 6815 12315 6841
rect 12435 6841 12537 6935
tri 12537 6841 12635 6939 sw
tri 12635 6841 12733 6939 ne
rect 12733 6935 13087 6939
rect 12733 6841 12865 6935
rect 12435 6815 12635 6841
rect 12213 6811 12635 6815
tri 12635 6811 12665 6841 sw
tri 12733 6811 12763 6841 ne
rect 12763 6815 12865 6841
rect 12985 6841 13087 6935
tri 13087 6841 13185 6939 sw
tri 13185 6841 13283 6939 ne
rect 13283 6935 13637 6939
rect 13283 6841 13415 6935
rect 12985 6815 13185 6841
rect 12763 6811 13185 6815
tri 13185 6811 13215 6841 sw
tri 13283 6811 13313 6841 ne
rect 13313 6815 13415 6841
rect 13535 6841 13637 6935
tri 13637 6841 13735 6939 sw
tri 13735 6841 13833 6939 ne
rect 13833 6935 14187 6939
rect 13833 6841 13965 6935
rect 13535 6815 13735 6841
rect 13313 6811 13735 6815
tri 13735 6811 13765 6841 sw
tri 13833 6811 13863 6841 ne
rect 13863 6815 13965 6841
rect 14085 6841 14187 6935
tri 14187 6841 14285 6939 sw
tri 14285 6841 14383 6939 ne
rect 14383 6935 14737 6939
rect 14383 6841 14515 6935
rect 14085 6815 14285 6841
rect 13863 6811 14285 6815
tri 14285 6811 14315 6841 sw
tri 14383 6811 14413 6841 ne
rect 14413 6815 14515 6841
rect 14635 6841 14737 6935
tri 14737 6841 14835 6939 sw
tri 14835 6841 14933 6939 ne
rect 14933 6935 15287 6939
rect 14933 6841 15065 6935
rect 14635 6815 14835 6841
rect 14413 6811 14835 6815
tri 14835 6811 14865 6841 sw
tri 14933 6811 14963 6841 ne
rect 14963 6815 15065 6841
rect 15185 6841 15287 6935
tri 15287 6841 15385 6939 sw
tri 15385 6841 15483 6939 ne
rect 15483 6935 15837 6939
rect 15483 6841 15615 6935
rect 15185 6815 15385 6841
rect 14963 6811 15385 6815
tri 15385 6811 15415 6841 sw
tri 15483 6811 15513 6841 ne
rect 15513 6815 15615 6841
rect 15735 6841 15837 6935
tri 15837 6841 15935 6939 sw
tri 15935 6841 16033 6939 ne
rect 16033 6935 16387 6939
rect 16033 6841 16165 6935
rect 15735 6815 15935 6841
rect 15513 6811 15935 6815
tri 15935 6811 15965 6841 sw
tri 16033 6811 16063 6841 ne
rect 16063 6815 16165 6841
rect 16285 6841 16387 6935
tri 16387 6841 16485 6939 sw
tri 16485 6841 16583 6939 ne
rect 16583 6935 16937 6939
rect 16583 6841 16715 6935
rect 16285 6815 16485 6841
rect 16063 6811 16485 6815
tri 16485 6811 16515 6841 sw
tri 16583 6811 16613 6841 ne
rect 16613 6815 16715 6841
rect 16835 6841 16937 6935
tri 16937 6841 17035 6939 sw
tri 17035 6841 17133 6939 ne
rect 17133 6935 17487 6939
rect 17133 6841 17265 6935
rect 16835 6815 17035 6841
rect 16613 6811 17035 6815
tri 17035 6811 17065 6841 sw
tri 17133 6811 17163 6841 ne
rect 17163 6815 17265 6841
rect 17385 6841 17487 6935
tri 17487 6841 17585 6939 sw
tri 17585 6841 17683 6939 ne
rect 17683 6935 18037 6939
rect 17683 6841 17815 6935
rect 17385 6815 17585 6841
rect 17163 6811 17585 6815
tri 17585 6811 17615 6841 sw
tri 17683 6811 17713 6841 ne
rect 17713 6815 17815 6841
rect 17935 6841 18037 6935
tri 18037 6841 18135 6939 sw
tri 18135 6841 18233 6939 ne
rect 18233 6935 18587 6939
rect 18233 6841 18365 6935
rect 17935 6815 18135 6841
rect 17713 6811 18135 6815
tri 18135 6811 18165 6841 sw
tri 18233 6811 18263 6841 ne
rect 18263 6815 18365 6841
rect 18485 6841 18587 6935
tri 18587 6841 18685 6939 sw
tri 18685 6841 18783 6939 ne
rect 18783 6935 19137 6939
rect 18783 6841 18915 6935
rect 18485 6815 18685 6841
rect 18263 6811 18685 6815
tri 18685 6811 18715 6841 sw
tri 18783 6811 18813 6841 ne
rect 18813 6815 18915 6841
rect 19035 6841 19137 6935
tri 19137 6841 19235 6939 sw
tri 19235 6841 19333 6939 ne
rect 19333 6935 20300 6939
rect 19333 6841 19465 6935
rect 19035 6815 19235 6841
rect 18813 6811 19235 6815
tri 19235 6811 19265 6841 sw
tri 19333 6811 19363 6841 ne
rect 19363 6815 19465 6841
rect 19585 6815 20300 6935
rect 19363 6811 20300 6815
tri 113 6713 211 6811 ne
rect 211 6713 565 6811
tri 565 6713 663 6811 sw
tri 663 6713 761 6811 ne
rect 761 6713 1115 6811
tri 1115 6713 1213 6811 sw
tri 1213 6713 1311 6811 ne
rect 1311 6713 1665 6811
tri 1665 6713 1763 6811 sw
tri 1763 6713 1861 6811 ne
rect 1861 6713 2215 6811
tri 2215 6713 2313 6811 sw
tri 2313 6713 2411 6811 ne
rect 2411 6713 2765 6811
tri 2765 6713 2863 6811 sw
tri 2863 6713 2961 6811 ne
rect 2961 6713 3315 6811
tri 3315 6713 3413 6811 sw
tri 3413 6713 3511 6811 ne
rect 3511 6713 3865 6811
tri 3865 6713 3963 6811 sw
tri 3963 6713 4061 6811 ne
rect 4061 6713 4415 6811
tri 4415 6713 4513 6811 sw
tri 4513 6713 4611 6811 ne
rect 4611 6713 4965 6811
tri 4965 6713 5063 6811 sw
tri 5063 6713 5161 6811 ne
rect 5161 6713 5515 6811
tri 5515 6713 5613 6811 sw
tri 5613 6713 5711 6811 ne
rect 5711 6713 6065 6811
tri 6065 6713 6163 6811 sw
tri 6163 6713 6261 6811 ne
rect 6261 6713 6615 6811
tri 6615 6713 6713 6811 sw
tri 6713 6713 6811 6811 ne
rect 6811 6713 7165 6811
tri 7165 6713 7263 6811 sw
tri 7263 6713 7361 6811 ne
rect 7361 6713 7715 6811
tri 7715 6713 7813 6811 sw
tri 7813 6713 7911 6811 ne
rect 7911 6713 8265 6811
tri 8265 6713 8363 6811 sw
tri 8363 6713 8461 6811 ne
rect 8461 6713 8815 6811
tri 8815 6713 8913 6811 sw
tri 8913 6713 9011 6811 ne
rect 9011 6713 9365 6811
tri 9365 6713 9463 6811 sw
tri 9463 6713 9561 6811 ne
rect 9561 6713 9915 6811
tri 9915 6713 10013 6811 sw
tri 10013 6713 10111 6811 ne
rect 10111 6713 10465 6811
tri 10465 6713 10563 6811 sw
tri 10563 6713 10661 6811 ne
rect 10661 6713 11015 6811
tri 11015 6713 11113 6811 sw
tri 11113 6713 11211 6811 ne
rect 11211 6713 11565 6811
tri 11565 6713 11663 6811 sw
tri 11663 6713 11761 6811 ne
rect 11761 6713 12115 6811
tri 12115 6713 12213 6811 sw
tri 12213 6713 12311 6811 ne
rect 12311 6713 12665 6811
tri 12665 6713 12763 6811 sw
tri 12763 6713 12861 6811 ne
rect 12861 6713 13215 6811
tri 13215 6713 13313 6811 sw
tri 13313 6713 13411 6811 ne
rect 13411 6713 13765 6811
tri 13765 6713 13863 6811 sw
tri 13863 6713 13961 6811 ne
rect 13961 6713 14315 6811
tri 14315 6713 14413 6811 sw
tri 14413 6713 14511 6811 ne
rect 14511 6713 14865 6811
tri 14865 6713 14963 6811 sw
tri 14963 6713 15061 6811 ne
rect 15061 6713 15415 6811
tri 15415 6713 15513 6811 sw
tri 15513 6713 15611 6811 ne
rect 15611 6713 15965 6811
tri 15965 6713 16063 6811 sw
tri 16063 6713 16161 6811 ne
rect 16161 6713 16515 6811
tri 16515 6713 16613 6811 sw
tri 16613 6713 16711 6811 ne
rect 16711 6713 17065 6811
tri 17065 6713 17163 6811 sw
tri 17163 6713 17261 6811 ne
rect 17261 6713 17615 6811
tri 17615 6713 17713 6811 sw
tri 17713 6713 17811 6811 ne
rect 17811 6713 18165 6811
tri 18165 6713 18263 6811 sw
tri 18263 6713 18361 6811 ne
rect 18361 6713 18715 6811
tri 18715 6713 18813 6811 sw
tri 18813 6713 18911 6811 ne
rect 18911 6713 19265 6811
tri 19265 6713 19363 6811 sw
tri 19363 6713 19461 6811 ne
rect 19461 6713 20300 6811
rect -2000 6683 113 6713
tri 113 6683 143 6713 sw
tri 211 6683 241 6713 ne
rect 241 6683 663 6713
tri 663 6683 693 6713 sw
tri 761 6683 791 6713 ne
rect 791 6683 1213 6713
tri 1213 6683 1243 6713 sw
tri 1311 6683 1341 6713 ne
rect 1341 6683 1763 6713
tri 1763 6683 1793 6713 sw
tri 1861 6683 1891 6713 ne
rect 1891 6683 2313 6713
tri 2313 6683 2343 6713 sw
tri 2411 6683 2441 6713 ne
rect 2441 6683 2863 6713
tri 2863 6683 2893 6713 sw
tri 2961 6683 2991 6713 ne
rect 2991 6683 3413 6713
tri 3413 6683 3443 6713 sw
tri 3511 6683 3541 6713 ne
rect 3541 6683 3963 6713
tri 3963 6683 3993 6713 sw
tri 4061 6683 4091 6713 ne
rect 4091 6683 4513 6713
tri 4513 6683 4543 6713 sw
tri 4611 6683 4641 6713 ne
rect 4641 6683 5063 6713
tri 5063 6683 5093 6713 sw
tri 5161 6683 5191 6713 ne
rect 5191 6683 5613 6713
tri 5613 6683 5643 6713 sw
tri 5711 6683 5741 6713 ne
rect 5741 6683 6163 6713
tri 6163 6683 6193 6713 sw
tri 6261 6683 6291 6713 ne
rect 6291 6683 6713 6713
tri 6713 6683 6743 6713 sw
tri 6811 6683 6841 6713 ne
rect 6841 6683 7263 6713
tri 7263 6683 7293 6713 sw
tri 7361 6683 7391 6713 ne
rect 7391 6683 7813 6713
tri 7813 6683 7843 6713 sw
tri 7911 6683 7941 6713 ne
rect 7941 6683 8363 6713
tri 8363 6683 8393 6713 sw
tri 8461 6683 8491 6713 ne
rect 8491 6683 8913 6713
tri 8913 6683 8943 6713 sw
tri 9011 6683 9041 6713 ne
rect 9041 6683 9463 6713
tri 9463 6683 9493 6713 sw
tri 9561 6683 9591 6713 ne
rect 9591 6683 10013 6713
tri 10013 6683 10043 6713 sw
tri 10111 6683 10141 6713 ne
rect 10141 6683 10563 6713
tri 10563 6683 10593 6713 sw
tri 10661 6683 10691 6713 ne
rect 10691 6683 11113 6713
tri 11113 6683 11143 6713 sw
tri 11211 6683 11241 6713 ne
rect 11241 6683 11663 6713
tri 11663 6683 11693 6713 sw
tri 11761 6683 11791 6713 ne
rect 11791 6683 12213 6713
tri 12213 6683 12243 6713 sw
tri 12311 6683 12341 6713 ne
rect 12341 6683 12763 6713
tri 12763 6683 12793 6713 sw
tri 12861 6683 12891 6713 ne
rect 12891 6683 13313 6713
tri 13313 6683 13343 6713 sw
tri 13411 6683 13441 6713 ne
rect 13441 6683 13863 6713
tri 13863 6683 13893 6713 sw
tri 13961 6683 13991 6713 ne
rect 13991 6683 14413 6713
tri 14413 6683 14443 6713 sw
tri 14511 6683 14541 6713 ne
rect 14541 6683 14963 6713
tri 14963 6683 14993 6713 sw
tri 15061 6683 15091 6713 ne
rect 15091 6683 15513 6713
tri 15513 6683 15543 6713 sw
tri 15611 6683 15641 6713 ne
rect 15641 6683 16063 6713
tri 16063 6683 16093 6713 sw
tri 16161 6683 16191 6713 ne
rect 16191 6683 16613 6713
tri 16613 6683 16643 6713 sw
tri 16711 6683 16741 6713 ne
rect 16741 6683 17163 6713
tri 17163 6683 17193 6713 sw
tri 17261 6683 17291 6713 ne
rect 17291 6683 17713 6713
tri 17713 6683 17743 6713 sw
tri 17811 6683 17841 6713 ne
rect 17841 6683 18263 6713
tri 18263 6683 18293 6713 sw
tri 18361 6683 18391 6713 ne
rect 18391 6683 18813 6713
tri 18813 6683 18843 6713 sw
tri 18911 6683 18941 6713 ne
rect 18941 6683 19363 6713
tri 19363 6683 19393 6713 sw
tri 19461 6683 19491 6713 ne
rect 19491 6683 20300 6713
rect -2000 6585 143 6683
tri 143 6585 241 6683 sw
tri 241 6585 339 6683 ne
rect 339 6585 693 6683
tri 693 6585 791 6683 sw
tri 791 6585 889 6683 ne
rect 889 6585 1243 6683
tri 1243 6585 1341 6683 sw
tri 1341 6585 1439 6683 ne
rect 1439 6585 1793 6683
tri 1793 6585 1891 6683 sw
tri 1891 6585 1989 6683 ne
rect 1989 6585 2343 6683
tri 2343 6585 2441 6683 sw
tri 2441 6585 2539 6683 ne
rect 2539 6585 2893 6683
tri 2893 6585 2991 6683 sw
tri 2991 6585 3089 6683 ne
rect 3089 6585 3443 6683
tri 3443 6585 3541 6683 sw
tri 3541 6585 3639 6683 ne
rect 3639 6585 3993 6683
tri 3993 6585 4091 6683 sw
tri 4091 6585 4189 6683 ne
rect 4189 6585 4543 6683
tri 4543 6585 4641 6683 sw
tri 4641 6585 4739 6683 ne
rect 4739 6585 5093 6683
tri 5093 6585 5191 6683 sw
tri 5191 6585 5289 6683 ne
rect 5289 6585 5643 6683
tri 5643 6585 5741 6683 sw
tri 5741 6585 5839 6683 ne
rect 5839 6585 6193 6683
tri 6193 6585 6291 6683 sw
tri 6291 6585 6389 6683 ne
rect 6389 6585 6743 6683
tri 6743 6585 6841 6683 sw
tri 6841 6585 6939 6683 ne
rect 6939 6585 7293 6683
tri 7293 6585 7391 6683 sw
tri 7391 6585 7489 6683 ne
rect 7489 6585 7843 6683
tri 7843 6585 7941 6683 sw
tri 7941 6585 8039 6683 ne
rect 8039 6585 8393 6683
tri 8393 6585 8491 6683 sw
tri 8491 6585 8589 6683 ne
rect 8589 6585 8943 6683
tri 8943 6585 9041 6683 sw
tri 9041 6585 9139 6683 ne
rect 9139 6585 9493 6683
tri 9493 6585 9591 6683 sw
tri 9591 6585 9689 6683 ne
rect 9689 6585 10043 6683
tri 10043 6585 10141 6683 sw
tri 10141 6585 10239 6683 ne
rect 10239 6585 10593 6683
tri 10593 6585 10691 6683 sw
tri 10691 6585 10789 6683 ne
rect 10789 6585 11143 6683
tri 11143 6585 11241 6683 sw
tri 11241 6585 11339 6683 ne
rect 11339 6585 11693 6683
tri 11693 6585 11791 6683 sw
tri 11791 6585 11889 6683 ne
rect 11889 6585 12243 6683
tri 12243 6585 12341 6683 sw
tri 12341 6585 12439 6683 ne
rect 12439 6585 12793 6683
tri 12793 6585 12891 6683 sw
tri 12891 6585 12989 6683 ne
rect 12989 6585 13343 6683
tri 13343 6585 13441 6683 sw
tri 13441 6585 13539 6683 ne
rect 13539 6585 13893 6683
tri 13893 6585 13991 6683 sw
tri 13991 6585 14089 6683 ne
rect 14089 6585 14443 6683
tri 14443 6585 14541 6683 sw
tri 14541 6585 14639 6683 ne
rect 14639 6585 14993 6683
tri 14993 6585 15091 6683 sw
tri 15091 6585 15189 6683 ne
rect 15189 6585 15543 6683
tri 15543 6585 15641 6683 sw
tri 15641 6585 15739 6683 ne
rect 15739 6585 16093 6683
tri 16093 6585 16191 6683 sw
tri 16191 6585 16289 6683 ne
rect 16289 6585 16643 6683
tri 16643 6585 16741 6683 sw
tri 16741 6585 16839 6683 ne
rect 16839 6585 17193 6683
tri 17193 6585 17291 6683 sw
tri 17291 6585 17389 6683 ne
rect 17389 6585 17743 6683
tri 17743 6585 17841 6683 sw
tri 17841 6585 17939 6683 ne
rect 17939 6585 18293 6683
tri 18293 6585 18391 6683 sw
tri 18391 6585 18489 6683 ne
rect 18489 6585 18843 6683
tri 18843 6585 18941 6683 sw
tri 18941 6585 19039 6683 ne
rect 19039 6585 19393 6683
tri 19393 6585 19491 6683 sw
tri 19491 6585 19589 6683 ne
rect 19589 6585 20300 6683
rect -2000 6487 241 6585
tri 241 6487 339 6585 sw
tri 339 6487 437 6585 ne
rect 437 6487 791 6585
tri 791 6487 889 6585 sw
tri 889 6487 987 6585 ne
rect 987 6487 1341 6585
tri 1341 6487 1439 6585 sw
tri 1439 6487 1537 6585 ne
rect 1537 6487 1891 6585
tri 1891 6487 1989 6585 sw
tri 1989 6487 2087 6585 ne
rect 2087 6487 2441 6585
tri 2441 6487 2539 6585 sw
tri 2539 6487 2637 6585 ne
rect 2637 6487 2991 6585
tri 2991 6487 3089 6585 sw
tri 3089 6487 3187 6585 ne
rect 3187 6487 3541 6585
tri 3541 6487 3639 6585 sw
tri 3639 6487 3737 6585 ne
rect 3737 6487 4091 6585
tri 4091 6487 4189 6585 sw
tri 4189 6487 4287 6585 ne
rect 4287 6487 4641 6585
tri 4641 6487 4739 6585 sw
tri 4739 6487 4837 6585 ne
rect 4837 6487 5191 6585
tri 5191 6487 5289 6585 sw
tri 5289 6487 5387 6585 ne
rect 5387 6487 5741 6585
tri 5741 6487 5839 6585 sw
tri 5839 6487 5937 6585 ne
rect 5937 6487 6291 6585
tri 6291 6487 6389 6585 sw
tri 6389 6487 6487 6585 ne
rect 6487 6487 6841 6585
tri 6841 6487 6939 6585 sw
tri 6939 6487 7037 6585 ne
rect 7037 6487 7391 6585
tri 7391 6487 7489 6585 sw
tri 7489 6487 7587 6585 ne
rect 7587 6487 7941 6585
tri 7941 6487 8039 6585 sw
tri 8039 6487 8137 6585 ne
rect 8137 6487 8491 6585
tri 8491 6487 8589 6585 sw
tri 8589 6487 8687 6585 ne
rect 8687 6487 9041 6585
tri 9041 6487 9139 6585 sw
tri 9139 6487 9237 6585 ne
rect 9237 6487 9591 6585
tri 9591 6487 9689 6585 sw
tri 9689 6487 9787 6585 ne
rect 9787 6487 10141 6585
tri 10141 6487 10239 6585 sw
tri 10239 6487 10337 6585 ne
rect 10337 6487 10691 6585
tri 10691 6487 10789 6585 sw
tri 10789 6487 10887 6585 ne
rect 10887 6487 11241 6585
tri 11241 6487 11339 6585 sw
tri 11339 6487 11437 6585 ne
rect 11437 6487 11791 6585
tri 11791 6487 11889 6585 sw
tri 11889 6487 11987 6585 ne
rect 11987 6487 12341 6585
tri 12341 6487 12439 6585 sw
tri 12439 6487 12537 6585 ne
rect 12537 6487 12891 6585
tri 12891 6487 12989 6585 sw
tri 12989 6487 13087 6585 ne
rect 13087 6487 13441 6585
tri 13441 6487 13539 6585 sw
tri 13539 6487 13637 6585 ne
rect 13637 6487 13991 6585
tri 13991 6487 14089 6585 sw
tri 14089 6487 14187 6585 ne
rect 14187 6487 14541 6585
tri 14541 6487 14639 6585 sw
tri 14639 6487 14737 6585 ne
rect 14737 6487 15091 6585
tri 15091 6487 15189 6585 sw
tri 15189 6487 15287 6585 ne
rect 15287 6487 15641 6585
tri 15641 6487 15739 6585 sw
tri 15739 6487 15837 6585 ne
rect 15837 6487 16191 6585
tri 16191 6487 16289 6585 sw
tri 16289 6487 16387 6585 ne
rect 16387 6487 16741 6585
tri 16741 6487 16839 6585 sw
tri 16839 6487 16937 6585 ne
rect 16937 6487 17291 6585
tri 17291 6487 17389 6585 sw
tri 17389 6487 17487 6585 ne
rect 17487 6487 17841 6585
tri 17841 6487 17939 6585 sw
tri 17939 6487 18037 6585 ne
rect 18037 6487 18391 6585
tri 18391 6487 18489 6585 sw
tri 18489 6487 18587 6585 ne
rect 18587 6487 18941 6585
tri 18941 6487 19039 6585 sw
tri 19039 6487 19137 6585 ne
rect 19137 6487 19491 6585
tri 19491 6487 19589 6585 sw
tri 19589 6487 19687 6585 ne
rect 19687 6487 20300 6585
rect -2000 6389 339 6487
tri 339 6389 437 6487 sw
tri 437 6389 535 6487 ne
rect 535 6389 889 6487
tri 889 6389 987 6487 sw
tri 987 6389 1085 6487 ne
rect 1085 6389 1439 6487
tri 1439 6389 1537 6487 sw
tri 1537 6389 1635 6487 ne
rect 1635 6389 1989 6487
tri 1989 6389 2087 6487 sw
tri 2087 6389 2185 6487 ne
rect 2185 6389 2539 6487
tri 2539 6389 2637 6487 sw
tri 2637 6389 2735 6487 ne
rect 2735 6389 3089 6487
tri 3089 6389 3187 6487 sw
tri 3187 6389 3285 6487 ne
rect 3285 6389 3639 6487
tri 3639 6389 3737 6487 sw
tri 3737 6389 3835 6487 ne
rect 3835 6389 4189 6487
tri 4189 6389 4287 6487 sw
tri 4287 6389 4385 6487 ne
rect 4385 6389 4739 6487
tri 4739 6389 4837 6487 sw
tri 4837 6389 4935 6487 ne
rect 4935 6389 5289 6487
tri 5289 6389 5387 6487 sw
tri 5387 6389 5485 6487 ne
rect 5485 6389 5839 6487
tri 5839 6389 5937 6487 sw
tri 5937 6389 6035 6487 ne
rect 6035 6389 6389 6487
tri 6389 6389 6487 6487 sw
tri 6487 6389 6585 6487 ne
rect 6585 6389 6939 6487
tri 6939 6389 7037 6487 sw
tri 7037 6389 7135 6487 ne
rect 7135 6389 7489 6487
tri 7489 6389 7587 6487 sw
tri 7587 6389 7685 6487 ne
rect 7685 6389 8039 6487
tri 8039 6389 8137 6487 sw
tri 8137 6389 8235 6487 ne
rect 8235 6389 8589 6487
tri 8589 6389 8687 6487 sw
tri 8687 6389 8785 6487 ne
rect 8785 6389 9139 6487
tri 9139 6389 9237 6487 sw
tri 9237 6389 9335 6487 ne
rect 9335 6389 9689 6487
tri 9689 6389 9787 6487 sw
tri 9787 6389 9885 6487 ne
rect 9885 6389 10239 6487
tri 10239 6389 10337 6487 sw
tri 10337 6389 10435 6487 ne
rect 10435 6389 10789 6487
tri 10789 6389 10887 6487 sw
tri 10887 6389 10985 6487 ne
rect 10985 6389 11339 6487
tri 11339 6389 11437 6487 sw
tri 11437 6389 11535 6487 ne
rect 11535 6389 11889 6487
tri 11889 6389 11987 6487 sw
tri 11987 6389 12085 6487 ne
rect 12085 6389 12439 6487
tri 12439 6389 12537 6487 sw
tri 12537 6389 12635 6487 ne
rect 12635 6389 12989 6487
tri 12989 6389 13087 6487 sw
tri 13087 6389 13185 6487 ne
rect 13185 6389 13539 6487
tri 13539 6389 13637 6487 sw
tri 13637 6389 13735 6487 ne
rect 13735 6389 14089 6487
tri 14089 6389 14187 6487 sw
tri 14187 6389 14285 6487 ne
rect 14285 6389 14639 6487
tri 14639 6389 14737 6487 sw
tri 14737 6389 14835 6487 ne
rect 14835 6389 15189 6487
tri 15189 6389 15287 6487 sw
tri 15287 6389 15385 6487 ne
rect 15385 6389 15739 6487
tri 15739 6389 15837 6487 sw
tri 15837 6389 15935 6487 ne
rect 15935 6389 16289 6487
tri 16289 6389 16387 6487 sw
tri 16387 6389 16485 6487 ne
rect 16485 6389 16839 6487
tri 16839 6389 16937 6487 sw
tri 16937 6389 17035 6487 ne
rect 17035 6389 17389 6487
tri 17389 6389 17487 6487 sw
tri 17487 6389 17585 6487 ne
rect 17585 6389 17939 6487
tri 17939 6389 18037 6487 sw
tri 18037 6389 18135 6487 ne
rect 18135 6389 18489 6487
tri 18489 6389 18587 6487 sw
tri 18587 6389 18685 6487 ne
rect 18685 6389 19039 6487
tri 19039 6389 19137 6487 sw
tri 19137 6389 19235 6487 ne
rect 19235 6389 19589 6487
tri 19589 6389 19687 6487 sw
rect 20800 6389 21800 7037
rect -2000 6385 437 6389
rect -2000 6265 215 6385
rect 335 6291 437 6385
tri 437 6291 535 6389 sw
tri 535 6291 633 6389 ne
rect 633 6385 987 6389
rect 633 6291 765 6385
rect 335 6265 535 6291
rect -2000 6261 535 6265
rect -2000 5613 -1000 6261
tri 113 6163 211 6261 ne
rect 211 6213 535 6261
tri 535 6213 613 6291 sw
tri 633 6213 711 6291 ne
rect 711 6265 765 6291
rect 885 6291 987 6385
tri 987 6291 1085 6389 sw
tri 1085 6291 1183 6389 ne
rect 1183 6385 1537 6389
rect 1183 6291 1315 6385
rect 885 6265 1085 6291
rect 711 6213 1085 6265
tri 1085 6213 1163 6291 sw
tri 1183 6213 1261 6291 ne
rect 1261 6265 1315 6291
rect 1435 6291 1537 6385
tri 1537 6291 1635 6389 sw
tri 1635 6291 1733 6389 ne
rect 1733 6385 2087 6389
rect 1733 6291 1865 6385
rect 1435 6265 1635 6291
rect 1261 6213 1635 6265
tri 1635 6213 1713 6291 sw
tri 1733 6213 1811 6291 ne
rect 1811 6265 1865 6291
rect 1985 6291 2087 6385
tri 2087 6291 2185 6389 sw
tri 2185 6291 2283 6389 ne
rect 2283 6385 2637 6389
rect 2283 6291 2415 6385
rect 1985 6265 2185 6291
rect 1811 6213 2185 6265
tri 2185 6213 2263 6291 sw
tri 2283 6213 2361 6291 ne
rect 2361 6265 2415 6291
rect 2535 6291 2637 6385
tri 2637 6291 2735 6389 sw
tri 2735 6291 2833 6389 ne
rect 2833 6385 3187 6389
rect 2833 6291 2965 6385
rect 2535 6265 2735 6291
rect 2361 6213 2735 6265
tri 2735 6213 2813 6291 sw
tri 2833 6213 2911 6291 ne
rect 2911 6265 2965 6291
rect 3085 6291 3187 6385
tri 3187 6291 3285 6389 sw
tri 3285 6291 3383 6389 ne
rect 3383 6385 3737 6389
rect 3383 6291 3515 6385
rect 3085 6265 3285 6291
rect 2911 6213 3285 6265
tri 3285 6213 3363 6291 sw
tri 3383 6213 3461 6291 ne
rect 3461 6265 3515 6291
rect 3635 6291 3737 6385
tri 3737 6291 3835 6389 sw
tri 3835 6291 3933 6389 ne
rect 3933 6385 4287 6389
rect 3933 6291 4065 6385
rect 3635 6265 3835 6291
rect 3461 6213 3835 6265
tri 3835 6213 3913 6291 sw
tri 3933 6213 4011 6291 ne
rect 4011 6265 4065 6291
rect 4185 6291 4287 6385
tri 4287 6291 4385 6389 sw
tri 4385 6291 4483 6389 ne
rect 4483 6385 4837 6389
rect 4483 6291 4615 6385
rect 4185 6265 4385 6291
rect 4011 6213 4385 6265
tri 4385 6213 4463 6291 sw
tri 4483 6213 4561 6291 ne
rect 4561 6265 4615 6291
rect 4735 6291 4837 6385
tri 4837 6291 4935 6389 sw
tri 4935 6291 5033 6389 ne
rect 5033 6385 5387 6389
rect 5033 6291 5165 6385
rect 4735 6265 4935 6291
rect 4561 6213 4935 6265
tri 4935 6213 5013 6291 sw
tri 5033 6213 5111 6291 ne
rect 5111 6265 5165 6291
rect 5285 6291 5387 6385
tri 5387 6291 5485 6389 sw
tri 5485 6291 5583 6389 ne
rect 5583 6385 5937 6389
rect 5583 6291 5715 6385
rect 5285 6265 5485 6291
rect 5111 6213 5485 6265
tri 5485 6213 5563 6291 sw
tri 5583 6213 5661 6291 ne
rect 5661 6265 5715 6291
rect 5835 6291 5937 6385
tri 5937 6291 6035 6389 sw
tri 6035 6291 6133 6389 ne
rect 6133 6385 6487 6389
rect 6133 6291 6265 6385
rect 5835 6265 6035 6291
rect 5661 6213 6035 6265
tri 6035 6213 6113 6291 sw
tri 6133 6213 6211 6291 ne
rect 6211 6265 6265 6291
rect 6385 6291 6487 6385
tri 6487 6291 6585 6389 sw
tri 6585 6291 6683 6389 ne
rect 6683 6385 7037 6389
rect 6683 6291 6815 6385
rect 6385 6265 6585 6291
rect 6211 6213 6585 6265
tri 6585 6213 6663 6291 sw
tri 6683 6213 6761 6291 ne
rect 6761 6265 6815 6291
rect 6935 6291 7037 6385
tri 7037 6291 7135 6389 sw
tri 7135 6291 7233 6389 ne
rect 7233 6385 7587 6389
rect 7233 6291 7365 6385
rect 6935 6265 7135 6291
rect 6761 6213 7135 6265
tri 7135 6213 7213 6291 sw
tri 7233 6213 7311 6291 ne
rect 7311 6265 7365 6291
rect 7485 6291 7587 6385
tri 7587 6291 7685 6389 sw
tri 7685 6291 7783 6389 ne
rect 7783 6385 8137 6389
rect 7783 6291 7915 6385
rect 7485 6265 7685 6291
rect 7311 6213 7685 6265
tri 7685 6213 7763 6291 sw
tri 7783 6213 7861 6291 ne
rect 7861 6265 7915 6291
rect 8035 6291 8137 6385
tri 8137 6291 8235 6389 sw
tri 8235 6291 8333 6389 ne
rect 8333 6385 8687 6389
rect 8333 6291 8465 6385
rect 8035 6265 8235 6291
rect 7861 6213 8235 6265
tri 8235 6213 8313 6291 sw
tri 8333 6213 8411 6291 ne
rect 8411 6265 8465 6291
rect 8585 6291 8687 6385
tri 8687 6291 8785 6389 sw
tri 8785 6291 8883 6389 ne
rect 8883 6385 9237 6389
rect 8883 6291 9015 6385
rect 8585 6265 8785 6291
rect 8411 6213 8785 6265
tri 8785 6213 8863 6291 sw
tri 8883 6213 8961 6291 ne
rect 8961 6265 9015 6291
rect 9135 6291 9237 6385
tri 9237 6291 9335 6389 sw
tri 9335 6291 9433 6389 ne
rect 9433 6385 9787 6389
rect 9433 6291 9565 6385
rect 9135 6265 9335 6291
rect 8961 6213 9335 6265
tri 9335 6213 9413 6291 sw
tri 9433 6213 9511 6291 ne
rect 9511 6265 9565 6291
rect 9685 6291 9787 6385
tri 9787 6291 9885 6389 sw
tri 9885 6291 9983 6389 ne
rect 9983 6385 10337 6389
rect 9983 6291 10115 6385
rect 9685 6265 9885 6291
rect 9511 6213 9885 6265
tri 9885 6213 9963 6291 sw
tri 9983 6213 10061 6291 ne
rect 10061 6265 10115 6291
rect 10235 6291 10337 6385
tri 10337 6291 10435 6389 sw
tri 10435 6291 10533 6389 ne
rect 10533 6385 10887 6389
rect 10533 6291 10665 6385
rect 10235 6265 10435 6291
rect 10061 6213 10435 6265
tri 10435 6213 10513 6291 sw
tri 10533 6213 10611 6291 ne
rect 10611 6265 10665 6291
rect 10785 6291 10887 6385
tri 10887 6291 10985 6389 sw
tri 10985 6291 11083 6389 ne
rect 11083 6385 11437 6389
rect 11083 6291 11215 6385
rect 10785 6265 10985 6291
rect 10611 6213 10985 6265
tri 10985 6213 11063 6291 sw
tri 11083 6213 11161 6291 ne
rect 11161 6265 11215 6291
rect 11335 6291 11437 6385
tri 11437 6291 11535 6389 sw
tri 11535 6291 11633 6389 ne
rect 11633 6385 11987 6389
rect 11633 6291 11765 6385
rect 11335 6265 11535 6291
rect 11161 6213 11535 6265
tri 11535 6213 11613 6291 sw
tri 11633 6213 11711 6291 ne
rect 11711 6265 11765 6291
rect 11885 6291 11987 6385
tri 11987 6291 12085 6389 sw
tri 12085 6291 12183 6389 ne
rect 12183 6385 12537 6389
rect 12183 6291 12315 6385
rect 11885 6265 12085 6291
rect 11711 6213 12085 6265
tri 12085 6213 12163 6291 sw
tri 12183 6213 12261 6291 ne
rect 12261 6265 12315 6291
rect 12435 6291 12537 6385
tri 12537 6291 12635 6389 sw
tri 12635 6291 12733 6389 ne
rect 12733 6385 13087 6389
rect 12733 6291 12865 6385
rect 12435 6265 12635 6291
rect 12261 6213 12635 6265
tri 12635 6213 12713 6291 sw
tri 12733 6213 12811 6291 ne
rect 12811 6265 12865 6291
rect 12985 6291 13087 6385
tri 13087 6291 13185 6389 sw
tri 13185 6291 13283 6389 ne
rect 13283 6385 13637 6389
rect 13283 6291 13415 6385
rect 12985 6265 13185 6291
rect 12811 6213 13185 6265
tri 13185 6213 13263 6291 sw
tri 13283 6213 13361 6291 ne
rect 13361 6265 13415 6291
rect 13535 6291 13637 6385
tri 13637 6291 13735 6389 sw
tri 13735 6291 13833 6389 ne
rect 13833 6385 14187 6389
rect 13833 6291 13965 6385
rect 13535 6265 13735 6291
rect 13361 6213 13735 6265
tri 13735 6213 13813 6291 sw
tri 13833 6213 13911 6291 ne
rect 13911 6265 13965 6291
rect 14085 6291 14187 6385
tri 14187 6291 14285 6389 sw
tri 14285 6291 14383 6389 ne
rect 14383 6385 14737 6389
rect 14383 6291 14515 6385
rect 14085 6265 14285 6291
rect 13911 6213 14285 6265
tri 14285 6213 14363 6291 sw
tri 14383 6213 14461 6291 ne
rect 14461 6265 14515 6291
rect 14635 6291 14737 6385
tri 14737 6291 14835 6389 sw
tri 14835 6291 14933 6389 ne
rect 14933 6385 15287 6389
rect 14933 6291 15065 6385
rect 14635 6265 14835 6291
rect 14461 6213 14835 6265
tri 14835 6213 14913 6291 sw
tri 14933 6213 15011 6291 ne
rect 15011 6265 15065 6291
rect 15185 6291 15287 6385
tri 15287 6291 15385 6389 sw
tri 15385 6291 15483 6389 ne
rect 15483 6385 15837 6389
rect 15483 6291 15615 6385
rect 15185 6265 15385 6291
rect 15011 6213 15385 6265
tri 15385 6213 15463 6291 sw
tri 15483 6213 15561 6291 ne
rect 15561 6265 15615 6291
rect 15735 6291 15837 6385
tri 15837 6291 15935 6389 sw
tri 15935 6291 16033 6389 ne
rect 16033 6385 16387 6389
rect 16033 6291 16165 6385
rect 15735 6265 15935 6291
rect 15561 6213 15935 6265
tri 15935 6213 16013 6291 sw
tri 16033 6213 16111 6291 ne
rect 16111 6265 16165 6291
rect 16285 6291 16387 6385
tri 16387 6291 16485 6389 sw
tri 16485 6291 16583 6389 ne
rect 16583 6385 16937 6389
rect 16583 6291 16715 6385
rect 16285 6265 16485 6291
rect 16111 6213 16485 6265
tri 16485 6213 16563 6291 sw
tri 16583 6213 16661 6291 ne
rect 16661 6265 16715 6291
rect 16835 6291 16937 6385
tri 16937 6291 17035 6389 sw
tri 17035 6291 17133 6389 ne
rect 17133 6385 17487 6389
rect 17133 6291 17265 6385
rect 16835 6265 17035 6291
rect 16661 6213 17035 6265
tri 17035 6213 17113 6291 sw
tri 17133 6213 17211 6291 ne
rect 17211 6265 17265 6291
rect 17385 6291 17487 6385
tri 17487 6291 17585 6389 sw
tri 17585 6291 17683 6389 ne
rect 17683 6385 18037 6389
rect 17683 6291 17815 6385
rect 17385 6265 17585 6291
rect 17211 6213 17585 6265
tri 17585 6213 17663 6291 sw
tri 17683 6213 17761 6291 ne
rect 17761 6265 17815 6291
rect 17935 6291 18037 6385
tri 18037 6291 18135 6389 sw
tri 18135 6291 18233 6389 ne
rect 18233 6385 18587 6389
rect 18233 6291 18365 6385
rect 17935 6265 18135 6291
rect 17761 6213 18135 6265
tri 18135 6213 18213 6291 sw
tri 18233 6213 18311 6291 ne
rect 18311 6265 18365 6291
rect 18485 6291 18587 6385
tri 18587 6291 18685 6389 sw
tri 18685 6291 18783 6389 ne
rect 18783 6385 19137 6389
rect 18783 6291 18915 6385
rect 18485 6265 18685 6291
rect 18311 6213 18685 6265
tri 18685 6213 18763 6291 sw
tri 18783 6213 18861 6291 ne
rect 18861 6265 18915 6291
rect 19035 6291 19137 6385
tri 19137 6291 19235 6389 sw
tri 19235 6291 19333 6389 ne
rect 19333 6385 21800 6389
rect 19333 6291 19465 6385
rect 19035 6265 19235 6291
rect 18861 6213 19235 6265
tri 19235 6213 19313 6291 sw
tri 19333 6213 19411 6291 ne
rect 19411 6265 19465 6291
rect 19585 6265 21800 6385
rect 19411 6213 21800 6265
rect 211 6163 613 6213
rect -500 6113 113 6163
tri 113 6113 163 6163 sw
tri 211 6113 261 6163 ne
rect 261 6133 613 6163
tri 613 6133 693 6213 sw
tri 711 6133 791 6213 ne
rect 791 6133 1163 6213
tri 1163 6133 1243 6213 sw
tri 1261 6133 1341 6213 ne
rect 1341 6133 1713 6213
tri 1713 6133 1793 6213 sw
tri 1811 6133 1891 6213 ne
rect 1891 6133 2263 6213
tri 2263 6133 2343 6213 sw
tri 2361 6133 2441 6213 ne
rect 2441 6133 2813 6213
tri 2813 6133 2893 6213 sw
tri 2911 6133 2991 6213 ne
rect 2991 6133 3363 6213
tri 3363 6133 3443 6213 sw
tri 3461 6133 3541 6213 ne
rect 3541 6133 3913 6213
tri 3913 6133 3993 6213 sw
tri 4011 6133 4091 6213 ne
rect 4091 6133 4463 6213
tri 4463 6133 4543 6213 sw
tri 4561 6133 4641 6213 ne
rect 4641 6133 5013 6213
tri 5013 6133 5093 6213 sw
tri 5111 6133 5191 6213 ne
rect 5191 6133 5563 6213
tri 5563 6133 5643 6213 sw
tri 5661 6133 5741 6213 ne
rect 5741 6133 6113 6213
tri 6113 6133 6193 6213 sw
tri 6211 6133 6291 6213 ne
rect 6291 6133 6663 6213
tri 6663 6133 6743 6213 sw
tri 6761 6133 6841 6213 ne
rect 6841 6133 7213 6213
tri 7213 6133 7293 6213 sw
tri 7311 6133 7391 6213 ne
rect 7391 6133 7763 6213
tri 7763 6133 7843 6213 sw
tri 7861 6133 7941 6213 ne
rect 7941 6133 8313 6213
tri 8313 6133 8393 6213 sw
tri 8411 6133 8491 6213 ne
rect 8491 6133 8863 6213
tri 8863 6133 8943 6213 sw
tri 8961 6133 9041 6213 ne
rect 9041 6133 9413 6213
tri 9413 6133 9493 6213 sw
tri 9511 6133 9591 6213 ne
rect 9591 6133 9963 6213
tri 9963 6133 10043 6213 sw
tri 10061 6133 10141 6213 ne
rect 10141 6133 10513 6213
tri 10513 6133 10593 6213 sw
tri 10611 6133 10691 6213 ne
rect 10691 6133 11063 6213
tri 11063 6133 11143 6213 sw
tri 11161 6133 11241 6213 ne
rect 11241 6133 11613 6213
tri 11613 6133 11693 6213 sw
tri 11711 6133 11791 6213 ne
rect 11791 6133 12163 6213
tri 12163 6133 12243 6213 sw
tri 12261 6133 12341 6213 ne
rect 12341 6133 12713 6213
tri 12713 6133 12793 6213 sw
tri 12811 6133 12891 6213 ne
rect 12891 6133 13263 6213
tri 13263 6133 13343 6213 sw
tri 13361 6133 13441 6213 ne
rect 13441 6133 13813 6213
tri 13813 6133 13893 6213 sw
tri 13911 6133 13991 6213 ne
rect 13991 6133 14363 6213
tri 14363 6133 14443 6213 sw
tri 14461 6133 14541 6213 ne
rect 14541 6133 14913 6213
tri 14913 6133 14993 6213 sw
tri 15011 6133 15091 6213 ne
rect 15091 6133 15463 6213
tri 15463 6133 15543 6213 sw
tri 15561 6133 15641 6213 ne
rect 15641 6133 16013 6213
tri 16013 6133 16093 6213 sw
tri 16111 6133 16191 6213 ne
rect 16191 6133 16563 6213
tri 16563 6133 16643 6213 sw
tri 16661 6133 16741 6213 ne
rect 16741 6133 17113 6213
tri 17113 6133 17193 6213 sw
tri 17211 6133 17291 6213 ne
rect 17291 6133 17663 6213
tri 17663 6133 17743 6213 sw
tri 17761 6133 17841 6213 ne
rect 17841 6133 18213 6213
tri 18213 6133 18293 6213 sw
tri 18311 6133 18391 6213 ne
rect 18391 6133 18763 6213
tri 18763 6133 18843 6213 sw
tri 18861 6133 18941 6213 ne
rect 18941 6133 19313 6213
tri 19313 6133 19393 6213 sw
tri 19411 6133 19491 6213 ne
rect 19491 6133 20100 6213
rect 261 6113 693 6133
rect -500 6035 163 6113
tri 163 6035 241 6113 sw
tri 261 6035 339 6113 ne
rect 339 6035 693 6113
tri 693 6035 791 6133 sw
tri 791 6035 889 6133 ne
rect 889 6035 1243 6133
tri 1243 6035 1341 6133 sw
tri 1341 6035 1439 6133 ne
rect 1439 6035 1793 6133
tri 1793 6035 1891 6133 sw
tri 1891 6035 1989 6133 ne
rect 1989 6035 2343 6133
tri 2343 6035 2441 6133 sw
tri 2441 6035 2539 6133 ne
rect 2539 6035 2893 6133
tri 2893 6035 2991 6133 sw
tri 2991 6035 3089 6133 ne
rect 3089 6035 3443 6133
tri 3443 6035 3541 6133 sw
tri 3541 6035 3639 6133 ne
rect 3639 6035 3993 6133
tri 3993 6035 4091 6133 sw
tri 4091 6035 4189 6133 ne
rect 4189 6035 4543 6133
tri 4543 6035 4641 6133 sw
tri 4641 6035 4739 6133 ne
rect 4739 6035 5093 6133
tri 5093 6035 5191 6133 sw
tri 5191 6035 5289 6133 ne
rect 5289 6035 5643 6133
tri 5643 6035 5741 6133 sw
tri 5741 6035 5839 6133 ne
rect 5839 6035 6193 6133
tri 6193 6035 6291 6133 sw
tri 6291 6035 6389 6133 ne
rect 6389 6035 6743 6133
tri 6743 6035 6841 6133 sw
tri 6841 6035 6939 6133 ne
rect 6939 6035 7293 6133
tri 7293 6035 7391 6133 sw
tri 7391 6035 7489 6133 ne
rect 7489 6035 7843 6133
tri 7843 6035 7941 6133 sw
tri 7941 6035 8039 6133 ne
rect 8039 6035 8393 6133
tri 8393 6035 8491 6133 sw
tri 8491 6035 8589 6133 ne
rect 8589 6035 8943 6133
tri 8943 6035 9041 6133 sw
tri 9041 6035 9139 6133 ne
rect 9139 6035 9493 6133
tri 9493 6035 9591 6133 sw
tri 9591 6035 9689 6133 ne
rect 9689 6035 10043 6133
tri 10043 6035 10141 6133 sw
tri 10141 6035 10239 6133 ne
rect 10239 6035 10593 6133
tri 10593 6035 10691 6133 sw
tri 10691 6035 10789 6133 ne
rect 10789 6035 11143 6133
tri 11143 6035 11241 6133 sw
tri 11241 6035 11339 6133 ne
rect 11339 6035 11693 6133
tri 11693 6035 11791 6133 sw
tri 11791 6035 11889 6133 ne
rect 11889 6035 12243 6133
tri 12243 6035 12341 6133 sw
tri 12341 6035 12439 6133 ne
rect 12439 6035 12793 6133
tri 12793 6035 12891 6133 sw
tri 12891 6035 12989 6133 ne
rect 12989 6035 13343 6133
tri 13343 6035 13441 6133 sw
tri 13441 6035 13539 6133 ne
rect 13539 6035 13893 6133
tri 13893 6035 13991 6133 sw
tri 13991 6035 14089 6133 ne
rect 14089 6035 14443 6133
tri 14443 6035 14541 6133 sw
tri 14541 6035 14639 6133 ne
rect 14639 6035 14993 6133
tri 14993 6035 15091 6133 sw
tri 15091 6035 15189 6133 ne
rect 15189 6035 15543 6133
tri 15543 6035 15641 6133 sw
tri 15641 6035 15739 6133 ne
rect 15739 6035 16093 6133
tri 16093 6035 16191 6133 sw
tri 16191 6035 16289 6133 ne
rect 16289 6035 16643 6133
tri 16643 6035 16741 6133 sw
tri 16741 6035 16839 6133 ne
rect 16839 6035 17193 6133
tri 17193 6035 17291 6133 sw
tri 17291 6035 17389 6133 ne
rect 17389 6035 17743 6133
tri 17743 6035 17841 6133 sw
tri 17841 6035 17939 6133 ne
rect 17939 6035 18293 6133
tri 18293 6035 18391 6133 sw
tri 18391 6035 18489 6133 ne
rect 18489 6035 18843 6133
tri 18843 6035 18941 6133 sw
tri 18941 6035 19039 6133 ne
rect 19039 6035 19393 6133
tri 19393 6035 19491 6133 sw
tri 19491 6035 19589 6133 ne
rect 19589 6113 20100 6133
rect 20200 6113 21800 6213
rect 19589 6035 21800 6113
rect -500 5987 241 6035
rect -500 5887 -400 5987
rect -300 5937 241 5987
tri 241 5937 339 6035 sw
tri 339 5937 437 6035 ne
rect 437 5937 791 6035
tri 791 5937 889 6035 sw
tri 889 5937 987 6035 ne
rect 987 5937 1341 6035
tri 1341 5937 1439 6035 sw
tri 1439 5937 1537 6035 ne
rect 1537 5937 1891 6035
tri 1891 5937 1989 6035 sw
tri 1989 5937 2087 6035 ne
rect 2087 5937 2441 6035
tri 2441 5937 2539 6035 sw
tri 2539 5937 2637 6035 ne
rect 2637 5937 2991 6035
tri 2991 5937 3089 6035 sw
tri 3089 5937 3187 6035 ne
rect 3187 5937 3541 6035
tri 3541 5937 3639 6035 sw
tri 3639 5937 3737 6035 ne
rect 3737 5937 4091 6035
tri 4091 5937 4189 6035 sw
tri 4189 5937 4287 6035 ne
rect 4287 5937 4641 6035
tri 4641 5937 4739 6035 sw
tri 4739 5937 4837 6035 ne
rect 4837 5937 5191 6035
tri 5191 5937 5289 6035 sw
tri 5289 5937 5387 6035 ne
rect 5387 5937 5741 6035
tri 5741 5937 5839 6035 sw
tri 5839 5937 5937 6035 ne
rect 5937 5937 6291 6035
tri 6291 5937 6389 6035 sw
tri 6389 5937 6487 6035 ne
rect 6487 5937 6841 6035
tri 6841 5937 6939 6035 sw
tri 6939 5937 7037 6035 ne
rect 7037 5937 7391 6035
tri 7391 5937 7489 6035 sw
tri 7489 5937 7587 6035 ne
rect 7587 5937 7941 6035
tri 7941 5937 8039 6035 sw
tri 8039 5937 8137 6035 ne
rect 8137 5937 8491 6035
tri 8491 5937 8589 6035 sw
tri 8589 5937 8687 6035 ne
rect 8687 5937 9041 6035
tri 9041 5937 9139 6035 sw
tri 9139 5937 9237 6035 ne
rect 9237 5937 9591 6035
tri 9591 5937 9689 6035 sw
tri 9689 5937 9787 6035 ne
rect 9787 5937 10141 6035
tri 10141 5937 10239 6035 sw
tri 10239 5937 10337 6035 ne
rect 10337 5937 10691 6035
tri 10691 5937 10789 6035 sw
tri 10789 5937 10887 6035 ne
rect 10887 5937 11241 6035
tri 11241 5937 11339 6035 sw
tri 11339 5937 11437 6035 ne
rect 11437 5937 11791 6035
tri 11791 5937 11889 6035 sw
tri 11889 5937 11987 6035 ne
rect 11987 5937 12341 6035
tri 12341 5937 12439 6035 sw
tri 12439 5937 12537 6035 ne
rect 12537 5937 12891 6035
tri 12891 5937 12989 6035 sw
tri 12989 5937 13087 6035 ne
rect 13087 5937 13441 6035
tri 13441 5937 13539 6035 sw
tri 13539 5937 13637 6035 ne
rect 13637 5937 13991 6035
tri 13991 5937 14089 6035 sw
tri 14089 5937 14187 6035 ne
rect 14187 5937 14541 6035
tri 14541 5937 14639 6035 sw
tri 14639 5937 14737 6035 ne
rect 14737 5937 15091 6035
tri 15091 5937 15189 6035 sw
tri 15189 5937 15287 6035 ne
rect 15287 5937 15641 6035
tri 15641 5937 15739 6035 sw
tri 15739 5937 15837 6035 ne
rect 15837 5937 16191 6035
tri 16191 5937 16289 6035 sw
tri 16289 5937 16387 6035 ne
rect 16387 5937 16741 6035
tri 16741 5937 16839 6035 sw
tri 16839 5937 16937 6035 ne
rect 16937 5937 17291 6035
tri 17291 5937 17389 6035 sw
tri 17389 5937 17487 6035 ne
rect 17487 5937 17841 6035
tri 17841 5937 17939 6035 sw
tri 17939 5937 18037 6035 ne
rect 18037 5937 18391 6035
tri 18391 5937 18489 6035 sw
tri 18489 5937 18587 6035 ne
rect 18587 5937 18941 6035
tri 18941 5937 19039 6035 sw
tri 19039 5937 19137 6035 ne
rect 19137 5937 19491 6035
tri 19491 5937 19589 6035 sw
tri 19589 5937 19687 6035 ne
rect 19687 5937 21800 6035
rect -300 5887 339 5937
rect -500 5839 339 5887
tri 339 5839 437 5937 sw
tri 437 5839 535 5937 ne
rect 535 5839 889 5937
tri 889 5839 987 5937 sw
tri 987 5839 1085 5937 ne
rect 1085 5839 1439 5937
tri 1439 5839 1537 5937 sw
tri 1537 5839 1635 5937 ne
rect 1635 5839 1989 5937
tri 1989 5839 2087 5937 sw
tri 2087 5839 2185 5937 ne
rect 2185 5839 2539 5937
tri 2539 5839 2637 5937 sw
tri 2637 5839 2735 5937 ne
rect 2735 5839 3089 5937
tri 3089 5839 3187 5937 sw
tri 3187 5839 3285 5937 ne
rect 3285 5839 3639 5937
tri 3639 5839 3737 5937 sw
tri 3737 5839 3835 5937 ne
rect 3835 5839 4189 5937
tri 4189 5839 4287 5937 sw
tri 4287 5839 4385 5937 ne
rect 4385 5839 4739 5937
tri 4739 5839 4837 5937 sw
tri 4837 5839 4935 5937 ne
rect 4935 5839 5289 5937
tri 5289 5839 5387 5937 sw
tri 5387 5839 5485 5937 ne
rect 5485 5839 5839 5937
tri 5839 5839 5937 5937 sw
tri 5937 5839 6035 5937 ne
rect 6035 5839 6389 5937
tri 6389 5839 6487 5937 sw
tri 6487 5839 6585 5937 ne
rect 6585 5839 6939 5937
tri 6939 5839 7037 5937 sw
tri 7037 5839 7135 5937 ne
rect 7135 5839 7489 5937
tri 7489 5839 7587 5937 sw
tri 7587 5839 7685 5937 ne
rect 7685 5839 8039 5937
tri 8039 5839 8137 5937 sw
tri 8137 5839 8235 5937 ne
rect 8235 5839 8589 5937
tri 8589 5839 8687 5937 sw
tri 8687 5839 8785 5937 ne
rect 8785 5839 9139 5937
tri 9139 5839 9237 5937 sw
tri 9237 5839 9335 5937 ne
rect 9335 5839 9689 5937
tri 9689 5839 9787 5937 sw
tri 9787 5839 9885 5937 ne
rect 9885 5839 10239 5937
tri 10239 5839 10337 5937 sw
tri 10337 5839 10435 5937 ne
rect 10435 5839 10789 5937
tri 10789 5839 10887 5937 sw
tri 10887 5839 10985 5937 ne
rect 10985 5839 11339 5937
tri 11339 5839 11437 5937 sw
tri 11437 5839 11535 5937 ne
rect 11535 5839 11889 5937
tri 11889 5839 11987 5937 sw
tri 11987 5839 12085 5937 ne
rect 12085 5839 12439 5937
tri 12439 5839 12537 5937 sw
tri 12537 5839 12635 5937 ne
rect 12635 5839 12989 5937
tri 12989 5839 13087 5937 sw
tri 13087 5839 13185 5937 ne
rect 13185 5839 13539 5937
tri 13539 5839 13637 5937 sw
tri 13637 5839 13735 5937 ne
rect 13735 5839 14089 5937
tri 14089 5839 14187 5937 sw
tri 14187 5839 14285 5937 ne
rect 14285 5839 14639 5937
tri 14639 5839 14737 5937 sw
tri 14737 5839 14835 5937 ne
rect 14835 5839 15189 5937
tri 15189 5839 15287 5937 sw
tri 15287 5839 15385 5937 ne
rect 15385 5839 15739 5937
tri 15739 5839 15837 5937 sw
tri 15837 5839 15935 5937 ne
rect 15935 5839 16289 5937
tri 16289 5839 16387 5937 sw
tri 16387 5839 16485 5937 ne
rect 16485 5839 16839 5937
tri 16839 5839 16937 5937 sw
tri 16937 5839 17035 5937 ne
rect 17035 5839 17389 5937
tri 17389 5839 17487 5937 sw
tri 17487 5839 17585 5937 ne
rect 17585 5839 17939 5937
tri 17939 5839 18037 5937 sw
tri 18037 5839 18135 5937 ne
rect 18135 5839 18489 5937
tri 18489 5839 18587 5937 sw
tri 18587 5839 18685 5937 ne
rect 18685 5839 19039 5937
tri 19039 5839 19137 5937 sw
tri 19137 5839 19235 5937 ne
rect 19235 5839 19589 5937
tri 19589 5839 19687 5937 sw
rect -500 5835 437 5839
rect -500 5715 215 5835
rect 335 5741 437 5835
tri 437 5741 535 5839 sw
tri 535 5741 633 5839 ne
rect 633 5835 987 5839
rect 633 5741 765 5835
rect 335 5715 535 5741
rect -500 5711 535 5715
tri 535 5711 565 5741 sw
tri 633 5711 663 5741 ne
rect 663 5715 765 5741
rect 885 5741 987 5835
tri 987 5741 1085 5839 sw
tri 1085 5741 1183 5839 ne
rect 1183 5835 1537 5839
rect 1183 5741 1315 5835
rect 885 5715 1085 5741
rect 663 5711 1085 5715
tri 1085 5711 1115 5741 sw
tri 1183 5711 1213 5741 ne
rect 1213 5715 1315 5741
rect 1435 5741 1537 5835
tri 1537 5741 1635 5839 sw
tri 1635 5741 1733 5839 ne
rect 1733 5835 2087 5839
rect 1733 5741 1865 5835
rect 1435 5715 1635 5741
rect 1213 5711 1635 5715
tri 1635 5711 1665 5741 sw
tri 1733 5711 1763 5741 ne
rect 1763 5715 1865 5741
rect 1985 5741 2087 5835
tri 2087 5741 2185 5839 sw
tri 2185 5741 2283 5839 ne
rect 2283 5835 2637 5839
rect 2283 5741 2415 5835
rect 1985 5715 2185 5741
rect 1763 5711 2185 5715
tri 2185 5711 2215 5741 sw
tri 2283 5711 2313 5741 ne
rect 2313 5715 2415 5741
rect 2535 5741 2637 5835
tri 2637 5741 2735 5839 sw
tri 2735 5741 2833 5839 ne
rect 2833 5835 3187 5839
rect 2833 5741 2965 5835
rect 2535 5715 2735 5741
rect 2313 5711 2735 5715
tri 2735 5711 2765 5741 sw
tri 2833 5711 2863 5741 ne
rect 2863 5715 2965 5741
rect 3085 5741 3187 5835
tri 3187 5741 3285 5839 sw
tri 3285 5741 3383 5839 ne
rect 3383 5835 3737 5839
rect 3383 5741 3515 5835
rect 3085 5715 3285 5741
rect 2863 5711 3285 5715
tri 3285 5711 3315 5741 sw
tri 3383 5711 3413 5741 ne
rect 3413 5715 3515 5741
rect 3635 5741 3737 5835
tri 3737 5741 3835 5839 sw
tri 3835 5741 3933 5839 ne
rect 3933 5835 4287 5839
rect 3933 5741 4065 5835
rect 3635 5715 3835 5741
rect 3413 5711 3835 5715
tri 3835 5711 3865 5741 sw
tri 3933 5711 3963 5741 ne
rect 3963 5715 4065 5741
rect 4185 5741 4287 5835
tri 4287 5741 4385 5839 sw
tri 4385 5741 4483 5839 ne
rect 4483 5835 4837 5839
rect 4483 5741 4615 5835
rect 4185 5715 4385 5741
rect 3963 5711 4385 5715
tri 4385 5711 4415 5741 sw
tri 4483 5711 4513 5741 ne
rect 4513 5715 4615 5741
rect 4735 5741 4837 5835
tri 4837 5741 4935 5839 sw
tri 4935 5741 5033 5839 ne
rect 5033 5835 5387 5839
rect 5033 5741 5165 5835
rect 4735 5715 4935 5741
rect 4513 5711 4935 5715
tri 4935 5711 4965 5741 sw
tri 5033 5711 5063 5741 ne
rect 5063 5715 5165 5741
rect 5285 5741 5387 5835
tri 5387 5741 5485 5839 sw
tri 5485 5741 5583 5839 ne
rect 5583 5835 5937 5839
rect 5583 5741 5715 5835
rect 5285 5715 5485 5741
rect 5063 5711 5485 5715
tri 5485 5711 5515 5741 sw
tri 5583 5711 5613 5741 ne
rect 5613 5715 5715 5741
rect 5835 5741 5937 5835
tri 5937 5741 6035 5839 sw
tri 6035 5741 6133 5839 ne
rect 6133 5835 6487 5839
rect 6133 5741 6265 5835
rect 5835 5715 6035 5741
rect 5613 5711 6035 5715
tri 6035 5711 6065 5741 sw
tri 6133 5711 6163 5741 ne
rect 6163 5715 6265 5741
rect 6385 5741 6487 5835
tri 6487 5741 6585 5839 sw
tri 6585 5741 6683 5839 ne
rect 6683 5835 7037 5839
rect 6683 5741 6815 5835
rect 6385 5715 6585 5741
rect 6163 5711 6585 5715
tri 6585 5711 6615 5741 sw
tri 6683 5711 6713 5741 ne
rect 6713 5715 6815 5741
rect 6935 5741 7037 5835
tri 7037 5741 7135 5839 sw
tri 7135 5741 7233 5839 ne
rect 7233 5835 7587 5839
rect 7233 5741 7365 5835
rect 6935 5715 7135 5741
rect 6713 5711 7135 5715
tri 7135 5711 7165 5741 sw
tri 7233 5711 7263 5741 ne
rect 7263 5715 7365 5741
rect 7485 5741 7587 5835
tri 7587 5741 7685 5839 sw
tri 7685 5741 7783 5839 ne
rect 7783 5835 8137 5839
rect 7783 5741 7915 5835
rect 7485 5715 7685 5741
rect 7263 5711 7685 5715
tri 7685 5711 7715 5741 sw
tri 7783 5711 7813 5741 ne
rect 7813 5715 7915 5741
rect 8035 5741 8137 5835
tri 8137 5741 8235 5839 sw
tri 8235 5741 8333 5839 ne
rect 8333 5835 8687 5839
rect 8333 5741 8465 5835
rect 8035 5715 8235 5741
rect 7813 5711 8235 5715
tri 8235 5711 8265 5741 sw
tri 8333 5711 8363 5741 ne
rect 8363 5715 8465 5741
rect 8585 5741 8687 5835
tri 8687 5741 8785 5839 sw
tri 8785 5741 8883 5839 ne
rect 8883 5835 9237 5839
rect 8883 5741 9015 5835
rect 8585 5715 8785 5741
rect 8363 5711 8785 5715
tri 8785 5711 8815 5741 sw
tri 8883 5711 8913 5741 ne
rect 8913 5715 9015 5741
rect 9135 5741 9237 5835
tri 9237 5741 9335 5839 sw
tri 9335 5741 9433 5839 ne
rect 9433 5835 9787 5839
rect 9433 5741 9565 5835
rect 9135 5715 9335 5741
rect 8913 5711 9335 5715
tri 9335 5711 9365 5741 sw
tri 9433 5711 9463 5741 ne
rect 9463 5715 9565 5741
rect 9685 5741 9787 5835
tri 9787 5741 9885 5839 sw
tri 9885 5741 9983 5839 ne
rect 9983 5835 10337 5839
rect 9983 5741 10115 5835
rect 9685 5715 9885 5741
rect 9463 5711 9885 5715
tri 9885 5711 9915 5741 sw
tri 9983 5711 10013 5741 ne
rect 10013 5715 10115 5741
rect 10235 5741 10337 5835
tri 10337 5741 10435 5839 sw
tri 10435 5741 10533 5839 ne
rect 10533 5835 10887 5839
rect 10533 5741 10665 5835
rect 10235 5715 10435 5741
rect 10013 5711 10435 5715
tri 10435 5711 10465 5741 sw
tri 10533 5711 10563 5741 ne
rect 10563 5715 10665 5741
rect 10785 5741 10887 5835
tri 10887 5741 10985 5839 sw
tri 10985 5741 11083 5839 ne
rect 11083 5835 11437 5839
rect 11083 5741 11215 5835
rect 10785 5715 10985 5741
rect 10563 5711 10985 5715
tri 10985 5711 11015 5741 sw
tri 11083 5711 11113 5741 ne
rect 11113 5715 11215 5741
rect 11335 5741 11437 5835
tri 11437 5741 11535 5839 sw
tri 11535 5741 11633 5839 ne
rect 11633 5835 11987 5839
rect 11633 5741 11765 5835
rect 11335 5715 11535 5741
rect 11113 5711 11535 5715
tri 11535 5711 11565 5741 sw
tri 11633 5711 11663 5741 ne
rect 11663 5715 11765 5741
rect 11885 5741 11987 5835
tri 11987 5741 12085 5839 sw
tri 12085 5741 12183 5839 ne
rect 12183 5835 12537 5839
rect 12183 5741 12315 5835
rect 11885 5715 12085 5741
rect 11663 5711 12085 5715
tri 12085 5711 12115 5741 sw
tri 12183 5711 12213 5741 ne
rect 12213 5715 12315 5741
rect 12435 5741 12537 5835
tri 12537 5741 12635 5839 sw
tri 12635 5741 12733 5839 ne
rect 12733 5835 13087 5839
rect 12733 5741 12865 5835
rect 12435 5715 12635 5741
rect 12213 5711 12635 5715
tri 12635 5711 12665 5741 sw
tri 12733 5711 12763 5741 ne
rect 12763 5715 12865 5741
rect 12985 5741 13087 5835
tri 13087 5741 13185 5839 sw
tri 13185 5741 13283 5839 ne
rect 13283 5835 13637 5839
rect 13283 5741 13415 5835
rect 12985 5715 13185 5741
rect 12763 5711 13185 5715
tri 13185 5711 13215 5741 sw
tri 13283 5711 13313 5741 ne
rect 13313 5715 13415 5741
rect 13535 5741 13637 5835
tri 13637 5741 13735 5839 sw
tri 13735 5741 13833 5839 ne
rect 13833 5835 14187 5839
rect 13833 5741 13965 5835
rect 13535 5715 13735 5741
rect 13313 5711 13735 5715
tri 13735 5711 13765 5741 sw
tri 13833 5711 13863 5741 ne
rect 13863 5715 13965 5741
rect 14085 5741 14187 5835
tri 14187 5741 14285 5839 sw
tri 14285 5741 14383 5839 ne
rect 14383 5835 14737 5839
rect 14383 5741 14515 5835
rect 14085 5715 14285 5741
rect 13863 5711 14285 5715
tri 14285 5711 14315 5741 sw
tri 14383 5711 14413 5741 ne
rect 14413 5715 14515 5741
rect 14635 5741 14737 5835
tri 14737 5741 14835 5839 sw
tri 14835 5741 14933 5839 ne
rect 14933 5835 15287 5839
rect 14933 5741 15065 5835
rect 14635 5715 14835 5741
rect 14413 5711 14835 5715
tri 14835 5711 14865 5741 sw
tri 14933 5711 14963 5741 ne
rect 14963 5715 15065 5741
rect 15185 5741 15287 5835
tri 15287 5741 15385 5839 sw
tri 15385 5741 15483 5839 ne
rect 15483 5835 15837 5839
rect 15483 5741 15615 5835
rect 15185 5715 15385 5741
rect 14963 5711 15385 5715
tri 15385 5711 15415 5741 sw
tri 15483 5711 15513 5741 ne
rect 15513 5715 15615 5741
rect 15735 5741 15837 5835
tri 15837 5741 15935 5839 sw
tri 15935 5741 16033 5839 ne
rect 16033 5835 16387 5839
rect 16033 5741 16165 5835
rect 15735 5715 15935 5741
rect 15513 5711 15935 5715
tri 15935 5711 15965 5741 sw
tri 16033 5711 16063 5741 ne
rect 16063 5715 16165 5741
rect 16285 5741 16387 5835
tri 16387 5741 16485 5839 sw
tri 16485 5741 16583 5839 ne
rect 16583 5835 16937 5839
rect 16583 5741 16715 5835
rect 16285 5715 16485 5741
rect 16063 5711 16485 5715
tri 16485 5711 16515 5741 sw
tri 16583 5711 16613 5741 ne
rect 16613 5715 16715 5741
rect 16835 5741 16937 5835
tri 16937 5741 17035 5839 sw
tri 17035 5741 17133 5839 ne
rect 17133 5835 17487 5839
rect 17133 5741 17265 5835
rect 16835 5715 17035 5741
rect 16613 5711 17035 5715
tri 17035 5711 17065 5741 sw
tri 17133 5711 17163 5741 ne
rect 17163 5715 17265 5741
rect 17385 5741 17487 5835
tri 17487 5741 17585 5839 sw
tri 17585 5741 17683 5839 ne
rect 17683 5835 18037 5839
rect 17683 5741 17815 5835
rect 17385 5715 17585 5741
rect 17163 5711 17585 5715
tri 17585 5711 17615 5741 sw
tri 17683 5711 17713 5741 ne
rect 17713 5715 17815 5741
rect 17935 5741 18037 5835
tri 18037 5741 18135 5839 sw
tri 18135 5741 18233 5839 ne
rect 18233 5835 18587 5839
rect 18233 5741 18365 5835
rect 17935 5715 18135 5741
rect 17713 5711 18135 5715
tri 18135 5711 18165 5741 sw
tri 18233 5711 18263 5741 ne
rect 18263 5715 18365 5741
rect 18485 5741 18587 5835
tri 18587 5741 18685 5839 sw
tri 18685 5741 18783 5839 ne
rect 18783 5835 19137 5839
rect 18783 5741 18915 5835
rect 18485 5715 18685 5741
rect 18263 5711 18685 5715
tri 18685 5711 18715 5741 sw
tri 18783 5711 18813 5741 ne
rect 18813 5715 18915 5741
rect 19035 5741 19137 5835
tri 19137 5741 19235 5839 sw
tri 19235 5741 19333 5839 ne
rect 19333 5835 20300 5839
rect 19333 5741 19465 5835
rect 19035 5715 19235 5741
rect 18813 5711 19235 5715
tri 19235 5711 19265 5741 sw
tri 19333 5711 19363 5741 ne
rect 19363 5715 19465 5741
rect 19585 5715 20300 5835
rect 19363 5711 20300 5715
tri 113 5613 211 5711 ne
rect 211 5613 565 5711
tri 565 5613 663 5711 sw
tri 663 5613 761 5711 ne
rect 761 5613 1115 5711
tri 1115 5613 1213 5711 sw
tri 1213 5613 1311 5711 ne
rect 1311 5613 1665 5711
tri 1665 5613 1763 5711 sw
tri 1763 5613 1861 5711 ne
rect 1861 5613 2215 5711
tri 2215 5613 2313 5711 sw
tri 2313 5613 2411 5711 ne
rect 2411 5613 2765 5711
tri 2765 5613 2863 5711 sw
tri 2863 5613 2961 5711 ne
rect 2961 5613 3315 5711
tri 3315 5613 3413 5711 sw
tri 3413 5613 3511 5711 ne
rect 3511 5613 3865 5711
tri 3865 5613 3963 5711 sw
tri 3963 5613 4061 5711 ne
rect 4061 5613 4415 5711
tri 4415 5613 4513 5711 sw
tri 4513 5613 4611 5711 ne
rect 4611 5613 4965 5711
tri 4965 5613 5063 5711 sw
tri 5063 5613 5161 5711 ne
rect 5161 5613 5515 5711
tri 5515 5613 5613 5711 sw
tri 5613 5613 5711 5711 ne
rect 5711 5613 6065 5711
tri 6065 5613 6163 5711 sw
tri 6163 5613 6261 5711 ne
rect 6261 5613 6615 5711
tri 6615 5613 6713 5711 sw
tri 6713 5613 6811 5711 ne
rect 6811 5613 7165 5711
tri 7165 5613 7263 5711 sw
tri 7263 5613 7361 5711 ne
rect 7361 5613 7715 5711
tri 7715 5613 7813 5711 sw
tri 7813 5613 7911 5711 ne
rect 7911 5613 8265 5711
tri 8265 5613 8363 5711 sw
tri 8363 5613 8461 5711 ne
rect 8461 5613 8815 5711
tri 8815 5613 8913 5711 sw
tri 8913 5613 9011 5711 ne
rect 9011 5613 9365 5711
tri 9365 5613 9463 5711 sw
tri 9463 5613 9561 5711 ne
rect 9561 5613 9915 5711
tri 9915 5613 10013 5711 sw
tri 10013 5613 10111 5711 ne
rect 10111 5613 10465 5711
tri 10465 5613 10563 5711 sw
tri 10563 5613 10661 5711 ne
rect 10661 5613 11015 5711
tri 11015 5613 11113 5711 sw
tri 11113 5613 11211 5711 ne
rect 11211 5613 11565 5711
tri 11565 5613 11663 5711 sw
tri 11663 5613 11761 5711 ne
rect 11761 5613 12115 5711
tri 12115 5613 12213 5711 sw
tri 12213 5613 12311 5711 ne
rect 12311 5613 12665 5711
tri 12665 5613 12763 5711 sw
tri 12763 5613 12861 5711 ne
rect 12861 5613 13215 5711
tri 13215 5613 13313 5711 sw
tri 13313 5613 13411 5711 ne
rect 13411 5613 13765 5711
tri 13765 5613 13863 5711 sw
tri 13863 5613 13961 5711 ne
rect 13961 5613 14315 5711
tri 14315 5613 14413 5711 sw
tri 14413 5613 14511 5711 ne
rect 14511 5613 14865 5711
tri 14865 5613 14963 5711 sw
tri 14963 5613 15061 5711 ne
rect 15061 5613 15415 5711
tri 15415 5613 15513 5711 sw
tri 15513 5613 15611 5711 ne
rect 15611 5613 15965 5711
tri 15965 5613 16063 5711 sw
tri 16063 5613 16161 5711 ne
rect 16161 5613 16515 5711
tri 16515 5613 16613 5711 sw
tri 16613 5613 16711 5711 ne
rect 16711 5613 17065 5711
tri 17065 5613 17163 5711 sw
tri 17163 5613 17261 5711 ne
rect 17261 5613 17615 5711
tri 17615 5613 17713 5711 sw
tri 17713 5613 17811 5711 ne
rect 17811 5613 18165 5711
tri 18165 5613 18263 5711 sw
tri 18263 5613 18361 5711 ne
rect 18361 5613 18715 5711
tri 18715 5613 18813 5711 sw
tri 18813 5613 18911 5711 ne
rect 18911 5613 19265 5711
tri 19265 5613 19363 5711 sw
tri 19363 5613 19461 5711 ne
rect 19461 5613 20300 5711
rect -2000 5583 113 5613
tri 113 5583 143 5613 sw
tri 211 5583 241 5613 ne
rect 241 5583 663 5613
tri 663 5583 693 5613 sw
tri 761 5583 791 5613 ne
rect 791 5583 1213 5613
tri 1213 5583 1243 5613 sw
tri 1311 5583 1341 5613 ne
rect 1341 5583 1763 5613
tri 1763 5583 1793 5613 sw
tri 1861 5583 1891 5613 ne
rect 1891 5583 2313 5613
tri 2313 5583 2343 5613 sw
tri 2411 5583 2441 5613 ne
rect 2441 5583 2863 5613
tri 2863 5583 2893 5613 sw
tri 2961 5583 2991 5613 ne
rect 2991 5583 3413 5613
tri 3413 5583 3443 5613 sw
tri 3511 5583 3541 5613 ne
rect 3541 5583 3963 5613
tri 3963 5583 3993 5613 sw
tri 4061 5583 4091 5613 ne
rect 4091 5583 4513 5613
tri 4513 5583 4543 5613 sw
tri 4611 5583 4641 5613 ne
rect 4641 5583 5063 5613
tri 5063 5583 5093 5613 sw
tri 5161 5583 5191 5613 ne
rect 5191 5583 5613 5613
tri 5613 5583 5643 5613 sw
tri 5711 5583 5741 5613 ne
rect 5741 5583 6163 5613
tri 6163 5583 6193 5613 sw
tri 6261 5583 6291 5613 ne
rect 6291 5583 6713 5613
tri 6713 5583 6743 5613 sw
tri 6811 5583 6841 5613 ne
rect 6841 5583 7263 5613
tri 7263 5583 7293 5613 sw
tri 7361 5583 7391 5613 ne
rect 7391 5583 7813 5613
tri 7813 5583 7843 5613 sw
tri 7911 5583 7941 5613 ne
rect 7941 5583 8363 5613
tri 8363 5583 8393 5613 sw
tri 8461 5583 8491 5613 ne
rect 8491 5583 8913 5613
tri 8913 5583 8943 5613 sw
tri 9011 5583 9041 5613 ne
rect 9041 5583 9463 5613
tri 9463 5583 9493 5613 sw
tri 9561 5583 9591 5613 ne
rect 9591 5583 10013 5613
tri 10013 5583 10043 5613 sw
tri 10111 5583 10141 5613 ne
rect 10141 5583 10563 5613
tri 10563 5583 10593 5613 sw
tri 10661 5583 10691 5613 ne
rect 10691 5583 11113 5613
tri 11113 5583 11143 5613 sw
tri 11211 5583 11241 5613 ne
rect 11241 5583 11663 5613
tri 11663 5583 11693 5613 sw
tri 11761 5583 11791 5613 ne
rect 11791 5583 12213 5613
tri 12213 5583 12243 5613 sw
tri 12311 5583 12341 5613 ne
rect 12341 5583 12763 5613
tri 12763 5583 12793 5613 sw
tri 12861 5583 12891 5613 ne
rect 12891 5583 13313 5613
tri 13313 5583 13343 5613 sw
tri 13411 5583 13441 5613 ne
rect 13441 5583 13863 5613
tri 13863 5583 13893 5613 sw
tri 13961 5583 13991 5613 ne
rect 13991 5583 14413 5613
tri 14413 5583 14443 5613 sw
tri 14511 5583 14541 5613 ne
rect 14541 5583 14963 5613
tri 14963 5583 14993 5613 sw
tri 15061 5583 15091 5613 ne
rect 15091 5583 15513 5613
tri 15513 5583 15543 5613 sw
tri 15611 5583 15641 5613 ne
rect 15641 5583 16063 5613
tri 16063 5583 16093 5613 sw
tri 16161 5583 16191 5613 ne
rect 16191 5583 16613 5613
tri 16613 5583 16643 5613 sw
tri 16711 5583 16741 5613 ne
rect 16741 5583 17163 5613
tri 17163 5583 17193 5613 sw
tri 17261 5583 17291 5613 ne
rect 17291 5583 17713 5613
tri 17713 5583 17743 5613 sw
tri 17811 5583 17841 5613 ne
rect 17841 5583 18263 5613
tri 18263 5583 18293 5613 sw
tri 18361 5583 18391 5613 ne
rect 18391 5583 18813 5613
tri 18813 5583 18843 5613 sw
tri 18911 5583 18941 5613 ne
rect 18941 5583 19363 5613
tri 19363 5583 19393 5613 sw
tri 19461 5583 19491 5613 ne
rect 19491 5583 20300 5613
rect -2000 5485 143 5583
tri 143 5485 241 5583 sw
tri 241 5485 339 5583 ne
rect 339 5485 693 5583
tri 693 5485 791 5583 sw
tri 791 5485 889 5583 ne
rect 889 5485 1243 5583
tri 1243 5485 1341 5583 sw
tri 1341 5485 1439 5583 ne
rect 1439 5485 1793 5583
tri 1793 5485 1891 5583 sw
tri 1891 5485 1989 5583 ne
rect 1989 5485 2343 5583
tri 2343 5485 2441 5583 sw
tri 2441 5485 2539 5583 ne
rect 2539 5485 2893 5583
tri 2893 5485 2991 5583 sw
tri 2991 5485 3089 5583 ne
rect 3089 5485 3443 5583
tri 3443 5485 3541 5583 sw
tri 3541 5485 3639 5583 ne
rect 3639 5485 3993 5583
tri 3993 5485 4091 5583 sw
tri 4091 5485 4189 5583 ne
rect 4189 5485 4543 5583
tri 4543 5485 4641 5583 sw
tri 4641 5485 4739 5583 ne
rect 4739 5485 5093 5583
tri 5093 5485 5191 5583 sw
tri 5191 5485 5289 5583 ne
rect 5289 5485 5643 5583
tri 5643 5485 5741 5583 sw
tri 5741 5485 5839 5583 ne
rect 5839 5485 6193 5583
tri 6193 5485 6291 5583 sw
tri 6291 5485 6389 5583 ne
rect 6389 5485 6743 5583
tri 6743 5485 6841 5583 sw
tri 6841 5485 6939 5583 ne
rect 6939 5485 7293 5583
tri 7293 5485 7391 5583 sw
tri 7391 5485 7489 5583 ne
rect 7489 5485 7843 5583
tri 7843 5485 7941 5583 sw
tri 7941 5485 8039 5583 ne
rect 8039 5485 8393 5583
tri 8393 5485 8491 5583 sw
tri 8491 5485 8589 5583 ne
rect 8589 5485 8943 5583
tri 8943 5485 9041 5583 sw
tri 9041 5485 9139 5583 ne
rect 9139 5485 9493 5583
tri 9493 5485 9591 5583 sw
tri 9591 5485 9689 5583 ne
rect 9689 5485 10043 5583
tri 10043 5485 10141 5583 sw
tri 10141 5485 10239 5583 ne
rect 10239 5485 10593 5583
tri 10593 5485 10691 5583 sw
tri 10691 5485 10789 5583 ne
rect 10789 5485 11143 5583
tri 11143 5485 11241 5583 sw
tri 11241 5485 11339 5583 ne
rect 11339 5485 11693 5583
tri 11693 5485 11791 5583 sw
tri 11791 5485 11889 5583 ne
rect 11889 5485 12243 5583
tri 12243 5485 12341 5583 sw
tri 12341 5485 12439 5583 ne
rect 12439 5485 12793 5583
tri 12793 5485 12891 5583 sw
tri 12891 5485 12989 5583 ne
rect 12989 5485 13343 5583
tri 13343 5485 13441 5583 sw
tri 13441 5485 13539 5583 ne
rect 13539 5485 13893 5583
tri 13893 5485 13991 5583 sw
tri 13991 5485 14089 5583 ne
rect 14089 5485 14443 5583
tri 14443 5485 14541 5583 sw
tri 14541 5485 14639 5583 ne
rect 14639 5485 14993 5583
tri 14993 5485 15091 5583 sw
tri 15091 5485 15189 5583 ne
rect 15189 5485 15543 5583
tri 15543 5485 15641 5583 sw
tri 15641 5485 15739 5583 ne
rect 15739 5485 16093 5583
tri 16093 5485 16191 5583 sw
tri 16191 5485 16289 5583 ne
rect 16289 5485 16643 5583
tri 16643 5485 16741 5583 sw
tri 16741 5485 16839 5583 ne
rect 16839 5485 17193 5583
tri 17193 5485 17291 5583 sw
tri 17291 5485 17389 5583 ne
rect 17389 5485 17743 5583
tri 17743 5485 17841 5583 sw
tri 17841 5485 17939 5583 ne
rect 17939 5485 18293 5583
tri 18293 5485 18391 5583 sw
tri 18391 5485 18489 5583 ne
rect 18489 5485 18843 5583
tri 18843 5485 18941 5583 sw
tri 18941 5485 19039 5583 ne
rect 19039 5485 19393 5583
tri 19393 5485 19491 5583 sw
tri 19491 5485 19589 5583 ne
rect 19589 5485 20300 5583
rect -2000 5387 241 5485
tri 241 5387 339 5485 sw
tri 339 5387 437 5485 ne
rect 437 5387 791 5485
tri 791 5387 889 5485 sw
tri 889 5387 987 5485 ne
rect 987 5387 1341 5485
tri 1341 5387 1439 5485 sw
tri 1439 5387 1537 5485 ne
rect 1537 5387 1891 5485
tri 1891 5387 1989 5485 sw
tri 1989 5387 2087 5485 ne
rect 2087 5387 2441 5485
tri 2441 5387 2539 5485 sw
tri 2539 5387 2637 5485 ne
rect 2637 5387 2991 5485
tri 2991 5387 3089 5485 sw
tri 3089 5387 3187 5485 ne
rect 3187 5387 3541 5485
tri 3541 5387 3639 5485 sw
tri 3639 5387 3737 5485 ne
rect 3737 5387 4091 5485
tri 4091 5387 4189 5485 sw
tri 4189 5387 4287 5485 ne
rect 4287 5387 4641 5485
tri 4641 5387 4739 5485 sw
tri 4739 5387 4837 5485 ne
rect 4837 5387 5191 5485
tri 5191 5387 5289 5485 sw
tri 5289 5387 5387 5485 ne
rect 5387 5387 5741 5485
tri 5741 5387 5839 5485 sw
tri 5839 5387 5937 5485 ne
rect 5937 5387 6291 5485
tri 6291 5387 6389 5485 sw
tri 6389 5387 6487 5485 ne
rect 6487 5387 6841 5485
tri 6841 5387 6939 5485 sw
tri 6939 5387 7037 5485 ne
rect 7037 5387 7391 5485
tri 7391 5387 7489 5485 sw
tri 7489 5387 7587 5485 ne
rect 7587 5387 7941 5485
tri 7941 5387 8039 5485 sw
tri 8039 5387 8137 5485 ne
rect 8137 5387 8491 5485
tri 8491 5387 8589 5485 sw
tri 8589 5387 8687 5485 ne
rect 8687 5387 9041 5485
tri 9041 5387 9139 5485 sw
tri 9139 5387 9237 5485 ne
rect 9237 5387 9591 5485
tri 9591 5387 9689 5485 sw
tri 9689 5387 9787 5485 ne
rect 9787 5387 10141 5485
tri 10141 5387 10239 5485 sw
tri 10239 5387 10337 5485 ne
rect 10337 5387 10691 5485
tri 10691 5387 10789 5485 sw
tri 10789 5387 10887 5485 ne
rect 10887 5387 11241 5485
tri 11241 5387 11339 5485 sw
tri 11339 5387 11437 5485 ne
rect 11437 5387 11791 5485
tri 11791 5387 11889 5485 sw
tri 11889 5387 11987 5485 ne
rect 11987 5387 12341 5485
tri 12341 5387 12439 5485 sw
tri 12439 5387 12537 5485 ne
rect 12537 5387 12891 5485
tri 12891 5387 12989 5485 sw
tri 12989 5387 13087 5485 ne
rect 13087 5387 13441 5485
tri 13441 5387 13539 5485 sw
tri 13539 5387 13637 5485 ne
rect 13637 5387 13991 5485
tri 13991 5387 14089 5485 sw
tri 14089 5387 14187 5485 ne
rect 14187 5387 14541 5485
tri 14541 5387 14639 5485 sw
tri 14639 5387 14737 5485 ne
rect 14737 5387 15091 5485
tri 15091 5387 15189 5485 sw
tri 15189 5387 15287 5485 ne
rect 15287 5387 15641 5485
tri 15641 5387 15739 5485 sw
tri 15739 5387 15837 5485 ne
rect 15837 5387 16191 5485
tri 16191 5387 16289 5485 sw
tri 16289 5387 16387 5485 ne
rect 16387 5387 16741 5485
tri 16741 5387 16839 5485 sw
tri 16839 5387 16937 5485 ne
rect 16937 5387 17291 5485
tri 17291 5387 17389 5485 sw
tri 17389 5387 17487 5485 ne
rect 17487 5387 17841 5485
tri 17841 5387 17939 5485 sw
tri 17939 5387 18037 5485 ne
rect 18037 5387 18391 5485
tri 18391 5387 18489 5485 sw
tri 18489 5387 18587 5485 ne
rect 18587 5387 18941 5485
tri 18941 5387 19039 5485 sw
tri 19039 5387 19137 5485 ne
rect 19137 5387 19491 5485
tri 19491 5387 19589 5485 sw
tri 19589 5387 19687 5485 ne
rect 19687 5387 20300 5485
rect -2000 5289 339 5387
tri 339 5289 437 5387 sw
tri 437 5289 535 5387 ne
rect 535 5289 889 5387
tri 889 5289 987 5387 sw
tri 987 5289 1085 5387 ne
rect 1085 5289 1439 5387
tri 1439 5289 1537 5387 sw
tri 1537 5289 1635 5387 ne
rect 1635 5289 1989 5387
tri 1989 5289 2087 5387 sw
tri 2087 5289 2185 5387 ne
rect 2185 5289 2539 5387
tri 2539 5289 2637 5387 sw
tri 2637 5289 2735 5387 ne
rect 2735 5289 3089 5387
tri 3089 5289 3187 5387 sw
tri 3187 5289 3285 5387 ne
rect 3285 5289 3639 5387
tri 3639 5289 3737 5387 sw
tri 3737 5289 3835 5387 ne
rect 3835 5289 4189 5387
tri 4189 5289 4287 5387 sw
tri 4287 5289 4385 5387 ne
rect 4385 5289 4739 5387
tri 4739 5289 4837 5387 sw
tri 4837 5289 4935 5387 ne
rect 4935 5289 5289 5387
tri 5289 5289 5387 5387 sw
tri 5387 5289 5485 5387 ne
rect 5485 5289 5839 5387
tri 5839 5289 5937 5387 sw
tri 5937 5289 6035 5387 ne
rect 6035 5289 6389 5387
tri 6389 5289 6487 5387 sw
tri 6487 5289 6585 5387 ne
rect 6585 5289 6939 5387
tri 6939 5289 7037 5387 sw
tri 7037 5289 7135 5387 ne
rect 7135 5289 7489 5387
tri 7489 5289 7587 5387 sw
tri 7587 5289 7685 5387 ne
rect 7685 5289 8039 5387
tri 8039 5289 8137 5387 sw
tri 8137 5289 8235 5387 ne
rect 8235 5289 8589 5387
tri 8589 5289 8687 5387 sw
tri 8687 5289 8785 5387 ne
rect 8785 5289 9139 5387
tri 9139 5289 9237 5387 sw
tri 9237 5289 9335 5387 ne
rect 9335 5289 9689 5387
tri 9689 5289 9787 5387 sw
tri 9787 5289 9885 5387 ne
rect 9885 5289 10239 5387
tri 10239 5289 10337 5387 sw
tri 10337 5289 10435 5387 ne
rect 10435 5289 10789 5387
tri 10789 5289 10887 5387 sw
tri 10887 5289 10985 5387 ne
rect 10985 5289 11339 5387
tri 11339 5289 11437 5387 sw
tri 11437 5289 11535 5387 ne
rect 11535 5289 11889 5387
tri 11889 5289 11987 5387 sw
tri 11987 5289 12085 5387 ne
rect 12085 5289 12439 5387
tri 12439 5289 12537 5387 sw
tri 12537 5289 12635 5387 ne
rect 12635 5289 12989 5387
tri 12989 5289 13087 5387 sw
tri 13087 5289 13185 5387 ne
rect 13185 5289 13539 5387
tri 13539 5289 13637 5387 sw
tri 13637 5289 13735 5387 ne
rect 13735 5289 14089 5387
tri 14089 5289 14187 5387 sw
tri 14187 5289 14285 5387 ne
rect 14285 5289 14639 5387
tri 14639 5289 14737 5387 sw
tri 14737 5289 14835 5387 ne
rect 14835 5289 15189 5387
tri 15189 5289 15287 5387 sw
tri 15287 5289 15385 5387 ne
rect 15385 5289 15739 5387
tri 15739 5289 15837 5387 sw
tri 15837 5289 15935 5387 ne
rect 15935 5289 16289 5387
tri 16289 5289 16387 5387 sw
tri 16387 5289 16485 5387 ne
rect 16485 5289 16839 5387
tri 16839 5289 16937 5387 sw
tri 16937 5289 17035 5387 ne
rect 17035 5289 17389 5387
tri 17389 5289 17487 5387 sw
tri 17487 5289 17585 5387 ne
rect 17585 5289 17939 5387
tri 17939 5289 18037 5387 sw
tri 18037 5289 18135 5387 ne
rect 18135 5289 18489 5387
tri 18489 5289 18587 5387 sw
tri 18587 5289 18685 5387 ne
rect 18685 5289 19039 5387
tri 19039 5289 19137 5387 sw
tri 19137 5289 19235 5387 ne
rect 19235 5289 19589 5387
tri 19589 5289 19687 5387 sw
rect 20800 5289 21800 5937
rect -2000 5285 437 5289
rect -2000 5165 215 5285
rect 335 5191 437 5285
tri 437 5191 535 5289 sw
tri 535 5191 633 5289 ne
rect 633 5285 987 5289
rect 633 5191 765 5285
rect 335 5165 535 5191
rect -2000 5161 535 5165
rect -2000 4513 -1000 5161
tri 113 5063 211 5161 ne
rect 211 5113 535 5161
tri 535 5113 613 5191 sw
tri 633 5113 711 5191 ne
rect 711 5165 765 5191
rect 885 5191 987 5285
tri 987 5191 1085 5289 sw
tri 1085 5191 1183 5289 ne
rect 1183 5285 1537 5289
rect 1183 5191 1315 5285
rect 885 5165 1085 5191
rect 711 5113 1085 5165
tri 1085 5113 1163 5191 sw
tri 1183 5113 1261 5191 ne
rect 1261 5165 1315 5191
rect 1435 5191 1537 5285
tri 1537 5191 1635 5289 sw
tri 1635 5191 1733 5289 ne
rect 1733 5285 2087 5289
rect 1733 5191 1865 5285
rect 1435 5165 1635 5191
rect 1261 5113 1635 5165
tri 1635 5113 1713 5191 sw
tri 1733 5113 1811 5191 ne
rect 1811 5165 1865 5191
rect 1985 5191 2087 5285
tri 2087 5191 2185 5289 sw
tri 2185 5191 2283 5289 ne
rect 2283 5285 2637 5289
rect 2283 5191 2415 5285
rect 1985 5165 2185 5191
rect 1811 5113 2185 5165
tri 2185 5113 2263 5191 sw
tri 2283 5113 2361 5191 ne
rect 2361 5165 2415 5191
rect 2535 5191 2637 5285
tri 2637 5191 2735 5289 sw
tri 2735 5191 2833 5289 ne
rect 2833 5285 3187 5289
rect 2833 5191 2965 5285
rect 2535 5165 2735 5191
rect 2361 5113 2735 5165
tri 2735 5113 2813 5191 sw
tri 2833 5113 2911 5191 ne
rect 2911 5165 2965 5191
rect 3085 5191 3187 5285
tri 3187 5191 3285 5289 sw
tri 3285 5191 3383 5289 ne
rect 3383 5285 3737 5289
rect 3383 5191 3515 5285
rect 3085 5165 3285 5191
rect 2911 5113 3285 5165
tri 3285 5113 3363 5191 sw
tri 3383 5113 3461 5191 ne
rect 3461 5165 3515 5191
rect 3635 5191 3737 5285
tri 3737 5191 3835 5289 sw
tri 3835 5191 3933 5289 ne
rect 3933 5285 4287 5289
rect 3933 5191 4065 5285
rect 3635 5165 3835 5191
rect 3461 5113 3835 5165
tri 3835 5113 3913 5191 sw
tri 3933 5113 4011 5191 ne
rect 4011 5165 4065 5191
rect 4185 5191 4287 5285
tri 4287 5191 4385 5289 sw
tri 4385 5191 4483 5289 ne
rect 4483 5285 4837 5289
rect 4483 5191 4615 5285
rect 4185 5165 4385 5191
rect 4011 5113 4385 5165
tri 4385 5113 4463 5191 sw
tri 4483 5113 4561 5191 ne
rect 4561 5165 4615 5191
rect 4735 5191 4837 5285
tri 4837 5191 4935 5289 sw
tri 4935 5191 5033 5289 ne
rect 5033 5285 5387 5289
rect 5033 5191 5165 5285
rect 4735 5165 4935 5191
rect 4561 5113 4935 5165
tri 4935 5113 5013 5191 sw
tri 5033 5113 5111 5191 ne
rect 5111 5165 5165 5191
rect 5285 5191 5387 5285
tri 5387 5191 5485 5289 sw
tri 5485 5191 5583 5289 ne
rect 5583 5285 5937 5289
rect 5583 5191 5715 5285
rect 5285 5165 5485 5191
rect 5111 5113 5485 5165
tri 5485 5113 5563 5191 sw
tri 5583 5113 5661 5191 ne
rect 5661 5165 5715 5191
rect 5835 5191 5937 5285
tri 5937 5191 6035 5289 sw
tri 6035 5191 6133 5289 ne
rect 6133 5285 6487 5289
rect 6133 5191 6265 5285
rect 5835 5165 6035 5191
rect 5661 5113 6035 5165
tri 6035 5113 6113 5191 sw
tri 6133 5113 6211 5191 ne
rect 6211 5165 6265 5191
rect 6385 5191 6487 5285
tri 6487 5191 6585 5289 sw
tri 6585 5191 6683 5289 ne
rect 6683 5285 7037 5289
rect 6683 5191 6815 5285
rect 6385 5165 6585 5191
rect 6211 5113 6585 5165
tri 6585 5113 6663 5191 sw
tri 6683 5113 6761 5191 ne
rect 6761 5165 6815 5191
rect 6935 5191 7037 5285
tri 7037 5191 7135 5289 sw
tri 7135 5191 7233 5289 ne
rect 7233 5285 7587 5289
rect 7233 5191 7365 5285
rect 6935 5165 7135 5191
rect 6761 5113 7135 5165
tri 7135 5113 7213 5191 sw
tri 7233 5113 7311 5191 ne
rect 7311 5165 7365 5191
rect 7485 5191 7587 5285
tri 7587 5191 7685 5289 sw
tri 7685 5191 7783 5289 ne
rect 7783 5285 8137 5289
rect 7783 5191 7915 5285
rect 7485 5165 7685 5191
rect 7311 5113 7685 5165
tri 7685 5113 7763 5191 sw
tri 7783 5113 7861 5191 ne
rect 7861 5165 7915 5191
rect 8035 5191 8137 5285
tri 8137 5191 8235 5289 sw
tri 8235 5191 8333 5289 ne
rect 8333 5285 8687 5289
rect 8333 5191 8465 5285
rect 8035 5165 8235 5191
rect 7861 5113 8235 5165
tri 8235 5113 8313 5191 sw
tri 8333 5113 8411 5191 ne
rect 8411 5165 8465 5191
rect 8585 5191 8687 5285
tri 8687 5191 8785 5289 sw
tri 8785 5191 8883 5289 ne
rect 8883 5285 9237 5289
rect 8883 5191 9015 5285
rect 8585 5165 8785 5191
rect 8411 5113 8785 5165
tri 8785 5113 8863 5191 sw
tri 8883 5113 8961 5191 ne
rect 8961 5165 9015 5191
rect 9135 5191 9237 5285
tri 9237 5191 9335 5289 sw
tri 9335 5191 9433 5289 ne
rect 9433 5285 9787 5289
rect 9433 5191 9565 5285
rect 9135 5165 9335 5191
rect 8961 5113 9335 5165
tri 9335 5113 9413 5191 sw
tri 9433 5113 9511 5191 ne
rect 9511 5165 9565 5191
rect 9685 5191 9787 5285
tri 9787 5191 9885 5289 sw
tri 9885 5191 9983 5289 ne
rect 9983 5285 10337 5289
rect 9983 5191 10115 5285
rect 9685 5165 9885 5191
rect 9511 5113 9885 5165
tri 9885 5113 9963 5191 sw
tri 9983 5113 10061 5191 ne
rect 10061 5165 10115 5191
rect 10235 5191 10337 5285
tri 10337 5191 10435 5289 sw
tri 10435 5191 10533 5289 ne
rect 10533 5285 10887 5289
rect 10533 5191 10665 5285
rect 10235 5165 10435 5191
rect 10061 5113 10435 5165
tri 10435 5113 10513 5191 sw
tri 10533 5113 10611 5191 ne
rect 10611 5165 10665 5191
rect 10785 5191 10887 5285
tri 10887 5191 10985 5289 sw
tri 10985 5191 11083 5289 ne
rect 11083 5285 11437 5289
rect 11083 5191 11215 5285
rect 10785 5165 10985 5191
rect 10611 5113 10985 5165
tri 10985 5113 11063 5191 sw
tri 11083 5113 11161 5191 ne
rect 11161 5165 11215 5191
rect 11335 5191 11437 5285
tri 11437 5191 11535 5289 sw
tri 11535 5191 11633 5289 ne
rect 11633 5285 11987 5289
rect 11633 5191 11765 5285
rect 11335 5165 11535 5191
rect 11161 5113 11535 5165
tri 11535 5113 11613 5191 sw
tri 11633 5113 11711 5191 ne
rect 11711 5165 11765 5191
rect 11885 5191 11987 5285
tri 11987 5191 12085 5289 sw
tri 12085 5191 12183 5289 ne
rect 12183 5285 12537 5289
rect 12183 5191 12315 5285
rect 11885 5165 12085 5191
rect 11711 5113 12085 5165
tri 12085 5113 12163 5191 sw
tri 12183 5113 12261 5191 ne
rect 12261 5165 12315 5191
rect 12435 5191 12537 5285
tri 12537 5191 12635 5289 sw
tri 12635 5191 12733 5289 ne
rect 12733 5285 13087 5289
rect 12733 5191 12865 5285
rect 12435 5165 12635 5191
rect 12261 5113 12635 5165
tri 12635 5113 12713 5191 sw
tri 12733 5113 12811 5191 ne
rect 12811 5165 12865 5191
rect 12985 5191 13087 5285
tri 13087 5191 13185 5289 sw
tri 13185 5191 13283 5289 ne
rect 13283 5285 13637 5289
rect 13283 5191 13415 5285
rect 12985 5165 13185 5191
rect 12811 5113 13185 5165
tri 13185 5113 13263 5191 sw
tri 13283 5113 13361 5191 ne
rect 13361 5165 13415 5191
rect 13535 5191 13637 5285
tri 13637 5191 13735 5289 sw
tri 13735 5191 13833 5289 ne
rect 13833 5285 14187 5289
rect 13833 5191 13965 5285
rect 13535 5165 13735 5191
rect 13361 5113 13735 5165
tri 13735 5113 13813 5191 sw
tri 13833 5113 13911 5191 ne
rect 13911 5165 13965 5191
rect 14085 5191 14187 5285
tri 14187 5191 14285 5289 sw
tri 14285 5191 14383 5289 ne
rect 14383 5285 14737 5289
rect 14383 5191 14515 5285
rect 14085 5165 14285 5191
rect 13911 5113 14285 5165
tri 14285 5113 14363 5191 sw
tri 14383 5113 14461 5191 ne
rect 14461 5165 14515 5191
rect 14635 5191 14737 5285
tri 14737 5191 14835 5289 sw
tri 14835 5191 14933 5289 ne
rect 14933 5285 15287 5289
rect 14933 5191 15065 5285
rect 14635 5165 14835 5191
rect 14461 5113 14835 5165
tri 14835 5113 14913 5191 sw
tri 14933 5113 15011 5191 ne
rect 15011 5165 15065 5191
rect 15185 5191 15287 5285
tri 15287 5191 15385 5289 sw
tri 15385 5191 15483 5289 ne
rect 15483 5285 15837 5289
rect 15483 5191 15615 5285
rect 15185 5165 15385 5191
rect 15011 5113 15385 5165
tri 15385 5113 15463 5191 sw
tri 15483 5113 15561 5191 ne
rect 15561 5165 15615 5191
rect 15735 5191 15837 5285
tri 15837 5191 15935 5289 sw
tri 15935 5191 16033 5289 ne
rect 16033 5285 16387 5289
rect 16033 5191 16165 5285
rect 15735 5165 15935 5191
rect 15561 5113 15935 5165
tri 15935 5113 16013 5191 sw
tri 16033 5113 16111 5191 ne
rect 16111 5165 16165 5191
rect 16285 5191 16387 5285
tri 16387 5191 16485 5289 sw
tri 16485 5191 16583 5289 ne
rect 16583 5285 16937 5289
rect 16583 5191 16715 5285
rect 16285 5165 16485 5191
rect 16111 5113 16485 5165
tri 16485 5113 16563 5191 sw
tri 16583 5113 16661 5191 ne
rect 16661 5165 16715 5191
rect 16835 5191 16937 5285
tri 16937 5191 17035 5289 sw
tri 17035 5191 17133 5289 ne
rect 17133 5285 17487 5289
rect 17133 5191 17265 5285
rect 16835 5165 17035 5191
rect 16661 5113 17035 5165
tri 17035 5113 17113 5191 sw
tri 17133 5113 17211 5191 ne
rect 17211 5165 17265 5191
rect 17385 5191 17487 5285
tri 17487 5191 17585 5289 sw
tri 17585 5191 17683 5289 ne
rect 17683 5285 18037 5289
rect 17683 5191 17815 5285
rect 17385 5165 17585 5191
rect 17211 5113 17585 5165
tri 17585 5113 17663 5191 sw
tri 17683 5113 17761 5191 ne
rect 17761 5165 17815 5191
rect 17935 5191 18037 5285
tri 18037 5191 18135 5289 sw
tri 18135 5191 18233 5289 ne
rect 18233 5285 18587 5289
rect 18233 5191 18365 5285
rect 17935 5165 18135 5191
rect 17761 5113 18135 5165
tri 18135 5113 18213 5191 sw
tri 18233 5113 18311 5191 ne
rect 18311 5165 18365 5191
rect 18485 5191 18587 5285
tri 18587 5191 18685 5289 sw
tri 18685 5191 18783 5289 ne
rect 18783 5285 19137 5289
rect 18783 5191 18915 5285
rect 18485 5165 18685 5191
rect 18311 5113 18685 5165
tri 18685 5113 18763 5191 sw
tri 18783 5113 18861 5191 ne
rect 18861 5165 18915 5191
rect 19035 5191 19137 5285
tri 19137 5191 19235 5289 sw
tri 19235 5191 19333 5289 ne
rect 19333 5285 21800 5289
rect 19333 5191 19465 5285
rect 19035 5165 19235 5191
rect 18861 5113 19235 5165
tri 19235 5113 19313 5191 sw
tri 19333 5113 19411 5191 ne
rect 19411 5165 19465 5191
rect 19585 5165 21800 5285
rect 19411 5113 21800 5165
rect 211 5063 613 5113
rect -500 5013 113 5063
tri 113 5013 163 5063 sw
tri 211 5013 261 5063 ne
rect 261 5033 613 5063
tri 613 5033 693 5113 sw
tri 711 5033 791 5113 ne
rect 791 5033 1163 5113
tri 1163 5033 1243 5113 sw
tri 1261 5033 1341 5113 ne
rect 1341 5033 1713 5113
tri 1713 5033 1793 5113 sw
tri 1811 5033 1891 5113 ne
rect 1891 5033 2263 5113
tri 2263 5033 2343 5113 sw
tri 2361 5033 2441 5113 ne
rect 2441 5033 2813 5113
tri 2813 5033 2893 5113 sw
tri 2911 5033 2991 5113 ne
rect 2991 5033 3363 5113
tri 3363 5033 3443 5113 sw
tri 3461 5033 3541 5113 ne
rect 3541 5033 3913 5113
tri 3913 5033 3993 5113 sw
tri 4011 5033 4091 5113 ne
rect 4091 5033 4463 5113
tri 4463 5033 4543 5113 sw
tri 4561 5033 4641 5113 ne
rect 4641 5033 5013 5113
tri 5013 5033 5093 5113 sw
tri 5111 5033 5191 5113 ne
rect 5191 5033 5563 5113
tri 5563 5033 5643 5113 sw
tri 5661 5033 5741 5113 ne
rect 5741 5033 6113 5113
tri 6113 5033 6193 5113 sw
tri 6211 5033 6291 5113 ne
rect 6291 5033 6663 5113
tri 6663 5033 6743 5113 sw
tri 6761 5033 6841 5113 ne
rect 6841 5033 7213 5113
tri 7213 5033 7293 5113 sw
tri 7311 5033 7391 5113 ne
rect 7391 5033 7763 5113
tri 7763 5033 7843 5113 sw
tri 7861 5033 7941 5113 ne
rect 7941 5033 8313 5113
tri 8313 5033 8393 5113 sw
tri 8411 5033 8491 5113 ne
rect 8491 5033 8863 5113
tri 8863 5033 8943 5113 sw
tri 8961 5033 9041 5113 ne
rect 9041 5033 9413 5113
tri 9413 5033 9493 5113 sw
tri 9511 5033 9591 5113 ne
rect 9591 5033 9963 5113
tri 9963 5033 10043 5113 sw
tri 10061 5033 10141 5113 ne
rect 10141 5033 10513 5113
tri 10513 5033 10593 5113 sw
tri 10611 5033 10691 5113 ne
rect 10691 5033 11063 5113
tri 11063 5033 11143 5113 sw
tri 11161 5033 11241 5113 ne
rect 11241 5033 11613 5113
tri 11613 5033 11693 5113 sw
tri 11711 5033 11791 5113 ne
rect 11791 5033 12163 5113
tri 12163 5033 12243 5113 sw
tri 12261 5033 12341 5113 ne
rect 12341 5033 12713 5113
tri 12713 5033 12793 5113 sw
tri 12811 5033 12891 5113 ne
rect 12891 5033 13263 5113
tri 13263 5033 13343 5113 sw
tri 13361 5033 13441 5113 ne
rect 13441 5033 13813 5113
tri 13813 5033 13893 5113 sw
tri 13911 5033 13991 5113 ne
rect 13991 5033 14363 5113
tri 14363 5033 14443 5113 sw
tri 14461 5033 14541 5113 ne
rect 14541 5033 14913 5113
tri 14913 5033 14993 5113 sw
tri 15011 5033 15091 5113 ne
rect 15091 5033 15463 5113
tri 15463 5033 15543 5113 sw
tri 15561 5033 15641 5113 ne
rect 15641 5033 16013 5113
tri 16013 5033 16093 5113 sw
tri 16111 5033 16191 5113 ne
rect 16191 5033 16563 5113
tri 16563 5033 16643 5113 sw
tri 16661 5033 16741 5113 ne
rect 16741 5033 17113 5113
tri 17113 5033 17193 5113 sw
tri 17211 5033 17291 5113 ne
rect 17291 5033 17663 5113
tri 17663 5033 17743 5113 sw
tri 17761 5033 17841 5113 ne
rect 17841 5033 18213 5113
tri 18213 5033 18293 5113 sw
tri 18311 5033 18391 5113 ne
rect 18391 5033 18763 5113
tri 18763 5033 18843 5113 sw
tri 18861 5033 18941 5113 ne
rect 18941 5033 19313 5113
tri 19313 5033 19393 5113 sw
tri 19411 5033 19491 5113 ne
rect 19491 5033 20100 5113
rect 261 5013 693 5033
rect -500 4935 163 5013
tri 163 4935 241 5013 sw
tri 261 4935 339 5013 ne
rect 339 4935 693 5013
tri 693 4935 791 5033 sw
tri 791 4935 889 5033 ne
rect 889 4935 1243 5033
tri 1243 4935 1341 5033 sw
tri 1341 4935 1439 5033 ne
rect 1439 4935 1793 5033
tri 1793 4935 1891 5033 sw
tri 1891 4935 1989 5033 ne
rect 1989 4935 2343 5033
tri 2343 4935 2441 5033 sw
tri 2441 4935 2539 5033 ne
rect 2539 4935 2893 5033
tri 2893 4935 2991 5033 sw
tri 2991 4935 3089 5033 ne
rect 3089 4935 3443 5033
tri 3443 4935 3541 5033 sw
tri 3541 4935 3639 5033 ne
rect 3639 4935 3993 5033
tri 3993 4935 4091 5033 sw
tri 4091 4935 4189 5033 ne
rect 4189 4935 4543 5033
tri 4543 4935 4641 5033 sw
tri 4641 4935 4739 5033 ne
rect 4739 4935 5093 5033
tri 5093 4935 5191 5033 sw
tri 5191 4935 5289 5033 ne
rect 5289 4935 5643 5033
tri 5643 4935 5741 5033 sw
tri 5741 4935 5839 5033 ne
rect 5839 4935 6193 5033
tri 6193 4935 6291 5033 sw
tri 6291 4935 6389 5033 ne
rect 6389 4935 6743 5033
tri 6743 4935 6841 5033 sw
tri 6841 4935 6939 5033 ne
rect 6939 4935 7293 5033
tri 7293 4935 7391 5033 sw
tri 7391 4935 7489 5033 ne
rect 7489 4935 7843 5033
tri 7843 4935 7941 5033 sw
tri 7941 4935 8039 5033 ne
rect 8039 4935 8393 5033
tri 8393 4935 8491 5033 sw
tri 8491 4935 8589 5033 ne
rect 8589 4935 8943 5033
tri 8943 4935 9041 5033 sw
tri 9041 4935 9139 5033 ne
rect 9139 4935 9493 5033
tri 9493 4935 9591 5033 sw
tri 9591 4935 9689 5033 ne
rect 9689 4935 10043 5033
tri 10043 4935 10141 5033 sw
tri 10141 4935 10239 5033 ne
rect 10239 4935 10593 5033
tri 10593 4935 10691 5033 sw
tri 10691 4935 10789 5033 ne
rect 10789 4935 11143 5033
tri 11143 4935 11241 5033 sw
tri 11241 4935 11339 5033 ne
rect 11339 4935 11693 5033
tri 11693 4935 11791 5033 sw
tri 11791 4935 11889 5033 ne
rect 11889 4935 12243 5033
tri 12243 4935 12341 5033 sw
tri 12341 4935 12439 5033 ne
rect 12439 4935 12793 5033
tri 12793 4935 12891 5033 sw
tri 12891 4935 12989 5033 ne
rect 12989 4935 13343 5033
tri 13343 4935 13441 5033 sw
tri 13441 4935 13539 5033 ne
rect 13539 4935 13893 5033
tri 13893 4935 13991 5033 sw
tri 13991 4935 14089 5033 ne
rect 14089 4935 14443 5033
tri 14443 4935 14541 5033 sw
tri 14541 4935 14639 5033 ne
rect 14639 4935 14993 5033
tri 14993 4935 15091 5033 sw
tri 15091 4935 15189 5033 ne
rect 15189 4935 15543 5033
tri 15543 4935 15641 5033 sw
tri 15641 4935 15739 5033 ne
rect 15739 4935 16093 5033
tri 16093 4935 16191 5033 sw
tri 16191 4935 16289 5033 ne
rect 16289 4935 16643 5033
tri 16643 4935 16741 5033 sw
tri 16741 4935 16839 5033 ne
rect 16839 4935 17193 5033
tri 17193 4935 17291 5033 sw
tri 17291 4935 17389 5033 ne
rect 17389 4935 17743 5033
tri 17743 4935 17841 5033 sw
tri 17841 4935 17939 5033 ne
rect 17939 4935 18293 5033
tri 18293 4935 18391 5033 sw
tri 18391 4935 18489 5033 ne
rect 18489 4935 18843 5033
tri 18843 4935 18941 5033 sw
tri 18941 4935 19039 5033 ne
rect 19039 4935 19393 5033
tri 19393 4935 19491 5033 sw
tri 19491 4935 19589 5033 ne
rect 19589 5013 20100 5033
rect 20200 5013 21800 5113
rect 19589 4935 21800 5013
rect -500 4887 241 4935
rect -500 4787 -400 4887
rect -300 4837 241 4887
tri 241 4837 339 4935 sw
tri 339 4837 437 4935 ne
rect 437 4837 791 4935
tri 791 4837 889 4935 sw
tri 889 4837 987 4935 ne
rect 987 4837 1341 4935
tri 1341 4837 1439 4935 sw
tri 1439 4837 1537 4935 ne
rect 1537 4837 1891 4935
tri 1891 4837 1989 4935 sw
tri 1989 4837 2087 4935 ne
rect 2087 4837 2441 4935
tri 2441 4837 2539 4935 sw
tri 2539 4837 2637 4935 ne
rect 2637 4837 2991 4935
tri 2991 4837 3089 4935 sw
tri 3089 4837 3187 4935 ne
rect 3187 4837 3541 4935
tri 3541 4837 3639 4935 sw
tri 3639 4837 3737 4935 ne
rect 3737 4837 4091 4935
tri 4091 4837 4189 4935 sw
tri 4189 4837 4287 4935 ne
rect 4287 4837 4641 4935
tri 4641 4837 4739 4935 sw
tri 4739 4837 4837 4935 ne
rect 4837 4837 5191 4935
tri 5191 4837 5289 4935 sw
tri 5289 4837 5387 4935 ne
rect 5387 4837 5741 4935
tri 5741 4837 5839 4935 sw
tri 5839 4837 5937 4935 ne
rect 5937 4837 6291 4935
tri 6291 4837 6389 4935 sw
tri 6389 4837 6487 4935 ne
rect 6487 4837 6841 4935
tri 6841 4837 6939 4935 sw
tri 6939 4837 7037 4935 ne
rect 7037 4837 7391 4935
tri 7391 4837 7489 4935 sw
tri 7489 4837 7587 4935 ne
rect 7587 4837 7941 4935
tri 7941 4837 8039 4935 sw
tri 8039 4837 8137 4935 ne
rect 8137 4837 8491 4935
tri 8491 4837 8589 4935 sw
tri 8589 4837 8687 4935 ne
rect 8687 4837 9041 4935
tri 9041 4837 9139 4935 sw
tri 9139 4837 9237 4935 ne
rect 9237 4837 9591 4935
tri 9591 4837 9689 4935 sw
tri 9689 4837 9787 4935 ne
rect 9787 4837 10141 4935
tri 10141 4837 10239 4935 sw
tri 10239 4837 10337 4935 ne
rect 10337 4837 10691 4935
tri 10691 4837 10789 4935 sw
tri 10789 4837 10887 4935 ne
rect 10887 4837 11241 4935
tri 11241 4837 11339 4935 sw
tri 11339 4837 11437 4935 ne
rect 11437 4837 11791 4935
tri 11791 4837 11889 4935 sw
tri 11889 4837 11987 4935 ne
rect 11987 4837 12341 4935
tri 12341 4837 12439 4935 sw
tri 12439 4837 12537 4935 ne
rect 12537 4837 12891 4935
tri 12891 4837 12989 4935 sw
tri 12989 4837 13087 4935 ne
rect 13087 4837 13441 4935
tri 13441 4837 13539 4935 sw
tri 13539 4837 13637 4935 ne
rect 13637 4837 13991 4935
tri 13991 4837 14089 4935 sw
tri 14089 4837 14187 4935 ne
rect 14187 4837 14541 4935
tri 14541 4837 14639 4935 sw
tri 14639 4837 14737 4935 ne
rect 14737 4837 15091 4935
tri 15091 4837 15189 4935 sw
tri 15189 4837 15287 4935 ne
rect 15287 4837 15641 4935
tri 15641 4837 15739 4935 sw
tri 15739 4837 15837 4935 ne
rect 15837 4837 16191 4935
tri 16191 4837 16289 4935 sw
tri 16289 4837 16387 4935 ne
rect 16387 4837 16741 4935
tri 16741 4837 16839 4935 sw
tri 16839 4837 16937 4935 ne
rect 16937 4837 17291 4935
tri 17291 4837 17389 4935 sw
tri 17389 4837 17487 4935 ne
rect 17487 4837 17841 4935
tri 17841 4837 17939 4935 sw
tri 17939 4837 18037 4935 ne
rect 18037 4837 18391 4935
tri 18391 4837 18489 4935 sw
tri 18489 4837 18587 4935 ne
rect 18587 4837 18941 4935
tri 18941 4837 19039 4935 sw
tri 19039 4837 19137 4935 ne
rect 19137 4837 19491 4935
tri 19491 4837 19589 4935 sw
tri 19589 4837 19687 4935 ne
rect 19687 4837 21800 4935
rect -300 4787 339 4837
rect -500 4739 339 4787
tri 339 4739 437 4837 sw
tri 437 4739 535 4837 ne
rect 535 4739 889 4837
tri 889 4739 987 4837 sw
tri 987 4739 1085 4837 ne
rect 1085 4739 1439 4837
tri 1439 4739 1537 4837 sw
tri 1537 4739 1635 4837 ne
rect 1635 4739 1989 4837
tri 1989 4739 2087 4837 sw
tri 2087 4739 2185 4837 ne
rect 2185 4739 2539 4837
tri 2539 4739 2637 4837 sw
tri 2637 4739 2735 4837 ne
rect 2735 4739 3089 4837
tri 3089 4739 3187 4837 sw
tri 3187 4739 3285 4837 ne
rect 3285 4739 3639 4837
tri 3639 4739 3737 4837 sw
tri 3737 4739 3835 4837 ne
rect 3835 4739 4189 4837
tri 4189 4739 4287 4837 sw
tri 4287 4739 4385 4837 ne
rect 4385 4739 4739 4837
tri 4739 4739 4837 4837 sw
tri 4837 4739 4935 4837 ne
rect 4935 4739 5289 4837
tri 5289 4739 5387 4837 sw
tri 5387 4739 5485 4837 ne
rect 5485 4739 5839 4837
tri 5839 4739 5937 4837 sw
tri 5937 4739 6035 4837 ne
rect 6035 4739 6389 4837
tri 6389 4739 6487 4837 sw
tri 6487 4739 6585 4837 ne
rect 6585 4739 6939 4837
tri 6939 4739 7037 4837 sw
tri 7037 4739 7135 4837 ne
rect 7135 4739 7489 4837
tri 7489 4739 7587 4837 sw
tri 7587 4739 7685 4837 ne
rect 7685 4739 8039 4837
tri 8039 4739 8137 4837 sw
tri 8137 4739 8235 4837 ne
rect 8235 4739 8589 4837
tri 8589 4739 8687 4837 sw
tri 8687 4739 8785 4837 ne
rect 8785 4739 9139 4837
tri 9139 4739 9237 4837 sw
tri 9237 4739 9335 4837 ne
rect 9335 4739 9689 4837
tri 9689 4739 9787 4837 sw
tri 9787 4739 9885 4837 ne
rect 9885 4739 10239 4837
tri 10239 4739 10337 4837 sw
tri 10337 4739 10435 4837 ne
rect 10435 4739 10789 4837
tri 10789 4739 10887 4837 sw
tri 10887 4739 10985 4837 ne
rect 10985 4739 11339 4837
tri 11339 4739 11437 4837 sw
tri 11437 4739 11535 4837 ne
rect 11535 4739 11889 4837
tri 11889 4739 11987 4837 sw
tri 11987 4739 12085 4837 ne
rect 12085 4739 12439 4837
tri 12439 4739 12537 4837 sw
tri 12537 4739 12635 4837 ne
rect 12635 4739 12989 4837
tri 12989 4739 13087 4837 sw
tri 13087 4739 13185 4837 ne
rect 13185 4739 13539 4837
tri 13539 4739 13637 4837 sw
tri 13637 4739 13735 4837 ne
rect 13735 4739 14089 4837
tri 14089 4739 14187 4837 sw
tri 14187 4739 14285 4837 ne
rect 14285 4739 14639 4837
tri 14639 4739 14737 4837 sw
tri 14737 4739 14835 4837 ne
rect 14835 4739 15189 4837
tri 15189 4739 15287 4837 sw
tri 15287 4739 15385 4837 ne
rect 15385 4739 15739 4837
tri 15739 4739 15837 4837 sw
tri 15837 4739 15935 4837 ne
rect 15935 4739 16289 4837
tri 16289 4739 16387 4837 sw
tri 16387 4739 16485 4837 ne
rect 16485 4739 16839 4837
tri 16839 4739 16937 4837 sw
tri 16937 4739 17035 4837 ne
rect 17035 4739 17389 4837
tri 17389 4739 17487 4837 sw
tri 17487 4739 17585 4837 ne
rect 17585 4739 17939 4837
tri 17939 4739 18037 4837 sw
tri 18037 4739 18135 4837 ne
rect 18135 4739 18489 4837
tri 18489 4739 18587 4837 sw
tri 18587 4739 18685 4837 ne
rect 18685 4739 19039 4837
tri 19039 4739 19137 4837 sw
tri 19137 4739 19235 4837 ne
rect 19235 4739 19589 4837
tri 19589 4739 19687 4837 sw
rect -500 4735 437 4739
rect -500 4615 215 4735
rect 335 4641 437 4735
tri 437 4641 535 4739 sw
tri 535 4641 633 4739 ne
rect 633 4735 987 4739
rect 633 4641 765 4735
rect 335 4615 535 4641
rect -500 4611 535 4615
tri 535 4611 565 4641 sw
tri 633 4611 663 4641 ne
rect 663 4615 765 4641
rect 885 4641 987 4735
tri 987 4641 1085 4739 sw
tri 1085 4641 1183 4739 ne
rect 1183 4735 1537 4739
rect 1183 4641 1315 4735
rect 885 4615 1085 4641
rect 663 4611 1085 4615
tri 1085 4611 1115 4641 sw
tri 1183 4611 1213 4641 ne
rect 1213 4615 1315 4641
rect 1435 4641 1537 4735
tri 1537 4641 1635 4739 sw
tri 1635 4641 1733 4739 ne
rect 1733 4735 2087 4739
rect 1733 4641 1865 4735
rect 1435 4615 1635 4641
rect 1213 4611 1635 4615
tri 1635 4611 1665 4641 sw
tri 1733 4611 1763 4641 ne
rect 1763 4615 1865 4641
rect 1985 4641 2087 4735
tri 2087 4641 2185 4739 sw
tri 2185 4641 2283 4739 ne
rect 2283 4735 2637 4739
rect 2283 4641 2415 4735
rect 1985 4615 2185 4641
rect 1763 4611 2185 4615
tri 2185 4611 2215 4641 sw
tri 2283 4611 2313 4641 ne
rect 2313 4615 2415 4641
rect 2535 4641 2637 4735
tri 2637 4641 2735 4739 sw
tri 2735 4641 2833 4739 ne
rect 2833 4735 3187 4739
rect 2833 4641 2965 4735
rect 2535 4615 2735 4641
rect 2313 4611 2735 4615
tri 2735 4611 2765 4641 sw
tri 2833 4611 2863 4641 ne
rect 2863 4615 2965 4641
rect 3085 4641 3187 4735
tri 3187 4641 3285 4739 sw
tri 3285 4641 3383 4739 ne
rect 3383 4735 3737 4739
rect 3383 4641 3515 4735
rect 3085 4615 3285 4641
rect 2863 4611 3285 4615
tri 3285 4611 3315 4641 sw
tri 3383 4611 3413 4641 ne
rect 3413 4615 3515 4641
rect 3635 4641 3737 4735
tri 3737 4641 3835 4739 sw
tri 3835 4641 3933 4739 ne
rect 3933 4735 4287 4739
rect 3933 4641 4065 4735
rect 3635 4615 3835 4641
rect 3413 4611 3835 4615
tri 3835 4611 3865 4641 sw
tri 3933 4611 3963 4641 ne
rect 3963 4615 4065 4641
rect 4185 4641 4287 4735
tri 4287 4641 4385 4739 sw
tri 4385 4641 4483 4739 ne
rect 4483 4735 4837 4739
rect 4483 4641 4615 4735
rect 4185 4615 4385 4641
rect 3963 4611 4385 4615
tri 4385 4611 4415 4641 sw
tri 4483 4611 4513 4641 ne
rect 4513 4615 4615 4641
rect 4735 4641 4837 4735
tri 4837 4641 4935 4739 sw
tri 4935 4641 5033 4739 ne
rect 5033 4735 5387 4739
rect 5033 4641 5165 4735
rect 4735 4615 4935 4641
rect 4513 4611 4935 4615
tri 4935 4611 4965 4641 sw
tri 5033 4611 5063 4641 ne
rect 5063 4615 5165 4641
rect 5285 4641 5387 4735
tri 5387 4641 5485 4739 sw
tri 5485 4641 5583 4739 ne
rect 5583 4735 5937 4739
rect 5583 4641 5715 4735
rect 5285 4615 5485 4641
rect 5063 4611 5485 4615
tri 5485 4611 5515 4641 sw
tri 5583 4611 5613 4641 ne
rect 5613 4615 5715 4641
rect 5835 4641 5937 4735
tri 5937 4641 6035 4739 sw
tri 6035 4641 6133 4739 ne
rect 6133 4735 6487 4739
rect 6133 4641 6265 4735
rect 5835 4615 6035 4641
rect 5613 4611 6035 4615
tri 6035 4611 6065 4641 sw
tri 6133 4611 6163 4641 ne
rect 6163 4615 6265 4641
rect 6385 4641 6487 4735
tri 6487 4641 6585 4739 sw
tri 6585 4641 6683 4739 ne
rect 6683 4735 7037 4739
rect 6683 4641 6815 4735
rect 6385 4615 6585 4641
rect 6163 4611 6585 4615
tri 6585 4611 6615 4641 sw
tri 6683 4611 6713 4641 ne
rect 6713 4615 6815 4641
rect 6935 4641 7037 4735
tri 7037 4641 7135 4739 sw
tri 7135 4641 7233 4739 ne
rect 7233 4735 7587 4739
rect 7233 4641 7365 4735
rect 6935 4615 7135 4641
rect 6713 4611 7135 4615
tri 7135 4611 7165 4641 sw
tri 7233 4611 7263 4641 ne
rect 7263 4615 7365 4641
rect 7485 4641 7587 4735
tri 7587 4641 7685 4739 sw
tri 7685 4641 7783 4739 ne
rect 7783 4735 8137 4739
rect 7783 4641 7915 4735
rect 7485 4615 7685 4641
rect 7263 4611 7685 4615
tri 7685 4611 7715 4641 sw
tri 7783 4611 7813 4641 ne
rect 7813 4615 7915 4641
rect 8035 4641 8137 4735
tri 8137 4641 8235 4739 sw
tri 8235 4641 8333 4739 ne
rect 8333 4735 8687 4739
rect 8333 4641 8465 4735
rect 8035 4615 8235 4641
rect 7813 4611 8235 4615
tri 8235 4611 8265 4641 sw
tri 8333 4611 8363 4641 ne
rect 8363 4615 8465 4641
rect 8585 4641 8687 4735
tri 8687 4641 8785 4739 sw
tri 8785 4641 8883 4739 ne
rect 8883 4735 9237 4739
rect 8883 4641 9015 4735
rect 8585 4615 8785 4641
rect 8363 4611 8785 4615
tri 8785 4611 8815 4641 sw
tri 8883 4611 8913 4641 ne
rect 8913 4615 9015 4641
rect 9135 4641 9237 4735
tri 9237 4641 9335 4739 sw
tri 9335 4641 9433 4739 ne
rect 9433 4735 9787 4739
rect 9433 4641 9565 4735
rect 9135 4615 9335 4641
rect 8913 4611 9335 4615
tri 9335 4611 9365 4641 sw
tri 9433 4611 9463 4641 ne
rect 9463 4615 9565 4641
rect 9685 4641 9787 4735
tri 9787 4641 9885 4739 sw
tri 9885 4641 9983 4739 ne
rect 9983 4735 10337 4739
rect 9983 4641 10115 4735
rect 9685 4615 9885 4641
rect 9463 4611 9885 4615
tri 9885 4611 9915 4641 sw
tri 9983 4611 10013 4641 ne
rect 10013 4615 10115 4641
rect 10235 4641 10337 4735
tri 10337 4641 10435 4739 sw
tri 10435 4641 10533 4739 ne
rect 10533 4735 10887 4739
rect 10533 4641 10665 4735
rect 10235 4615 10435 4641
rect 10013 4611 10435 4615
tri 10435 4611 10465 4641 sw
tri 10533 4611 10563 4641 ne
rect 10563 4615 10665 4641
rect 10785 4641 10887 4735
tri 10887 4641 10985 4739 sw
tri 10985 4641 11083 4739 ne
rect 11083 4735 11437 4739
rect 11083 4641 11215 4735
rect 10785 4615 10985 4641
rect 10563 4611 10985 4615
tri 10985 4611 11015 4641 sw
tri 11083 4611 11113 4641 ne
rect 11113 4615 11215 4641
rect 11335 4641 11437 4735
tri 11437 4641 11535 4739 sw
tri 11535 4641 11633 4739 ne
rect 11633 4735 11987 4739
rect 11633 4641 11765 4735
rect 11335 4615 11535 4641
rect 11113 4611 11535 4615
tri 11535 4611 11565 4641 sw
tri 11633 4611 11663 4641 ne
rect 11663 4615 11765 4641
rect 11885 4641 11987 4735
tri 11987 4641 12085 4739 sw
tri 12085 4641 12183 4739 ne
rect 12183 4735 12537 4739
rect 12183 4641 12315 4735
rect 11885 4615 12085 4641
rect 11663 4611 12085 4615
tri 12085 4611 12115 4641 sw
tri 12183 4611 12213 4641 ne
rect 12213 4615 12315 4641
rect 12435 4641 12537 4735
tri 12537 4641 12635 4739 sw
tri 12635 4641 12733 4739 ne
rect 12733 4735 13087 4739
rect 12733 4641 12865 4735
rect 12435 4615 12635 4641
rect 12213 4611 12635 4615
tri 12635 4611 12665 4641 sw
tri 12733 4611 12763 4641 ne
rect 12763 4615 12865 4641
rect 12985 4641 13087 4735
tri 13087 4641 13185 4739 sw
tri 13185 4641 13283 4739 ne
rect 13283 4735 13637 4739
rect 13283 4641 13415 4735
rect 12985 4615 13185 4641
rect 12763 4611 13185 4615
tri 13185 4611 13215 4641 sw
tri 13283 4611 13313 4641 ne
rect 13313 4615 13415 4641
rect 13535 4641 13637 4735
tri 13637 4641 13735 4739 sw
tri 13735 4641 13833 4739 ne
rect 13833 4735 14187 4739
rect 13833 4641 13965 4735
rect 13535 4615 13735 4641
rect 13313 4611 13735 4615
tri 13735 4611 13765 4641 sw
tri 13833 4611 13863 4641 ne
rect 13863 4615 13965 4641
rect 14085 4641 14187 4735
tri 14187 4641 14285 4739 sw
tri 14285 4641 14383 4739 ne
rect 14383 4735 14737 4739
rect 14383 4641 14515 4735
rect 14085 4615 14285 4641
rect 13863 4611 14285 4615
tri 14285 4611 14315 4641 sw
tri 14383 4611 14413 4641 ne
rect 14413 4615 14515 4641
rect 14635 4641 14737 4735
tri 14737 4641 14835 4739 sw
tri 14835 4641 14933 4739 ne
rect 14933 4735 15287 4739
rect 14933 4641 15065 4735
rect 14635 4615 14835 4641
rect 14413 4611 14835 4615
tri 14835 4611 14865 4641 sw
tri 14933 4611 14963 4641 ne
rect 14963 4615 15065 4641
rect 15185 4641 15287 4735
tri 15287 4641 15385 4739 sw
tri 15385 4641 15483 4739 ne
rect 15483 4735 15837 4739
rect 15483 4641 15615 4735
rect 15185 4615 15385 4641
rect 14963 4611 15385 4615
tri 15385 4611 15415 4641 sw
tri 15483 4611 15513 4641 ne
rect 15513 4615 15615 4641
rect 15735 4641 15837 4735
tri 15837 4641 15935 4739 sw
tri 15935 4641 16033 4739 ne
rect 16033 4735 16387 4739
rect 16033 4641 16165 4735
rect 15735 4615 15935 4641
rect 15513 4611 15935 4615
tri 15935 4611 15965 4641 sw
tri 16033 4611 16063 4641 ne
rect 16063 4615 16165 4641
rect 16285 4641 16387 4735
tri 16387 4641 16485 4739 sw
tri 16485 4641 16583 4739 ne
rect 16583 4735 16937 4739
rect 16583 4641 16715 4735
rect 16285 4615 16485 4641
rect 16063 4611 16485 4615
tri 16485 4611 16515 4641 sw
tri 16583 4611 16613 4641 ne
rect 16613 4615 16715 4641
rect 16835 4641 16937 4735
tri 16937 4641 17035 4739 sw
tri 17035 4641 17133 4739 ne
rect 17133 4735 17487 4739
rect 17133 4641 17265 4735
rect 16835 4615 17035 4641
rect 16613 4611 17035 4615
tri 17035 4611 17065 4641 sw
tri 17133 4611 17163 4641 ne
rect 17163 4615 17265 4641
rect 17385 4641 17487 4735
tri 17487 4641 17585 4739 sw
tri 17585 4641 17683 4739 ne
rect 17683 4735 18037 4739
rect 17683 4641 17815 4735
rect 17385 4615 17585 4641
rect 17163 4611 17585 4615
tri 17585 4611 17615 4641 sw
tri 17683 4611 17713 4641 ne
rect 17713 4615 17815 4641
rect 17935 4641 18037 4735
tri 18037 4641 18135 4739 sw
tri 18135 4641 18233 4739 ne
rect 18233 4735 18587 4739
rect 18233 4641 18365 4735
rect 17935 4615 18135 4641
rect 17713 4611 18135 4615
tri 18135 4611 18165 4641 sw
tri 18233 4611 18263 4641 ne
rect 18263 4615 18365 4641
rect 18485 4641 18587 4735
tri 18587 4641 18685 4739 sw
tri 18685 4641 18783 4739 ne
rect 18783 4735 19137 4739
rect 18783 4641 18915 4735
rect 18485 4615 18685 4641
rect 18263 4611 18685 4615
tri 18685 4611 18715 4641 sw
tri 18783 4611 18813 4641 ne
rect 18813 4615 18915 4641
rect 19035 4641 19137 4735
tri 19137 4641 19235 4739 sw
tri 19235 4641 19333 4739 ne
rect 19333 4735 20300 4739
rect 19333 4641 19465 4735
rect 19035 4615 19235 4641
rect 18813 4611 19235 4615
tri 19235 4611 19265 4641 sw
tri 19333 4611 19363 4641 ne
rect 19363 4615 19465 4641
rect 19585 4615 20300 4735
rect 19363 4611 20300 4615
tri 113 4513 211 4611 ne
rect 211 4513 565 4611
tri 565 4513 663 4611 sw
tri 663 4513 761 4611 ne
rect 761 4513 1115 4611
tri 1115 4513 1213 4611 sw
tri 1213 4513 1311 4611 ne
rect 1311 4513 1665 4611
tri 1665 4513 1763 4611 sw
tri 1763 4513 1861 4611 ne
rect 1861 4513 2215 4611
tri 2215 4513 2313 4611 sw
tri 2313 4513 2411 4611 ne
rect 2411 4513 2765 4611
tri 2765 4513 2863 4611 sw
tri 2863 4513 2961 4611 ne
rect 2961 4513 3315 4611
tri 3315 4513 3413 4611 sw
tri 3413 4513 3511 4611 ne
rect 3511 4513 3865 4611
tri 3865 4513 3963 4611 sw
tri 3963 4513 4061 4611 ne
rect 4061 4513 4415 4611
tri 4415 4513 4513 4611 sw
tri 4513 4513 4611 4611 ne
rect 4611 4513 4965 4611
tri 4965 4513 5063 4611 sw
tri 5063 4513 5161 4611 ne
rect 5161 4513 5515 4611
tri 5515 4513 5613 4611 sw
tri 5613 4513 5711 4611 ne
rect 5711 4513 6065 4611
tri 6065 4513 6163 4611 sw
tri 6163 4513 6261 4611 ne
rect 6261 4513 6615 4611
tri 6615 4513 6713 4611 sw
tri 6713 4513 6811 4611 ne
rect 6811 4513 7165 4611
tri 7165 4513 7263 4611 sw
tri 7263 4513 7361 4611 ne
rect 7361 4513 7715 4611
tri 7715 4513 7813 4611 sw
tri 7813 4513 7911 4611 ne
rect 7911 4513 8265 4611
tri 8265 4513 8363 4611 sw
tri 8363 4513 8461 4611 ne
rect 8461 4513 8815 4611
tri 8815 4513 8913 4611 sw
tri 8913 4513 9011 4611 ne
rect 9011 4513 9365 4611
tri 9365 4513 9463 4611 sw
tri 9463 4513 9561 4611 ne
rect 9561 4513 9915 4611
tri 9915 4513 10013 4611 sw
tri 10013 4513 10111 4611 ne
rect 10111 4513 10465 4611
tri 10465 4513 10563 4611 sw
tri 10563 4513 10661 4611 ne
rect 10661 4513 11015 4611
tri 11015 4513 11113 4611 sw
tri 11113 4513 11211 4611 ne
rect 11211 4513 11565 4611
tri 11565 4513 11663 4611 sw
tri 11663 4513 11761 4611 ne
rect 11761 4513 12115 4611
tri 12115 4513 12213 4611 sw
tri 12213 4513 12311 4611 ne
rect 12311 4513 12665 4611
tri 12665 4513 12763 4611 sw
tri 12763 4513 12861 4611 ne
rect 12861 4513 13215 4611
tri 13215 4513 13313 4611 sw
tri 13313 4513 13411 4611 ne
rect 13411 4513 13765 4611
tri 13765 4513 13863 4611 sw
tri 13863 4513 13961 4611 ne
rect 13961 4513 14315 4611
tri 14315 4513 14413 4611 sw
tri 14413 4513 14511 4611 ne
rect 14511 4513 14865 4611
tri 14865 4513 14963 4611 sw
tri 14963 4513 15061 4611 ne
rect 15061 4513 15415 4611
tri 15415 4513 15513 4611 sw
tri 15513 4513 15611 4611 ne
rect 15611 4513 15965 4611
tri 15965 4513 16063 4611 sw
tri 16063 4513 16161 4611 ne
rect 16161 4513 16515 4611
tri 16515 4513 16613 4611 sw
tri 16613 4513 16711 4611 ne
rect 16711 4513 17065 4611
tri 17065 4513 17163 4611 sw
tri 17163 4513 17261 4611 ne
rect 17261 4513 17615 4611
tri 17615 4513 17713 4611 sw
tri 17713 4513 17811 4611 ne
rect 17811 4513 18165 4611
tri 18165 4513 18263 4611 sw
tri 18263 4513 18361 4611 ne
rect 18361 4513 18715 4611
tri 18715 4513 18813 4611 sw
tri 18813 4513 18911 4611 ne
rect 18911 4513 19265 4611
tri 19265 4513 19363 4611 sw
tri 19363 4513 19461 4611 ne
rect 19461 4513 20300 4611
rect -2000 4483 113 4513
tri 113 4483 143 4513 sw
tri 211 4483 241 4513 ne
rect 241 4483 663 4513
tri 663 4483 693 4513 sw
tri 761 4483 791 4513 ne
rect 791 4483 1213 4513
tri 1213 4483 1243 4513 sw
tri 1311 4483 1341 4513 ne
rect 1341 4483 1763 4513
tri 1763 4483 1793 4513 sw
tri 1861 4483 1891 4513 ne
rect 1891 4483 2313 4513
tri 2313 4483 2343 4513 sw
tri 2411 4483 2441 4513 ne
rect 2441 4483 2863 4513
tri 2863 4483 2893 4513 sw
tri 2961 4483 2991 4513 ne
rect 2991 4483 3413 4513
tri 3413 4483 3443 4513 sw
tri 3511 4483 3541 4513 ne
rect 3541 4483 3963 4513
tri 3963 4483 3993 4513 sw
tri 4061 4483 4091 4513 ne
rect 4091 4483 4513 4513
tri 4513 4483 4543 4513 sw
tri 4611 4483 4641 4513 ne
rect 4641 4483 5063 4513
tri 5063 4483 5093 4513 sw
tri 5161 4483 5191 4513 ne
rect 5191 4483 5613 4513
tri 5613 4483 5643 4513 sw
tri 5711 4483 5741 4513 ne
rect 5741 4483 6163 4513
tri 6163 4483 6193 4513 sw
tri 6261 4483 6291 4513 ne
rect 6291 4483 6713 4513
tri 6713 4483 6743 4513 sw
tri 6811 4483 6841 4513 ne
rect 6841 4483 7263 4513
tri 7263 4483 7293 4513 sw
tri 7361 4483 7391 4513 ne
rect 7391 4483 7813 4513
tri 7813 4483 7843 4513 sw
tri 7911 4483 7941 4513 ne
rect 7941 4483 8363 4513
tri 8363 4483 8393 4513 sw
tri 8461 4483 8491 4513 ne
rect 8491 4483 8913 4513
tri 8913 4483 8943 4513 sw
tri 9011 4483 9041 4513 ne
rect 9041 4483 9463 4513
tri 9463 4483 9493 4513 sw
tri 9561 4483 9591 4513 ne
rect 9591 4483 10013 4513
tri 10013 4483 10043 4513 sw
tri 10111 4483 10141 4513 ne
rect 10141 4483 10563 4513
tri 10563 4483 10593 4513 sw
tri 10661 4483 10691 4513 ne
rect 10691 4483 11113 4513
tri 11113 4483 11143 4513 sw
tri 11211 4483 11241 4513 ne
rect 11241 4483 11663 4513
tri 11663 4483 11693 4513 sw
tri 11761 4483 11791 4513 ne
rect 11791 4483 12213 4513
tri 12213 4483 12243 4513 sw
tri 12311 4483 12341 4513 ne
rect 12341 4483 12763 4513
tri 12763 4483 12793 4513 sw
tri 12861 4483 12891 4513 ne
rect 12891 4483 13313 4513
tri 13313 4483 13343 4513 sw
tri 13411 4483 13441 4513 ne
rect 13441 4483 13863 4513
tri 13863 4483 13893 4513 sw
tri 13961 4483 13991 4513 ne
rect 13991 4483 14413 4513
tri 14413 4483 14443 4513 sw
tri 14511 4483 14541 4513 ne
rect 14541 4483 14963 4513
tri 14963 4483 14993 4513 sw
tri 15061 4483 15091 4513 ne
rect 15091 4483 15513 4513
tri 15513 4483 15543 4513 sw
tri 15611 4483 15641 4513 ne
rect 15641 4483 16063 4513
tri 16063 4483 16093 4513 sw
tri 16161 4483 16191 4513 ne
rect 16191 4483 16613 4513
tri 16613 4483 16643 4513 sw
tri 16711 4483 16741 4513 ne
rect 16741 4483 17163 4513
tri 17163 4483 17193 4513 sw
tri 17261 4483 17291 4513 ne
rect 17291 4483 17713 4513
tri 17713 4483 17743 4513 sw
tri 17811 4483 17841 4513 ne
rect 17841 4483 18263 4513
tri 18263 4483 18293 4513 sw
tri 18361 4483 18391 4513 ne
rect 18391 4483 18813 4513
tri 18813 4483 18843 4513 sw
tri 18911 4483 18941 4513 ne
rect 18941 4483 19363 4513
tri 19363 4483 19393 4513 sw
tri 19461 4483 19491 4513 ne
rect 19491 4483 20300 4513
rect -2000 4385 143 4483
tri 143 4385 241 4483 sw
tri 241 4385 339 4483 ne
rect 339 4385 693 4483
tri 693 4385 791 4483 sw
tri 791 4385 889 4483 ne
rect 889 4385 1243 4483
tri 1243 4385 1341 4483 sw
tri 1341 4385 1439 4483 ne
rect 1439 4385 1793 4483
tri 1793 4385 1891 4483 sw
tri 1891 4385 1989 4483 ne
rect 1989 4385 2343 4483
tri 2343 4385 2441 4483 sw
tri 2441 4385 2539 4483 ne
rect 2539 4385 2893 4483
tri 2893 4385 2991 4483 sw
tri 2991 4385 3089 4483 ne
rect 3089 4385 3443 4483
tri 3443 4385 3541 4483 sw
tri 3541 4385 3639 4483 ne
rect 3639 4385 3993 4483
tri 3993 4385 4091 4483 sw
tri 4091 4385 4189 4483 ne
rect 4189 4385 4543 4483
tri 4543 4385 4641 4483 sw
tri 4641 4385 4739 4483 ne
rect 4739 4385 5093 4483
tri 5093 4385 5191 4483 sw
tri 5191 4385 5289 4483 ne
rect 5289 4385 5643 4483
tri 5643 4385 5741 4483 sw
tri 5741 4385 5839 4483 ne
rect 5839 4385 6193 4483
tri 6193 4385 6291 4483 sw
tri 6291 4385 6389 4483 ne
rect 6389 4385 6743 4483
tri 6743 4385 6841 4483 sw
tri 6841 4385 6939 4483 ne
rect 6939 4385 7293 4483
tri 7293 4385 7391 4483 sw
tri 7391 4385 7489 4483 ne
rect 7489 4385 7843 4483
tri 7843 4385 7941 4483 sw
tri 7941 4385 8039 4483 ne
rect 8039 4385 8393 4483
tri 8393 4385 8491 4483 sw
tri 8491 4385 8589 4483 ne
rect 8589 4385 8943 4483
tri 8943 4385 9041 4483 sw
tri 9041 4385 9139 4483 ne
rect 9139 4385 9493 4483
tri 9493 4385 9591 4483 sw
tri 9591 4385 9689 4483 ne
rect 9689 4385 10043 4483
tri 10043 4385 10141 4483 sw
tri 10141 4385 10239 4483 ne
rect 10239 4385 10593 4483
tri 10593 4385 10691 4483 sw
tri 10691 4385 10789 4483 ne
rect 10789 4385 11143 4483
tri 11143 4385 11241 4483 sw
tri 11241 4385 11339 4483 ne
rect 11339 4385 11693 4483
tri 11693 4385 11791 4483 sw
tri 11791 4385 11889 4483 ne
rect 11889 4385 12243 4483
tri 12243 4385 12341 4483 sw
tri 12341 4385 12439 4483 ne
rect 12439 4385 12793 4483
tri 12793 4385 12891 4483 sw
tri 12891 4385 12989 4483 ne
rect 12989 4385 13343 4483
tri 13343 4385 13441 4483 sw
tri 13441 4385 13539 4483 ne
rect 13539 4385 13893 4483
tri 13893 4385 13991 4483 sw
tri 13991 4385 14089 4483 ne
rect 14089 4385 14443 4483
tri 14443 4385 14541 4483 sw
tri 14541 4385 14639 4483 ne
rect 14639 4385 14993 4483
tri 14993 4385 15091 4483 sw
tri 15091 4385 15189 4483 ne
rect 15189 4385 15543 4483
tri 15543 4385 15641 4483 sw
tri 15641 4385 15739 4483 ne
rect 15739 4385 16093 4483
tri 16093 4385 16191 4483 sw
tri 16191 4385 16289 4483 ne
rect 16289 4385 16643 4483
tri 16643 4385 16741 4483 sw
tri 16741 4385 16839 4483 ne
rect 16839 4385 17193 4483
tri 17193 4385 17291 4483 sw
tri 17291 4385 17389 4483 ne
rect 17389 4385 17743 4483
tri 17743 4385 17841 4483 sw
tri 17841 4385 17939 4483 ne
rect 17939 4385 18293 4483
tri 18293 4385 18391 4483 sw
tri 18391 4385 18489 4483 ne
rect 18489 4385 18843 4483
tri 18843 4385 18941 4483 sw
tri 18941 4385 19039 4483 ne
rect 19039 4385 19393 4483
tri 19393 4385 19491 4483 sw
tri 19491 4385 19589 4483 ne
rect 19589 4385 20300 4483
rect -2000 4287 241 4385
tri 241 4287 339 4385 sw
tri 339 4287 437 4385 ne
rect 437 4287 791 4385
tri 791 4287 889 4385 sw
tri 889 4287 987 4385 ne
rect 987 4287 1341 4385
tri 1341 4287 1439 4385 sw
tri 1439 4287 1537 4385 ne
rect 1537 4287 1891 4385
tri 1891 4287 1989 4385 sw
tri 1989 4287 2087 4385 ne
rect 2087 4287 2441 4385
tri 2441 4287 2539 4385 sw
tri 2539 4287 2637 4385 ne
rect 2637 4287 2991 4385
tri 2991 4287 3089 4385 sw
tri 3089 4287 3187 4385 ne
rect 3187 4287 3541 4385
tri 3541 4287 3639 4385 sw
tri 3639 4287 3737 4385 ne
rect 3737 4287 4091 4385
tri 4091 4287 4189 4385 sw
tri 4189 4287 4287 4385 ne
rect 4287 4287 4641 4385
tri 4641 4287 4739 4385 sw
tri 4739 4287 4837 4385 ne
rect 4837 4287 5191 4385
tri 5191 4287 5289 4385 sw
tri 5289 4287 5387 4385 ne
rect 5387 4287 5741 4385
tri 5741 4287 5839 4385 sw
tri 5839 4287 5937 4385 ne
rect 5937 4287 6291 4385
tri 6291 4287 6389 4385 sw
tri 6389 4287 6487 4385 ne
rect 6487 4287 6841 4385
tri 6841 4287 6939 4385 sw
tri 6939 4287 7037 4385 ne
rect 7037 4287 7391 4385
tri 7391 4287 7489 4385 sw
tri 7489 4287 7587 4385 ne
rect 7587 4287 7941 4385
tri 7941 4287 8039 4385 sw
tri 8039 4287 8137 4385 ne
rect 8137 4287 8491 4385
tri 8491 4287 8589 4385 sw
tri 8589 4287 8687 4385 ne
rect 8687 4287 9041 4385
tri 9041 4287 9139 4385 sw
tri 9139 4287 9237 4385 ne
rect 9237 4287 9591 4385
tri 9591 4287 9689 4385 sw
tri 9689 4287 9787 4385 ne
rect 9787 4287 10141 4385
tri 10141 4287 10239 4385 sw
tri 10239 4287 10337 4385 ne
rect 10337 4287 10691 4385
tri 10691 4287 10789 4385 sw
tri 10789 4287 10887 4385 ne
rect 10887 4287 11241 4385
tri 11241 4287 11339 4385 sw
tri 11339 4287 11437 4385 ne
rect 11437 4287 11791 4385
tri 11791 4287 11889 4385 sw
tri 11889 4287 11987 4385 ne
rect 11987 4287 12341 4385
tri 12341 4287 12439 4385 sw
tri 12439 4287 12537 4385 ne
rect 12537 4287 12891 4385
tri 12891 4287 12989 4385 sw
tri 12989 4287 13087 4385 ne
rect 13087 4287 13441 4385
tri 13441 4287 13539 4385 sw
tri 13539 4287 13637 4385 ne
rect 13637 4287 13991 4385
tri 13991 4287 14089 4385 sw
tri 14089 4287 14187 4385 ne
rect 14187 4287 14541 4385
tri 14541 4287 14639 4385 sw
tri 14639 4287 14737 4385 ne
rect 14737 4287 15091 4385
tri 15091 4287 15189 4385 sw
tri 15189 4287 15287 4385 ne
rect 15287 4287 15641 4385
tri 15641 4287 15739 4385 sw
tri 15739 4287 15837 4385 ne
rect 15837 4287 16191 4385
tri 16191 4287 16289 4385 sw
tri 16289 4287 16387 4385 ne
rect 16387 4287 16741 4385
tri 16741 4287 16839 4385 sw
tri 16839 4287 16937 4385 ne
rect 16937 4287 17291 4385
tri 17291 4287 17389 4385 sw
tri 17389 4287 17487 4385 ne
rect 17487 4287 17841 4385
tri 17841 4287 17939 4385 sw
tri 17939 4287 18037 4385 ne
rect 18037 4287 18391 4385
tri 18391 4287 18489 4385 sw
tri 18489 4287 18587 4385 ne
rect 18587 4287 18941 4385
tri 18941 4287 19039 4385 sw
tri 19039 4287 19137 4385 ne
rect 19137 4287 19491 4385
tri 19491 4287 19589 4385 sw
tri 19589 4287 19687 4385 ne
rect 19687 4287 20300 4385
rect -2000 4189 339 4287
tri 339 4189 437 4287 sw
tri 437 4189 535 4287 ne
rect 535 4189 889 4287
tri 889 4189 987 4287 sw
tri 987 4189 1085 4287 ne
rect 1085 4189 1439 4287
tri 1439 4189 1537 4287 sw
tri 1537 4189 1635 4287 ne
rect 1635 4189 1989 4287
tri 1989 4189 2087 4287 sw
tri 2087 4189 2185 4287 ne
rect 2185 4189 2539 4287
tri 2539 4189 2637 4287 sw
tri 2637 4189 2735 4287 ne
rect 2735 4189 3089 4287
tri 3089 4189 3187 4287 sw
tri 3187 4189 3285 4287 ne
rect 3285 4189 3639 4287
tri 3639 4189 3737 4287 sw
tri 3737 4189 3835 4287 ne
rect 3835 4189 4189 4287
tri 4189 4189 4287 4287 sw
tri 4287 4189 4385 4287 ne
rect 4385 4189 4739 4287
tri 4739 4189 4837 4287 sw
tri 4837 4189 4935 4287 ne
rect 4935 4189 5289 4287
tri 5289 4189 5387 4287 sw
tri 5387 4189 5485 4287 ne
rect 5485 4189 5839 4287
tri 5839 4189 5937 4287 sw
tri 5937 4189 6035 4287 ne
rect 6035 4189 6389 4287
tri 6389 4189 6487 4287 sw
tri 6487 4189 6585 4287 ne
rect 6585 4189 6939 4287
tri 6939 4189 7037 4287 sw
tri 7037 4189 7135 4287 ne
rect 7135 4189 7489 4287
tri 7489 4189 7587 4287 sw
tri 7587 4189 7685 4287 ne
rect 7685 4189 8039 4287
tri 8039 4189 8137 4287 sw
tri 8137 4189 8235 4287 ne
rect 8235 4189 8589 4287
tri 8589 4189 8687 4287 sw
tri 8687 4189 8785 4287 ne
rect 8785 4189 9139 4287
tri 9139 4189 9237 4287 sw
tri 9237 4189 9335 4287 ne
rect 9335 4189 9689 4287
tri 9689 4189 9787 4287 sw
tri 9787 4189 9885 4287 ne
rect 9885 4189 10239 4287
tri 10239 4189 10337 4287 sw
tri 10337 4189 10435 4287 ne
rect 10435 4189 10789 4287
tri 10789 4189 10887 4287 sw
tri 10887 4189 10985 4287 ne
rect 10985 4189 11339 4287
tri 11339 4189 11437 4287 sw
tri 11437 4189 11535 4287 ne
rect 11535 4189 11889 4287
tri 11889 4189 11987 4287 sw
tri 11987 4189 12085 4287 ne
rect 12085 4189 12439 4287
tri 12439 4189 12537 4287 sw
tri 12537 4189 12635 4287 ne
rect 12635 4189 12989 4287
tri 12989 4189 13087 4287 sw
tri 13087 4189 13185 4287 ne
rect 13185 4189 13539 4287
tri 13539 4189 13637 4287 sw
tri 13637 4189 13735 4287 ne
rect 13735 4189 14089 4287
tri 14089 4189 14187 4287 sw
tri 14187 4189 14285 4287 ne
rect 14285 4189 14639 4287
tri 14639 4189 14737 4287 sw
tri 14737 4189 14835 4287 ne
rect 14835 4189 15189 4287
tri 15189 4189 15287 4287 sw
tri 15287 4189 15385 4287 ne
rect 15385 4189 15739 4287
tri 15739 4189 15837 4287 sw
tri 15837 4189 15935 4287 ne
rect 15935 4189 16289 4287
tri 16289 4189 16387 4287 sw
tri 16387 4189 16485 4287 ne
rect 16485 4189 16839 4287
tri 16839 4189 16937 4287 sw
tri 16937 4189 17035 4287 ne
rect 17035 4189 17389 4287
tri 17389 4189 17487 4287 sw
tri 17487 4189 17585 4287 ne
rect 17585 4189 17939 4287
tri 17939 4189 18037 4287 sw
tri 18037 4189 18135 4287 ne
rect 18135 4189 18489 4287
tri 18489 4189 18587 4287 sw
tri 18587 4189 18685 4287 ne
rect 18685 4189 19039 4287
tri 19039 4189 19137 4287 sw
tri 19137 4189 19235 4287 ne
rect 19235 4189 19589 4287
tri 19589 4189 19687 4287 sw
rect 20800 4189 21800 4837
rect -2000 4185 437 4189
rect -2000 4065 215 4185
rect 335 4091 437 4185
tri 437 4091 535 4189 sw
tri 535 4091 633 4189 ne
rect 633 4185 987 4189
rect 633 4091 765 4185
rect 335 4065 535 4091
rect -2000 4061 535 4065
rect -2000 3413 -1000 4061
tri 113 3963 211 4061 ne
rect 211 4013 535 4061
tri 535 4013 613 4091 sw
tri 633 4013 711 4091 ne
rect 711 4065 765 4091
rect 885 4091 987 4185
tri 987 4091 1085 4189 sw
tri 1085 4091 1183 4189 ne
rect 1183 4185 1537 4189
rect 1183 4091 1315 4185
rect 885 4065 1085 4091
rect 711 4013 1085 4065
tri 1085 4013 1163 4091 sw
tri 1183 4013 1261 4091 ne
rect 1261 4065 1315 4091
rect 1435 4091 1537 4185
tri 1537 4091 1635 4189 sw
tri 1635 4091 1733 4189 ne
rect 1733 4185 2087 4189
rect 1733 4091 1865 4185
rect 1435 4065 1635 4091
rect 1261 4013 1635 4065
tri 1635 4013 1713 4091 sw
tri 1733 4013 1811 4091 ne
rect 1811 4065 1865 4091
rect 1985 4091 2087 4185
tri 2087 4091 2185 4189 sw
tri 2185 4091 2283 4189 ne
rect 2283 4185 2637 4189
rect 2283 4091 2415 4185
rect 1985 4065 2185 4091
rect 1811 4013 2185 4065
tri 2185 4013 2263 4091 sw
tri 2283 4013 2361 4091 ne
rect 2361 4065 2415 4091
rect 2535 4091 2637 4185
tri 2637 4091 2735 4189 sw
tri 2735 4091 2833 4189 ne
rect 2833 4185 3187 4189
rect 2833 4091 2965 4185
rect 2535 4065 2735 4091
rect 2361 4013 2735 4065
tri 2735 4013 2813 4091 sw
tri 2833 4013 2911 4091 ne
rect 2911 4065 2965 4091
rect 3085 4091 3187 4185
tri 3187 4091 3285 4189 sw
tri 3285 4091 3383 4189 ne
rect 3383 4185 3737 4189
rect 3383 4091 3515 4185
rect 3085 4065 3285 4091
rect 2911 4013 3285 4065
tri 3285 4013 3363 4091 sw
tri 3383 4013 3461 4091 ne
rect 3461 4065 3515 4091
rect 3635 4091 3737 4185
tri 3737 4091 3835 4189 sw
tri 3835 4091 3933 4189 ne
rect 3933 4185 4287 4189
rect 3933 4091 4065 4185
rect 3635 4065 3835 4091
rect 3461 4013 3835 4065
tri 3835 4013 3913 4091 sw
tri 3933 4013 4011 4091 ne
rect 4011 4065 4065 4091
rect 4185 4091 4287 4185
tri 4287 4091 4385 4189 sw
tri 4385 4091 4483 4189 ne
rect 4483 4185 4837 4189
rect 4483 4091 4615 4185
rect 4185 4065 4385 4091
rect 4011 4013 4385 4065
tri 4385 4013 4463 4091 sw
tri 4483 4013 4561 4091 ne
rect 4561 4065 4615 4091
rect 4735 4091 4837 4185
tri 4837 4091 4935 4189 sw
tri 4935 4091 5033 4189 ne
rect 5033 4185 5387 4189
rect 5033 4091 5165 4185
rect 4735 4065 4935 4091
rect 4561 4013 4935 4065
tri 4935 4013 5013 4091 sw
tri 5033 4013 5111 4091 ne
rect 5111 4065 5165 4091
rect 5285 4091 5387 4185
tri 5387 4091 5485 4189 sw
tri 5485 4091 5583 4189 ne
rect 5583 4185 5937 4189
rect 5583 4091 5715 4185
rect 5285 4065 5485 4091
rect 5111 4013 5485 4065
tri 5485 4013 5563 4091 sw
tri 5583 4013 5661 4091 ne
rect 5661 4065 5715 4091
rect 5835 4091 5937 4185
tri 5937 4091 6035 4189 sw
tri 6035 4091 6133 4189 ne
rect 6133 4185 6487 4189
rect 6133 4091 6265 4185
rect 5835 4065 6035 4091
rect 5661 4013 6035 4065
tri 6035 4013 6113 4091 sw
tri 6133 4013 6211 4091 ne
rect 6211 4065 6265 4091
rect 6385 4091 6487 4185
tri 6487 4091 6585 4189 sw
tri 6585 4091 6683 4189 ne
rect 6683 4185 7037 4189
rect 6683 4091 6815 4185
rect 6385 4065 6585 4091
rect 6211 4013 6585 4065
tri 6585 4013 6663 4091 sw
tri 6683 4013 6761 4091 ne
rect 6761 4065 6815 4091
rect 6935 4091 7037 4185
tri 7037 4091 7135 4189 sw
tri 7135 4091 7233 4189 ne
rect 7233 4185 7587 4189
rect 7233 4091 7365 4185
rect 6935 4065 7135 4091
rect 6761 4013 7135 4065
tri 7135 4013 7213 4091 sw
tri 7233 4013 7311 4091 ne
rect 7311 4065 7365 4091
rect 7485 4091 7587 4185
tri 7587 4091 7685 4189 sw
tri 7685 4091 7783 4189 ne
rect 7783 4185 8137 4189
rect 7783 4091 7915 4185
rect 7485 4065 7685 4091
rect 7311 4013 7685 4065
tri 7685 4013 7763 4091 sw
tri 7783 4013 7861 4091 ne
rect 7861 4065 7915 4091
rect 8035 4091 8137 4185
tri 8137 4091 8235 4189 sw
tri 8235 4091 8333 4189 ne
rect 8333 4185 8687 4189
rect 8333 4091 8465 4185
rect 8035 4065 8235 4091
rect 7861 4013 8235 4065
tri 8235 4013 8313 4091 sw
tri 8333 4013 8411 4091 ne
rect 8411 4065 8465 4091
rect 8585 4091 8687 4185
tri 8687 4091 8785 4189 sw
tri 8785 4091 8883 4189 ne
rect 8883 4185 9237 4189
rect 8883 4091 9015 4185
rect 8585 4065 8785 4091
rect 8411 4013 8785 4065
tri 8785 4013 8863 4091 sw
tri 8883 4013 8961 4091 ne
rect 8961 4065 9015 4091
rect 9135 4091 9237 4185
tri 9237 4091 9335 4189 sw
tri 9335 4091 9433 4189 ne
rect 9433 4185 9787 4189
rect 9433 4091 9565 4185
rect 9135 4065 9335 4091
rect 8961 4013 9335 4065
tri 9335 4013 9413 4091 sw
tri 9433 4013 9511 4091 ne
rect 9511 4065 9565 4091
rect 9685 4091 9787 4185
tri 9787 4091 9885 4189 sw
tri 9885 4091 9983 4189 ne
rect 9983 4185 10337 4189
rect 9983 4091 10115 4185
rect 9685 4065 9885 4091
rect 9511 4013 9885 4065
tri 9885 4013 9963 4091 sw
tri 9983 4013 10061 4091 ne
rect 10061 4065 10115 4091
rect 10235 4091 10337 4185
tri 10337 4091 10435 4189 sw
tri 10435 4091 10533 4189 ne
rect 10533 4185 10887 4189
rect 10533 4091 10665 4185
rect 10235 4065 10435 4091
rect 10061 4013 10435 4065
tri 10435 4013 10513 4091 sw
tri 10533 4013 10611 4091 ne
rect 10611 4065 10665 4091
rect 10785 4091 10887 4185
tri 10887 4091 10985 4189 sw
tri 10985 4091 11083 4189 ne
rect 11083 4185 11437 4189
rect 11083 4091 11215 4185
rect 10785 4065 10985 4091
rect 10611 4013 10985 4065
tri 10985 4013 11063 4091 sw
tri 11083 4013 11161 4091 ne
rect 11161 4065 11215 4091
rect 11335 4091 11437 4185
tri 11437 4091 11535 4189 sw
tri 11535 4091 11633 4189 ne
rect 11633 4185 11987 4189
rect 11633 4091 11765 4185
rect 11335 4065 11535 4091
rect 11161 4013 11535 4065
tri 11535 4013 11613 4091 sw
tri 11633 4013 11711 4091 ne
rect 11711 4065 11765 4091
rect 11885 4091 11987 4185
tri 11987 4091 12085 4189 sw
tri 12085 4091 12183 4189 ne
rect 12183 4185 12537 4189
rect 12183 4091 12315 4185
rect 11885 4065 12085 4091
rect 11711 4013 12085 4065
tri 12085 4013 12163 4091 sw
tri 12183 4013 12261 4091 ne
rect 12261 4065 12315 4091
rect 12435 4091 12537 4185
tri 12537 4091 12635 4189 sw
tri 12635 4091 12733 4189 ne
rect 12733 4185 13087 4189
rect 12733 4091 12865 4185
rect 12435 4065 12635 4091
rect 12261 4013 12635 4065
tri 12635 4013 12713 4091 sw
tri 12733 4013 12811 4091 ne
rect 12811 4065 12865 4091
rect 12985 4091 13087 4185
tri 13087 4091 13185 4189 sw
tri 13185 4091 13283 4189 ne
rect 13283 4185 13637 4189
rect 13283 4091 13415 4185
rect 12985 4065 13185 4091
rect 12811 4013 13185 4065
tri 13185 4013 13263 4091 sw
tri 13283 4013 13361 4091 ne
rect 13361 4065 13415 4091
rect 13535 4091 13637 4185
tri 13637 4091 13735 4189 sw
tri 13735 4091 13833 4189 ne
rect 13833 4185 14187 4189
rect 13833 4091 13965 4185
rect 13535 4065 13735 4091
rect 13361 4013 13735 4065
tri 13735 4013 13813 4091 sw
tri 13833 4013 13911 4091 ne
rect 13911 4065 13965 4091
rect 14085 4091 14187 4185
tri 14187 4091 14285 4189 sw
tri 14285 4091 14383 4189 ne
rect 14383 4185 14737 4189
rect 14383 4091 14515 4185
rect 14085 4065 14285 4091
rect 13911 4013 14285 4065
tri 14285 4013 14363 4091 sw
tri 14383 4013 14461 4091 ne
rect 14461 4065 14515 4091
rect 14635 4091 14737 4185
tri 14737 4091 14835 4189 sw
tri 14835 4091 14933 4189 ne
rect 14933 4185 15287 4189
rect 14933 4091 15065 4185
rect 14635 4065 14835 4091
rect 14461 4013 14835 4065
tri 14835 4013 14913 4091 sw
tri 14933 4013 15011 4091 ne
rect 15011 4065 15065 4091
rect 15185 4091 15287 4185
tri 15287 4091 15385 4189 sw
tri 15385 4091 15483 4189 ne
rect 15483 4185 15837 4189
rect 15483 4091 15615 4185
rect 15185 4065 15385 4091
rect 15011 4013 15385 4065
tri 15385 4013 15463 4091 sw
tri 15483 4013 15561 4091 ne
rect 15561 4065 15615 4091
rect 15735 4091 15837 4185
tri 15837 4091 15935 4189 sw
tri 15935 4091 16033 4189 ne
rect 16033 4185 16387 4189
rect 16033 4091 16165 4185
rect 15735 4065 15935 4091
rect 15561 4013 15935 4065
tri 15935 4013 16013 4091 sw
tri 16033 4013 16111 4091 ne
rect 16111 4065 16165 4091
rect 16285 4091 16387 4185
tri 16387 4091 16485 4189 sw
tri 16485 4091 16583 4189 ne
rect 16583 4185 16937 4189
rect 16583 4091 16715 4185
rect 16285 4065 16485 4091
rect 16111 4013 16485 4065
tri 16485 4013 16563 4091 sw
tri 16583 4013 16661 4091 ne
rect 16661 4065 16715 4091
rect 16835 4091 16937 4185
tri 16937 4091 17035 4189 sw
tri 17035 4091 17133 4189 ne
rect 17133 4185 17487 4189
rect 17133 4091 17265 4185
rect 16835 4065 17035 4091
rect 16661 4013 17035 4065
tri 17035 4013 17113 4091 sw
tri 17133 4013 17211 4091 ne
rect 17211 4065 17265 4091
rect 17385 4091 17487 4185
tri 17487 4091 17585 4189 sw
tri 17585 4091 17683 4189 ne
rect 17683 4185 18037 4189
rect 17683 4091 17815 4185
rect 17385 4065 17585 4091
rect 17211 4013 17585 4065
tri 17585 4013 17663 4091 sw
tri 17683 4013 17761 4091 ne
rect 17761 4065 17815 4091
rect 17935 4091 18037 4185
tri 18037 4091 18135 4189 sw
tri 18135 4091 18233 4189 ne
rect 18233 4185 18587 4189
rect 18233 4091 18365 4185
rect 17935 4065 18135 4091
rect 17761 4013 18135 4065
tri 18135 4013 18213 4091 sw
tri 18233 4013 18311 4091 ne
rect 18311 4065 18365 4091
rect 18485 4091 18587 4185
tri 18587 4091 18685 4189 sw
tri 18685 4091 18783 4189 ne
rect 18783 4185 19137 4189
rect 18783 4091 18915 4185
rect 18485 4065 18685 4091
rect 18311 4013 18685 4065
tri 18685 4013 18763 4091 sw
tri 18783 4013 18861 4091 ne
rect 18861 4065 18915 4091
rect 19035 4091 19137 4185
tri 19137 4091 19235 4189 sw
tri 19235 4091 19333 4189 ne
rect 19333 4185 21800 4189
rect 19333 4091 19465 4185
rect 19035 4065 19235 4091
rect 18861 4013 19235 4065
tri 19235 4013 19313 4091 sw
tri 19333 4013 19411 4091 ne
rect 19411 4065 19465 4091
rect 19585 4065 21800 4185
rect 19411 4013 21800 4065
rect 211 3963 613 4013
rect -500 3913 113 3963
tri 113 3913 163 3963 sw
tri 211 3913 261 3963 ne
rect 261 3933 613 3963
tri 613 3933 693 4013 sw
tri 711 3933 791 4013 ne
rect 791 3933 1163 4013
tri 1163 3933 1243 4013 sw
tri 1261 3933 1341 4013 ne
rect 1341 3933 1713 4013
tri 1713 3933 1793 4013 sw
tri 1811 3933 1891 4013 ne
rect 1891 3933 2263 4013
tri 2263 3933 2343 4013 sw
tri 2361 3933 2441 4013 ne
rect 2441 3933 2813 4013
tri 2813 3933 2893 4013 sw
tri 2911 3933 2991 4013 ne
rect 2991 3933 3363 4013
tri 3363 3933 3443 4013 sw
tri 3461 3933 3541 4013 ne
rect 3541 3933 3913 4013
tri 3913 3933 3993 4013 sw
tri 4011 3933 4091 4013 ne
rect 4091 3933 4463 4013
tri 4463 3933 4543 4013 sw
tri 4561 3933 4641 4013 ne
rect 4641 3933 5013 4013
tri 5013 3933 5093 4013 sw
tri 5111 3933 5191 4013 ne
rect 5191 3933 5563 4013
tri 5563 3933 5643 4013 sw
tri 5661 3933 5741 4013 ne
rect 5741 3933 6113 4013
tri 6113 3933 6193 4013 sw
tri 6211 3933 6291 4013 ne
rect 6291 3933 6663 4013
tri 6663 3933 6743 4013 sw
tri 6761 3933 6841 4013 ne
rect 6841 3933 7213 4013
tri 7213 3933 7293 4013 sw
tri 7311 3933 7391 4013 ne
rect 7391 3933 7763 4013
tri 7763 3933 7843 4013 sw
tri 7861 3933 7941 4013 ne
rect 7941 3933 8313 4013
tri 8313 3933 8393 4013 sw
tri 8411 3933 8491 4013 ne
rect 8491 3933 8863 4013
tri 8863 3933 8943 4013 sw
tri 8961 3933 9041 4013 ne
rect 9041 3933 9413 4013
tri 9413 3933 9493 4013 sw
tri 9511 3933 9591 4013 ne
rect 9591 3933 9963 4013
tri 9963 3933 10043 4013 sw
tri 10061 3933 10141 4013 ne
rect 10141 3933 10513 4013
tri 10513 3933 10593 4013 sw
tri 10611 3933 10691 4013 ne
rect 10691 3933 11063 4013
tri 11063 3933 11143 4013 sw
tri 11161 3933 11241 4013 ne
rect 11241 3933 11613 4013
tri 11613 3933 11693 4013 sw
tri 11711 3933 11791 4013 ne
rect 11791 3933 12163 4013
tri 12163 3933 12243 4013 sw
tri 12261 3933 12341 4013 ne
rect 12341 3933 12713 4013
tri 12713 3933 12793 4013 sw
tri 12811 3933 12891 4013 ne
rect 12891 3933 13263 4013
tri 13263 3933 13343 4013 sw
tri 13361 3933 13441 4013 ne
rect 13441 3933 13813 4013
tri 13813 3933 13893 4013 sw
tri 13911 3933 13991 4013 ne
rect 13991 3933 14363 4013
tri 14363 3933 14443 4013 sw
tri 14461 3933 14541 4013 ne
rect 14541 3933 14913 4013
tri 14913 3933 14993 4013 sw
tri 15011 3933 15091 4013 ne
rect 15091 3933 15463 4013
tri 15463 3933 15543 4013 sw
tri 15561 3933 15641 4013 ne
rect 15641 3933 16013 4013
tri 16013 3933 16093 4013 sw
tri 16111 3933 16191 4013 ne
rect 16191 3933 16563 4013
tri 16563 3933 16643 4013 sw
tri 16661 3933 16741 4013 ne
rect 16741 3933 17113 4013
tri 17113 3933 17193 4013 sw
tri 17211 3933 17291 4013 ne
rect 17291 3933 17663 4013
tri 17663 3933 17743 4013 sw
tri 17761 3933 17841 4013 ne
rect 17841 3933 18213 4013
tri 18213 3933 18293 4013 sw
tri 18311 3933 18391 4013 ne
rect 18391 3933 18763 4013
tri 18763 3933 18843 4013 sw
tri 18861 3933 18941 4013 ne
rect 18941 3933 19313 4013
tri 19313 3933 19393 4013 sw
tri 19411 3933 19491 4013 ne
rect 19491 3933 20100 4013
rect 261 3913 693 3933
rect -500 3835 163 3913
tri 163 3835 241 3913 sw
tri 261 3835 339 3913 ne
rect 339 3835 693 3913
tri 693 3835 791 3933 sw
tri 791 3835 889 3933 ne
rect 889 3835 1243 3933
tri 1243 3835 1341 3933 sw
tri 1341 3835 1439 3933 ne
rect 1439 3835 1793 3933
tri 1793 3835 1891 3933 sw
tri 1891 3835 1989 3933 ne
rect 1989 3835 2343 3933
tri 2343 3835 2441 3933 sw
tri 2441 3835 2539 3933 ne
rect 2539 3835 2893 3933
tri 2893 3835 2991 3933 sw
tri 2991 3835 3089 3933 ne
rect 3089 3835 3443 3933
tri 3443 3835 3541 3933 sw
tri 3541 3835 3639 3933 ne
rect 3639 3835 3993 3933
tri 3993 3835 4091 3933 sw
tri 4091 3835 4189 3933 ne
rect 4189 3835 4543 3933
tri 4543 3835 4641 3933 sw
tri 4641 3835 4739 3933 ne
rect 4739 3835 5093 3933
tri 5093 3835 5191 3933 sw
tri 5191 3835 5289 3933 ne
rect 5289 3835 5643 3933
tri 5643 3835 5741 3933 sw
tri 5741 3835 5839 3933 ne
rect 5839 3835 6193 3933
tri 6193 3835 6291 3933 sw
tri 6291 3835 6389 3933 ne
rect 6389 3835 6743 3933
tri 6743 3835 6841 3933 sw
tri 6841 3835 6939 3933 ne
rect 6939 3835 7293 3933
tri 7293 3835 7391 3933 sw
tri 7391 3835 7489 3933 ne
rect 7489 3835 7843 3933
tri 7843 3835 7941 3933 sw
tri 7941 3835 8039 3933 ne
rect 8039 3835 8393 3933
tri 8393 3835 8491 3933 sw
tri 8491 3835 8589 3933 ne
rect 8589 3835 8943 3933
tri 8943 3835 9041 3933 sw
tri 9041 3835 9139 3933 ne
rect 9139 3835 9493 3933
tri 9493 3835 9591 3933 sw
tri 9591 3835 9689 3933 ne
rect 9689 3835 10043 3933
tri 10043 3835 10141 3933 sw
tri 10141 3835 10239 3933 ne
rect 10239 3835 10593 3933
tri 10593 3835 10691 3933 sw
tri 10691 3835 10789 3933 ne
rect 10789 3835 11143 3933
tri 11143 3835 11241 3933 sw
tri 11241 3835 11339 3933 ne
rect 11339 3835 11693 3933
tri 11693 3835 11791 3933 sw
tri 11791 3835 11889 3933 ne
rect 11889 3835 12243 3933
tri 12243 3835 12341 3933 sw
tri 12341 3835 12439 3933 ne
rect 12439 3835 12793 3933
tri 12793 3835 12891 3933 sw
tri 12891 3835 12989 3933 ne
rect 12989 3835 13343 3933
tri 13343 3835 13441 3933 sw
tri 13441 3835 13539 3933 ne
rect 13539 3835 13893 3933
tri 13893 3835 13991 3933 sw
tri 13991 3835 14089 3933 ne
rect 14089 3835 14443 3933
tri 14443 3835 14541 3933 sw
tri 14541 3835 14639 3933 ne
rect 14639 3835 14993 3933
tri 14993 3835 15091 3933 sw
tri 15091 3835 15189 3933 ne
rect 15189 3835 15543 3933
tri 15543 3835 15641 3933 sw
tri 15641 3835 15739 3933 ne
rect 15739 3835 16093 3933
tri 16093 3835 16191 3933 sw
tri 16191 3835 16289 3933 ne
rect 16289 3835 16643 3933
tri 16643 3835 16741 3933 sw
tri 16741 3835 16839 3933 ne
rect 16839 3835 17193 3933
tri 17193 3835 17291 3933 sw
tri 17291 3835 17389 3933 ne
rect 17389 3835 17743 3933
tri 17743 3835 17841 3933 sw
tri 17841 3835 17939 3933 ne
rect 17939 3835 18293 3933
tri 18293 3835 18391 3933 sw
tri 18391 3835 18489 3933 ne
rect 18489 3835 18843 3933
tri 18843 3835 18941 3933 sw
tri 18941 3835 19039 3933 ne
rect 19039 3835 19393 3933
tri 19393 3835 19491 3933 sw
tri 19491 3835 19589 3933 ne
rect 19589 3913 20100 3933
rect 20200 3913 21800 4013
rect 19589 3835 21800 3913
rect -500 3787 241 3835
rect -500 3687 -400 3787
rect -300 3737 241 3787
tri 241 3737 339 3835 sw
tri 339 3737 437 3835 ne
rect 437 3737 791 3835
tri 791 3737 889 3835 sw
tri 889 3737 987 3835 ne
rect 987 3737 1341 3835
tri 1341 3737 1439 3835 sw
tri 1439 3737 1537 3835 ne
rect 1537 3737 1891 3835
tri 1891 3737 1989 3835 sw
tri 1989 3737 2087 3835 ne
rect 2087 3737 2441 3835
tri 2441 3737 2539 3835 sw
tri 2539 3737 2637 3835 ne
rect 2637 3737 2991 3835
tri 2991 3737 3089 3835 sw
tri 3089 3737 3187 3835 ne
rect 3187 3737 3541 3835
tri 3541 3737 3639 3835 sw
tri 3639 3737 3737 3835 ne
rect 3737 3737 4091 3835
tri 4091 3737 4189 3835 sw
tri 4189 3737 4287 3835 ne
rect 4287 3737 4641 3835
tri 4641 3737 4739 3835 sw
tri 4739 3737 4837 3835 ne
rect 4837 3737 5191 3835
tri 5191 3737 5289 3835 sw
tri 5289 3737 5387 3835 ne
rect 5387 3737 5741 3835
tri 5741 3737 5839 3835 sw
tri 5839 3737 5937 3835 ne
rect 5937 3737 6291 3835
tri 6291 3737 6389 3835 sw
tri 6389 3737 6487 3835 ne
rect 6487 3737 6841 3835
tri 6841 3737 6939 3835 sw
tri 6939 3737 7037 3835 ne
rect 7037 3737 7391 3835
tri 7391 3737 7489 3835 sw
tri 7489 3737 7587 3835 ne
rect 7587 3737 7941 3835
tri 7941 3737 8039 3835 sw
tri 8039 3737 8137 3835 ne
rect 8137 3737 8491 3835
tri 8491 3737 8589 3835 sw
tri 8589 3737 8687 3835 ne
rect 8687 3737 9041 3835
tri 9041 3737 9139 3835 sw
tri 9139 3737 9237 3835 ne
rect 9237 3737 9591 3835
tri 9591 3737 9689 3835 sw
tri 9689 3737 9787 3835 ne
rect 9787 3737 10141 3835
tri 10141 3737 10239 3835 sw
tri 10239 3737 10337 3835 ne
rect 10337 3737 10691 3835
tri 10691 3737 10789 3835 sw
tri 10789 3737 10887 3835 ne
rect 10887 3737 11241 3835
tri 11241 3737 11339 3835 sw
tri 11339 3737 11437 3835 ne
rect 11437 3737 11791 3835
tri 11791 3737 11889 3835 sw
tri 11889 3737 11987 3835 ne
rect 11987 3737 12341 3835
tri 12341 3737 12439 3835 sw
tri 12439 3737 12537 3835 ne
rect 12537 3737 12891 3835
tri 12891 3737 12989 3835 sw
tri 12989 3737 13087 3835 ne
rect 13087 3737 13441 3835
tri 13441 3737 13539 3835 sw
tri 13539 3737 13637 3835 ne
rect 13637 3737 13991 3835
tri 13991 3737 14089 3835 sw
tri 14089 3737 14187 3835 ne
rect 14187 3737 14541 3835
tri 14541 3737 14639 3835 sw
tri 14639 3737 14737 3835 ne
rect 14737 3737 15091 3835
tri 15091 3737 15189 3835 sw
tri 15189 3737 15287 3835 ne
rect 15287 3737 15641 3835
tri 15641 3737 15739 3835 sw
tri 15739 3737 15837 3835 ne
rect 15837 3737 16191 3835
tri 16191 3737 16289 3835 sw
tri 16289 3737 16387 3835 ne
rect 16387 3737 16741 3835
tri 16741 3737 16839 3835 sw
tri 16839 3737 16937 3835 ne
rect 16937 3737 17291 3835
tri 17291 3737 17389 3835 sw
tri 17389 3737 17487 3835 ne
rect 17487 3737 17841 3835
tri 17841 3737 17939 3835 sw
tri 17939 3737 18037 3835 ne
rect 18037 3737 18391 3835
tri 18391 3737 18489 3835 sw
tri 18489 3737 18587 3835 ne
rect 18587 3737 18941 3835
tri 18941 3737 19039 3835 sw
tri 19039 3737 19137 3835 ne
rect 19137 3737 19491 3835
tri 19491 3737 19589 3835 sw
tri 19589 3737 19687 3835 ne
rect 19687 3737 21800 3835
rect -300 3687 339 3737
rect -500 3639 339 3687
tri 339 3639 437 3737 sw
tri 437 3639 535 3737 ne
rect 535 3639 889 3737
tri 889 3639 987 3737 sw
tri 987 3639 1085 3737 ne
rect 1085 3639 1439 3737
tri 1439 3639 1537 3737 sw
tri 1537 3639 1635 3737 ne
rect 1635 3639 1989 3737
tri 1989 3639 2087 3737 sw
tri 2087 3639 2185 3737 ne
rect 2185 3639 2539 3737
tri 2539 3639 2637 3737 sw
tri 2637 3639 2735 3737 ne
rect 2735 3639 3089 3737
tri 3089 3639 3187 3737 sw
tri 3187 3639 3285 3737 ne
rect 3285 3639 3639 3737
tri 3639 3639 3737 3737 sw
tri 3737 3639 3835 3737 ne
rect 3835 3639 4189 3737
tri 4189 3639 4287 3737 sw
tri 4287 3639 4385 3737 ne
rect 4385 3639 4739 3737
tri 4739 3639 4837 3737 sw
tri 4837 3639 4935 3737 ne
rect 4935 3639 5289 3737
tri 5289 3639 5387 3737 sw
tri 5387 3639 5485 3737 ne
rect 5485 3639 5839 3737
tri 5839 3639 5937 3737 sw
tri 5937 3639 6035 3737 ne
rect 6035 3639 6389 3737
tri 6389 3639 6487 3737 sw
tri 6487 3639 6585 3737 ne
rect 6585 3639 6939 3737
tri 6939 3639 7037 3737 sw
tri 7037 3639 7135 3737 ne
rect 7135 3639 7489 3737
tri 7489 3639 7587 3737 sw
tri 7587 3639 7685 3737 ne
rect 7685 3639 8039 3737
tri 8039 3639 8137 3737 sw
tri 8137 3639 8235 3737 ne
rect 8235 3639 8589 3737
tri 8589 3639 8687 3737 sw
tri 8687 3639 8785 3737 ne
rect 8785 3639 9139 3737
tri 9139 3639 9237 3737 sw
tri 9237 3639 9335 3737 ne
rect 9335 3639 9689 3737
tri 9689 3639 9787 3737 sw
tri 9787 3639 9885 3737 ne
rect 9885 3639 10239 3737
tri 10239 3639 10337 3737 sw
tri 10337 3639 10435 3737 ne
rect 10435 3639 10789 3737
tri 10789 3639 10887 3737 sw
tri 10887 3639 10985 3737 ne
rect 10985 3639 11339 3737
tri 11339 3639 11437 3737 sw
tri 11437 3639 11535 3737 ne
rect 11535 3639 11889 3737
tri 11889 3639 11987 3737 sw
tri 11987 3639 12085 3737 ne
rect 12085 3639 12439 3737
tri 12439 3639 12537 3737 sw
tri 12537 3639 12635 3737 ne
rect 12635 3639 12989 3737
tri 12989 3639 13087 3737 sw
tri 13087 3639 13185 3737 ne
rect 13185 3639 13539 3737
tri 13539 3639 13637 3737 sw
tri 13637 3639 13735 3737 ne
rect 13735 3639 14089 3737
tri 14089 3639 14187 3737 sw
tri 14187 3639 14285 3737 ne
rect 14285 3639 14639 3737
tri 14639 3639 14737 3737 sw
tri 14737 3639 14835 3737 ne
rect 14835 3639 15189 3737
tri 15189 3639 15287 3737 sw
tri 15287 3639 15385 3737 ne
rect 15385 3639 15739 3737
tri 15739 3639 15837 3737 sw
tri 15837 3639 15935 3737 ne
rect 15935 3639 16289 3737
tri 16289 3639 16387 3737 sw
tri 16387 3639 16485 3737 ne
rect 16485 3639 16839 3737
tri 16839 3639 16937 3737 sw
tri 16937 3639 17035 3737 ne
rect 17035 3639 17389 3737
tri 17389 3639 17487 3737 sw
tri 17487 3639 17585 3737 ne
rect 17585 3639 17939 3737
tri 17939 3639 18037 3737 sw
tri 18037 3639 18135 3737 ne
rect 18135 3639 18489 3737
tri 18489 3639 18587 3737 sw
tri 18587 3639 18685 3737 ne
rect 18685 3639 19039 3737
tri 19039 3639 19137 3737 sw
tri 19137 3639 19235 3737 ne
rect 19235 3639 19589 3737
tri 19589 3639 19687 3737 sw
rect -500 3635 437 3639
rect -500 3515 215 3635
rect 335 3541 437 3635
tri 437 3541 535 3639 sw
tri 535 3541 633 3639 ne
rect 633 3635 987 3639
rect 633 3541 765 3635
rect 335 3515 535 3541
rect -500 3511 535 3515
tri 535 3511 565 3541 sw
tri 633 3511 663 3541 ne
rect 663 3515 765 3541
rect 885 3541 987 3635
tri 987 3541 1085 3639 sw
tri 1085 3541 1183 3639 ne
rect 1183 3635 1537 3639
rect 1183 3541 1315 3635
rect 885 3515 1085 3541
rect 663 3511 1085 3515
tri 1085 3511 1115 3541 sw
tri 1183 3511 1213 3541 ne
rect 1213 3515 1315 3541
rect 1435 3541 1537 3635
tri 1537 3541 1635 3639 sw
tri 1635 3541 1733 3639 ne
rect 1733 3635 2087 3639
rect 1733 3541 1865 3635
rect 1435 3515 1635 3541
rect 1213 3511 1635 3515
tri 1635 3511 1665 3541 sw
tri 1733 3511 1763 3541 ne
rect 1763 3515 1865 3541
rect 1985 3541 2087 3635
tri 2087 3541 2185 3639 sw
tri 2185 3541 2283 3639 ne
rect 2283 3635 2637 3639
rect 2283 3541 2415 3635
rect 1985 3515 2185 3541
rect 1763 3511 2185 3515
tri 2185 3511 2215 3541 sw
tri 2283 3511 2313 3541 ne
rect 2313 3515 2415 3541
rect 2535 3541 2637 3635
tri 2637 3541 2735 3639 sw
tri 2735 3541 2833 3639 ne
rect 2833 3635 3187 3639
rect 2833 3541 2965 3635
rect 2535 3515 2735 3541
rect 2313 3511 2735 3515
tri 2735 3511 2765 3541 sw
tri 2833 3511 2863 3541 ne
rect 2863 3515 2965 3541
rect 3085 3541 3187 3635
tri 3187 3541 3285 3639 sw
tri 3285 3541 3383 3639 ne
rect 3383 3635 3737 3639
rect 3383 3541 3515 3635
rect 3085 3515 3285 3541
rect 2863 3511 3285 3515
tri 3285 3511 3315 3541 sw
tri 3383 3511 3413 3541 ne
rect 3413 3515 3515 3541
rect 3635 3541 3737 3635
tri 3737 3541 3835 3639 sw
tri 3835 3541 3933 3639 ne
rect 3933 3635 4287 3639
rect 3933 3541 4065 3635
rect 3635 3515 3835 3541
rect 3413 3511 3835 3515
tri 3835 3511 3865 3541 sw
tri 3933 3511 3963 3541 ne
rect 3963 3515 4065 3541
rect 4185 3541 4287 3635
tri 4287 3541 4385 3639 sw
tri 4385 3541 4483 3639 ne
rect 4483 3635 4837 3639
rect 4483 3541 4615 3635
rect 4185 3515 4385 3541
rect 3963 3511 4385 3515
tri 4385 3511 4415 3541 sw
tri 4483 3511 4513 3541 ne
rect 4513 3515 4615 3541
rect 4735 3541 4837 3635
tri 4837 3541 4935 3639 sw
tri 4935 3541 5033 3639 ne
rect 5033 3635 5387 3639
rect 5033 3541 5165 3635
rect 4735 3515 4935 3541
rect 4513 3511 4935 3515
tri 4935 3511 4965 3541 sw
tri 5033 3511 5063 3541 ne
rect 5063 3515 5165 3541
rect 5285 3541 5387 3635
tri 5387 3541 5485 3639 sw
tri 5485 3541 5583 3639 ne
rect 5583 3635 5937 3639
rect 5583 3541 5715 3635
rect 5285 3515 5485 3541
rect 5063 3511 5485 3515
tri 5485 3511 5515 3541 sw
tri 5583 3511 5613 3541 ne
rect 5613 3515 5715 3541
rect 5835 3541 5937 3635
tri 5937 3541 6035 3639 sw
tri 6035 3541 6133 3639 ne
rect 6133 3635 6487 3639
rect 6133 3541 6265 3635
rect 5835 3515 6035 3541
rect 5613 3511 6035 3515
tri 6035 3511 6065 3541 sw
tri 6133 3511 6163 3541 ne
rect 6163 3515 6265 3541
rect 6385 3541 6487 3635
tri 6487 3541 6585 3639 sw
tri 6585 3541 6683 3639 ne
rect 6683 3635 7037 3639
rect 6683 3541 6815 3635
rect 6385 3515 6585 3541
rect 6163 3511 6585 3515
tri 6585 3511 6615 3541 sw
tri 6683 3511 6713 3541 ne
rect 6713 3515 6815 3541
rect 6935 3541 7037 3635
tri 7037 3541 7135 3639 sw
tri 7135 3541 7233 3639 ne
rect 7233 3635 7587 3639
rect 7233 3541 7365 3635
rect 6935 3515 7135 3541
rect 6713 3511 7135 3515
tri 7135 3511 7165 3541 sw
tri 7233 3511 7263 3541 ne
rect 7263 3515 7365 3541
rect 7485 3541 7587 3635
tri 7587 3541 7685 3639 sw
tri 7685 3541 7783 3639 ne
rect 7783 3635 8137 3639
rect 7783 3541 7915 3635
rect 7485 3515 7685 3541
rect 7263 3511 7685 3515
tri 7685 3511 7715 3541 sw
tri 7783 3511 7813 3541 ne
rect 7813 3515 7915 3541
rect 8035 3541 8137 3635
tri 8137 3541 8235 3639 sw
tri 8235 3541 8333 3639 ne
rect 8333 3635 8687 3639
rect 8333 3541 8465 3635
rect 8035 3515 8235 3541
rect 7813 3511 8235 3515
tri 8235 3511 8265 3541 sw
tri 8333 3511 8363 3541 ne
rect 8363 3515 8465 3541
rect 8585 3541 8687 3635
tri 8687 3541 8785 3639 sw
tri 8785 3541 8883 3639 ne
rect 8883 3635 9237 3639
rect 8883 3541 9015 3635
rect 8585 3515 8785 3541
rect 8363 3511 8785 3515
tri 8785 3511 8815 3541 sw
tri 8883 3511 8913 3541 ne
rect 8913 3515 9015 3541
rect 9135 3541 9237 3635
tri 9237 3541 9335 3639 sw
tri 9335 3541 9433 3639 ne
rect 9433 3635 9787 3639
rect 9433 3541 9565 3635
rect 9135 3515 9335 3541
rect 8913 3511 9335 3515
tri 9335 3511 9365 3541 sw
tri 9433 3511 9463 3541 ne
rect 9463 3515 9565 3541
rect 9685 3541 9787 3635
tri 9787 3541 9885 3639 sw
tri 9885 3541 9983 3639 ne
rect 9983 3635 10337 3639
rect 9983 3541 10115 3635
rect 9685 3515 9885 3541
rect 9463 3511 9885 3515
tri 9885 3511 9915 3541 sw
tri 9983 3511 10013 3541 ne
rect 10013 3515 10115 3541
rect 10235 3541 10337 3635
tri 10337 3541 10435 3639 sw
tri 10435 3541 10533 3639 ne
rect 10533 3635 10887 3639
rect 10533 3541 10665 3635
rect 10235 3515 10435 3541
rect 10013 3511 10435 3515
tri 10435 3511 10465 3541 sw
tri 10533 3511 10563 3541 ne
rect 10563 3515 10665 3541
rect 10785 3541 10887 3635
tri 10887 3541 10985 3639 sw
tri 10985 3541 11083 3639 ne
rect 11083 3635 11437 3639
rect 11083 3541 11215 3635
rect 10785 3515 10985 3541
rect 10563 3511 10985 3515
tri 10985 3511 11015 3541 sw
tri 11083 3511 11113 3541 ne
rect 11113 3515 11215 3541
rect 11335 3541 11437 3635
tri 11437 3541 11535 3639 sw
tri 11535 3541 11633 3639 ne
rect 11633 3635 11987 3639
rect 11633 3541 11765 3635
rect 11335 3515 11535 3541
rect 11113 3511 11535 3515
tri 11535 3511 11565 3541 sw
tri 11633 3511 11663 3541 ne
rect 11663 3515 11765 3541
rect 11885 3541 11987 3635
tri 11987 3541 12085 3639 sw
tri 12085 3541 12183 3639 ne
rect 12183 3635 12537 3639
rect 12183 3541 12315 3635
rect 11885 3515 12085 3541
rect 11663 3511 12085 3515
tri 12085 3511 12115 3541 sw
tri 12183 3511 12213 3541 ne
rect 12213 3515 12315 3541
rect 12435 3541 12537 3635
tri 12537 3541 12635 3639 sw
tri 12635 3541 12733 3639 ne
rect 12733 3635 13087 3639
rect 12733 3541 12865 3635
rect 12435 3515 12635 3541
rect 12213 3511 12635 3515
tri 12635 3511 12665 3541 sw
tri 12733 3511 12763 3541 ne
rect 12763 3515 12865 3541
rect 12985 3541 13087 3635
tri 13087 3541 13185 3639 sw
tri 13185 3541 13283 3639 ne
rect 13283 3635 13637 3639
rect 13283 3541 13415 3635
rect 12985 3515 13185 3541
rect 12763 3511 13185 3515
tri 13185 3511 13215 3541 sw
tri 13283 3511 13313 3541 ne
rect 13313 3515 13415 3541
rect 13535 3541 13637 3635
tri 13637 3541 13735 3639 sw
tri 13735 3541 13833 3639 ne
rect 13833 3635 14187 3639
rect 13833 3541 13965 3635
rect 13535 3515 13735 3541
rect 13313 3511 13735 3515
tri 13735 3511 13765 3541 sw
tri 13833 3511 13863 3541 ne
rect 13863 3515 13965 3541
rect 14085 3541 14187 3635
tri 14187 3541 14285 3639 sw
tri 14285 3541 14383 3639 ne
rect 14383 3635 14737 3639
rect 14383 3541 14515 3635
rect 14085 3515 14285 3541
rect 13863 3511 14285 3515
tri 14285 3511 14315 3541 sw
tri 14383 3511 14413 3541 ne
rect 14413 3515 14515 3541
rect 14635 3541 14737 3635
tri 14737 3541 14835 3639 sw
tri 14835 3541 14933 3639 ne
rect 14933 3635 15287 3639
rect 14933 3541 15065 3635
rect 14635 3515 14835 3541
rect 14413 3511 14835 3515
tri 14835 3511 14865 3541 sw
tri 14933 3511 14963 3541 ne
rect 14963 3515 15065 3541
rect 15185 3541 15287 3635
tri 15287 3541 15385 3639 sw
tri 15385 3541 15483 3639 ne
rect 15483 3635 15837 3639
rect 15483 3541 15615 3635
rect 15185 3515 15385 3541
rect 14963 3511 15385 3515
tri 15385 3511 15415 3541 sw
tri 15483 3511 15513 3541 ne
rect 15513 3515 15615 3541
rect 15735 3541 15837 3635
tri 15837 3541 15935 3639 sw
tri 15935 3541 16033 3639 ne
rect 16033 3635 16387 3639
rect 16033 3541 16165 3635
rect 15735 3515 15935 3541
rect 15513 3511 15935 3515
tri 15935 3511 15965 3541 sw
tri 16033 3511 16063 3541 ne
rect 16063 3515 16165 3541
rect 16285 3541 16387 3635
tri 16387 3541 16485 3639 sw
tri 16485 3541 16583 3639 ne
rect 16583 3635 16937 3639
rect 16583 3541 16715 3635
rect 16285 3515 16485 3541
rect 16063 3511 16485 3515
tri 16485 3511 16515 3541 sw
tri 16583 3511 16613 3541 ne
rect 16613 3515 16715 3541
rect 16835 3541 16937 3635
tri 16937 3541 17035 3639 sw
tri 17035 3541 17133 3639 ne
rect 17133 3635 17487 3639
rect 17133 3541 17265 3635
rect 16835 3515 17035 3541
rect 16613 3511 17035 3515
tri 17035 3511 17065 3541 sw
tri 17133 3511 17163 3541 ne
rect 17163 3515 17265 3541
rect 17385 3541 17487 3635
tri 17487 3541 17585 3639 sw
tri 17585 3541 17683 3639 ne
rect 17683 3635 18037 3639
rect 17683 3541 17815 3635
rect 17385 3515 17585 3541
rect 17163 3511 17585 3515
tri 17585 3511 17615 3541 sw
tri 17683 3511 17713 3541 ne
rect 17713 3515 17815 3541
rect 17935 3541 18037 3635
tri 18037 3541 18135 3639 sw
tri 18135 3541 18233 3639 ne
rect 18233 3635 18587 3639
rect 18233 3541 18365 3635
rect 17935 3515 18135 3541
rect 17713 3511 18135 3515
tri 18135 3511 18165 3541 sw
tri 18233 3511 18263 3541 ne
rect 18263 3515 18365 3541
rect 18485 3541 18587 3635
tri 18587 3541 18685 3639 sw
tri 18685 3541 18783 3639 ne
rect 18783 3635 19137 3639
rect 18783 3541 18915 3635
rect 18485 3515 18685 3541
rect 18263 3511 18685 3515
tri 18685 3511 18715 3541 sw
tri 18783 3511 18813 3541 ne
rect 18813 3515 18915 3541
rect 19035 3541 19137 3635
tri 19137 3541 19235 3639 sw
tri 19235 3541 19333 3639 ne
rect 19333 3635 20300 3639
rect 19333 3541 19465 3635
rect 19035 3515 19235 3541
rect 18813 3511 19235 3515
tri 19235 3511 19265 3541 sw
tri 19333 3511 19363 3541 ne
rect 19363 3515 19465 3541
rect 19585 3515 20300 3635
rect 19363 3511 20300 3515
tri 113 3413 211 3511 ne
rect 211 3413 565 3511
tri 565 3413 663 3511 sw
tri 663 3413 761 3511 ne
rect 761 3413 1115 3511
tri 1115 3413 1213 3511 sw
tri 1213 3413 1311 3511 ne
rect 1311 3413 1665 3511
tri 1665 3413 1763 3511 sw
tri 1763 3413 1861 3511 ne
rect 1861 3413 2215 3511
tri 2215 3413 2313 3511 sw
tri 2313 3413 2411 3511 ne
rect 2411 3413 2765 3511
tri 2765 3413 2863 3511 sw
tri 2863 3413 2961 3511 ne
rect 2961 3413 3315 3511
tri 3315 3413 3413 3511 sw
tri 3413 3413 3511 3511 ne
rect 3511 3413 3865 3511
tri 3865 3413 3963 3511 sw
tri 3963 3413 4061 3511 ne
rect 4061 3413 4415 3511
tri 4415 3413 4513 3511 sw
tri 4513 3413 4611 3511 ne
rect 4611 3413 4965 3511
tri 4965 3413 5063 3511 sw
tri 5063 3413 5161 3511 ne
rect 5161 3413 5515 3511
tri 5515 3413 5613 3511 sw
tri 5613 3413 5711 3511 ne
rect 5711 3413 6065 3511
tri 6065 3413 6163 3511 sw
tri 6163 3413 6261 3511 ne
rect 6261 3413 6615 3511
tri 6615 3413 6713 3511 sw
tri 6713 3413 6811 3511 ne
rect 6811 3413 7165 3511
tri 7165 3413 7263 3511 sw
tri 7263 3413 7361 3511 ne
rect 7361 3413 7715 3511
tri 7715 3413 7813 3511 sw
tri 7813 3413 7911 3511 ne
rect 7911 3413 8265 3511
tri 8265 3413 8363 3511 sw
tri 8363 3413 8461 3511 ne
rect 8461 3413 8815 3511
tri 8815 3413 8913 3511 sw
tri 8913 3413 9011 3511 ne
rect 9011 3413 9365 3511
tri 9365 3413 9463 3511 sw
tri 9463 3413 9561 3511 ne
rect 9561 3413 9915 3511
tri 9915 3413 10013 3511 sw
tri 10013 3413 10111 3511 ne
rect 10111 3413 10465 3511
tri 10465 3413 10563 3511 sw
tri 10563 3413 10661 3511 ne
rect 10661 3413 11015 3511
tri 11015 3413 11113 3511 sw
tri 11113 3413 11211 3511 ne
rect 11211 3413 11565 3511
tri 11565 3413 11663 3511 sw
tri 11663 3413 11761 3511 ne
rect 11761 3413 12115 3511
tri 12115 3413 12213 3511 sw
tri 12213 3413 12311 3511 ne
rect 12311 3413 12665 3511
tri 12665 3413 12763 3511 sw
tri 12763 3413 12861 3511 ne
rect 12861 3413 13215 3511
tri 13215 3413 13313 3511 sw
tri 13313 3413 13411 3511 ne
rect 13411 3413 13765 3511
tri 13765 3413 13863 3511 sw
tri 13863 3413 13961 3511 ne
rect 13961 3413 14315 3511
tri 14315 3413 14413 3511 sw
tri 14413 3413 14511 3511 ne
rect 14511 3413 14865 3511
tri 14865 3413 14963 3511 sw
tri 14963 3413 15061 3511 ne
rect 15061 3413 15415 3511
tri 15415 3413 15513 3511 sw
tri 15513 3413 15611 3511 ne
rect 15611 3413 15965 3511
tri 15965 3413 16063 3511 sw
tri 16063 3413 16161 3511 ne
rect 16161 3413 16515 3511
tri 16515 3413 16613 3511 sw
tri 16613 3413 16711 3511 ne
rect 16711 3413 17065 3511
tri 17065 3413 17163 3511 sw
tri 17163 3413 17261 3511 ne
rect 17261 3413 17615 3511
tri 17615 3413 17713 3511 sw
tri 17713 3413 17811 3511 ne
rect 17811 3413 18165 3511
tri 18165 3413 18263 3511 sw
tri 18263 3413 18361 3511 ne
rect 18361 3413 18715 3511
tri 18715 3413 18813 3511 sw
tri 18813 3413 18911 3511 ne
rect 18911 3413 19265 3511
tri 19265 3413 19363 3511 sw
tri 19363 3413 19461 3511 ne
rect 19461 3413 20300 3511
rect -2000 3383 113 3413
tri 113 3383 143 3413 sw
tri 211 3383 241 3413 ne
rect 241 3383 663 3413
tri 663 3383 693 3413 sw
tri 761 3383 791 3413 ne
rect 791 3383 1213 3413
tri 1213 3383 1243 3413 sw
tri 1311 3383 1341 3413 ne
rect 1341 3383 1763 3413
tri 1763 3383 1793 3413 sw
tri 1861 3383 1891 3413 ne
rect 1891 3383 2313 3413
tri 2313 3383 2343 3413 sw
tri 2411 3383 2441 3413 ne
rect 2441 3383 2863 3413
tri 2863 3383 2893 3413 sw
tri 2961 3383 2991 3413 ne
rect 2991 3383 3413 3413
tri 3413 3383 3443 3413 sw
tri 3511 3383 3541 3413 ne
rect 3541 3383 3963 3413
tri 3963 3383 3993 3413 sw
tri 4061 3383 4091 3413 ne
rect 4091 3383 4513 3413
tri 4513 3383 4543 3413 sw
tri 4611 3383 4641 3413 ne
rect 4641 3383 5063 3413
tri 5063 3383 5093 3413 sw
tri 5161 3383 5191 3413 ne
rect 5191 3383 5613 3413
tri 5613 3383 5643 3413 sw
tri 5711 3383 5741 3413 ne
rect 5741 3383 6163 3413
tri 6163 3383 6193 3413 sw
tri 6261 3383 6291 3413 ne
rect 6291 3383 6713 3413
tri 6713 3383 6743 3413 sw
tri 6811 3383 6841 3413 ne
rect 6841 3383 7263 3413
tri 7263 3383 7293 3413 sw
tri 7361 3383 7391 3413 ne
rect 7391 3383 7813 3413
tri 7813 3383 7843 3413 sw
tri 7911 3383 7941 3413 ne
rect 7941 3383 8363 3413
tri 8363 3383 8393 3413 sw
tri 8461 3383 8491 3413 ne
rect 8491 3383 8913 3413
tri 8913 3383 8943 3413 sw
tri 9011 3383 9041 3413 ne
rect 9041 3383 9463 3413
tri 9463 3383 9493 3413 sw
tri 9561 3383 9591 3413 ne
rect 9591 3383 10013 3413
tri 10013 3383 10043 3413 sw
tri 10111 3383 10141 3413 ne
rect 10141 3383 10563 3413
tri 10563 3383 10593 3413 sw
tri 10661 3383 10691 3413 ne
rect 10691 3383 11113 3413
tri 11113 3383 11143 3413 sw
tri 11211 3383 11241 3413 ne
rect 11241 3383 11663 3413
tri 11663 3383 11693 3413 sw
tri 11761 3383 11791 3413 ne
rect 11791 3383 12213 3413
tri 12213 3383 12243 3413 sw
tri 12311 3383 12341 3413 ne
rect 12341 3383 12763 3413
tri 12763 3383 12793 3413 sw
tri 12861 3383 12891 3413 ne
rect 12891 3383 13313 3413
tri 13313 3383 13343 3413 sw
tri 13411 3383 13441 3413 ne
rect 13441 3383 13863 3413
tri 13863 3383 13893 3413 sw
tri 13961 3383 13991 3413 ne
rect 13991 3383 14413 3413
tri 14413 3383 14443 3413 sw
tri 14511 3383 14541 3413 ne
rect 14541 3383 14963 3413
tri 14963 3383 14993 3413 sw
tri 15061 3383 15091 3413 ne
rect 15091 3383 15513 3413
tri 15513 3383 15543 3413 sw
tri 15611 3383 15641 3413 ne
rect 15641 3383 16063 3413
tri 16063 3383 16093 3413 sw
tri 16161 3383 16191 3413 ne
rect 16191 3383 16613 3413
tri 16613 3383 16643 3413 sw
tri 16711 3383 16741 3413 ne
rect 16741 3383 17163 3413
tri 17163 3383 17193 3413 sw
tri 17261 3383 17291 3413 ne
rect 17291 3383 17713 3413
tri 17713 3383 17743 3413 sw
tri 17811 3383 17841 3413 ne
rect 17841 3383 18263 3413
tri 18263 3383 18293 3413 sw
tri 18361 3383 18391 3413 ne
rect 18391 3383 18813 3413
tri 18813 3383 18843 3413 sw
tri 18911 3383 18941 3413 ne
rect 18941 3383 19363 3413
tri 19363 3383 19393 3413 sw
tri 19461 3383 19491 3413 ne
rect 19491 3383 20300 3413
rect -2000 3285 143 3383
tri 143 3285 241 3383 sw
tri 241 3285 339 3383 ne
rect 339 3285 693 3383
tri 693 3285 791 3383 sw
tri 791 3285 889 3383 ne
rect 889 3285 1243 3383
tri 1243 3285 1341 3383 sw
tri 1341 3285 1439 3383 ne
rect 1439 3285 1793 3383
tri 1793 3285 1891 3383 sw
tri 1891 3285 1989 3383 ne
rect 1989 3285 2343 3383
tri 2343 3285 2441 3383 sw
tri 2441 3285 2539 3383 ne
rect 2539 3285 2893 3383
tri 2893 3285 2991 3383 sw
tri 2991 3285 3089 3383 ne
rect 3089 3285 3443 3383
tri 3443 3285 3541 3383 sw
tri 3541 3285 3639 3383 ne
rect 3639 3285 3993 3383
tri 3993 3285 4091 3383 sw
tri 4091 3285 4189 3383 ne
rect 4189 3285 4543 3383
tri 4543 3285 4641 3383 sw
tri 4641 3285 4739 3383 ne
rect 4739 3285 5093 3383
tri 5093 3285 5191 3383 sw
tri 5191 3285 5289 3383 ne
rect 5289 3285 5643 3383
tri 5643 3285 5741 3383 sw
tri 5741 3285 5839 3383 ne
rect 5839 3285 6193 3383
tri 6193 3285 6291 3383 sw
tri 6291 3285 6389 3383 ne
rect 6389 3285 6743 3383
tri 6743 3285 6841 3383 sw
tri 6841 3285 6939 3383 ne
rect 6939 3285 7293 3383
tri 7293 3285 7391 3383 sw
tri 7391 3285 7489 3383 ne
rect 7489 3285 7843 3383
tri 7843 3285 7941 3383 sw
tri 7941 3285 8039 3383 ne
rect 8039 3285 8393 3383
tri 8393 3285 8491 3383 sw
tri 8491 3285 8589 3383 ne
rect 8589 3285 8943 3383
tri 8943 3285 9041 3383 sw
tri 9041 3285 9139 3383 ne
rect 9139 3285 9493 3383
tri 9493 3285 9591 3383 sw
tri 9591 3285 9689 3383 ne
rect 9689 3285 10043 3383
tri 10043 3285 10141 3383 sw
tri 10141 3285 10239 3383 ne
rect 10239 3285 10593 3383
tri 10593 3285 10691 3383 sw
tri 10691 3285 10789 3383 ne
rect 10789 3285 11143 3383
tri 11143 3285 11241 3383 sw
tri 11241 3285 11339 3383 ne
rect 11339 3285 11693 3383
tri 11693 3285 11791 3383 sw
tri 11791 3285 11889 3383 ne
rect 11889 3285 12243 3383
tri 12243 3285 12341 3383 sw
tri 12341 3285 12439 3383 ne
rect 12439 3285 12793 3383
tri 12793 3285 12891 3383 sw
tri 12891 3285 12989 3383 ne
rect 12989 3285 13343 3383
tri 13343 3285 13441 3383 sw
tri 13441 3285 13539 3383 ne
rect 13539 3285 13893 3383
tri 13893 3285 13991 3383 sw
tri 13991 3285 14089 3383 ne
rect 14089 3285 14443 3383
tri 14443 3285 14541 3383 sw
tri 14541 3285 14639 3383 ne
rect 14639 3285 14993 3383
tri 14993 3285 15091 3383 sw
tri 15091 3285 15189 3383 ne
rect 15189 3285 15543 3383
tri 15543 3285 15641 3383 sw
tri 15641 3285 15739 3383 ne
rect 15739 3285 16093 3383
tri 16093 3285 16191 3383 sw
tri 16191 3285 16289 3383 ne
rect 16289 3285 16643 3383
tri 16643 3285 16741 3383 sw
tri 16741 3285 16839 3383 ne
rect 16839 3285 17193 3383
tri 17193 3285 17291 3383 sw
tri 17291 3285 17389 3383 ne
rect 17389 3285 17743 3383
tri 17743 3285 17841 3383 sw
tri 17841 3285 17939 3383 ne
rect 17939 3285 18293 3383
tri 18293 3285 18391 3383 sw
tri 18391 3285 18489 3383 ne
rect 18489 3285 18843 3383
tri 18843 3285 18941 3383 sw
tri 18941 3285 19039 3383 ne
rect 19039 3285 19393 3383
tri 19393 3285 19491 3383 sw
tri 19491 3285 19589 3383 ne
rect 19589 3285 20300 3383
rect -2000 3187 241 3285
tri 241 3187 339 3285 sw
tri 339 3187 437 3285 ne
rect 437 3187 791 3285
tri 791 3187 889 3285 sw
tri 889 3187 987 3285 ne
rect 987 3187 1341 3285
tri 1341 3187 1439 3285 sw
tri 1439 3187 1537 3285 ne
rect 1537 3187 1891 3285
tri 1891 3187 1989 3285 sw
tri 1989 3187 2087 3285 ne
rect 2087 3187 2441 3285
tri 2441 3187 2539 3285 sw
tri 2539 3187 2637 3285 ne
rect 2637 3187 2991 3285
tri 2991 3187 3089 3285 sw
tri 3089 3187 3187 3285 ne
rect 3187 3187 3541 3285
tri 3541 3187 3639 3285 sw
tri 3639 3187 3737 3285 ne
rect 3737 3187 4091 3285
tri 4091 3187 4189 3285 sw
tri 4189 3187 4287 3285 ne
rect 4287 3187 4641 3285
tri 4641 3187 4739 3285 sw
tri 4739 3187 4837 3285 ne
rect 4837 3187 5191 3285
tri 5191 3187 5289 3285 sw
tri 5289 3187 5387 3285 ne
rect 5387 3187 5741 3285
tri 5741 3187 5839 3285 sw
tri 5839 3187 5937 3285 ne
rect 5937 3187 6291 3285
tri 6291 3187 6389 3285 sw
tri 6389 3187 6487 3285 ne
rect 6487 3187 6841 3285
tri 6841 3187 6939 3285 sw
tri 6939 3187 7037 3285 ne
rect 7037 3187 7391 3285
tri 7391 3187 7489 3285 sw
tri 7489 3187 7587 3285 ne
rect 7587 3187 7941 3285
tri 7941 3187 8039 3285 sw
tri 8039 3187 8137 3285 ne
rect 8137 3187 8491 3285
tri 8491 3187 8589 3285 sw
tri 8589 3187 8687 3285 ne
rect 8687 3187 9041 3285
tri 9041 3187 9139 3285 sw
tri 9139 3187 9237 3285 ne
rect 9237 3187 9591 3285
tri 9591 3187 9689 3285 sw
tri 9689 3187 9787 3285 ne
rect 9787 3187 10141 3285
tri 10141 3187 10239 3285 sw
tri 10239 3187 10337 3285 ne
rect 10337 3187 10691 3285
tri 10691 3187 10789 3285 sw
tri 10789 3187 10887 3285 ne
rect 10887 3187 11241 3285
tri 11241 3187 11339 3285 sw
tri 11339 3187 11437 3285 ne
rect 11437 3187 11791 3285
tri 11791 3187 11889 3285 sw
tri 11889 3187 11987 3285 ne
rect 11987 3187 12341 3285
tri 12341 3187 12439 3285 sw
tri 12439 3187 12537 3285 ne
rect 12537 3187 12891 3285
tri 12891 3187 12989 3285 sw
tri 12989 3187 13087 3285 ne
rect 13087 3187 13441 3285
tri 13441 3187 13539 3285 sw
tri 13539 3187 13637 3285 ne
rect 13637 3187 13991 3285
tri 13991 3187 14089 3285 sw
tri 14089 3187 14187 3285 ne
rect 14187 3187 14541 3285
tri 14541 3187 14639 3285 sw
tri 14639 3187 14737 3285 ne
rect 14737 3187 15091 3285
tri 15091 3187 15189 3285 sw
tri 15189 3187 15287 3285 ne
rect 15287 3187 15641 3285
tri 15641 3187 15739 3285 sw
tri 15739 3187 15837 3285 ne
rect 15837 3187 16191 3285
tri 16191 3187 16289 3285 sw
tri 16289 3187 16387 3285 ne
rect 16387 3187 16741 3285
tri 16741 3187 16839 3285 sw
tri 16839 3187 16937 3285 ne
rect 16937 3187 17291 3285
tri 17291 3187 17389 3285 sw
tri 17389 3187 17487 3285 ne
rect 17487 3187 17841 3285
tri 17841 3187 17939 3285 sw
tri 17939 3187 18037 3285 ne
rect 18037 3187 18391 3285
tri 18391 3187 18489 3285 sw
tri 18489 3187 18587 3285 ne
rect 18587 3187 18941 3285
tri 18941 3187 19039 3285 sw
tri 19039 3187 19137 3285 ne
rect 19137 3187 19491 3285
tri 19491 3187 19589 3285 sw
tri 19589 3187 19687 3285 ne
rect 19687 3187 20300 3285
rect -2000 3089 339 3187
tri 339 3089 437 3187 sw
tri 437 3089 535 3187 ne
rect 535 3089 889 3187
tri 889 3089 987 3187 sw
tri 987 3089 1085 3187 ne
rect 1085 3089 1439 3187
tri 1439 3089 1537 3187 sw
tri 1537 3089 1635 3187 ne
rect 1635 3089 1989 3187
tri 1989 3089 2087 3187 sw
tri 2087 3089 2185 3187 ne
rect 2185 3089 2539 3187
tri 2539 3089 2637 3187 sw
tri 2637 3089 2735 3187 ne
rect 2735 3089 3089 3187
tri 3089 3089 3187 3187 sw
tri 3187 3089 3285 3187 ne
rect 3285 3089 3639 3187
tri 3639 3089 3737 3187 sw
tri 3737 3089 3835 3187 ne
rect 3835 3089 4189 3187
tri 4189 3089 4287 3187 sw
tri 4287 3089 4385 3187 ne
rect 4385 3089 4739 3187
tri 4739 3089 4837 3187 sw
tri 4837 3089 4935 3187 ne
rect 4935 3089 5289 3187
tri 5289 3089 5387 3187 sw
tri 5387 3089 5485 3187 ne
rect 5485 3089 5839 3187
tri 5839 3089 5937 3187 sw
tri 5937 3089 6035 3187 ne
rect 6035 3089 6389 3187
tri 6389 3089 6487 3187 sw
tri 6487 3089 6585 3187 ne
rect 6585 3089 6939 3187
tri 6939 3089 7037 3187 sw
tri 7037 3089 7135 3187 ne
rect 7135 3089 7489 3187
tri 7489 3089 7587 3187 sw
tri 7587 3089 7685 3187 ne
rect 7685 3089 8039 3187
tri 8039 3089 8137 3187 sw
tri 8137 3089 8235 3187 ne
rect 8235 3089 8589 3187
tri 8589 3089 8687 3187 sw
tri 8687 3089 8785 3187 ne
rect 8785 3089 9139 3187
tri 9139 3089 9237 3187 sw
tri 9237 3089 9335 3187 ne
rect 9335 3089 9689 3187
tri 9689 3089 9787 3187 sw
tri 9787 3089 9885 3187 ne
rect 9885 3089 10239 3187
tri 10239 3089 10337 3187 sw
tri 10337 3089 10435 3187 ne
rect 10435 3089 10789 3187
tri 10789 3089 10887 3187 sw
tri 10887 3089 10985 3187 ne
rect 10985 3089 11339 3187
tri 11339 3089 11437 3187 sw
tri 11437 3089 11535 3187 ne
rect 11535 3089 11889 3187
tri 11889 3089 11987 3187 sw
tri 11987 3089 12085 3187 ne
rect 12085 3089 12439 3187
tri 12439 3089 12537 3187 sw
tri 12537 3089 12635 3187 ne
rect 12635 3089 12989 3187
tri 12989 3089 13087 3187 sw
tri 13087 3089 13185 3187 ne
rect 13185 3089 13539 3187
tri 13539 3089 13637 3187 sw
tri 13637 3089 13735 3187 ne
rect 13735 3089 14089 3187
tri 14089 3089 14187 3187 sw
tri 14187 3089 14285 3187 ne
rect 14285 3089 14639 3187
tri 14639 3089 14737 3187 sw
tri 14737 3089 14835 3187 ne
rect 14835 3089 15189 3187
tri 15189 3089 15287 3187 sw
tri 15287 3089 15385 3187 ne
rect 15385 3089 15739 3187
tri 15739 3089 15837 3187 sw
tri 15837 3089 15935 3187 ne
rect 15935 3089 16289 3187
tri 16289 3089 16387 3187 sw
tri 16387 3089 16485 3187 ne
rect 16485 3089 16839 3187
tri 16839 3089 16937 3187 sw
tri 16937 3089 17035 3187 ne
rect 17035 3089 17389 3187
tri 17389 3089 17487 3187 sw
tri 17487 3089 17585 3187 ne
rect 17585 3089 17939 3187
tri 17939 3089 18037 3187 sw
tri 18037 3089 18135 3187 ne
rect 18135 3089 18489 3187
tri 18489 3089 18587 3187 sw
tri 18587 3089 18685 3187 ne
rect 18685 3089 19039 3187
tri 19039 3089 19137 3187 sw
tri 19137 3089 19235 3187 ne
rect 19235 3089 19589 3187
tri 19589 3089 19687 3187 sw
rect 20800 3089 21800 3737
rect -2000 3085 437 3089
rect -2000 2965 215 3085
rect 335 2991 437 3085
tri 437 2991 535 3089 sw
tri 535 2991 633 3089 ne
rect 633 3085 987 3089
rect 633 2991 765 3085
rect 335 2965 535 2991
rect -2000 2961 535 2965
rect -2000 2313 -1000 2961
tri 113 2863 211 2961 ne
rect 211 2913 535 2961
tri 535 2913 613 2991 sw
tri 633 2913 711 2991 ne
rect 711 2965 765 2991
rect 885 2991 987 3085
tri 987 2991 1085 3089 sw
tri 1085 2991 1183 3089 ne
rect 1183 3085 1537 3089
rect 1183 2991 1315 3085
rect 885 2965 1085 2991
rect 711 2913 1085 2965
tri 1085 2913 1163 2991 sw
tri 1183 2913 1261 2991 ne
rect 1261 2965 1315 2991
rect 1435 2991 1537 3085
tri 1537 2991 1635 3089 sw
tri 1635 2991 1733 3089 ne
rect 1733 3085 2087 3089
rect 1733 2991 1865 3085
rect 1435 2965 1635 2991
rect 1261 2913 1635 2965
tri 1635 2913 1713 2991 sw
tri 1733 2913 1811 2991 ne
rect 1811 2965 1865 2991
rect 1985 2991 2087 3085
tri 2087 2991 2185 3089 sw
tri 2185 2991 2283 3089 ne
rect 2283 3085 2637 3089
rect 2283 2991 2415 3085
rect 1985 2965 2185 2991
rect 1811 2913 2185 2965
tri 2185 2913 2263 2991 sw
tri 2283 2913 2361 2991 ne
rect 2361 2965 2415 2991
rect 2535 2991 2637 3085
tri 2637 2991 2735 3089 sw
tri 2735 2991 2833 3089 ne
rect 2833 3085 3187 3089
rect 2833 2991 2965 3085
rect 2535 2965 2735 2991
rect 2361 2913 2735 2965
tri 2735 2913 2813 2991 sw
tri 2833 2913 2911 2991 ne
rect 2911 2965 2965 2991
rect 3085 2991 3187 3085
tri 3187 2991 3285 3089 sw
tri 3285 2991 3383 3089 ne
rect 3383 3085 3737 3089
rect 3383 2991 3515 3085
rect 3085 2965 3285 2991
rect 2911 2913 3285 2965
tri 3285 2913 3363 2991 sw
tri 3383 2913 3461 2991 ne
rect 3461 2965 3515 2991
rect 3635 2991 3737 3085
tri 3737 2991 3835 3089 sw
tri 3835 2991 3933 3089 ne
rect 3933 3085 4287 3089
rect 3933 2991 4065 3085
rect 3635 2965 3835 2991
rect 3461 2913 3835 2965
tri 3835 2913 3913 2991 sw
tri 3933 2913 4011 2991 ne
rect 4011 2965 4065 2991
rect 4185 2991 4287 3085
tri 4287 2991 4385 3089 sw
tri 4385 2991 4483 3089 ne
rect 4483 3085 4837 3089
rect 4483 2991 4615 3085
rect 4185 2965 4385 2991
rect 4011 2913 4385 2965
tri 4385 2913 4463 2991 sw
tri 4483 2913 4561 2991 ne
rect 4561 2965 4615 2991
rect 4735 2991 4837 3085
tri 4837 2991 4935 3089 sw
tri 4935 2991 5033 3089 ne
rect 5033 3085 5387 3089
rect 5033 2991 5165 3085
rect 4735 2965 4935 2991
rect 4561 2913 4935 2965
tri 4935 2913 5013 2991 sw
tri 5033 2913 5111 2991 ne
rect 5111 2965 5165 2991
rect 5285 2991 5387 3085
tri 5387 2991 5485 3089 sw
tri 5485 2991 5583 3089 ne
rect 5583 3085 5937 3089
rect 5583 2991 5715 3085
rect 5285 2965 5485 2991
rect 5111 2913 5485 2965
tri 5485 2913 5563 2991 sw
tri 5583 2913 5661 2991 ne
rect 5661 2965 5715 2991
rect 5835 2991 5937 3085
tri 5937 2991 6035 3089 sw
tri 6035 2991 6133 3089 ne
rect 6133 3085 6487 3089
rect 6133 2991 6265 3085
rect 5835 2965 6035 2991
rect 5661 2913 6035 2965
tri 6035 2913 6113 2991 sw
tri 6133 2913 6211 2991 ne
rect 6211 2965 6265 2991
rect 6385 2991 6487 3085
tri 6487 2991 6585 3089 sw
tri 6585 2991 6683 3089 ne
rect 6683 3085 7037 3089
rect 6683 2991 6815 3085
rect 6385 2965 6585 2991
rect 6211 2913 6585 2965
tri 6585 2913 6663 2991 sw
tri 6683 2913 6761 2991 ne
rect 6761 2965 6815 2991
rect 6935 2991 7037 3085
tri 7037 2991 7135 3089 sw
tri 7135 2991 7233 3089 ne
rect 7233 3085 7587 3089
rect 7233 2991 7365 3085
rect 6935 2965 7135 2991
rect 6761 2913 7135 2965
tri 7135 2913 7213 2991 sw
tri 7233 2913 7311 2991 ne
rect 7311 2965 7365 2991
rect 7485 2991 7587 3085
tri 7587 2991 7685 3089 sw
tri 7685 2991 7783 3089 ne
rect 7783 3085 8137 3089
rect 7783 2991 7915 3085
rect 7485 2965 7685 2991
rect 7311 2913 7685 2965
tri 7685 2913 7763 2991 sw
tri 7783 2913 7861 2991 ne
rect 7861 2965 7915 2991
rect 8035 2991 8137 3085
tri 8137 2991 8235 3089 sw
tri 8235 2991 8333 3089 ne
rect 8333 3085 8687 3089
rect 8333 2991 8465 3085
rect 8035 2965 8235 2991
rect 7861 2913 8235 2965
tri 8235 2913 8313 2991 sw
tri 8333 2913 8411 2991 ne
rect 8411 2965 8465 2991
rect 8585 2991 8687 3085
tri 8687 2991 8785 3089 sw
tri 8785 2991 8883 3089 ne
rect 8883 3085 9237 3089
rect 8883 2991 9015 3085
rect 8585 2965 8785 2991
rect 8411 2913 8785 2965
tri 8785 2913 8863 2991 sw
tri 8883 2913 8961 2991 ne
rect 8961 2965 9015 2991
rect 9135 2991 9237 3085
tri 9237 2991 9335 3089 sw
tri 9335 2991 9433 3089 ne
rect 9433 3085 9787 3089
rect 9433 2991 9565 3085
rect 9135 2965 9335 2991
rect 8961 2913 9335 2965
tri 9335 2913 9413 2991 sw
tri 9433 2913 9511 2991 ne
rect 9511 2965 9565 2991
rect 9685 2991 9787 3085
tri 9787 2991 9885 3089 sw
tri 9885 2991 9983 3089 ne
rect 9983 3085 10337 3089
rect 9983 2991 10115 3085
rect 9685 2965 9885 2991
rect 9511 2913 9885 2965
tri 9885 2913 9963 2991 sw
tri 9983 2913 10061 2991 ne
rect 10061 2965 10115 2991
rect 10235 2991 10337 3085
tri 10337 2991 10435 3089 sw
tri 10435 2991 10533 3089 ne
rect 10533 3085 10887 3089
rect 10533 2991 10665 3085
rect 10235 2965 10435 2991
rect 10061 2913 10435 2965
tri 10435 2913 10513 2991 sw
tri 10533 2913 10611 2991 ne
rect 10611 2965 10665 2991
rect 10785 2991 10887 3085
tri 10887 2991 10985 3089 sw
tri 10985 2991 11083 3089 ne
rect 11083 3085 11437 3089
rect 11083 2991 11215 3085
rect 10785 2965 10985 2991
rect 10611 2913 10985 2965
tri 10985 2913 11063 2991 sw
tri 11083 2913 11161 2991 ne
rect 11161 2965 11215 2991
rect 11335 2991 11437 3085
tri 11437 2991 11535 3089 sw
tri 11535 2991 11633 3089 ne
rect 11633 3085 11987 3089
rect 11633 2991 11765 3085
rect 11335 2965 11535 2991
rect 11161 2913 11535 2965
tri 11535 2913 11613 2991 sw
tri 11633 2913 11711 2991 ne
rect 11711 2965 11765 2991
rect 11885 2991 11987 3085
tri 11987 2991 12085 3089 sw
tri 12085 2991 12183 3089 ne
rect 12183 3085 12537 3089
rect 12183 2991 12315 3085
rect 11885 2965 12085 2991
rect 11711 2913 12085 2965
tri 12085 2913 12163 2991 sw
tri 12183 2913 12261 2991 ne
rect 12261 2965 12315 2991
rect 12435 2991 12537 3085
tri 12537 2991 12635 3089 sw
tri 12635 2991 12733 3089 ne
rect 12733 3085 13087 3089
rect 12733 2991 12865 3085
rect 12435 2965 12635 2991
rect 12261 2913 12635 2965
tri 12635 2913 12713 2991 sw
tri 12733 2913 12811 2991 ne
rect 12811 2965 12865 2991
rect 12985 2991 13087 3085
tri 13087 2991 13185 3089 sw
tri 13185 2991 13283 3089 ne
rect 13283 3085 13637 3089
rect 13283 2991 13415 3085
rect 12985 2965 13185 2991
rect 12811 2913 13185 2965
tri 13185 2913 13263 2991 sw
tri 13283 2913 13361 2991 ne
rect 13361 2965 13415 2991
rect 13535 2991 13637 3085
tri 13637 2991 13735 3089 sw
tri 13735 2991 13833 3089 ne
rect 13833 3085 14187 3089
rect 13833 2991 13965 3085
rect 13535 2965 13735 2991
rect 13361 2913 13735 2965
tri 13735 2913 13813 2991 sw
tri 13833 2913 13911 2991 ne
rect 13911 2965 13965 2991
rect 14085 2991 14187 3085
tri 14187 2991 14285 3089 sw
tri 14285 2991 14383 3089 ne
rect 14383 3085 14737 3089
rect 14383 2991 14515 3085
rect 14085 2965 14285 2991
rect 13911 2913 14285 2965
tri 14285 2913 14363 2991 sw
tri 14383 2913 14461 2991 ne
rect 14461 2965 14515 2991
rect 14635 2991 14737 3085
tri 14737 2991 14835 3089 sw
tri 14835 2991 14933 3089 ne
rect 14933 3085 15287 3089
rect 14933 2991 15065 3085
rect 14635 2965 14835 2991
rect 14461 2913 14835 2965
tri 14835 2913 14913 2991 sw
tri 14933 2913 15011 2991 ne
rect 15011 2965 15065 2991
rect 15185 2991 15287 3085
tri 15287 2991 15385 3089 sw
tri 15385 2991 15483 3089 ne
rect 15483 3085 15837 3089
rect 15483 2991 15615 3085
rect 15185 2965 15385 2991
rect 15011 2913 15385 2965
tri 15385 2913 15463 2991 sw
tri 15483 2913 15561 2991 ne
rect 15561 2965 15615 2991
rect 15735 2991 15837 3085
tri 15837 2991 15935 3089 sw
tri 15935 2991 16033 3089 ne
rect 16033 3085 16387 3089
rect 16033 2991 16165 3085
rect 15735 2965 15935 2991
rect 15561 2913 15935 2965
tri 15935 2913 16013 2991 sw
tri 16033 2913 16111 2991 ne
rect 16111 2965 16165 2991
rect 16285 2991 16387 3085
tri 16387 2991 16485 3089 sw
tri 16485 2991 16583 3089 ne
rect 16583 3085 16937 3089
rect 16583 2991 16715 3085
rect 16285 2965 16485 2991
rect 16111 2913 16485 2965
tri 16485 2913 16563 2991 sw
tri 16583 2913 16661 2991 ne
rect 16661 2965 16715 2991
rect 16835 2991 16937 3085
tri 16937 2991 17035 3089 sw
tri 17035 2991 17133 3089 ne
rect 17133 3085 17487 3089
rect 17133 2991 17265 3085
rect 16835 2965 17035 2991
rect 16661 2913 17035 2965
tri 17035 2913 17113 2991 sw
tri 17133 2913 17211 2991 ne
rect 17211 2965 17265 2991
rect 17385 2991 17487 3085
tri 17487 2991 17585 3089 sw
tri 17585 2991 17683 3089 ne
rect 17683 3085 18037 3089
rect 17683 2991 17815 3085
rect 17385 2965 17585 2991
rect 17211 2913 17585 2965
tri 17585 2913 17663 2991 sw
tri 17683 2913 17761 2991 ne
rect 17761 2965 17815 2991
rect 17935 2991 18037 3085
tri 18037 2991 18135 3089 sw
tri 18135 2991 18233 3089 ne
rect 18233 3085 18587 3089
rect 18233 2991 18365 3085
rect 17935 2965 18135 2991
rect 17761 2913 18135 2965
tri 18135 2913 18213 2991 sw
tri 18233 2913 18311 2991 ne
rect 18311 2965 18365 2991
rect 18485 2991 18587 3085
tri 18587 2991 18685 3089 sw
tri 18685 2991 18783 3089 ne
rect 18783 3085 19137 3089
rect 18783 2991 18915 3085
rect 18485 2965 18685 2991
rect 18311 2913 18685 2965
tri 18685 2913 18763 2991 sw
tri 18783 2913 18861 2991 ne
rect 18861 2965 18915 2991
rect 19035 2991 19137 3085
tri 19137 2991 19235 3089 sw
tri 19235 2991 19333 3089 ne
rect 19333 3085 21800 3089
rect 19333 2991 19465 3085
rect 19035 2965 19235 2991
rect 18861 2913 19235 2965
tri 19235 2913 19313 2991 sw
tri 19333 2913 19411 2991 ne
rect 19411 2965 19465 2991
rect 19585 2965 21800 3085
rect 19411 2913 21800 2965
rect 211 2863 613 2913
rect -500 2813 113 2863
tri 113 2813 163 2863 sw
tri 211 2813 261 2863 ne
rect 261 2833 613 2863
tri 613 2833 693 2913 sw
tri 711 2833 791 2913 ne
rect 791 2833 1163 2913
tri 1163 2833 1243 2913 sw
tri 1261 2833 1341 2913 ne
rect 1341 2833 1713 2913
tri 1713 2833 1793 2913 sw
tri 1811 2833 1891 2913 ne
rect 1891 2833 2263 2913
tri 2263 2833 2343 2913 sw
tri 2361 2833 2441 2913 ne
rect 2441 2833 2813 2913
tri 2813 2833 2893 2913 sw
tri 2911 2833 2991 2913 ne
rect 2991 2833 3363 2913
tri 3363 2833 3443 2913 sw
tri 3461 2833 3541 2913 ne
rect 3541 2833 3913 2913
tri 3913 2833 3993 2913 sw
tri 4011 2833 4091 2913 ne
rect 4091 2833 4463 2913
tri 4463 2833 4543 2913 sw
tri 4561 2833 4641 2913 ne
rect 4641 2833 5013 2913
tri 5013 2833 5093 2913 sw
tri 5111 2833 5191 2913 ne
rect 5191 2833 5563 2913
tri 5563 2833 5643 2913 sw
tri 5661 2833 5741 2913 ne
rect 5741 2833 6113 2913
tri 6113 2833 6193 2913 sw
tri 6211 2833 6291 2913 ne
rect 6291 2833 6663 2913
tri 6663 2833 6743 2913 sw
tri 6761 2833 6841 2913 ne
rect 6841 2833 7213 2913
tri 7213 2833 7293 2913 sw
tri 7311 2833 7391 2913 ne
rect 7391 2833 7763 2913
tri 7763 2833 7843 2913 sw
tri 7861 2833 7941 2913 ne
rect 7941 2833 8313 2913
tri 8313 2833 8393 2913 sw
tri 8411 2833 8491 2913 ne
rect 8491 2833 8863 2913
tri 8863 2833 8943 2913 sw
tri 8961 2833 9041 2913 ne
rect 9041 2833 9413 2913
tri 9413 2833 9493 2913 sw
tri 9511 2833 9591 2913 ne
rect 9591 2833 9963 2913
tri 9963 2833 10043 2913 sw
tri 10061 2833 10141 2913 ne
rect 10141 2833 10513 2913
tri 10513 2833 10593 2913 sw
tri 10611 2833 10691 2913 ne
rect 10691 2833 11063 2913
tri 11063 2833 11143 2913 sw
tri 11161 2833 11241 2913 ne
rect 11241 2833 11613 2913
tri 11613 2833 11693 2913 sw
tri 11711 2833 11791 2913 ne
rect 11791 2833 12163 2913
tri 12163 2833 12243 2913 sw
tri 12261 2833 12341 2913 ne
rect 12341 2833 12713 2913
tri 12713 2833 12793 2913 sw
tri 12811 2833 12891 2913 ne
rect 12891 2833 13263 2913
tri 13263 2833 13343 2913 sw
tri 13361 2833 13441 2913 ne
rect 13441 2833 13813 2913
tri 13813 2833 13893 2913 sw
tri 13911 2833 13991 2913 ne
rect 13991 2833 14363 2913
tri 14363 2833 14443 2913 sw
tri 14461 2833 14541 2913 ne
rect 14541 2833 14913 2913
tri 14913 2833 14993 2913 sw
tri 15011 2833 15091 2913 ne
rect 15091 2833 15463 2913
tri 15463 2833 15543 2913 sw
tri 15561 2833 15641 2913 ne
rect 15641 2833 16013 2913
tri 16013 2833 16093 2913 sw
tri 16111 2833 16191 2913 ne
rect 16191 2833 16563 2913
tri 16563 2833 16643 2913 sw
tri 16661 2833 16741 2913 ne
rect 16741 2833 17113 2913
tri 17113 2833 17193 2913 sw
tri 17211 2833 17291 2913 ne
rect 17291 2833 17663 2913
tri 17663 2833 17743 2913 sw
tri 17761 2833 17841 2913 ne
rect 17841 2833 18213 2913
tri 18213 2833 18293 2913 sw
tri 18311 2833 18391 2913 ne
rect 18391 2833 18763 2913
tri 18763 2833 18843 2913 sw
tri 18861 2833 18941 2913 ne
rect 18941 2833 19313 2913
tri 19313 2833 19393 2913 sw
tri 19411 2833 19491 2913 ne
rect 19491 2833 20100 2913
rect 261 2813 693 2833
rect -500 2735 163 2813
tri 163 2735 241 2813 sw
tri 261 2735 339 2813 ne
rect 339 2735 693 2813
tri 693 2735 791 2833 sw
tri 791 2735 889 2833 ne
rect 889 2735 1243 2833
tri 1243 2735 1341 2833 sw
tri 1341 2735 1439 2833 ne
rect 1439 2735 1793 2833
tri 1793 2735 1891 2833 sw
tri 1891 2735 1989 2833 ne
rect 1989 2735 2343 2833
tri 2343 2735 2441 2833 sw
tri 2441 2735 2539 2833 ne
rect 2539 2735 2893 2833
tri 2893 2735 2991 2833 sw
tri 2991 2735 3089 2833 ne
rect 3089 2735 3443 2833
tri 3443 2735 3541 2833 sw
tri 3541 2735 3639 2833 ne
rect 3639 2735 3993 2833
tri 3993 2735 4091 2833 sw
tri 4091 2735 4189 2833 ne
rect 4189 2735 4543 2833
tri 4543 2735 4641 2833 sw
tri 4641 2735 4739 2833 ne
rect 4739 2735 5093 2833
tri 5093 2735 5191 2833 sw
tri 5191 2735 5289 2833 ne
rect 5289 2735 5643 2833
tri 5643 2735 5741 2833 sw
tri 5741 2735 5839 2833 ne
rect 5839 2735 6193 2833
tri 6193 2735 6291 2833 sw
tri 6291 2735 6389 2833 ne
rect 6389 2735 6743 2833
tri 6743 2735 6841 2833 sw
tri 6841 2735 6939 2833 ne
rect 6939 2735 7293 2833
tri 7293 2735 7391 2833 sw
tri 7391 2735 7489 2833 ne
rect 7489 2735 7843 2833
tri 7843 2735 7941 2833 sw
tri 7941 2735 8039 2833 ne
rect 8039 2735 8393 2833
tri 8393 2735 8491 2833 sw
tri 8491 2735 8589 2833 ne
rect 8589 2735 8943 2833
tri 8943 2735 9041 2833 sw
tri 9041 2735 9139 2833 ne
rect 9139 2735 9493 2833
tri 9493 2735 9591 2833 sw
tri 9591 2735 9689 2833 ne
rect 9689 2735 10043 2833
tri 10043 2735 10141 2833 sw
tri 10141 2735 10239 2833 ne
rect 10239 2735 10593 2833
tri 10593 2735 10691 2833 sw
tri 10691 2735 10789 2833 ne
rect 10789 2735 11143 2833
tri 11143 2735 11241 2833 sw
tri 11241 2735 11339 2833 ne
rect 11339 2735 11693 2833
tri 11693 2735 11791 2833 sw
tri 11791 2735 11889 2833 ne
rect 11889 2735 12243 2833
tri 12243 2735 12341 2833 sw
tri 12341 2735 12439 2833 ne
rect 12439 2735 12793 2833
tri 12793 2735 12891 2833 sw
tri 12891 2735 12989 2833 ne
rect 12989 2735 13343 2833
tri 13343 2735 13441 2833 sw
tri 13441 2735 13539 2833 ne
rect 13539 2735 13893 2833
tri 13893 2735 13991 2833 sw
tri 13991 2735 14089 2833 ne
rect 14089 2735 14443 2833
tri 14443 2735 14541 2833 sw
tri 14541 2735 14639 2833 ne
rect 14639 2735 14993 2833
tri 14993 2735 15091 2833 sw
tri 15091 2735 15189 2833 ne
rect 15189 2735 15543 2833
tri 15543 2735 15641 2833 sw
tri 15641 2735 15739 2833 ne
rect 15739 2735 16093 2833
tri 16093 2735 16191 2833 sw
tri 16191 2735 16289 2833 ne
rect 16289 2735 16643 2833
tri 16643 2735 16741 2833 sw
tri 16741 2735 16839 2833 ne
rect 16839 2735 17193 2833
tri 17193 2735 17291 2833 sw
tri 17291 2735 17389 2833 ne
rect 17389 2735 17743 2833
tri 17743 2735 17841 2833 sw
tri 17841 2735 17939 2833 ne
rect 17939 2735 18293 2833
tri 18293 2735 18391 2833 sw
tri 18391 2735 18489 2833 ne
rect 18489 2735 18843 2833
tri 18843 2735 18941 2833 sw
tri 18941 2735 19039 2833 ne
rect 19039 2735 19393 2833
tri 19393 2735 19491 2833 sw
tri 19491 2735 19589 2833 ne
rect 19589 2813 20100 2833
rect 20200 2813 21800 2913
rect 19589 2735 21800 2813
rect -500 2687 241 2735
rect -500 2587 -400 2687
rect -300 2637 241 2687
tri 241 2637 339 2735 sw
tri 339 2637 437 2735 ne
rect 437 2637 791 2735
tri 791 2637 889 2735 sw
tri 889 2637 987 2735 ne
rect 987 2637 1341 2735
tri 1341 2637 1439 2735 sw
tri 1439 2637 1537 2735 ne
rect 1537 2637 1891 2735
tri 1891 2637 1989 2735 sw
tri 1989 2637 2087 2735 ne
rect 2087 2637 2441 2735
tri 2441 2637 2539 2735 sw
tri 2539 2637 2637 2735 ne
rect 2637 2637 2991 2735
tri 2991 2637 3089 2735 sw
tri 3089 2637 3187 2735 ne
rect 3187 2637 3541 2735
tri 3541 2637 3639 2735 sw
tri 3639 2637 3737 2735 ne
rect 3737 2637 4091 2735
tri 4091 2637 4189 2735 sw
tri 4189 2637 4287 2735 ne
rect 4287 2637 4641 2735
tri 4641 2637 4739 2735 sw
tri 4739 2637 4837 2735 ne
rect 4837 2637 5191 2735
tri 5191 2637 5289 2735 sw
tri 5289 2637 5387 2735 ne
rect 5387 2637 5741 2735
tri 5741 2637 5839 2735 sw
tri 5839 2637 5937 2735 ne
rect 5937 2637 6291 2735
tri 6291 2637 6389 2735 sw
tri 6389 2637 6487 2735 ne
rect 6487 2637 6841 2735
tri 6841 2637 6939 2735 sw
tri 6939 2637 7037 2735 ne
rect 7037 2637 7391 2735
tri 7391 2637 7489 2735 sw
tri 7489 2637 7587 2735 ne
rect 7587 2637 7941 2735
tri 7941 2637 8039 2735 sw
tri 8039 2637 8137 2735 ne
rect 8137 2637 8491 2735
tri 8491 2637 8589 2735 sw
tri 8589 2637 8687 2735 ne
rect 8687 2637 9041 2735
tri 9041 2637 9139 2735 sw
tri 9139 2637 9237 2735 ne
rect 9237 2637 9591 2735
tri 9591 2637 9689 2735 sw
tri 9689 2637 9787 2735 ne
rect 9787 2637 10141 2735
tri 10141 2637 10239 2735 sw
tri 10239 2637 10337 2735 ne
rect 10337 2637 10691 2735
tri 10691 2637 10789 2735 sw
tri 10789 2637 10887 2735 ne
rect 10887 2637 11241 2735
tri 11241 2637 11339 2735 sw
tri 11339 2637 11437 2735 ne
rect 11437 2637 11791 2735
tri 11791 2637 11889 2735 sw
tri 11889 2637 11987 2735 ne
rect 11987 2637 12341 2735
tri 12341 2637 12439 2735 sw
tri 12439 2637 12537 2735 ne
rect 12537 2637 12891 2735
tri 12891 2637 12989 2735 sw
tri 12989 2637 13087 2735 ne
rect 13087 2637 13441 2735
tri 13441 2637 13539 2735 sw
tri 13539 2637 13637 2735 ne
rect 13637 2637 13991 2735
tri 13991 2637 14089 2735 sw
tri 14089 2637 14187 2735 ne
rect 14187 2637 14541 2735
tri 14541 2637 14639 2735 sw
tri 14639 2637 14737 2735 ne
rect 14737 2637 15091 2735
tri 15091 2637 15189 2735 sw
tri 15189 2637 15287 2735 ne
rect 15287 2637 15641 2735
tri 15641 2637 15739 2735 sw
tri 15739 2637 15837 2735 ne
rect 15837 2637 16191 2735
tri 16191 2637 16289 2735 sw
tri 16289 2637 16387 2735 ne
rect 16387 2637 16741 2735
tri 16741 2637 16839 2735 sw
tri 16839 2637 16937 2735 ne
rect 16937 2637 17291 2735
tri 17291 2637 17389 2735 sw
tri 17389 2637 17487 2735 ne
rect 17487 2637 17841 2735
tri 17841 2637 17939 2735 sw
tri 17939 2637 18037 2735 ne
rect 18037 2637 18391 2735
tri 18391 2637 18489 2735 sw
tri 18489 2637 18587 2735 ne
rect 18587 2637 18941 2735
tri 18941 2637 19039 2735 sw
tri 19039 2637 19137 2735 ne
rect 19137 2637 19491 2735
tri 19491 2637 19589 2735 sw
tri 19589 2637 19687 2735 ne
rect 19687 2637 21800 2735
rect -300 2587 339 2637
rect -500 2539 339 2587
tri 339 2539 437 2637 sw
tri 437 2539 535 2637 ne
rect 535 2539 889 2637
tri 889 2539 987 2637 sw
tri 987 2539 1085 2637 ne
rect 1085 2539 1439 2637
tri 1439 2539 1537 2637 sw
tri 1537 2539 1635 2637 ne
rect 1635 2539 1989 2637
tri 1989 2539 2087 2637 sw
tri 2087 2539 2185 2637 ne
rect 2185 2539 2539 2637
tri 2539 2539 2637 2637 sw
tri 2637 2539 2735 2637 ne
rect 2735 2539 3089 2637
tri 3089 2539 3187 2637 sw
tri 3187 2539 3285 2637 ne
rect 3285 2539 3639 2637
tri 3639 2539 3737 2637 sw
tri 3737 2539 3835 2637 ne
rect 3835 2539 4189 2637
tri 4189 2539 4287 2637 sw
tri 4287 2539 4385 2637 ne
rect 4385 2539 4739 2637
tri 4739 2539 4837 2637 sw
tri 4837 2539 4935 2637 ne
rect 4935 2539 5289 2637
tri 5289 2539 5387 2637 sw
tri 5387 2539 5485 2637 ne
rect 5485 2539 5839 2637
tri 5839 2539 5937 2637 sw
tri 5937 2539 6035 2637 ne
rect 6035 2539 6389 2637
tri 6389 2539 6487 2637 sw
tri 6487 2539 6585 2637 ne
rect 6585 2539 6939 2637
tri 6939 2539 7037 2637 sw
tri 7037 2539 7135 2637 ne
rect 7135 2539 7489 2637
tri 7489 2539 7587 2637 sw
tri 7587 2539 7685 2637 ne
rect 7685 2539 8039 2637
tri 8039 2539 8137 2637 sw
tri 8137 2539 8235 2637 ne
rect 8235 2539 8589 2637
tri 8589 2539 8687 2637 sw
tri 8687 2539 8785 2637 ne
rect 8785 2539 9139 2637
tri 9139 2539 9237 2637 sw
tri 9237 2539 9335 2637 ne
rect 9335 2539 9689 2637
tri 9689 2539 9787 2637 sw
tri 9787 2539 9885 2637 ne
rect 9885 2539 10239 2637
tri 10239 2539 10337 2637 sw
tri 10337 2539 10435 2637 ne
rect 10435 2539 10789 2637
tri 10789 2539 10887 2637 sw
tri 10887 2539 10985 2637 ne
rect 10985 2539 11339 2637
tri 11339 2539 11437 2637 sw
tri 11437 2539 11535 2637 ne
rect 11535 2539 11889 2637
tri 11889 2539 11987 2637 sw
tri 11987 2539 12085 2637 ne
rect 12085 2539 12439 2637
tri 12439 2539 12537 2637 sw
tri 12537 2539 12635 2637 ne
rect 12635 2539 12989 2637
tri 12989 2539 13087 2637 sw
tri 13087 2539 13185 2637 ne
rect 13185 2539 13539 2637
tri 13539 2539 13637 2637 sw
tri 13637 2539 13735 2637 ne
rect 13735 2539 14089 2637
tri 14089 2539 14187 2637 sw
tri 14187 2539 14285 2637 ne
rect 14285 2539 14639 2637
tri 14639 2539 14737 2637 sw
tri 14737 2539 14835 2637 ne
rect 14835 2539 15189 2637
tri 15189 2539 15287 2637 sw
tri 15287 2539 15385 2637 ne
rect 15385 2539 15739 2637
tri 15739 2539 15837 2637 sw
tri 15837 2539 15935 2637 ne
rect 15935 2539 16289 2637
tri 16289 2539 16387 2637 sw
tri 16387 2539 16485 2637 ne
rect 16485 2539 16839 2637
tri 16839 2539 16937 2637 sw
tri 16937 2539 17035 2637 ne
rect 17035 2539 17389 2637
tri 17389 2539 17487 2637 sw
tri 17487 2539 17585 2637 ne
rect 17585 2539 17939 2637
tri 17939 2539 18037 2637 sw
tri 18037 2539 18135 2637 ne
rect 18135 2539 18489 2637
tri 18489 2539 18587 2637 sw
tri 18587 2539 18685 2637 ne
rect 18685 2539 19039 2637
tri 19039 2539 19137 2637 sw
tri 19137 2539 19235 2637 ne
rect 19235 2539 19589 2637
tri 19589 2539 19687 2637 sw
rect -500 2535 437 2539
rect -500 2415 215 2535
rect 335 2441 437 2535
tri 437 2441 535 2539 sw
tri 535 2441 633 2539 ne
rect 633 2535 987 2539
rect 633 2441 765 2535
rect 335 2415 535 2441
rect -500 2411 535 2415
tri 535 2411 565 2441 sw
tri 633 2411 663 2441 ne
rect 663 2415 765 2441
rect 885 2441 987 2535
tri 987 2441 1085 2539 sw
tri 1085 2441 1183 2539 ne
rect 1183 2535 1537 2539
rect 1183 2441 1315 2535
rect 885 2415 1085 2441
rect 663 2411 1085 2415
tri 1085 2411 1115 2441 sw
tri 1183 2411 1213 2441 ne
rect 1213 2415 1315 2441
rect 1435 2441 1537 2535
tri 1537 2441 1635 2539 sw
tri 1635 2441 1733 2539 ne
rect 1733 2535 2087 2539
rect 1733 2441 1865 2535
rect 1435 2415 1635 2441
rect 1213 2411 1635 2415
tri 1635 2411 1665 2441 sw
tri 1733 2411 1763 2441 ne
rect 1763 2415 1865 2441
rect 1985 2441 2087 2535
tri 2087 2441 2185 2539 sw
tri 2185 2441 2283 2539 ne
rect 2283 2535 2637 2539
rect 2283 2441 2415 2535
rect 1985 2415 2185 2441
rect 1763 2411 2185 2415
tri 2185 2411 2215 2441 sw
tri 2283 2411 2313 2441 ne
rect 2313 2415 2415 2441
rect 2535 2441 2637 2535
tri 2637 2441 2735 2539 sw
tri 2735 2441 2833 2539 ne
rect 2833 2535 3187 2539
rect 2833 2441 2965 2535
rect 2535 2415 2735 2441
rect 2313 2411 2735 2415
tri 2735 2411 2765 2441 sw
tri 2833 2411 2863 2441 ne
rect 2863 2415 2965 2441
rect 3085 2441 3187 2535
tri 3187 2441 3285 2539 sw
tri 3285 2441 3383 2539 ne
rect 3383 2535 3737 2539
rect 3383 2441 3515 2535
rect 3085 2415 3285 2441
rect 2863 2411 3285 2415
tri 3285 2411 3315 2441 sw
tri 3383 2411 3413 2441 ne
rect 3413 2415 3515 2441
rect 3635 2441 3737 2535
tri 3737 2441 3835 2539 sw
tri 3835 2441 3933 2539 ne
rect 3933 2535 4287 2539
rect 3933 2441 4065 2535
rect 3635 2415 3835 2441
rect 3413 2411 3835 2415
tri 3835 2411 3865 2441 sw
tri 3933 2411 3963 2441 ne
rect 3963 2415 4065 2441
rect 4185 2441 4287 2535
tri 4287 2441 4385 2539 sw
tri 4385 2441 4483 2539 ne
rect 4483 2535 4837 2539
rect 4483 2441 4615 2535
rect 4185 2415 4385 2441
rect 3963 2411 4385 2415
tri 4385 2411 4415 2441 sw
tri 4483 2411 4513 2441 ne
rect 4513 2415 4615 2441
rect 4735 2441 4837 2535
tri 4837 2441 4935 2539 sw
tri 4935 2441 5033 2539 ne
rect 5033 2535 5387 2539
rect 5033 2441 5165 2535
rect 4735 2415 4935 2441
rect 4513 2411 4935 2415
tri 4935 2411 4965 2441 sw
tri 5033 2411 5063 2441 ne
rect 5063 2415 5165 2441
rect 5285 2441 5387 2535
tri 5387 2441 5485 2539 sw
tri 5485 2441 5583 2539 ne
rect 5583 2535 5937 2539
rect 5583 2441 5715 2535
rect 5285 2415 5485 2441
rect 5063 2411 5485 2415
tri 5485 2411 5515 2441 sw
tri 5583 2411 5613 2441 ne
rect 5613 2415 5715 2441
rect 5835 2441 5937 2535
tri 5937 2441 6035 2539 sw
tri 6035 2441 6133 2539 ne
rect 6133 2535 6487 2539
rect 6133 2441 6265 2535
rect 5835 2415 6035 2441
rect 5613 2411 6035 2415
tri 6035 2411 6065 2441 sw
tri 6133 2411 6163 2441 ne
rect 6163 2415 6265 2441
rect 6385 2441 6487 2535
tri 6487 2441 6585 2539 sw
tri 6585 2441 6683 2539 ne
rect 6683 2535 7037 2539
rect 6683 2441 6815 2535
rect 6385 2415 6585 2441
rect 6163 2411 6585 2415
tri 6585 2411 6615 2441 sw
tri 6683 2411 6713 2441 ne
rect 6713 2415 6815 2441
rect 6935 2441 7037 2535
tri 7037 2441 7135 2539 sw
tri 7135 2441 7233 2539 ne
rect 7233 2535 7587 2539
rect 7233 2441 7365 2535
rect 6935 2415 7135 2441
rect 6713 2411 7135 2415
tri 7135 2411 7165 2441 sw
tri 7233 2411 7263 2441 ne
rect 7263 2415 7365 2441
rect 7485 2441 7587 2535
tri 7587 2441 7685 2539 sw
tri 7685 2441 7783 2539 ne
rect 7783 2535 8137 2539
rect 7783 2441 7915 2535
rect 7485 2415 7685 2441
rect 7263 2411 7685 2415
tri 7685 2411 7715 2441 sw
tri 7783 2411 7813 2441 ne
rect 7813 2415 7915 2441
rect 8035 2441 8137 2535
tri 8137 2441 8235 2539 sw
tri 8235 2441 8333 2539 ne
rect 8333 2535 8687 2539
rect 8333 2441 8465 2535
rect 8035 2415 8235 2441
rect 7813 2411 8235 2415
tri 8235 2411 8265 2441 sw
tri 8333 2411 8363 2441 ne
rect 8363 2415 8465 2441
rect 8585 2441 8687 2535
tri 8687 2441 8785 2539 sw
tri 8785 2441 8883 2539 ne
rect 8883 2535 9237 2539
rect 8883 2441 9015 2535
rect 8585 2415 8785 2441
rect 8363 2411 8785 2415
tri 8785 2411 8815 2441 sw
tri 8883 2411 8913 2441 ne
rect 8913 2415 9015 2441
rect 9135 2441 9237 2535
tri 9237 2441 9335 2539 sw
tri 9335 2441 9433 2539 ne
rect 9433 2535 9787 2539
rect 9433 2441 9565 2535
rect 9135 2415 9335 2441
rect 8913 2411 9335 2415
tri 9335 2411 9365 2441 sw
tri 9433 2411 9463 2441 ne
rect 9463 2415 9565 2441
rect 9685 2441 9787 2535
tri 9787 2441 9885 2539 sw
tri 9885 2441 9983 2539 ne
rect 9983 2535 10337 2539
rect 9983 2441 10115 2535
rect 9685 2415 9885 2441
rect 9463 2411 9885 2415
tri 9885 2411 9915 2441 sw
tri 9983 2411 10013 2441 ne
rect 10013 2415 10115 2441
rect 10235 2441 10337 2535
tri 10337 2441 10435 2539 sw
tri 10435 2441 10533 2539 ne
rect 10533 2535 10887 2539
rect 10533 2441 10665 2535
rect 10235 2415 10435 2441
rect 10013 2411 10435 2415
tri 10435 2411 10465 2441 sw
tri 10533 2411 10563 2441 ne
rect 10563 2415 10665 2441
rect 10785 2441 10887 2535
tri 10887 2441 10985 2539 sw
tri 10985 2441 11083 2539 ne
rect 11083 2535 11437 2539
rect 11083 2441 11215 2535
rect 10785 2415 10985 2441
rect 10563 2411 10985 2415
tri 10985 2411 11015 2441 sw
tri 11083 2411 11113 2441 ne
rect 11113 2415 11215 2441
rect 11335 2441 11437 2535
tri 11437 2441 11535 2539 sw
tri 11535 2441 11633 2539 ne
rect 11633 2535 11987 2539
rect 11633 2441 11765 2535
rect 11335 2415 11535 2441
rect 11113 2411 11535 2415
tri 11535 2411 11565 2441 sw
tri 11633 2411 11663 2441 ne
rect 11663 2415 11765 2441
rect 11885 2441 11987 2535
tri 11987 2441 12085 2539 sw
tri 12085 2441 12183 2539 ne
rect 12183 2535 12537 2539
rect 12183 2441 12315 2535
rect 11885 2415 12085 2441
rect 11663 2411 12085 2415
tri 12085 2411 12115 2441 sw
tri 12183 2411 12213 2441 ne
rect 12213 2415 12315 2441
rect 12435 2441 12537 2535
tri 12537 2441 12635 2539 sw
tri 12635 2441 12733 2539 ne
rect 12733 2535 13087 2539
rect 12733 2441 12865 2535
rect 12435 2415 12635 2441
rect 12213 2411 12635 2415
tri 12635 2411 12665 2441 sw
tri 12733 2411 12763 2441 ne
rect 12763 2415 12865 2441
rect 12985 2441 13087 2535
tri 13087 2441 13185 2539 sw
tri 13185 2441 13283 2539 ne
rect 13283 2535 13637 2539
rect 13283 2441 13415 2535
rect 12985 2415 13185 2441
rect 12763 2411 13185 2415
tri 13185 2411 13215 2441 sw
tri 13283 2411 13313 2441 ne
rect 13313 2415 13415 2441
rect 13535 2441 13637 2535
tri 13637 2441 13735 2539 sw
tri 13735 2441 13833 2539 ne
rect 13833 2535 14187 2539
rect 13833 2441 13965 2535
rect 13535 2415 13735 2441
rect 13313 2411 13735 2415
tri 13735 2411 13765 2441 sw
tri 13833 2411 13863 2441 ne
rect 13863 2415 13965 2441
rect 14085 2441 14187 2535
tri 14187 2441 14285 2539 sw
tri 14285 2441 14383 2539 ne
rect 14383 2535 14737 2539
rect 14383 2441 14515 2535
rect 14085 2415 14285 2441
rect 13863 2411 14285 2415
tri 14285 2411 14315 2441 sw
tri 14383 2411 14413 2441 ne
rect 14413 2415 14515 2441
rect 14635 2441 14737 2535
tri 14737 2441 14835 2539 sw
tri 14835 2441 14933 2539 ne
rect 14933 2535 15287 2539
rect 14933 2441 15065 2535
rect 14635 2415 14835 2441
rect 14413 2411 14835 2415
tri 14835 2411 14865 2441 sw
tri 14933 2411 14963 2441 ne
rect 14963 2415 15065 2441
rect 15185 2441 15287 2535
tri 15287 2441 15385 2539 sw
tri 15385 2441 15483 2539 ne
rect 15483 2535 15837 2539
rect 15483 2441 15615 2535
rect 15185 2415 15385 2441
rect 14963 2411 15385 2415
tri 15385 2411 15415 2441 sw
tri 15483 2411 15513 2441 ne
rect 15513 2415 15615 2441
rect 15735 2441 15837 2535
tri 15837 2441 15935 2539 sw
tri 15935 2441 16033 2539 ne
rect 16033 2535 16387 2539
rect 16033 2441 16165 2535
rect 15735 2415 15935 2441
rect 15513 2411 15935 2415
tri 15935 2411 15965 2441 sw
tri 16033 2411 16063 2441 ne
rect 16063 2415 16165 2441
rect 16285 2441 16387 2535
tri 16387 2441 16485 2539 sw
tri 16485 2441 16583 2539 ne
rect 16583 2535 16937 2539
rect 16583 2441 16715 2535
rect 16285 2415 16485 2441
rect 16063 2411 16485 2415
tri 16485 2411 16515 2441 sw
tri 16583 2411 16613 2441 ne
rect 16613 2415 16715 2441
rect 16835 2441 16937 2535
tri 16937 2441 17035 2539 sw
tri 17035 2441 17133 2539 ne
rect 17133 2535 17487 2539
rect 17133 2441 17265 2535
rect 16835 2415 17035 2441
rect 16613 2411 17035 2415
tri 17035 2411 17065 2441 sw
tri 17133 2411 17163 2441 ne
rect 17163 2415 17265 2441
rect 17385 2441 17487 2535
tri 17487 2441 17585 2539 sw
tri 17585 2441 17683 2539 ne
rect 17683 2535 18037 2539
rect 17683 2441 17815 2535
rect 17385 2415 17585 2441
rect 17163 2411 17585 2415
tri 17585 2411 17615 2441 sw
tri 17683 2411 17713 2441 ne
rect 17713 2415 17815 2441
rect 17935 2441 18037 2535
tri 18037 2441 18135 2539 sw
tri 18135 2441 18233 2539 ne
rect 18233 2535 18587 2539
rect 18233 2441 18365 2535
rect 17935 2415 18135 2441
rect 17713 2411 18135 2415
tri 18135 2411 18165 2441 sw
tri 18233 2411 18263 2441 ne
rect 18263 2415 18365 2441
rect 18485 2441 18587 2535
tri 18587 2441 18685 2539 sw
tri 18685 2441 18783 2539 ne
rect 18783 2535 19137 2539
rect 18783 2441 18915 2535
rect 18485 2415 18685 2441
rect 18263 2411 18685 2415
tri 18685 2411 18715 2441 sw
tri 18783 2411 18813 2441 ne
rect 18813 2415 18915 2441
rect 19035 2441 19137 2535
tri 19137 2441 19235 2539 sw
tri 19235 2441 19333 2539 ne
rect 19333 2535 20300 2539
rect 19333 2441 19465 2535
rect 19035 2415 19235 2441
rect 18813 2411 19235 2415
tri 19235 2411 19265 2441 sw
tri 19333 2411 19363 2441 ne
rect 19363 2415 19465 2441
rect 19585 2415 20300 2535
rect 19363 2411 20300 2415
tri 113 2313 211 2411 ne
rect 211 2313 565 2411
tri 565 2313 663 2411 sw
tri 663 2313 761 2411 ne
rect 761 2313 1115 2411
tri 1115 2313 1213 2411 sw
tri 1213 2313 1311 2411 ne
rect 1311 2313 1665 2411
tri 1665 2313 1763 2411 sw
tri 1763 2313 1861 2411 ne
rect 1861 2313 2215 2411
tri 2215 2313 2313 2411 sw
tri 2313 2313 2411 2411 ne
rect 2411 2313 2765 2411
tri 2765 2313 2863 2411 sw
tri 2863 2313 2961 2411 ne
rect 2961 2313 3315 2411
tri 3315 2313 3413 2411 sw
tri 3413 2313 3511 2411 ne
rect 3511 2313 3865 2411
tri 3865 2313 3963 2411 sw
tri 3963 2313 4061 2411 ne
rect 4061 2313 4415 2411
tri 4415 2313 4513 2411 sw
tri 4513 2313 4611 2411 ne
rect 4611 2313 4965 2411
tri 4965 2313 5063 2411 sw
tri 5063 2313 5161 2411 ne
rect 5161 2313 5515 2411
tri 5515 2313 5613 2411 sw
tri 5613 2313 5711 2411 ne
rect 5711 2313 6065 2411
tri 6065 2313 6163 2411 sw
tri 6163 2313 6261 2411 ne
rect 6261 2313 6615 2411
tri 6615 2313 6713 2411 sw
tri 6713 2313 6811 2411 ne
rect 6811 2313 7165 2411
tri 7165 2313 7263 2411 sw
tri 7263 2313 7361 2411 ne
rect 7361 2313 7715 2411
tri 7715 2313 7813 2411 sw
tri 7813 2313 7911 2411 ne
rect 7911 2313 8265 2411
tri 8265 2313 8363 2411 sw
tri 8363 2313 8461 2411 ne
rect 8461 2313 8815 2411
tri 8815 2313 8913 2411 sw
tri 8913 2313 9011 2411 ne
rect 9011 2313 9365 2411
tri 9365 2313 9463 2411 sw
tri 9463 2313 9561 2411 ne
rect 9561 2313 9915 2411
tri 9915 2313 10013 2411 sw
tri 10013 2313 10111 2411 ne
rect 10111 2313 10465 2411
tri 10465 2313 10563 2411 sw
tri 10563 2313 10661 2411 ne
rect 10661 2313 11015 2411
tri 11015 2313 11113 2411 sw
tri 11113 2313 11211 2411 ne
rect 11211 2313 11565 2411
tri 11565 2313 11663 2411 sw
tri 11663 2313 11761 2411 ne
rect 11761 2313 12115 2411
tri 12115 2313 12213 2411 sw
tri 12213 2313 12311 2411 ne
rect 12311 2313 12665 2411
tri 12665 2313 12763 2411 sw
tri 12763 2313 12861 2411 ne
rect 12861 2313 13215 2411
tri 13215 2313 13313 2411 sw
tri 13313 2313 13411 2411 ne
rect 13411 2313 13765 2411
tri 13765 2313 13863 2411 sw
tri 13863 2313 13961 2411 ne
rect 13961 2313 14315 2411
tri 14315 2313 14413 2411 sw
tri 14413 2313 14511 2411 ne
rect 14511 2313 14865 2411
tri 14865 2313 14963 2411 sw
tri 14963 2313 15061 2411 ne
rect 15061 2313 15415 2411
tri 15415 2313 15513 2411 sw
tri 15513 2313 15611 2411 ne
rect 15611 2313 15965 2411
tri 15965 2313 16063 2411 sw
tri 16063 2313 16161 2411 ne
rect 16161 2313 16515 2411
tri 16515 2313 16613 2411 sw
tri 16613 2313 16711 2411 ne
rect 16711 2313 17065 2411
tri 17065 2313 17163 2411 sw
tri 17163 2313 17261 2411 ne
rect 17261 2313 17615 2411
tri 17615 2313 17713 2411 sw
tri 17713 2313 17811 2411 ne
rect 17811 2313 18165 2411
tri 18165 2313 18263 2411 sw
tri 18263 2313 18361 2411 ne
rect 18361 2313 18715 2411
tri 18715 2313 18813 2411 sw
tri 18813 2313 18911 2411 ne
rect 18911 2313 19265 2411
tri 19265 2313 19363 2411 sw
tri 19363 2313 19461 2411 ne
rect 19461 2313 20300 2411
rect -2000 2283 113 2313
tri 113 2283 143 2313 sw
tri 211 2283 241 2313 ne
rect 241 2283 663 2313
tri 663 2283 693 2313 sw
tri 761 2283 791 2313 ne
rect 791 2283 1213 2313
tri 1213 2283 1243 2313 sw
tri 1311 2283 1341 2313 ne
rect 1341 2283 1763 2313
tri 1763 2283 1793 2313 sw
tri 1861 2283 1891 2313 ne
rect 1891 2283 2313 2313
tri 2313 2283 2343 2313 sw
tri 2411 2283 2441 2313 ne
rect 2441 2283 2863 2313
tri 2863 2283 2893 2313 sw
tri 2961 2283 2991 2313 ne
rect 2991 2283 3413 2313
tri 3413 2283 3443 2313 sw
tri 3511 2283 3541 2313 ne
rect 3541 2283 3963 2313
tri 3963 2283 3993 2313 sw
tri 4061 2283 4091 2313 ne
rect 4091 2283 4513 2313
tri 4513 2283 4543 2313 sw
tri 4611 2283 4641 2313 ne
rect 4641 2283 5063 2313
tri 5063 2283 5093 2313 sw
tri 5161 2283 5191 2313 ne
rect 5191 2283 5613 2313
tri 5613 2283 5643 2313 sw
tri 5711 2283 5741 2313 ne
rect 5741 2283 6163 2313
tri 6163 2283 6193 2313 sw
tri 6261 2283 6291 2313 ne
rect 6291 2283 6713 2313
tri 6713 2283 6743 2313 sw
tri 6811 2283 6841 2313 ne
rect 6841 2283 7263 2313
tri 7263 2283 7293 2313 sw
tri 7361 2283 7391 2313 ne
rect 7391 2283 7813 2313
tri 7813 2283 7843 2313 sw
tri 7911 2283 7941 2313 ne
rect 7941 2283 8363 2313
tri 8363 2283 8393 2313 sw
tri 8461 2283 8491 2313 ne
rect 8491 2283 8913 2313
tri 8913 2283 8943 2313 sw
tri 9011 2283 9041 2313 ne
rect 9041 2283 9463 2313
tri 9463 2283 9493 2313 sw
tri 9561 2283 9591 2313 ne
rect 9591 2283 10013 2313
tri 10013 2283 10043 2313 sw
tri 10111 2283 10141 2313 ne
rect 10141 2283 10563 2313
tri 10563 2283 10593 2313 sw
tri 10661 2283 10691 2313 ne
rect 10691 2283 11113 2313
tri 11113 2283 11143 2313 sw
tri 11211 2283 11241 2313 ne
rect 11241 2283 11663 2313
tri 11663 2283 11693 2313 sw
tri 11761 2283 11791 2313 ne
rect 11791 2283 12213 2313
tri 12213 2283 12243 2313 sw
tri 12311 2283 12341 2313 ne
rect 12341 2283 12763 2313
tri 12763 2283 12793 2313 sw
tri 12861 2283 12891 2313 ne
rect 12891 2283 13313 2313
tri 13313 2283 13343 2313 sw
tri 13411 2283 13441 2313 ne
rect 13441 2283 13863 2313
tri 13863 2283 13893 2313 sw
tri 13961 2283 13991 2313 ne
rect 13991 2283 14413 2313
tri 14413 2283 14443 2313 sw
tri 14511 2283 14541 2313 ne
rect 14541 2283 14963 2313
tri 14963 2283 14993 2313 sw
tri 15061 2283 15091 2313 ne
rect 15091 2283 15513 2313
tri 15513 2283 15543 2313 sw
tri 15611 2283 15641 2313 ne
rect 15641 2283 16063 2313
tri 16063 2283 16093 2313 sw
tri 16161 2283 16191 2313 ne
rect 16191 2283 16613 2313
tri 16613 2283 16643 2313 sw
tri 16711 2283 16741 2313 ne
rect 16741 2283 17163 2313
tri 17163 2283 17193 2313 sw
tri 17261 2283 17291 2313 ne
rect 17291 2283 17713 2313
tri 17713 2283 17743 2313 sw
tri 17811 2283 17841 2313 ne
rect 17841 2283 18263 2313
tri 18263 2283 18293 2313 sw
tri 18361 2283 18391 2313 ne
rect 18391 2283 18813 2313
tri 18813 2283 18843 2313 sw
tri 18911 2283 18941 2313 ne
rect 18941 2283 19363 2313
tri 19363 2283 19393 2313 sw
tri 19461 2283 19491 2313 ne
rect 19491 2283 20300 2313
rect -2000 2185 143 2283
tri 143 2185 241 2283 sw
tri 241 2185 339 2283 ne
rect 339 2185 693 2283
tri 693 2185 791 2283 sw
tri 791 2185 889 2283 ne
rect 889 2185 1243 2283
tri 1243 2185 1341 2283 sw
tri 1341 2185 1439 2283 ne
rect 1439 2185 1793 2283
tri 1793 2185 1891 2283 sw
tri 1891 2185 1989 2283 ne
rect 1989 2185 2343 2283
tri 2343 2185 2441 2283 sw
tri 2441 2185 2539 2283 ne
rect 2539 2185 2893 2283
tri 2893 2185 2991 2283 sw
tri 2991 2185 3089 2283 ne
rect 3089 2185 3443 2283
tri 3443 2185 3541 2283 sw
tri 3541 2185 3639 2283 ne
rect 3639 2185 3993 2283
tri 3993 2185 4091 2283 sw
tri 4091 2185 4189 2283 ne
rect 4189 2185 4543 2283
tri 4543 2185 4641 2283 sw
tri 4641 2185 4739 2283 ne
rect 4739 2185 5093 2283
tri 5093 2185 5191 2283 sw
tri 5191 2185 5289 2283 ne
rect 5289 2185 5643 2283
tri 5643 2185 5741 2283 sw
tri 5741 2185 5839 2283 ne
rect 5839 2185 6193 2283
tri 6193 2185 6291 2283 sw
tri 6291 2185 6389 2283 ne
rect 6389 2185 6743 2283
tri 6743 2185 6841 2283 sw
tri 6841 2185 6939 2283 ne
rect 6939 2185 7293 2283
tri 7293 2185 7391 2283 sw
tri 7391 2185 7489 2283 ne
rect 7489 2185 7843 2283
tri 7843 2185 7941 2283 sw
tri 7941 2185 8039 2283 ne
rect 8039 2185 8393 2283
tri 8393 2185 8491 2283 sw
tri 8491 2185 8589 2283 ne
rect 8589 2185 8943 2283
tri 8943 2185 9041 2283 sw
tri 9041 2185 9139 2283 ne
rect 9139 2185 9493 2283
tri 9493 2185 9591 2283 sw
tri 9591 2185 9689 2283 ne
rect 9689 2185 10043 2283
tri 10043 2185 10141 2283 sw
tri 10141 2185 10239 2283 ne
rect 10239 2185 10593 2283
tri 10593 2185 10691 2283 sw
tri 10691 2185 10789 2283 ne
rect 10789 2185 11143 2283
tri 11143 2185 11241 2283 sw
tri 11241 2185 11339 2283 ne
rect 11339 2185 11693 2283
tri 11693 2185 11791 2283 sw
tri 11791 2185 11889 2283 ne
rect 11889 2185 12243 2283
tri 12243 2185 12341 2283 sw
tri 12341 2185 12439 2283 ne
rect 12439 2185 12793 2283
tri 12793 2185 12891 2283 sw
tri 12891 2185 12989 2283 ne
rect 12989 2185 13343 2283
tri 13343 2185 13441 2283 sw
tri 13441 2185 13539 2283 ne
rect 13539 2185 13893 2283
tri 13893 2185 13991 2283 sw
tri 13991 2185 14089 2283 ne
rect 14089 2185 14443 2283
tri 14443 2185 14541 2283 sw
tri 14541 2185 14639 2283 ne
rect 14639 2185 14993 2283
tri 14993 2185 15091 2283 sw
tri 15091 2185 15189 2283 ne
rect 15189 2185 15543 2283
tri 15543 2185 15641 2283 sw
tri 15641 2185 15739 2283 ne
rect 15739 2185 16093 2283
tri 16093 2185 16191 2283 sw
tri 16191 2185 16289 2283 ne
rect 16289 2185 16643 2283
tri 16643 2185 16741 2283 sw
tri 16741 2185 16839 2283 ne
rect 16839 2185 17193 2283
tri 17193 2185 17291 2283 sw
tri 17291 2185 17389 2283 ne
rect 17389 2185 17743 2283
tri 17743 2185 17841 2283 sw
tri 17841 2185 17939 2283 ne
rect 17939 2185 18293 2283
tri 18293 2185 18391 2283 sw
tri 18391 2185 18489 2283 ne
rect 18489 2185 18843 2283
tri 18843 2185 18941 2283 sw
tri 18941 2185 19039 2283 ne
rect 19039 2185 19393 2283
tri 19393 2185 19491 2283 sw
tri 19491 2185 19589 2283 ne
rect 19589 2185 20300 2283
rect -2000 2087 241 2185
tri 241 2087 339 2185 sw
tri 339 2087 437 2185 ne
rect 437 2087 791 2185
tri 791 2087 889 2185 sw
tri 889 2087 987 2185 ne
rect 987 2087 1341 2185
tri 1341 2087 1439 2185 sw
tri 1439 2087 1537 2185 ne
rect 1537 2087 1891 2185
tri 1891 2087 1989 2185 sw
tri 1989 2087 2087 2185 ne
rect 2087 2087 2441 2185
tri 2441 2087 2539 2185 sw
tri 2539 2087 2637 2185 ne
rect 2637 2087 2991 2185
tri 2991 2087 3089 2185 sw
tri 3089 2087 3187 2185 ne
rect 3187 2087 3541 2185
tri 3541 2087 3639 2185 sw
tri 3639 2087 3737 2185 ne
rect 3737 2087 4091 2185
tri 4091 2087 4189 2185 sw
tri 4189 2087 4287 2185 ne
rect 4287 2087 4641 2185
tri 4641 2087 4739 2185 sw
tri 4739 2087 4837 2185 ne
rect 4837 2087 5191 2185
tri 5191 2087 5289 2185 sw
tri 5289 2087 5387 2185 ne
rect 5387 2087 5741 2185
tri 5741 2087 5839 2185 sw
tri 5839 2087 5937 2185 ne
rect 5937 2087 6291 2185
tri 6291 2087 6389 2185 sw
tri 6389 2087 6487 2185 ne
rect 6487 2087 6841 2185
tri 6841 2087 6939 2185 sw
tri 6939 2087 7037 2185 ne
rect 7037 2087 7391 2185
tri 7391 2087 7489 2185 sw
tri 7489 2087 7587 2185 ne
rect 7587 2087 7941 2185
tri 7941 2087 8039 2185 sw
tri 8039 2087 8137 2185 ne
rect 8137 2087 8491 2185
tri 8491 2087 8589 2185 sw
tri 8589 2087 8687 2185 ne
rect 8687 2087 9041 2185
tri 9041 2087 9139 2185 sw
tri 9139 2087 9237 2185 ne
rect 9237 2087 9591 2185
tri 9591 2087 9689 2185 sw
tri 9689 2087 9787 2185 ne
rect 9787 2087 10141 2185
tri 10141 2087 10239 2185 sw
tri 10239 2087 10337 2185 ne
rect 10337 2087 10691 2185
tri 10691 2087 10789 2185 sw
tri 10789 2087 10887 2185 ne
rect 10887 2087 11241 2185
tri 11241 2087 11339 2185 sw
tri 11339 2087 11437 2185 ne
rect 11437 2087 11791 2185
tri 11791 2087 11889 2185 sw
tri 11889 2087 11987 2185 ne
rect 11987 2087 12341 2185
tri 12341 2087 12439 2185 sw
tri 12439 2087 12537 2185 ne
rect 12537 2087 12891 2185
tri 12891 2087 12989 2185 sw
tri 12989 2087 13087 2185 ne
rect 13087 2087 13441 2185
tri 13441 2087 13539 2185 sw
tri 13539 2087 13637 2185 ne
rect 13637 2087 13991 2185
tri 13991 2087 14089 2185 sw
tri 14089 2087 14187 2185 ne
rect 14187 2087 14541 2185
tri 14541 2087 14639 2185 sw
tri 14639 2087 14737 2185 ne
rect 14737 2087 15091 2185
tri 15091 2087 15189 2185 sw
tri 15189 2087 15287 2185 ne
rect 15287 2087 15641 2185
tri 15641 2087 15739 2185 sw
tri 15739 2087 15837 2185 ne
rect 15837 2087 16191 2185
tri 16191 2087 16289 2185 sw
tri 16289 2087 16387 2185 ne
rect 16387 2087 16741 2185
tri 16741 2087 16839 2185 sw
tri 16839 2087 16937 2185 ne
rect 16937 2087 17291 2185
tri 17291 2087 17389 2185 sw
tri 17389 2087 17487 2185 ne
rect 17487 2087 17841 2185
tri 17841 2087 17939 2185 sw
tri 17939 2087 18037 2185 ne
rect 18037 2087 18391 2185
tri 18391 2087 18489 2185 sw
tri 18489 2087 18587 2185 ne
rect 18587 2087 18941 2185
tri 18941 2087 19039 2185 sw
tri 19039 2087 19137 2185 ne
rect 19137 2087 19491 2185
tri 19491 2087 19589 2185 sw
tri 19589 2087 19687 2185 ne
rect 19687 2087 20300 2185
rect -2000 1989 339 2087
tri 339 1989 437 2087 sw
tri 437 1989 535 2087 ne
rect 535 1989 889 2087
tri 889 1989 987 2087 sw
tri 987 1989 1085 2087 ne
rect 1085 1989 1439 2087
tri 1439 1989 1537 2087 sw
tri 1537 1989 1635 2087 ne
rect 1635 1989 1989 2087
tri 1989 1989 2087 2087 sw
tri 2087 1989 2185 2087 ne
rect 2185 1989 2539 2087
tri 2539 1989 2637 2087 sw
tri 2637 1989 2735 2087 ne
rect 2735 1989 3089 2087
tri 3089 1989 3187 2087 sw
tri 3187 1989 3285 2087 ne
rect 3285 1989 3639 2087
tri 3639 1989 3737 2087 sw
tri 3737 1989 3835 2087 ne
rect 3835 1989 4189 2087
tri 4189 1989 4287 2087 sw
tri 4287 1989 4385 2087 ne
rect 4385 1989 4739 2087
tri 4739 1989 4837 2087 sw
tri 4837 1989 4935 2087 ne
rect 4935 1989 5289 2087
tri 5289 1989 5387 2087 sw
tri 5387 1989 5485 2087 ne
rect 5485 1989 5839 2087
tri 5839 1989 5937 2087 sw
tri 5937 1989 6035 2087 ne
rect 6035 1989 6389 2087
tri 6389 1989 6487 2087 sw
tri 6487 1989 6585 2087 ne
rect 6585 1989 6939 2087
tri 6939 1989 7037 2087 sw
tri 7037 1989 7135 2087 ne
rect 7135 1989 7489 2087
tri 7489 1989 7587 2087 sw
tri 7587 1989 7685 2087 ne
rect 7685 1989 8039 2087
tri 8039 1989 8137 2087 sw
tri 8137 1989 8235 2087 ne
rect 8235 1989 8589 2087
tri 8589 1989 8687 2087 sw
tri 8687 1989 8785 2087 ne
rect 8785 1989 9139 2087
tri 9139 1989 9237 2087 sw
tri 9237 1989 9335 2087 ne
rect 9335 1989 9689 2087
tri 9689 1989 9787 2087 sw
tri 9787 1989 9885 2087 ne
rect 9885 1989 10239 2087
tri 10239 1989 10337 2087 sw
tri 10337 1989 10435 2087 ne
rect 10435 1989 10789 2087
tri 10789 1989 10887 2087 sw
tri 10887 1989 10985 2087 ne
rect 10985 1989 11339 2087
tri 11339 1989 11437 2087 sw
tri 11437 1989 11535 2087 ne
rect 11535 1989 11889 2087
tri 11889 1989 11987 2087 sw
tri 11987 1989 12085 2087 ne
rect 12085 1989 12439 2087
tri 12439 1989 12537 2087 sw
tri 12537 1989 12635 2087 ne
rect 12635 1989 12989 2087
tri 12989 1989 13087 2087 sw
tri 13087 1989 13185 2087 ne
rect 13185 1989 13539 2087
tri 13539 1989 13637 2087 sw
tri 13637 1989 13735 2087 ne
rect 13735 1989 14089 2087
tri 14089 1989 14187 2087 sw
tri 14187 1989 14285 2087 ne
rect 14285 1989 14639 2087
tri 14639 1989 14737 2087 sw
tri 14737 1989 14835 2087 ne
rect 14835 1989 15189 2087
tri 15189 1989 15287 2087 sw
tri 15287 1989 15385 2087 ne
rect 15385 1989 15739 2087
tri 15739 1989 15837 2087 sw
tri 15837 1989 15935 2087 ne
rect 15935 1989 16289 2087
tri 16289 1989 16387 2087 sw
tri 16387 1989 16485 2087 ne
rect 16485 1989 16839 2087
tri 16839 1989 16937 2087 sw
tri 16937 1989 17035 2087 ne
rect 17035 1989 17389 2087
tri 17389 1989 17487 2087 sw
tri 17487 1989 17585 2087 ne
rect 17585 1989 17939 2087
tri 17939 1989 18037 2087 sw
tri 18037 1989 18135 2087 ne
rect 18135 1989 18489 2087
tri 18489 1989 18587 2087 sw
tri 18587 1989 18685 2087 ne
rect 18685 1989 19039 2087
tri 19039 1989 19137 2087 sw
tri 19137 1989 19235 2087 ne
rect 19235 1989 19589 2087
tri 19589 1989 19687 2087 sw
rect 20800 1989 21800 2637
rect -2000 1985 437 1989
rect -2000 1865 215 1985
rect 335 1891 437 1985
tri 437 1891 535 1989 sw
tri 535 1891 633 1989 ne
rect 633 1985 987 1989
rect 633 1891 765 1985
rect 335 1865 535 1891
rect -2000 1861 535 1865
rect -2000 1650 -1000 1861
tri 113 1763 211 1861 ne
rect 211 1813 535 1861
tri 535 1813 613 1891 sw
tri 633 1813 711 1891 ne
rect 711 1865 765 1891
rect 885 1891 987 1985
tri 987 1891 1085 1989 sw
tri 1085 1891 1183 1989 ne
rect 1183 1985 1537 1989
rect 1183 1891 1315 1985
rect 885 1865 1085 1891
rect 711 1813 1085 1865
tri 1085 1813 1163 1891 sw
tri 1183 1813 1261 1891 ne
rect 1261 1865 1315 1891
rect 1435 1891 1537 1985
tri 1537 1891 1635 1989 sw
tri 1635 1891 1733 1989 ne
rect 1733 1985 2087 1989
rect 1733 1891 1865 1985
rect 1435 1865 1635 1891
rect 1261 1813 1635 1865
tri 1635 1813 1713 1891 sw
tri 1733 1813 1811 1891 ne
rect 1811 1865 1865 1891
rect 1985 1891 2087 1985
tri 2087 1891 2185 1989 sw
tri 2185 1891 2283 1989 ne
rect 2283 1985 2637 1989
rect 2283 1891 2415 1985
rect 1985 1865 2185 1891
rect 1811 1813 2185 1865
tri 2185 1813 2263 1891 sw
tri 2283 1813 2361 1891 ne
rect 2361 1865 2415 1891
rect 2535 1891 2637 1985
tri 2637 1891 2735 1989 sw
tri 2735 1891 2833 1989 ne
rect 2833 1985 3187 1989
rect 2833 1891 2965 1985
rect 2535 1865 2735 1891
rect 2361 1813 2735 1865
tri 2735 1813 2813 1891 sw
tri 2833 1813 2911 1891 ne
rect 2911 1865 2965 1891
rect 3085 1891 3187 1985
tri 3187 1891 3285 1989 sw
tri 3285 1891 3383 1989 ne
rect 3383 1985 3737 1989
rect 3383 1891 3515 1985
rect 3085 1865 3285 1891
rect 2911 1813 3285 1865
tri 3285 1813 3363 1891 sw
tri 3383 1813 3461 1891 ne
rect 3461 1865 3515 1891
rect 3635 1891 3737 1985
tri 3737 1891 3835 1989 sw
tri 3835 1891 3933 1989 ne
rect 3933 1985 4287 1989
rect 3933 1891 4065 1985
rect 3635 1865 3835 1891
rect 3461 1813 3835 1865
tri 3835 1813 3913 1891 sw
tri 3933 1813 4011 1891 ne
rect 4011 1865 4065 1891
rect 4185 1891 4287 1985
tri 4287 1891 4385 1989 sw
tri 4385 1891 4483 1989 ne
rect 4483 1985 4837 1989
rect 4483 1891 4615 1985
rect 4185 1865 4385 1891
rect 4011 1813 4385 1865
tri 4385 1813 4463 1891 sw
tri 4483 1813 4561 1891 ne
rect 4561 1865 4615 1891
rect 4735 1891 4837 1985
tri 4837 1891 4935 1989 sw
tri 4935 1891 5033 1989 ne
rect 5033 1985 5387 1989
rect 5033 1891 5165 1985
rect 4735 1865 4935 1891
rect 4561 1813 4935 1865
tri 4935 1813 5013 1891 sw
tri 5033 1813 5111 1891 ne
rect 5111 1865 5165 1891
rect 5285 1891 5387 1985
tri 5387 1891 5485 1989 sw
tri 5485 1891 5583 1989 ne
rect 5583 1985 5937 1989
rect 5583 1891 5715 1985
rect 5285 1865 5485 1891
rect 5111 1813 5485 1865
tri 5485 1813 5563 1891 sw
tri 5583 1813 5661 1891 ne
rect 5661 1865 5715 1891
rect 5835 1891 5937 1985
tri 5937 1891 6035 1989 sw
tri 6035 1891 6133 1989 ne
rect 6133 1985 6487 1989
rect 6133 1891 6265 1985
rect 5835 1865 6035 1891
rect 5661 1813 6035 1865
tri 6035 1813 6113 1891 sw
tri 6133 1813 6211 1891 ne
rect 6211 1865 6265 1891
rect 6385 1891 6487 1985
tri 6487 1891 6585 1989 sw
tri 6585 1891 6683 1989 ne
rect 6683 1985 7037 1989
rect 6683 1891 6815 1985
rect 6385 1865 6585 1891
rect 6211 1813 6585 1865
tri 6585 1813 6663 1891 sw
tri 6683 1813 6761 1891 ne
rect 6761 1865 6815 1891
rect 6935 1891 7037 1985
tri 7037 1891 7135 1989 sw
tri 7135 1891 7233 1989 ne
rect 7233 1985 7587 1989
rect 7233 1891 7365 1985
rect 6935 1865 7135 1891
rect 6761 1813 7135 1865
tri 7135 1813 7213 1891 sw
tri 7233 1813 7311 1891 ne
rect 7311 1865 7365 1891
rect 7485 1891 7587 1985
tri 7587 1891 7685 1989 sw
tri 7685 1891 7783 1989 ne
rect 7783 1985 8137 1989
rect 7783 1891 7915 1985
rect 7485 1865 7685 1891
rect 7311 1813 7685 1865
tri 7685 1813 7763 1891 sw
tri 7783 1813 7861 1891 ne
rect 7861 1865 7915 1891
rect 8035 1891 8137 1985
tri 8137 1891 8235 1989 sw
tri 8235 1891 8333 1989 ne
rect 8333 1985 8687 1989
rect 8333 1891 8465 1985
rect 8035 1865 8235 1891
rect 7861 1813 8235 1865
tri 8235 1813 8313 1891 sw
tri 8333 1813 8411 1891 ne
rect 8411 1865 8465 1891
rect 8585 1891 8687 1985
tri 8687 1891 8785 1989 sw
tri 8785 1891 8883 1989 ne
rect 8883 1985 9237 1989
rect 8883 1891 9015 1985
rect 8585 1865 8785 1891
rect 8411 1813 8785 1865
tri 8785 1813 8863 1891 sw
tri 8883 1813 8961 1891 ne
rect 8961 1865 9015 1891
rect 9135 1891 9237 1985
tri 9237 1891 9335 1989 sw
tri 9335 1891 9433 1989 ne
rect 9433 1985 9787 1989
rect 9433 1891 9565 1985
rect 9135 1865 9335 1891
rect 8961 1813 9335 1865
tri 9335 1813 9413 1891 sw
tri 9433 1813 9511 1891 ne
rect 9511 1865 9565 1891
rect 9685 1891 9787 1985
tri 9787 1891 9885 1989 sw
tri 9885 1891 9983 1989 ne
rect 9983 1985 10337 1989
rect 9983 1891 10115 1985
rect 9685 1865 9885 1891
rect 9511 1813 9885 1865
tri 9885 1813 9963 1891 sw
tri 9983 1813 10061 1891 ne
rect 10061 1865 10115 1891
rect 10235 1891 10337 1985
tri 10337 1891 10435 1989 sw
tri 10435 1891 10533 1989 ne
rect 10533 1985 10887 1989
rect 10533 1891 10665 1985
rect 10235 1865 10435 1891
rect 10061 1813 10435 1865
tri 10435 1813 10513 1891 sw
tri 10533 1813 10611 1891 ne
rect 10611 1865 10665 1891
rect 10785 1891 10887 1985
tri 10887 1891 10985 1989 sw
tri 10985 1891 11083 1989 ne
rect 11083 1985 11437 1989
rect 11083 1891 11215 1985
rect 10785 1865 10985 1891
rect 10611 1813 10985 1865
tri 10985 1813 11063 1891 sw
tri 11083 1813 11161 1891 ne
rect 11161 1865 11215 1891
rect 11335 1891 11437 1985
tri 11437 1891 11535 1989 sw
tri 11535 1891 11633 1989 ne
rect 11633 1985 11987 1989
rect 11633 1891 11765 1985
rect 11335 1865 11535 1891
rect 11161 1813 11535 1865
tri 11535 1813 11613 1891 sw
tri 11633 1813 11711 1891 ne
rect 11711 1865 11765 1891
rect 11885 1891 11987 1985
tri 11987 1891 12085 1989 sw
tri 12085 1891 12183 1989 ne
rect 12183 1985 12537 1989
rect 12183 1891 12315 1985
rect 11885 1865 12085 1891
rect 11711 1813 12085 1865
tri 12085 1813 12163 1891 sw
tri 12183 1813 12261 1891 ne
rect 12261 1865 12315 1891
rect 12435 1891 12537 1985
tri 12537 1891 12635 1989 sw
tri 12635 1891 12733 1989 ne
rect 12733 1985 13087 1989
rect 12733 1891 12865 1985
rect 12435 1865 12635 1891
rect 12261 1813 12635 1865
tri 12635 1813 12713 1891 sw
tri 12733 1813 12811 1891 ne
rect 12811 1865 12865 1891
rect 12985 1891 13087 1985
tri 13087 1891 13185 1989 sw
tri 13185 1891 13283 1989 ne
rect 13283 1985 13637 1989
rect 13283 1891 13415 1985
rect 12985 1865 13185 1891
rect 12811 1813 13185 1865
tri 13185 1813 13263 1891 sw
tri 13283 1813 13361 1891 ne
rect 13361 1865 13415 1891
rect 13535 1891 13637 1985
tri 13637 1891 13735 1989 sw
tri 13735 1891 13833 1989 ne
rect 13833 1985 14187 1989
rect 13833 1891 13965 1985
rect 13535 1865 13735 1891
rect 13361 1813 13735 1865
tri 13735 1813 13813 1891 sw
tri 13833 1813 13911 1891 ne
rect 13911 1865 13965 1891
rect 14085 1891 14187 1985
tri 14187 1891 14285 1989 sw
tri 14285 1891 14383 1989 ne
rect 14383 1985 14737 1989
rect 14383 1891 14515 1985
rect 14085 1865 14285 1891
rect 13911 1813 14285 1865
tri 14285 1813 14363 1891 sw
tri 14383 1813 14461 1891 ne
rect 14461 1865 14515 1891
rect 14635 1891 14737 1985
tri 14737 1891 14835 1989 sw
tri 14835 1891 14933 1989 ne
rect 14933 1985 15287 1989
rect 14933 1891 15065 1985
rect 14635 1865 14835 1891
rect 14461 1813 14835 1865
tri 14835 1813 14913 1891 sw
tri 14933 1813 15011 1891 ne
rect 15011 1865 15065 1891
rect 15185 1891 15287 1985
tri 15287 1891 15385 1989 sw
tri 15385 1891 15483 1989 ne
rect 15483 1985 15837 1989
rect 15483 1891 15615 1985
rect 15185 1865 15385 1891
rect 15011 1813 15385 1865
tri 15385 1813 15463 1891 sw
tri 15483 1813 15561 1891 ne
rect 15561 1865 15615 1891
rect 15735 1891 15837 1985
tri 15837 1891 15935 1989 sw
tri 15935 1891 16033 1989 ne
rect 16033 1985 16387 1989
rect 16033 1891 16165 1985
rect 15735 1865 15935 1891
rect 15561 1813 15935 1865
tri 15935 1813 16013 1891 sw
tri 16033 1813 16111 1891 ne
rect 16111 1865 16165 1891
rect 16285 1891 16387 1985
tri 16387 1891 16485 1989 sw
tri 16485 1891 16583 1989 ne
rect 16583 1985 16937 1989
rect 16583 1891 16715 1985
rect 16285 1865 16485 1891
rect 16111 1813 16485 1865
tri 16485 1813 16563 1891 sw
tri 16583 1813 16661 1891 ne
rect 16661 1865 16715 1891
rect 16835 1891 16937 1985
tri 16937 1891 17035 1989 sw
tri 17035 1891 17133 1989 ne
rect 17133 1985 17487 1989
rect 17133 1891 17265 1985
rect 16835 1865 17035 1891
rect 16661 1813 17035 1865
tri 17035 1813 17113 1891 sw
tri 17133 1813 17211 1891 ne
rect 17211 1865 17265 1891
rect 17385 1891 17487 1985
tri 17487 1891 17585 1989 sw
tri 17585 1891 17683 1989 ne
rect 17683 1985 18037 1989
rect 17683 1891 17815 1985
rect 17385 1865 17585 1891
rect 17211 1813 17585 1865
tri 17585 1813 17663 1891 sw
tri 17683 1813 17761 1891 ne
rect 17761 1865 17815 1891
rect 17935 1891 18037 1985
tri 18037 1891 18135 1989 sw
tri 18135 1891 18233 1989 ne
rect 18233 1985 18587 1989
rect 18233 1891 18365 1985
rect 17935 1865 18135 1891
rect 17761 1813 18135 1865
tri 18135 1813 18213 1891 sw
tri 18233 1813 18311 1891 ne
rect 18311 1865 18365 1891
rect 18485 1891 18587 1985
tri 18587 1891 18685 1989 sw
tri 18685 1891 18783 1989 ne
rect 18783 1985 19137 1989
rect 18783 1891 18915 1985
rect 18485 1865 18685 1891
rect 18311 1813 18685 1865
tri 18685 1813 18763 1891 sw
tri 18783 1813 18861 1891 ne
rect 18861 1865 18915 1891
rect 19035 1891 19137 1985
tri 19137 1891 19235 1989 sw
tri 19235 1891 19333 1989 ne
rect 19333 1985 21800 1989
rect 19333 1891 19465 1985
rect 19035 1865 19235 1891
rect 18861 1813 19235 1865
tri 19235 1813 19313 1891 sw
tri 19333 1813 19411 1891 ne
rect 19411 1865 19465 1891
rect 19585 1865 21800 1985
rect 19411 1813 21800 1865
rect 211 1763 613 1813
rect -500 1713 113 1763
tri 113 1713 163 1763 sw
tri 211 1713 261 1763 ne
rect 261 1733 613 1763
tri 613 1733 693 1813 sw
tri 711 1733 791 1813 ne
rect 791 1733 1163 1813
tri 1163 1733 1243 1813 sw
tri 1261 1733 1341 1813 ne
rect 1341 1733 1713 1813
tri 1713 1733 1793 1813 sw
tri 1811 1733 1891 1813 ne
rect 1891 1733 2263 1813
tri 2263 1733 2343 1813 sw
tri 2361 1733 2441 1813 ne
rect 2441 1733 2813 1813
tri 2813 1733 2893 1813 sw
tri 2911 1733 2991 1813 ne
rect 2991 1733 3363 1813
tri 3363 1733 3443 1813 sw
tri 3461 1733 3541 1813 ne
rect 3541 1733 3913 1813
tri 3913 1733 3993 1813 sw
tri 4011 1733 4091 1813 ne
rect 4091 1733 4463 1813
tri 4463 1733 4543 1813 sw
tri 4561 1733 4641 1813 ne
rect 4641 1733 5013 1813
tri 5013 1733 5093 1813 sw
tri 5111 1733 5191 1813 ne
rect 5191 1733 5563 1813
tri 5563 1733 5643 1813 sw
tri 5661 1733 5741 1813 ne
rect 5741 1733 6113 1813
tri 6113 1733 6193 1813 sw
tri 6211 1733 6291 1813 ne
rect 6291 1733 6663 1813
tri 6663 1733 6743 1813 sw
tri 6761 1733 6841 1813 ne
rect 6841 1733 7213 1813
tri 7213 1733 7293 1813 sw
tri 7311 1733 7391 1813 ne
rect 7391 1733 7763 1813
tri 7763 1733 7843 1813 sw
tri 7861 1733 7941 1813 ne
rect 7941 1733 8313 1813
tri 8313 1733 8393 1813 sw
tri 8411 1733 8491 1813 ne
rect 8491 1733 8863 1813
tri 8863 1733 8943 1813 sw
tri 8961 1733 9041 1813 ne
rect 9041 1733 9413 1813
tri 9413 1733 9493 1813 sw
tri 9511 1733 9591 1813 ne
rect 9591 1733 9963 1813
tri 9963 1733 10043 1813 sw
tri 10061 1733 10141 1813 ne
rect 10141 1733 10513 1813
tri 10513 1733 10593 1813 sw
tri 10611 1733 10691 1813 ne
rect 10691 1733 11063 1813
tri 11063 1733 11143 1813 sw
tri 11161 1733 11241 1813 ne
rect 11241 1733 11613 1813
tri 11613 1733 11693 1813 sw
tri 11711 1733 11791 1813 ne
rect 11791 1733 12163 1813
tri 12163 1733 12243 1813 sw
tri 12261 1733 12341 1813 ne
rect 12341 1733 12713 1813
tri 12713 1733 12793 1813 sw
tri 12811 1733 12891 1813 ne
rect 12891 1733 13263 1813
tri 13263 1733 13343 1813 sw
tri 13361 1733 13441 1813 ne
rect 13441 1733 13813 1813
tri 13813 1733 13893 1813 sw
tri 13911 1733 13991 1813 ne
rect 13991 1733 14363 1813
tri 14363 1733 14443 1813 sw
tri 14461 1733 14541 1813 ne
rect 14541 1733 14913 1813
tri 14913 1733 14993 1813 sw
tri 15011 1733 15091 1813 ne
rect 15091 1733 15463 1813
tri 15463 1733 15543 1813 sw
tri 15561 1733 15641 1813 ne
rect 15641 1733 16013 1813
tri 16013 1733 16093 1813 sw
tri 16111 1733 16191 1813 ne
rect 16191 1733 16563 1813
tri 16563 1733 16643 1813 sw
tri 16661 1733 16741 1813 ne
rect 16741 1733 17113 1813
tri 17113 1733 17193 1813 sw
tri 17211 1733 17291 1813 ne
rect 17291 1733 17663 1813
tri 17663 1733 17743 1813 sw
tri 17761 1733 17841 1813 ne
rect 17841 1733 18213 1813
tri 18213 1733 18293 1813 sw
tri 18311 1733 18391 1813 ne
rect 18391 1733 18763 1813
tri 18763 1733 18843 1813 sw
tri 18861 1733 18941 1813 ne
rect 18941 1733 19313 1813
tri 19313 1733 19393 1813 sw
tri 19411 1733 19491 1813 ne
rect 19491 1733 20100 1813
rect 261 1713 693 1733
rect -500 1635 163 1713
tri 163 1635 241 1713 sw
tri 261 1635 339 1713 ne
rect 339 1635 693 1713
tri 693 1635 791 1733 sw
tri 791 1635 889 1733 ne
rect 889 1635 1243 1733
tri 1243 1635 1341 1733 sw
tri 1341 1635 1439 1733 ne
rect 1439 1635 1793 1733
tri 1793 1635 1891 1733 sw
tri 1891 1635 1989 1733 ne
rect 1989 1635 2343 1733
tri 2343 1635 2441 1733 sw
tri 2441 1635 2539 1733 ne
rect 2539 1635 2893 1733
tri 2893 1635 2991 1733 sw
tri 2991 1635 3089 1733 ne
rect 3089 1635 3443 1733
tri 3443 1635 3541 1733 sw
tri 3541 1635 3639 1733 ne
rect 3639 1635 3993 1733
tri 3993 1635 4091 1733 sw
tri 4091 1635 4189 1733 ne
rect 4189 1635 4543 1733
tri 4543 1635 4641 1733 sw
tri 4641 1635 4739 1733 ne
rect 4739 1635 5093 1733
tri 5093 1635 5191 1733 sw
tri 5191 1635 5289 1733 ne
rect 5289 1635 5643 1733
tri 5643 1635 5741 1733 sw
tri 5741 1635 5839 1733 ne
rect 5839 1635 6193 1733
tri 6193 1635 6291 1733 sw
tri 6291 1635 6389 1733 ne
rect 6389 1635 6743 1733
tri 6743 1635 6841 1733 sw
tri 6841 1635 6939 1733 ne
rect 6939 1635 7293 1733
tri 7293 1635 7391 1733 sw
tri 7391 1635 7489 1733 ne
rect 7489 1635 7843 1733
tri 7843 1635 7941 1733 sw
tri 7941 1635 8039 1733 ne
rect 8039 1635 8393 1733
tri 8393 1635 8491 1733 sw
tri 8491 1635 8589 1733 ne
rect 8589 1635 8943 1733
tri 8943 1635 9041 1733 sw
tri 9041 1635 9139 1733 ne
rect 9139 1635 9493 1733
tri 9493 1635 9591 1733 sw
tri 9591 1635 9689 1733 ne
rect 9689 1635 10043 1733
tri 10043 1635 10141 1733 sw
tri 10141 1635 10239 1733 ne
rect 10239 1635 10593 1733
tri 10593 1635 10691 1733 sw
tri 10691 1635 10789 1733 ne
rect 10789 1635 11143 1733
tri 11143 1635 11241 1733 sw
tri 11241 1635 11339 1733 ne
rect 11339 1635 11693 1733
tri 11693 1635 11791 1733 sw
tri 11791 1635 11889 1733 ne
rect 11889 1635 12243 1733
tri 12243 1635 12341 1733 sw
tri 12341 1635 12439 1733 ne
rect 12439 1635 12793 1733
tri 12793 1635 12891 1733 sw
tri 12891 1635 12989 1733 ne
rect 12989 1635 13343 1733
tri 13343 1635 13441 1733 sw
tri 13441 1635 13539 1733 ne
rect 13539 1635 13893 1733
tri 13893 1635 13991 1733 sw
tri 13991 1635 14089 1733 ne
rect 14089 1635 14443 1733
tri 14443 1635 14541 1733 sw
tri 14541 1635 14639 1733 ne
rect 14639 1635 14993 1733
tri 14993 1635 15091 1733 sw
tri 15091 1635 15189 1733 ne
rect 15189 1635 15543 1733
tri 15543 1635 15641 1733 sw
tri 15641 1635 15739 1733 ne
rect 15739 1635 16093 1733
tri 16093 1635 16191 1733 sw
tri 16191 1635 16289 1733 ne
rect 16289 1635 16643 1733
tri 16643 1635 16741 1733 sw
tri 16741 1635 16839 1733 ne
rect 16839 1635 17193 1733
tri 17193 1635 17291 1733 sw
tri 17291 1635 17389 1733 ne
rect 17389 1635 17743 1733
tri 17743 1635 17841 1733 sw
tri 17841 1635 17939 1733 ne
rect 17939 1635 18293 1733
tri 18293 1635 18391 1733 sw
tri 18391 1635 18489 1733 ne
rect 18489 1635 18843 1733
tri 18843 1635 18941 1733 sw
tri 18941 1635 19039 1733 ne
rect 19039 1635 19393 1733
tri 19393 1635 19491 1733 sw
tri 19491 1635 19589 1733 ne
rect 19589 1713 20100 1733
rect 20200 1713 21800 1813
rect 19589 1635 21800 1713
rect -500 1587 241 1635
rect -500 1487 -400 1587
rect -300 1537 241 1587
tri 241 1537 339 1635 sw
tri 339 1537 437 1635 ne
rect 437 1537 791 1635
tri 791 1537 889 1635 sw
tri 889 1537 987 1635 ne
rect 987 1537 1341 1635
tri 1341 1537 1439 1635 sw
tri 1439 1537 1537 1635 ne
rect 1537 1537 1891 1635
tri 1891 1537 1989 1635 sw
tri 1989 1537 2087 1635 ne
rect 2087 1537 2441 1635
tri 2441 1537 2539 1635 sw
tri 2539 1537 2637 1635 ne
rect 2637 1537 2991 1635
tri 2991 1537 3089 1635 sw
tri 3089 1537 3187 1635 ne
rect 3187 1537 3541 1635
tri 3541 1537 3639 1635 sw
tri 3639 1537 3737 1635 ne
rect 3737 1537 4091 1635
tri 4091 1537 4189 1635 sw
tri 4189 1537 4287 1635 ne
rect 4287 1537 4641 1635
tri 4641 1537 4739 1635 sw
tri 4739 1537 4837 1635 ne
rect 4837 1537 5191 1635
tri 5191 1537 5289 1635 sw
tri 5289 1537 5387 1635 ne
rect 5387 1537 5741 1635
tri 5741 1537 5839 1635 sw
tri 5839 1537 5937 1635 ne
rect 5937 1537 6291 1635
tri 6291 1537 6389 1635 sw
tri 6389 1537 6487 1635 ne
rect 6487 1537 6841 1635
tri 6841 1537 6939 1635 sw
tri 6939 1537 7037 1635 ne
rect 7037 1537 7391 1635
tri 7391 1537 7489 1635 sw
tri 7489 1537 7587 1635 ne
rect 7587 1537 7941 1635
tri 7941 1537 8039 1635 sw
tri 8039 1537 8137 1635 ne
rect 8137 1537 8491 1635
tri 8491 1537 8589 1635 sw
tri 8589 1537 8687 1635 ne
rect 8687 1537 9041 1635
tri 9041 1537 9139 1635 sw
tri 9139 1537 9237 1635 ne
rect 9237 1537 9591 1635
tri 9591 1537 9689 1635 sw
tri 9689 1537 9787 1635 ne
rect 9787 1537 10141 1635
tri 10141 1537 10239 1635 sw
tri 10239 1537 10337 1635 ne
rect 10337 1537 10691 1635
tri 10691 1537 10789 1635 sw
tri 10789 1537 10887 1635 ne
rect 10887 1537 11241 1635
tri 11241 1537 11339 1635 sw
tri 11339 1537 11437 1635 ne
rect 11437 1537 11791 1635
tri 11791 1537 11889 1635 sw
tri 11889 1537 11987 1635 ne
rect 11987 1537 12341 1635
tri 12341 1537 12439 1635 sw
tri 12439 1537 12537 1635 ne
rect 12537 1537 12891 1635
tri 12891 1537 12989 1635 sw
tri 12989 1537 13087 1635 ne
rect 13087 1537 13441 1635
tri 13441 1537 13539 1635 sw
tri 13539 1537 13637 1635 ne
rect 13637 1537 13991 1635
tri 13991 1537 14089 1635 sw
tri 14089 1537 14187 1635 ne
rect 14187 1537 14541 1635
tri 14541 1537 14639 1635 sw
tri 14639 1537 14737 1635 ne
rect 14737 1537 15091 1635
tri 15091 1537 15189 1635 sw
tri 15189 1537 15287 1635 ne
rect 15287 1537 15641 1635
tri 15641 1537 15739 1635 sw
tri 15739 1537 15837 1635 ne
rect 15837 1537 16191 1635
tri 16191 1537 16289 1635 sw
tri 16289 1537 16387 1635 ne
rect 16387 1537 16741 1635
tri 16741 1537 16839 1635 sw
tri 16839 1537 16937 1635 ne
rect 16937 1537 17291 1635
tri 17291 1537 17389 1635 sw
tri 17389 1537 17487 1635 ne
rect 17487 1537 17841 1635
tri 17841 1537 17939 1635 sw
tri 17939 1537 18037 1635 ne
rect 18037 1537 18391 1635
tri 18391 1537 18489 1635 sw
tri 18489 1537 18587 1635 ne
rect 18587 1537 18941 1635
tri 18941 1537 19039 1635 sw
tri 19039 1537 19137 1635 ne
rect 19137 1537 19491 1635
tri 19491 1537 19589 1635 sw
tri 19589 1537 19687 1635 ne
rect 19687 1537 21800 1635
rect -300 1487 339 1537
rect -500 1439 339 1487
tri 339 1439 437 1537 sw
tri 437 1439 535 1537 ne
rect 535 1439 889 1537
tri 889 1439 987 1537 sw
tri 987 1439 1085 1537 ne
rect 1085 1439 1439 1537
tri 1439 1439 1537 1537 sw
tri 1537 1439 1635 1537 ne
rect 1635 1439 1989 1537
tri 1989 1439 2087 1537 sw
tri 2087 1439 2185 1537 ne
rect 2185 1439 2539 1537
tri 2539 1439 2637 1537 sw
tri 2637 1439 2735 1537 ne
rect 2735 1439 3089 1537
tri 3089 1439 3187 1537 sw
tri 3187 1439 3285 1537 ne
rect 3285 1439 3639 1537
tri 3639 1439 3737 1537 sw
tri 3737 1439 3835 1537 ne
rect 3835 1439 4189 1537
tri 4189 1439 4287 1537 sw
tri 4287 1439 4385 1537 ne
rect 4385 1439 4739 1537
tri 4739 1439 4837 1537 sw
tri 4837 1439 4935 1537 ne
rect 4935 1439 5289 1537
tri 5289 1439 5387 1537 sw
tri 5387 1439 5485 1537 ne
rect 5485 1439 5839 1537
tri 5839 1439 5937 1537 sw
tri 5937 1439 6035 1537 ne
rect 6035 1439 6389 1537
tri 6389 1439 6487 1537 sw
tri 6487 1439 6585 1537 ne
rect 6585 1439 6939 1537
tri 6939 1439 7037 1537 sw
tri 7037 1439 7135 1537 ne
rect 7135 1439 7489 1537
tri 7489 1439 7587 1537 sw
tri 7587 1439 7685 1537 ne
rect 7685 1439 8039 1537
tri 8039 1439 8137 1537 sw
tri 8137 1439 8235 1537 ne
rect 8235 1439 8589 1537
tri 8589 1439 8687 1537 sw
tri 8687 1439 8785 1537 ne
rect 8785 1439 9139 1537
tri 9139 1439 9237 1537 sw
tri 9237 1439 9335 1537 ne
rect 9335 1439 9689 1537
tri 9689 1439 9787 1537 sw
tri 9787 1439 9885 1537 ne
rect 9885 1439 10239 1537
tri 10239 1439 10337 1537 sw
tri 10337 1439 10435 1537 ne
rect 10435 1439 10789 1537
tri 10789 1439 10887 1537 sw
tri 10887 1439 10985 1537 ne
rect 10985 1439 11339 1537
tri 11339 1439 11437 1537 sw
tri 11437 1439 11535 1537 ne
rect 11535 1439 11889 1537
tri 11889 1439 11987 1537 sw
tri 11987 1439 12085 1537 ne
rect 12085 1439 12439 1537
tri 12439 1439 12537 1537 sw
tri 12537 1439 12635 1537 ne
rect 12635 1439 12989 1537
tri 12989 1439 13087 1537 sw
tri 13087 1439 13185 1537 ne
rect 13185 1439 13539 1537
tri 13539 1439 13637 1537 sw
tri 13637 1439 13735 1537 ne
rect 13735 1439 14089 1537
tri 14089 1439 14187 1537 sw
tri 14187 1439 14285 1537 ne
rect 14285 1439 14639 1537
tri 14639 1439 14737 1537 sw
tri 14737 1439 14835 1537 ne
rect 14835 1439 15189 1537
tri 15189 1439 15287 1537 sw
tri 15287 1439 15385 1537 ne
rect 15385 1439 15739 1537
tri 15739 1439 15837 1537 sw
tri 15837 1439 15935 1537 ne
rect 15935 1439 16289 1537
tri 16289 1439 16387 1537 sw
tri 16387 1439 16485 1537 ne
rect 16485 1439 16839 1537
tri 16839 1439 16937 1537 sw
tri 16937 1439 17035 1537 ne
rect 17035 1439 17389 1537
tri 17389 1439 17487 1537 sw
tri 17487 1439 17585 1537 ne
rect 17585 1439 17939 1537
tri 17939 1439 18037 1537 sw
tri 18037 1439 18135 1537 ne
rect 18135 1439 18489 1537
tri 18489 1439 18587 1537 sw
tri 18587 1439 18685 1537 ne
rect 18685 1439 19039 1537
tri 19039 1439 19137 1537 sw
tri 19137 1439 19235 1537 ne
rect 19235 1439 19589 1537
tri 19589 1439 19687 1537 sw
rect -500 1435 437 1439
rect -500 1315 215 1435
rect 335 1341 437 1435
tri 437 1341 535 1439 sw
tri 535 1341 633 1439 ne
rect 633 1435 987 1439
rect 633 1341 765 1435
rect 335 1315 535 1341
rect -500 1311 535 1315
tri 535 1311 565 1341 sw
tri 633 1311 663 1341 ne
rect 663 1315 765 1341
rect 885 1341 987 1435
tri 987 1341 1085 1439 sw
tri 1085 1341 1183 1439 ne
rect 1183 1435 1537 1439
rect 1183 1341 1315 1435
rect 885 1315 1085 1341
rect 663 1311 1085 1315
tri 1085 1311 1115 1341 sw
tri 1183 1311 1213 1341 ne
rect 1213 1315 1315 1341
rect 1435 1341 1537 1435
tri 1537 1341 1635 1439 sw
tri 1635 1341 1733 1439 ne
rect 1733 1435 2087 1439
rect 1733 1341 1865 1435
rect 1435 1315 1635 1341
rect 1213 1311 1635 1315
tri 1635 1311 1665 1341 sw
tri 1733 1311 1763 1341 ne
rect 1763 1315 1865 1341
rect 1985 1341 2087 1435
tri 2087 1341 2185 1439 sw
tri 2185 1341 2283 1439 ne
rect 2283 1435 2637 1439
rect 2283 1341 2415 1435
rect 1985 1315 2185 1341
rect 1763 1311 2185 1315
tri 2185 1311 2215 1341 sw
tri 2283 1311 2313 1341 ne
rect 2313 1315 2415 1341
rect 2535 1341 2637 1435
tri 2637 1341 2735 1439 sw
tri 2735 1341 2833 1439 ne
rect 2833 1435 3187 1439
rect 2833 1341 2965 1435
rect 2535 1315 2735 1341
rect 2313 1311 2735 1315
tri 2735 1311 2765 1341 sw
tri 2833 1311 2863 1341 ne
rect 2863 1315 2965 1341
rect 3085 1341 3187 1435
tri 3187 1341 3285 1439 sw
tri 3285 1341 3383 1439 ne
rect 3383 1435 3737 1439
rect 3383 1341 3515 1435
rect 3085 1315 3285 1341
rect 2863 1311 3285 1315
tri 3285 1311 3315 1341 sw
tri 3383 1311 3413 1341 ne
rect 3413 1315 3515 1341
rect 3635 1341 3737 1435
tri 3737 1341 3835 1439 sw
tri 3835 1341 3933 1439 ne
rect 3933 1435 4287 1439
rect 3933 1341 4065 1435
rect 3635 1315 3835 1341
rect 3413 1311 3835 1315
tri 3835 1311 3865 1341 sw
tri 3933 1311 3963 1341 ne
rect 3963 1315 4065 1341
rect 4185 1341 4287 1435
tri 4287 1341 4385 1439 sw
tri 4385 1341 4483 1439 ne
rect 4483 1435 4837 1439
rect 4483 1341 4615 1435
rect 4185 1315 4385 1341
rect 3963 1311 4385 1315
tri 4385 1311 4415 1341 sw
tri 4483 1311 4513 1341 ne
rect 4513 1315 4615 1341
rect 4735 1341 4837 1435
tri 4837 1341 4935 1439 sw
tri 4935 1341 5033 1439 ne
rect 5033 1435 5387 1439
rect 5033 1341 5165 1435
rect 4735 1315 4935 1341
rect 4513 1311 4935 1315
tri 4935 1311 4965 1341 sw
tri 5033 1311 5063 1341 ne
rect 5063 1315 5165 1341
rect 5285 1341 5387 1435
tri 5387 1341 5485 1439 sw
tri 5485 1341 5583 1439 ne
rect 5583 1435 5937 1439
rect 5583 1341 5715 1435
rect 5285 1315 5485 1341
rect 5063 1311 5485 1315
tri 5485 1311 5515 1341 sw
tri 5583 1311 5613 1341 ne
rect 5613 1315 5715 1341
rect 5835 1341 5937 1435
tri 5937 1341 6035 1439 sw
tri 6035 1341 6133 1439 ne
rect 6133 1435 6487 1439
rect 6133 1341 6265 1435
rect 5835 1315 6035 1341
rect 5613 1311 6035 1315
tri 6035 1311 6065 1341 sw
tri 6133 1311 6163 1341 ne
rect 6163 1315 6265 1341
rect 6385 1341 6487 1435
tri 6487 1341 6585 1439 sw
tri 6585 1341 6683 1439 ne
rect 6683 1435 7037 1439
rect 6683 1341 6815 1435
rect 6385 1315 6585 1341
rect 6163 1311 6585 1315
tri 6585 1311 6615 1341 sw
tri 6683 1311 6713 1341 ne
rect 6713 1315 6815 1341
rect 6935 1341 7037 1435
tri 7037 1341 7135 1439 sw
tri 7135 1341 7233 1439 ne
rect 7233 1435 7587 1439
rect 7233 1341 7365 1435
rect 6935 1315 7135 1341
rect 6713 1311 7135 1315
tri 7135 1311 7165 1341 sw
tri 7233 1311 7263 1341 ne
rect 7263 1315 7365 1341
rect 7485 1341 7587 1435
tri 7587 1341 7685 1439 sw
tri 7685 1341 7783 1439 ne
rect 7783 1435 8137 1439
rect 7783 1341 7915 1435
rect 7485 1315 7685 1341
rect 7263 1311 7685 1315
tri 7685 1311 7715 1341 sw
tri 7783 1311 7813 1341 ne
rect 7813 1315 7915 1341
rect 8035 1341 8137 1435
tri 8137 1341 8235 1439 sw
tri 8235 1341 8333 1439 ne
rect 8333 1435 8687 1439
rect 8333 1341 8465 1435
rect 8035 1315 8235 1341
rect 7813 1311 8235 1315
tri 8235 1311 8265 1341 sw
tri 8333 1311 8363 1341 ne
rect 8363 1315 8465 1341
rect 8585 1341 8687 1435
tri 8687 1341 8785 1439 sw
tri 8785 1341 8883 1439 ne
rect 8883 1435 9237 1439
rect 8883 1341 9015 1435
rect 8585 1315 8785 1341
rect 8363 1311 8785 1315
tri 8785 1311 8815 1341 sw
tri 8883 1311 8913 1341 ne
rect 8913 1315 9015 1341
rect 9135 1341 9237 1435
tri 9237 1341 9335 1439 sw
tri 9335 1341 9433 1439 ne
rect 9433 1435 9787 1439
rect 9433 1341 9565 1435
rect 9135 1315 9335 1341
rect 8913 1311 9335 1315
tri 9335 1311 9365 1341 sw
tri 9433 1311 9463 1341 ne
rect 9463 1315 9565 1341
rect 9685 1341 9787 1435
tri 9787 1341 9885 1439 sw
tri 9885 1341 9983 1439 ne
rect 9983 1435 10337 1439
rect 9983 1341 10115 1435
rect 9685 1315 9885 1341
rect 9463 1311 9885 1315
tri 9885 1311 9915 1341 sw
tri 9983 1311 10013 1341 ne
rect 10013 1315 10115 1341
rect 10235 1341 10337 1435
tri 10337 1341 10435 1439 sw
tri 10435 1341 10533 1439 ne
rect 10533 1435 10887 1439
rect 10533 1341 10665 1435
rect 10235 1315 10435 1341
rect 10013 1311 10435 1315
tri 10435 1311 10465 1341 sw
tri 10533 1311 10563 1341 ne
rect 10563 1315 10665 1341
rect 10785 1341 10887 1435
tri 10887 1341 10985 1439 sw
tri 10985 1341 11083 1439 ne
rect 11083 1435 11437 1439
rect 11083 1341 11215 1435
rect 10785 1315 10985 1341
rect 10563 1311 10985 1315
tri 10985 1311 11015 1341 sw
tri 11083 1311 11113 1341 ne
rect 11113 1315 11215 1341
rect 11335 1341 11437 1435
tri 11437 1341 11535 1439 sw
tri 11535 1341 11633 1439 ne
rect 11633 1435 11987 1439
rect 11633 1341 11765 1435
rect 11335 1315 11535 1341
rect 11113 1311 11535 1315
tri 11535 1311 11565 1341 sw
tri 11633 1311 11663 1341 ne
rect 11663 1315 11765 1341
rect 11885 1341 11987 1435
tri 11987 1341 12085 1439 sw
tri 12085 1341 12183 1439 ne
rect 12183 1435 12537 1439
rect 12183 1341 12315 1435
rect 11885 1315 12085 1341
rect 11663 1311 12085 1315
tri 12085 1311 12115 1341 sw
tri 12183 1311 12213 1341 ne
rect 12213 1315 12315 1341
rect 12435 1341 12537 1435
tri 12537 1341 12635 1439 sw
tri 12635 1341 12733 1439 ne
rect 12733 1435 13087 1439
rect 12733 1341 12865 1435
rect 12435 1315 12635 1341
rect 12213 1311 12635 1315
tri 12635 1311 12665 1341 sw
tri 12733 1311 12763 1341 ne
rect 12763 1315 12865 1341
rect 12985 1341 13087 1435
tri 13087 1341 13185 1439 sw
tri 13185 1341 13283 1439 ne
rect 13283 1435 13637 1439
rect 13283 1341 13415 1435
rect 12985 1315 13185 1341
rect 12763 1311 13185 1315
tri 13185 1311 13215 1341 sw
tri 13283 1311 13313 1341 ne
rect 13313 1315 13415 1341
rect 13535 1341 13637 1435
tri 13637 1341 13735 1439 sw
tri 13735 1341 13833 1439 ne
rect 13833 1435 14187 1439
rect 13833 1341 13965 1435
rect 13535 1315 13735 1341
rect 13313 1311 13735 1315
tri 13735 1311 13765 1341 sw
tri 13833 1311 13863 1341 ne
rect 13863 1315 13965 1341
rect 14085 1341 14187 1435
tri 14187 1341 14285 1439 sw
tri 14285 1341 14383 1439 ne
rect 14383 1435 14737 1439
rect 14383 1341 14515 1435
rect 14085 1315 14285 1341
rect 13863 1311 14285 1315
tri 14285 1311 14315 1341 sw
tri 14383 1311 14413 1341 ne
rect 14413 1315 14515 1341
rect 14635 1341 14737 1435
tri 14737 1341 14835 1439 sw
tri 14835 1341 14933 1439 ne
rect 14933 1435 15287 1439
rect 14933 1341 15065 1435
rect 14635 1315 14835 1341
rect 14413 1311 14835 1315
tri 14835 1311 14865 1341 sw
tri 14933 1311 14963 1341 ne
rect 14963 1315 15065 1341
rect 15185 1341 15287 1435
tri 15287 1341 15385 1439 sw
tri 15385 1341 15483 1439 ne
rect 15483 1435 15837 1439
rect 15483 1341 15615 1435
rect 15185 1315 15385 1341
rect 14963 1311 15385 1315
tri 15385 1311 15415 1341 sw
tri 15483 1311 15513 1341 ne
rect 15513 1315 15615 1341
rect 15735 1341 15837 1435
tri 15837 1341 15935 1439 sw
tri 15935 1341 16033 1439 ne
rect 16033 1435 16387 1439
rect 16033 1341 16165 1435
rect 15735 1315 15935 1341
rect 15513 1311 15935 1315
tri 15935 1311 15965 1341 sw
tri 16033 1311 16063 1341 ne
rect 16063 1315 16165 1341
rect 16285 1341 16387 1435
tri 16387 1341 16485 1439 sw
tri 16485 1341 16583 1439 ne
rect 16583 1435 16937 1439
rect 16583 1341 16715 1435
rect 16285 1315 16485 1341
rect 16063 1311 16485 1315
tri 16485 1311 16515 1341 sw
tri 16583 1311 16613 1341 ne
rect 16613 1315 16715 1341
rect 16835 1341 16937 1435
tri 16937 1341 17035 1439 sw
tri 17035 1341 17133 1439 ne
rect 17133 1435 17487 1439
rect 17133 1341 17265 1435
rect 16835 1315 17035 1341
rect 16613 1311 17035 1315
tri 17035 1311 17065 1341 sw
tri 17133 1311 17163 1341 ne
rect 17163 1315 17265 1341
rect 17385 1341 17487 1435
tri 17487 1341 17585 1439 sw
tri 17585 1341 17683 1439 ne
rect 17683 1435 18037 1439
rect 17683 1341 17815 1435
rect 17385 1315 17585 1341
rect 17163 1311 17585 1315
tri 17585 1311 17615 1341 sw
tri 17683 1311 17713 1341 ne
rect 17713 1315 17815 1341
rect 17935 1341 18037 1435
tri 18037 1341 18135 1439 sw
tri 18135 1341 18233 1439 ne
rect 18233 1435 18587 1439
rect 18233 1341 18365 1435
rect 17935 1315 18135 1341
rect 17713 1311 18135 1315
tri 18135 1311 18165 1341 sw
tri 18233 1311 18263 1341 ne
rect 18263 1315 18365 1341
rect 18485 1341 18587 1435
tri 18587 1341 18685 1439 sw
tri 18685 1341 18783 1439 ne
rect 18783 1435 19137 1439
rect 18783 1341 18915 1435
rect 18485 1315 18685 1341
rect 18263 1311 18685 1315
tri 18685 1311 18715 1341 sw
tri 18783 1311 18813 1341 ne
rect 18813 1315 18915 1341
rect 19035 1341 19137 1435
tri 19137 1341 19235 1439 sw
tri 19235 1341 19333 1439 ne
rect 19333 1435 20300 1439
rect 19333 1341 19465 1435
rect 19035 1315 19235 1341
rect 18813 1311 19235 1315
tri 19235 1311 19265 1341 sw
tri 19333 1311 19363 1341 ne
rect 19363 1315 19465 1341
rect 19585 1315 20300 1435
rect 19363 1311 20300 1315
tri 113 1213 211 1311 ne
rect 211 1213 565 1311
tri 565 1213 663 1311 sw
tri 663 1213 761 1311 ne
rect 761 1213 1115 1311
tri 1115 1213 1213 1311 sw
tri 1213 1213 1311 1311 ne
rect 1311 1213 1665 1311
tri 1665 1213 1763 1311 sw
tri 1763 1213 1861 1311 ne
rect 1861 1213 2215 1311
tri 2215 1213 2313 1311 sw
tri 2313 1213 2411 1311 ne
rect 2411 1213 2765 1311
tri 2765 1213 2863 1311 sw
tri 2863 1213 2961 1311 ne
rect 2961 1213 3315 1311
tri 3315 1213 3413 1311 sw
tri 3413 1213 3511 1311 ne
rect 3511 1213 3865 1311
tri 3865 1213 3963 1311 sw
tri 3963 1213 4061 1311 ne
rect 4061 1213 4415 1311
tri 4415 1213 4513 1311 sw
tri 4513 1213 4611 1311 ne
rect 4611 1213 4965 1311
tri 4965 1213 5063 1311 sw
tri 5063 1213 5161 1311 ne
rect 5161 1213 5515 1311
tri 5515 1213 5613 1311 sw
tri 5613 1213 5711 1311 ne
rect 5711 1213 6065 1311
tri 6065 1213 6163 1311 sw
tri 6163 1213 6261 1311 ne
rect 6261 1213 6615 1311
tri 6615 1213 6713 1311 sw
tri 6713 1213 6811 1311 ne
rect 6811 1213 7165 1311
tri 7165 1213 7263 1311 sw
tri 7263 1213 7361 1311 ne
rect 7361 1213 7715 1311
tri 7715 1213 7813 1311 sw
tri 7813 1213 7911 1311 ne
rect 7911 1213 8265 1311
tri 8265 1213 8363 1311 sw
tri 8363 1213 8461 1311 ne
rect 8461 1213 8815 1311
tri 8815 1213 8913 1311 sw
tri 8913 1213 9011 1311 ne
rect 9011 1213 9365 1311
tri 9365 1213 9463 1311 sw
tri 9463 1213 9561 1311 ne
rect 9561 1213 9915 1311
tri 9915 1213 10013 1311 sw
tri 10013 1213 10111 1311 ne
rect 10111 1213 10465 1311
tri 10465 1213 10563 1311 sw
tri 10563 1213 10661 1311 ne
rect 10661 1213 11015 1311
tri 11015 1213 11113 1311 sw
tri 11113 1213 11211 1311 ne
rect 11211 1213 11565 1311
tri 11565 1213 11663 1311 sw
tri 11663 1213 11761 1311 ne
rect 11761 1213 12115 1311
tri 12115 1213 12213 1311 sw
tri 12213 1213 12311 1311 ne
rect 12311 1213 12665 1311
tri 12665 1213 12763 1311 sw
tri 12763 1213 12861 1311 ne
rect 12861 1213 13215 1311
tri 13215 1213 13313 1311 sw
tri 13313 1213 13411 1311 ne
rect 13411 1213 13765 1311
tri 13765 1213 13863 1311 sw
tri 13863 1213 13961 1311 ne
rect 13961 1213 14315 1311
tri 14315 1213 14413 1311 sw
tri 14413 1213 14511 1311 ne
rect 14511 1213 14865 1311
tri 14865 1213 14963 1311 sw
tri 14963 1213 15061 1311 ne
rect 15061 1213 15415 1311
tri 15415 1213 15513 1311 sw
tri 15513 1213 15611 1311 ne
rect 15611 1213 15965 1311
tri 15965 1213 16063 1311 sw
tri 16063 1213 16161 1311 ne
rect 16161 1213 16515 1311
tri 16515 1213 16613 1311 sw
tri 16613 1213 16711 1311 ne
rect 16711 1213 17065 1311
tri 17065 1213 17163 1311 sw
tri 17163 1213 17261 1311 ne
rect 17261 1213 17615 1311
tri 17615 1213 17713 1311 sw
tri 17713 1213 17811 1311 ne
rect 17811 1213 18165 1311
tri 18165 1213 18263 1311 sw
tri 18263 1213 18361 1311 ne
rect 18361 1213 18715 1311
tri 18715 1213 18813 1311 sw
tri 18813 1213 18911 1311 ne
rect 18911 1213 19265 1311
tri 19265 1213 19363 1311 sw
tri 19363 1213 19461 1311 ne
rect 19461 1213 20300 1311
rect -1000 1183 113 1213
tri 113 1183 143 1213 sw
tri 211 1183 241 1213 ne
rect 241 1183 663 1213
tri 663 1183 693 1213 sw
tri 761 1183 791 1213 ne
rect 791 1183 1213 1213
tri 1213 1183 1243 1213 sw
tri 1311 1183 1341 1213 ne
rect 1341 1183 1763 1213
tri 1763 1183 1793 1213 sw
tri 1861 1183 1891 1213 ne
rect 1891 1183 2313 1213
tri 2313 1183 2343 1213 sw
tri 2411 1183 2441 1213 ne
rect 2441 1183 2863 1213
tri 2863 1183 2893 1213 sw
tri 2961 1183 2991 1213 ne
rect 2991 1183 3413 1213
tri 3413 1183 3443 1213 sw
tri 3511 1183 3541 1213 ne
rect 3541 1183 3963 1213
tri 3963 1183 3993 1213 sw
tri 4061 1183 4091 1213 ne
rect 4091 1183 4513 1213
tri 4513 1183 4543 1213 sw
tri 4611 1183 4641 1213 ne
rect 4641 1183 5063 1213
tri 5063 1183 5093 1213 sw
tri 5161 1183 5191 1213 ne
rect 5191 1183 5613 1213
tri 5613 1183 5643 1213 sw
tri 5711 1183 5741 1213 ne
rect 5741 1183 6163 1213
tri 6163 1183 6193 1213 sw
tri 6261 1183 6291 1213 ne
rect 6291 1183 6713 1213
tri 6713 1183 6743 1213 sw
tri 6811 1183 6841 1213 ne
rect 6841 1183 7263 1213
tri 7263 1183 7293 1213 sw
tri 7361 1183 7391 1213 ne
rect 7391 1183 7813 1213
tri 7813 1183 7843 1213 sw
tri 7911 1183 7941 1213 ne
rect 7941 1183 8363 1213
tri 8363 1183 8393 1213 sw
tri 8461 1183 8491 1213 ne
rect 8491 1183 8913 1213
tri 8913 1183 8943 1213 sw
tri 9011 1183 9041 1213 ne
rect 9041 1183 9463 1213
tri 9463 1183 9493 1213 sw
tri 9561 1183 9591 1213 ne
rect 9591 1183 10013 1213
tri 10013 1183 10043 1213 sw
tri 10111 1183 10141 1213 ne
rect 10141 1183 10563 1213
tri 10563 1183 10593 1213 sw
tri 10661 1183 10691 1213 ne
rect 10691 1183 11113 1213
tri 11113 1183 11143 1213 sw
tri 11211 1183 11241 1213 ne
rect 11241 1183 11663 1213
tri 11663 1183 11693 1213 sw
tri 11761 1183 11791 1213 ne
rect 11791 1183 12213 1213
tri 12213 1183 12243 1213 sw
tri 12311 1183 12341 1213 ne
rect 12341 1183 12763 1213
tri 12763 1183 12793 1213 sw
tri 12861 1183 12891 1213 ne
rect 12891 1183 13313 1213
tri 13313 1183 13343 1213 sw
tri 13411 1183 13441 1213 ne
rect 13441 1183 13863 1213
tri 13863 1183 13893 1213 sw
tri 13961 1183 13991 1213 ne
rect 13991 1183 14413 1213
tri 14413 1183 14443 1213 sw
tri 14511 1183 14541 1213 ne
rect 14541 1183 14963 1213
tri 14963 1183 14993 1213 sw
tri 15061 1183 15091 1213 ne
rect 15091 1183 15513 1213
tri 15513 1183 15543 1213 sw
tri 15611 1183 15641 1213 ne
rect 15641 1183 16063 1213
tri 16063 1183 16093 1213 sw
tri 16161 1183 16191 1213 ne
rect 16191 1183 16613 1213
tri 16613 1183 16643 1213 sw
tri 16711 1183 16741 1213 ne
rect 16741 1183 17163 1213
tri 17163 1183 17193 1213 sw
tri 17261 1183 17291 1213 ne
rect 17291 1183 17713 1213
tri 17713 1183 17743 1213 sw
tri 17811 1183 17841 1213 ne
rect 17841 1183 18263 1213
tri 18263 1183 18293 1213 sw
tri 18361 1183 18391 1213 ne
rect 18391 1183 18813 1213
tri 18813 1183 18843 1213 sw
tri 18911 1183 18941 1213 ne
rect 18941 1183 19363 1213
tri 19363 1183 19393 1213 sw
tri 19461 1183 19491 1213 ne
rect 19491 1183 20300 1213
rect -1000 1085 143 1183
tri 143 1085 241 1183 sw
tri 241 1085 339 1183 ne
rect 339 1085 693 1183
tri 693 1085 791 1183 sw
tri 791 1085 889 1183 ne
rect 889 1085 1243 1183
tri 1243 1085 1341 1183 sw
tri 1341 1085 1439 1183 ne
rect 1439 1085 1793 1183
tri 1793 1085 1891 1183 sw
tri 1891 1085 1989 1183 ne
rect 1989 1085 2343 1183
tri 2343 1085 2441 1183 sw
tri 2441 1085 2539 1183 ne
rect 2539 1085 2893 1183
tri 2893 1085 2991 1183 sw
tri 2991 1085 3089 1183 ne
rect 3089 1085 3443 1183
tri 3443 1085 3541 1183 sw
tri 3541 1085 3639 1183 ne
rect 3639 1085 3993 1183
tri 3993 1085 4091 1183 sw
tri 4091 1085 4189 1183 ne
rect 4189 1085 4543 1183
tri 4543 1085 4641 1183 sw
tri 4641 1085 4739 1183 ne
rect 4739 1085 5093 1183
tri 5093 1085 5191 1183 sw
tri 5191 1085 5289 1183 ne
rect 5289 1085 5643 1183
tri 5643 1085 5741 1183 sw
tri 5741 1085 5839 1183 ne
rect 5839 1085 6193 1183
tri 6193 1085 6291 1183 sw
tri 6291 1085 6389 1183 ne
rect 6389 1085 6743 1183
tri 6743 1085 6841 1183 sw
tri 6841 1085 6939 1183 ne
rect 6939 1085 7293 1183
tri 7293 1085 7391 1183 sw
tri 7391 1085 7489 1183 ne
rect 7489 1085 7843 1183
tri 7843 1085 7941 1183 sw
tri 7941 1085 8039 1183 ne
rect 8039 1085 8393 1183
tri 8393 1085 8491 1183 sw
tri 8491 1085 8589 1183 ne
rect 8589 1085 8943 1183
tri 8943 1085 9041 1183 sw
tri 9041 1085 9139 1183 ne
rect 9139 1085 9493 1183
tri 9493 1085 9591 1183 sw
tri 9591 1085 9689 1183 ne
rect 9689 1085 10043 1183
tri 10043 1085 10141 1183 sw
tri 10141 1085 10239 1183 ne
rect 10239 1085 10593 1183
tri 10593 1085 10691 1183 sw
tri 10691 1085 10789 1183 ne
rect 10789 1085 11143 1183
tri 11143 1085 11241 1183 sw
tri 11241 1085 11339 1183 ne
rect 11339 1085 11693 1183
tri 11693 1085 11791 1183 sw
tri 11791 1085 11889 1183 ne
rect 11889 1085 12243 1183
tri 12243 1085 12341 1183 sw
tri 12341 1085 12439 1183 ne
rect 12439 1085 12793 1183
tri 12793 1085 12891 1183 sw
tri 12891 1085 12989 1183 ne
rect 12989 1085 13343 1183
tri 13343 1085 13441 1183 sw
tri 13441 1085 13539 1183 ne
rect 13539 1085 13893 1183
tri 13893 1085 13991 1183 sw
tri 13991 1085 14089 1183 ne
rect 14089 1085 14443 1183
tri 14443 1085 14541 1183 sw
tri 14541 1085 14639 1183 ne
rect 14639 1085 14993 1183
tri 14993 1085 15091 1183 sw
tri 15091 1085 15189 1183 ne
rect 15189 1085 15543 1183
tri 15543 1085 15641 1183 sw
tri 15641 1085 15739 1183 ne
rect 15739 1085 16093 1183
tri 16093 1085 16191 1183 sw
tri 16191 1085 16289 1183 ne
rect 16289 1085 16643 1183
tri 16643 1085 16741 1183 sw
tri 16741 1085 16839 1183 ne
rect 16839 1085 17193 1183
tri 17193 1085 17291 1183 sw
tri 17291 1085 17389 1183 ne
rect 17389 1085 17743 1183
tri 17743 1085 17841 1183 sw
tri 17841 1085 17939 1183 ne
rect 17939 1085 18293 1183
tri 18293 1085 18391 1183 sw
tri 18391 1085 18489 1183 ne
rect 18489 1085 18843 1183
tri 18843 1085 18941 1183 sw
tri 18941 1085 19039 1183 ne
rect 19039 1085 19393 1183
tri 19393 1085 19491 1183 sw
tri 19491 1085 19589 1183 ne
rect 19589 1085 20300 1183
rect -1000 987 241 1085
tri 241 987 339 1085 sw
tri 339 987 437 1085 ne
rect 437 987 791 1085
tri 791 987 889 1085 sw
tri 889 987 987 1085 ne
rect 987 987 1341 1085
tri 1341 987 1439 1085 sw
tri 1439 987 1537 1085 ne
rect 1537 987 1891 1085
tri 1891 987 1989 1085 sw
tri 1989 987 2087 1085 ne
rect 2087 987 2441 1085
tri 2441 987 2539 1085 sw
tri 2539 987 2637 1085 ne
rect 2637 987 2991 1085
tri 2991 987 3089 1085 sw
tri 3089 987 3187 1085 ne
rect 3187 987 3541 1085
tri 3541 987 3639 1085 sw
tri 3639 987 3737 1085 ne
rect 3737 987 4091 1085
tri 4091 987 4189 1085 sw
tri 4189 987 4287 1085 ne
rect 4287 987 4641 1085
tri 4641 987 4739 1085 sw
tri 4739 987 4837 1085 ne
rect 4837 987 5191 1085
tri 5191 987 5289 1085 sw
tri 5289 987 5387 1085 ne
rect 5387 987 5741 1085
tri 5741 987 5839 1085 sw
tri 5839 987 5937 1085 ne
rect 5937 987 6291 1085
tri 6291 987 6389 1085 sw
tri 6389 987 6487 1085 ne
rect 6487 987 6841 1085
tri 6841 987 6939 1085 sw
tri 6939 987 7037 1085 ne
rect 7037 987 7391 1085
tri 7391 987 7489 1085 sw
tri 7489 987 7587 1085 ne
rect 7587 987 7941 1085
tri 7941 987 8039 1085 sw
tri 8039 987 8137 1085 ne
rect 8137 987 8491 1085
tri 8491 987 8589 1085 sw
tri 8589 987 8687 1085 ne
rect 8687 987 9041 1085
tri 9041 987 9139 1085 sw
tri 9139 987 9237 1085 ne
rect 9237 987 9591 1085
tri 9591 987 9689 1085 sw
tri 9689 987 9787 1085 ne
rect 9787 987 10141 1085
tri 10141 987 10239 1085 sw
tri 10239 987 10337 1085 ne
rect 10337 987 10691 1085
tri 10691 987 10789 1085 sw
tri 10789 987 10887 1085 ne
rect 10887 987 11241 1085
tri 11241 987 11339 1085 sw
tri 11339 987 11437 1085 ne
rect 11437 987 11791 1085
tri 11791 987 11889 1085 sw
tri 11889 987 11987 1085 ne
rect 11987 987 12341 1085
tri 12341 987 12439 1085 sw
tri 12439 987 12537 1085 ne
rect 12537 987 12891 1085
tri 12891 987 12989 1085 sw
tri 12989 987 13087 1085 ne
rect 13087 987 13441 1085
tri 13441 987 13539 1085 sw
tri 13539 987 13637 1085 ne
rect 13637 987 13991 1085
tri 13991 987 14089 1085 sw
tri 14089 987 14187 1085 ne
rect 14187 987 14541 1085
tri 14541 987 14639 1085 sw
tri 14639 987 14737 1085 ne
rect 14737 987 15091 1085
tri 15091 987 15189 1085 sw
tri 15189 987 15287 1085 ne
rect 15287 987 15641 1085
tri 15641 987 15739 1085 sw
tri 15739 987 15837 1085 ne
rect 15837 987 16191 1085
tri 16191 987 16289 1085 sw
tri 16289 987 16387 1085 ne
rect 16387 987 16741 1085
tri 16741 987 16839 1085 sw
tri 16839 987 16937 1085 ne
rect 16937 987 17291 1085
tri 17291 987 17389 1085 sw
tri 17389 987 17487 1085 ne
rect 17487 987 17841 1085
tri 17841 987 17939 1085 sw
tri 17939 987 18037 1085 ne
rect 18037 987 18391 1085
tri 18391 987 18489 1085 sw
tri 18489 987 18587 1085 ne
rect 18587 987 18941 1085
tri 18941 987 19039 1085 sw
tri 19039 987 19137 1085 ne
rect 19137 987 19491 1085
tri 19491 987 19589 1085 sw
tri 19589 987 19687 1085 ne
rect 19687 987 20300 1085
rect -1000 889 339 987
tri 339 889 437 987 sw
tri 437 889 535 987 ne
rect 535 889 889 987
tri 889 889 987 987 sw
tri 987 889 1085 987 ne
rect 1085 889 1439 987
tri 1439 889 1537 987 sw
tri 1537 889 1635 987 ne
rect 1635 889 1989 987
tri 1989 889 2087 987 sw
tri 2087 889 2185 987 ne
rect 2185 889 2539 987
tri 2539 889 2637 987 sw
tri 2637 889 2735 987 ne
rect 2735 889 3089 987
tri 3089 889 3187 987 sw
tri 3187 889 3285 987 ne
rect 3285 889 3639 987
tri 3639 889 3737 987 sw
tri 3737 889 3835 987 ne
rect 3835 889 4189 987
tri 4189 889 4287 987 sw
tri 4287 889 4385 987 ne
rect 4385 889 4739 987
tri 4739 889 4837 987 sw
tri 4837 889 4935 987 ne
rect 4935 889 5289 987
tri 5289 889 5387 987 sw
tri 5387 889 5485 987 ne
rect 5485 889 5839 987
tri 5839 889 5937 987 sw
tri 5937 889 6035 987 ne
rect 6035 889 6389 987
tri 6389 889 6487 987 sw
tri 6487 889 6585 987 ne
rect 6585 889 6939 987
tri 6939 889 7037 987 sw
tri 7037 889 7135 987 ne
rect 7135 889 7489 987
tri 7489 889 7587 987 sw
tri 7587 889 7685 987 ne
rect 7685 889 8039 987
tri 8039 889 8137 987 sw
tri 8137 889 8235 987 ne
rect 8235 889 8589 987
tri 8589 889 8687 987 sw
tri 8687 889 8785 987 ne
rect 8785 889 9139 987
tri 9139 889 9237 987 sw
tri 9237 889 9335 987 ne
rect 9335 889 9689 987
tri 9689 889 9787 987 sw
tri 9787 889 9885 987 ne
rect 9885 889 10239 987
tri 10239 889 10337 987 sw
tri 10337 889 10435 987 ne
rect 10435 889 10789 987
tri 10789 889 10887 987 sw
tri 10887 889 10985 987 ne
rect 10985 889 11339 987
tri 11339 889 11437 987 sw
tri 11437 889 11535 987 ne
rect 11535 889 11889 987
tri 11889 889 11987 987 sw
tri 11987 889 12085 987 ne
rect 12085 889 12439 987
tri 12439 889 12537 987 sw
tri 12537 889 12635 987 ne
rect 12635 889 12989 987
tri 12989 889 13087 987 sw
tri 13087 889 13185 987 ne
rect 13185 889 13539 987
tri 13539 889 13637 987 sw
tri 13637 889 13735 987 ne
rect 13735 889 14089 987
tri 14089 889 14187 987 sw
tri 14187 889 14285 987 ne
rect 14285 889 14639 987
tri 14639 889 14737 987 sw
tri 14737 889 14835 987 ne
rect 14835 889 15189 987
tri 15189 889 15287 987 sw
tri 15287 889 15385 987 ne
rect 15385 889 15739 987
tri 15739 889 15837 987 sw
tri 15837 889 15935 987 ne
rect 15935 889 16289 987
tri 16289 889 16387 987 sw
tri 16387 889 16485 987 ne
rect 16485 889 16839 987
tri 16839 889 16937 987 sw
tri 16937 889 17035 987 ne
rect 17035 889 17389 987
tri 17389 889 17487 987 sw
tri 17487 889 17585 987 ne
rect 17585 889 17939 987
tri 17939 889 18037 987 sw
tri 18037 889 18135 987 ne
rect 18135 889 18489 987
tri 18489 889 18587 987 sw
tri 18587 889 18685 987 ne
rect 18685 889 19039 987
tri 19039 889 19137 987 sw
tri 19137 889 19235 987 ne
rect 19235 889 19589 987
tri 19589 889 19687 987 sw
rect 20800 889 21800 1537
rect -1000 885 437 889
rect -1000 765 215 885
rect 335 791 437 885
tri 437 791 535 889 sw
tri 535 791 633 889 ne
rect 633 885 987 889
rect 633 791 765 885
rect 335 765 535 791
rect -1000 761 535 765
tri 113 663 211 761 ne
rect 211 713 535 761
tri 535 713 613 791 sw
tri 633 713 711 791 ne
rect 711 765 765 791
rect 885 791 987 885
tri 987 791 1085 889 sw
tri 1085 791 1183 889 ne
rect 1183 885 1537 889
rect 1183 791 1315 885
rect 885 765 1085 791
rect 711 713 1085 765
tri 1085 713 1163 791 sw
tri 1183 713 1261 791 ne
rect 1261 765 1315 791
rect 1435 791 1537 885
tri 1537 791 1635 889 sw
tri 1635 791 1733 889 ne
rect 1733 885 2087 889
rect 1733 791 1865 885
rect 1435 765 1635 791
rect 1261 713 1635 765
tri 1635 713 1713 791 sw
tri 1733 713 1811 791 ne
rect 1811 765 1865 791
rect 1985 791 2087 885
tri 2087 791 2185 889 sw
tri 2185 791 2283 889 ne
rect 2283 885 2637 889
rect 2283 791 2415 885
rect 1985 765 2185 791
rect 1811 713 2185 765
tri 2185 713 2263 791 sw
tri 2283 713 2361 791 ne
rect 2361 765 2415 791
rect 2535 791 2637 885
tri 2637 791 2735 889 sw
tri 2735 791 2833 889 ne
rect 2833 885 3187 889
rect 2833 791 2965 885
rect 2535 765 2735 791
rect 2361 713 2735 765
tri 2735 713 2813 791 sw
tri 2833 713 2911 791 ne
rect 2911 765 2965 791
rect 3085 791 3187 885
tri 3187 791 3285 889 sw
tri 3285 791 3383 889 ne
rect 3383 885 3737 889
rect 3383 791 3515 885
rect 3085 765 3285 791
rect 2911 713 3285 765
tri 3285 713 3363 791 sw
tri 3383 713 3461 791 ne
rect 3461 765 3515 791
rect 3635 791 3737 885
tri 3737 791 3835 889 sw
tri 3835 791 3933 889 ne
rect 3933 885 4287 889
rect 3933 791 4065 885
rect 3635 765 3835 791
rect 3461 713 3835 765
tri 3835 713 3913 791 sw
tri 3933 713 4011 791 ne
rect 4011 765 4065 791
rect 4185 791 4287 885
tri 4287 791 4385 889 sw
tri 4385 791 4483 889 ne
rect 4483 885 4837 889
rect 4483 791 4615 885
rect 4185 765 4385 791
rect 4011 713 4385 765
tri 4385 713 4463 791 sw
tri 4483 713 4561 791 ne
rect 4561 765 4615 791
rect 4735 791 4837 885
tri 4837 791 4935 889 sw
tri 4935 791 5033 889 ne
rect 5033 885 5387 889
rect 5033 791 5165 885
rect 4735 765 4935 791
rect 4561 713 4935 765
tri 4935 713 5013 791 sw
tri 5033 713 5111 791 ne
rect 5111 765 5165 791
rect 5285 791 5387 885
tri 5387 791 5485 889 sw
tri 5485 791 5583 889 ne
rect 5583 885 5937 889
rect 5583 791 5715 885
rect 5285 765 5485 791
rect 5111 713 5485 765
tri 5485 713 5563 791 sw
tri 5583 713 5661 791 ne
rect 5661 765 5715 791
rect 5835 791 5937 885
tri 5937 791 6035 889 sw
tri 6035 791 6133 889 ne
rect 6133 885 6487 889
rect 6133 791 6265 885
rect 5835 765 6035 791
rect 5661 713 6035 765
tri 6035 713 6113 791 sw
tri 6133 713 6211 791 ne
rect 6211 765 6265 791
rect 6385 791 6487 885
tri 6487 791 6585 889 sw
tri 6585 791 6683 889 ne
rect 6683 885 7037 889
rect 6683 791 6815 885
rect 6385 765 6585 791
rect 6211 713 6585 765
tri 6585 713 6663 791 sw
tri 6683 713 6761 791 ne
rect 6761 765 6815 791
rect 6935 791 7037 885
tri 7037 791 7135 889 sw
tri 7135 791 7233 889 ne
rect 7233 885 7587 889
rect 7233 791 7365 885
rect 6935 765 7135 791
rect 6761 713 7135 765
tri 7135 713 7213 791 sw
tri 7233 713 7311 791 ne
rect 7311 765 7365 791
rect 7485 791 7587 885
tri 7587 791 7685 889 sw
tri 7685 791 7783 889 ne
rect 7783 885 8137 889
rect 7783 791 7915 885
rect 7485 765 7685 791
rect 7311 713 7685 765
tri 7685 713 7763 791 sw
tri 7783 713 7861 791 ne
rect 7861 765 7915 791
rect 8035 791 8137 885
tri 8137 791 8235 889 sw
tri 8235 791 8333 889 ne
rect 8333 885 8687 889
rect 8333 791 8465 885
rect 8035 765 8235 791
rect 7861 713 8235 765
tri 8235 713 8313 791 sw
tri 8333 713 8411 791 ne
rect 8411 765 8465 791
rect 8585 791 8687 885
tri 8687 791 8785 889 sw
tri 8785 791 8883 889 ne
rect 8883 885 9237 889
rect 8883 791 9015 885
rect 8585 765 8785 791
rect 8411 713 8785 765
tri 8785 713 8863 791 sw
tri 8883 713 8961 791 ne
rect 8961 765 9015 791
rect 9135 791 9237 885
tri 9237 791 9335 889 sw
tri 9335 791 9433 889 ne
rect 9433 885 9787 889
rect 9433 791 9565 885
rect 9135 765 9335 791
rect 8961 713 9335 765
tri 9335 713 9413 791 sw
tri 9433 713 9511 791 ne
rect 9511 765 9565 791
rect 9685 791 9787 885
tri 9787 791 9885 889 sw
tri 9885 791 9983 889 ne
rect 9983 885 10337 889
rect 9983 791 10115 885
rect 9685 765 9885 791
rect 9511 713 9885 765
tri 9885 713 9963 791 sw
tri 9983 713 10061 791 ne
rect 10061 765 10115 791
rect 10235 791 10337 885
tri 10337 791 10435 889 sw
tri 10435 791 10533 889 ne
rect 10533 885 10887 889
rect 10533 791 10665 885
rect 10235 765 10435 791
rect 10061 713 10435 765
tri 10435 713 10513 791 sw
tri 10533 713 10611 791 ne
rect 10611 765 10665 791
rect 10785 791 10887 885
tri 10887 791 10985 889 sw
tri 10985 791 11083 889 ne
rect 11083 885 11437 889
rect 11083 791 11215 885
rect 10785 765 10985 791
rect 10611 713 10985 765
tri 10985 713 11063 791 sw
tri 11083 713 11161 791 ne
rect 11161 765 11215 791
rect 11335 791 11437 885
tri 11437 791 11535 889 sw
tri 11535 791 11633 889 ne
rect 11633 885 11987 889
rect 11633 791 11765 885
rect 11335 765 11535 791
rect 11161 713 11535 765
tri 11535 713 11613 791 sw
tri 11633 713 11711 791 ne
rect 11711 765 11765 791
rect 11885 791 11987 885
tri 11987 791 12085 889 sw
tri 12085 791 12183 889 ne
rect 12183 885 12537 889
rect 12183 791 12315 885
rect 11885 765 12085 791
rect 11711 713 12085 765
tri 12085 713 12163 791 sw
tri 12183 713 12261 791 ne
rect 12261 765 12315 791
rect 12435 791 12537 885
tri 12537 791 12635 889 sw
tri 12635 791 12733 889 ne
rect 12733 885 13087 889
rect 12733 791 12865 885
rect 12435 765 12635 791
rect 12261 713 12635 765
tri 12635 713 12713 791 sw
tri 12733 713 12811 791 ne
rect 12811 765 12865 791
rect 12985 791 13087 885
tri 13087 791 13185 889 sw
tri 13185 791 13283 889 ne
rect 13283 885 13637 889
rect 13283 791 13415 885
rect 12985 765 13185 791
rect 12811 713 13185 765
tri 13185 713 13263 791 sw
tri 13283 713 13361 791 ne
rect 13361 765 13415 791
rect 13535 791 13637 885
tri 13637 791 13735 889 sw
tri 13735 791 13833 889 ne
rect 13833 885 14187 889
rect 13833 791 13965 885
rect 13535 765 13735 791
rect 13361 713 13735 765
tri 13735 713 13813 791 sw
tri 13833 713 13911 791 ne
rect 13911 765 13965 791
rect 14085 791 14187 885
tri 14187 791 14285 889 sw
tri 14285 791 14383 889 ne
rect 14383 885 14737 889
rect 14383 791 14515 885
rect 14085 765 14285 791
rect 13911 713 14285 765
tri 14285 713 14363 791 sw
tri 14383 713 14461 791 ne
rect 14461 765 14515 791
rect 14635 791 14737 885
tri 14737 791 14835 889 sw
tri 14835 791 14933 889 ne
rect 14933 885 15287 889
rect 14933 791 15065 885
rect 14635 765 14835 791
rect 14461 713 14835 765
tri 14835 713 14913 791 sw
tri 14933 713 15011 791 ne
rect 15011 765 15065 791
rect 15185 791 15287 885
tri 15287 791 15385 889 sw
tri 15385 791 15483 889 ne
rect 15483 885 15837 889
rect 15483 791 15615 885
rect 15185 765 15385 791
rect 15011 713 15385 765
tri 15385 713 15463 791 sw
tri 15483 713 15561 791 ne
rect 15561 765 15615 791
rect 15735 791 15837 885
tri 15837 791 15935 889 sw
tri 15935 791 16033 889 ne
rect 16033 885 16387 889
rect 16033 791 16165 885
rect 15735 765 15935 791
rect 15561 713 15935 765
tri 15935 713 16013 791 sw
tri 16033 713 16111 791 ne
rect 16111 765 16165 791
rect 16285 791 16387 885
tri 16387 791 16485 889 sw
tri 16485 791 16583 889 ne
rect 16583 885 16937 889
rect 16583 791 16715 885
rect 16285 765 16485 791
rect 16111 713 16485 765
tri 16485 713 16563 791 sw
tri 16583 713 16661 791 ne
rect 16661 765 16715 791
rect 16835 791 16937 885
tri 16937 791 17035 889 sw
tri 17035 791 17133 889 ne
rect 17133 885 17487 889
rect 17133 791 17265 885
rect 16835 765 17035 791
rect 16661 713 17035 765
tri 17035 713 17113 791 sw
tri 17133 713 17211 791 ne
rect 17211 765 17265 791
rect 17385 791 17487 885
tri 17487 791 17585 889 sw
tri 17585 791 17683 889 ne
rect 17683 885 18037 889
rect 17683 791 17815 885
rect 17385 765 17585 791
rect 17211 713 17585 765
tri 17585 713 17663 791 sw
tri 17683 713 17761 791 ne
rect 17761 765 17815 791
rect 17935 791 18037 885
tri 18037 791 18135 889 sw
tri 18135 791 18233 889 ne
rect 18233 885 18587 889
rect 18233 791 18365 885
rect 17935 765 18135 791
rect 17761 713 18135 765
tri 18135 713 18213 791 sw
tri 18233 713 18311 791 ne
rect 18311 765 18365 791
rect 18485 791 18587 885
tri 18587 791 18685 889 sw
tri 18685 791 18783 889 ne
rect 18783 885 19137 889
rect 18783 791 18915 885
rect 18485 765 18685 791
rect 18311 713 18685 765
tri 18685 713 18763 791 sw
tri 18783 713 18861 791 ne
rect 18861 765 18915 791
rect 19035 791 19137 885
tri 19137 791 19235 889 sw
tri 19235 791 19333 889 ne
rect 19333 885 21800 889
rect 19333 791 19465 885
rect 19035 765 19235 791
rect 18861 713 19235 765
tri 19235 713 19313 791 sw
tri 19333 713 19411 791 ne
rect 19411 765 19465 791
rect 19585 765 21800 885
rect 19411 713 21800 765
rect 211 663 613 713
rect -500 613 113 663
tri 113 613 163 663 sw
tri 211 613 261 663 ne
rect 261 633 613 663
tri 613 633 693 713 sw
tri 711 633 791 713 ne
rect 791 633 1163 713
tri 1163 633 1243 713 sw
tri 1261 633 1341 713 ne
rect 1341 633 1713 713
tri 1713 633 1793 713 sw
tri 1811 633 1891 713 ne
rect 1891 633 2263 713
tri 2263 633 2343 713 sw
tri 2361 633 2441 713 ne
rect 2441 633 2813 713
tri 2813 633 2893 713 sw
tri 2911 633 2991 713 ne
rect 2991 633 3363 713
tri 3363 633 3443 713 sw
tri 3461 633 3541 713 ne
rect 3541 633 3913 713
tri 3913 633 3993 713 sw
tri 4011 633 4091 713 ne
rect 4091 633 4463 713
tri 4463 633 4543 713 sw
tri 4561 633 4641 713 ne
rect 4641 633 5013 713
tri 5013 633 5093 713 sw
tri 5111 633 5191 713 ne
rect 5191 633 5563 713
tri 5563 633 5643 713 sw
tri 5661 633 5741 713 ne
rect 5741 633 6113 713
tri 6113 633 6193 713 sw
tri 6211 633 6291 713 ne
rect 6291 633 6663 713
tri 6663 633 6743 713 sw
tri 6761 633 6841 713 ne
rect 6841 633 7213 713
tri 7213 633 7293 713 sw
tri 7311 633 7391 713 ne
rect 7391 633 7763 713
tri 7763 633 7843 713 sw
tri 7861 633 7941 713 ne
rect 7941 633 8313 713
tri 8313 633 8393 713 sw
tri 8411 633 8491 713 ne
rect 8491 633 8863 713
tri 8863 633 8943 713 sw
tri 8961 633 9041 713 ne
rect 9041 633 9413 713
tri 9413 633 9493 713 sw
tri 9511 633 9591 713 ne
rect 9591 633 9963 713
tri 9963 633 10043 713 sw
tri 10061 633 10141 713 ne
rect 10141 633 10513 713
tri 10513 633 10593 713 sw
tri 10611 633 10691 713 ne
rect 10691 633 11063 713
tri 11063 633 11143 713 sw
tri 11161 633 11241 713 ne
rect 11241 633 11613 713
tri 11613 633 11693 713 sw
tri 11711 633 11791 713 ne
rect 11791 633 12163 713
tri 12163 633 12243 713 sw
tri 12261 633 12341 713 ne
rect 12341 633 12713 713
tri 12713 633 12793 713 sw
tri 12811 633 12891 713 ne
rect 12891 633 13263 713
tri 13263 633 13343 713 sw
tri 13361 633 13441 713 ne
rect 13441 633 13813 713
tri 13813 633 13893 713 sw
tri 13911 633 13991 713 ne
rect 13991 633 14363 713
tri 14363 633 14443 713 sw
tri 14461 633 14541 713 ne
rect 14541 633 14913 713
tri 14913 633 14993 713 sw
tri 15011 633 15091 713 ne
rect 15091 633 15463 713
tri 15463 633 15543 713 sw
tri 15561 633 15641 713 ne
rect 15641 633 16013 713
tri 16013 633 16093 713 sw
tri 16111 633 16191 713 ne
rect 16191 633 16563 713
tri 16563 633 16643 713 sw
tri 16661 633 16741 713 ne
rect 16741 633 17113 713
tri 17113 633 17193 713 sw
tri 17211 633 17291 713 ne
rect 17291 633 17663 713
tri 17663 633 17743 713 sw
tri 17761 633 17841 713 ne
rect 17841 633 18213 713
tri 18213 633 18293 713 sw
tri 18311 633 18391 713 ne
rect 18391 633 18763 713
tri 18763 633 18843 713 sw
tri 18861 633 18941 713 ne
rect 18941 633 19313 713
tri 19313 633 19393 713 sw
tri 19411 633 19491 713 ne
rect 19491 633 20100 713
rect 261 613 693 633
rect -500 535 163 613
tri 163 535 241 613 sw
tri 261 535 339 613 ne
rect 339 535 693 613
tri 693 535 791 633 sw
tri 791 535 889 633 ne
rect 889 535 1243 633
tri 1243 535 1341 633 sw
tri 1341 535 1439 633 ne
rect 1439 535 1793 633
tri 1793 535 1891 633 sw
tri 1891 535 1989 633 ne
rect 1989 535 2343 633
tri 2343 535 2441 633 sw
tri 2441 535 2539 633 ne
rect 2539 535 2893 633
tri 2893 535 2991 633 sw
tri 2991 535 3089 633 ne
rect 3089 535 3443 633
tri 3443 535 3541 633 sw
tri 3541 535 3639 633 ne
rect 3639 535 3993 633
tri 3993 535 4091 633 sw
tri 4091 535 4189 633 ne
rect 4189 535 4543 633
tri 4543 535 4641 633 sw
tri 4641 535 4739 633 ne
rect 4739 535 5093 633
tri 5093 535 5191 633 sw
tri 5191 535 5289 633 ne
rect 5289 535 5643 633
tri 5643 535 5741 633 sw
tri 5741 535 5839 633 ne
rect 5839 535 6193 633
tri 6193 535 6291 633 sw
tri 6291 535 6389 633 ne
rect 6389 535 6743 633
tri 6743 535 6841 633 sw
tri 6841 535 6939 633 ne
rect 6939 535 7293 633
tri 7293 535 7391 633 sw
tri 7391 535 7489 633 ne
rect 7489 535 7843 633
tri 7843 535 7941 633 sw
tri 7941 535 8039 633 ne
rect 8039 535 8393 633
tri 8393 535 8491 633 sw
tri 8491 535 8589 633 ne
rect 8589 535 8943 633
tri 8943 535 9041 633 sw
tri 9041 535 9139 633 ne
rect 9139 535 9493 633
tri 9493 535 9591 633 sw
tri 9591 535 9689 633 ne
rect 9689 535 10043 633
tri 10043 535 10141 633 sw
tri 10141 535 10239 633 ne
rect 10239 535 10593 633
tri 10593 535 10691 633 sw
tri 10691 535 10789 633 ne
rect 10789 535 11143 633
tri 11143 535 11241 633 sw
tri 11241 535 11339 633 ne
rect 11339 535 11693 633
tri 11693 535 11791 633 sw
tri 11791 535 11889 633 ne
rect 11889 535 12243 633
tri 12243 535 12341 633 sw
tri 12341 535 12439 633 ne
rect 12439 535 12793 633
tri 12793 535 12891 633 sw
tri 12891 535 12989 633 ne
rect 12989 535 13343 633
tri 13343 535 13441 633 sw
tri 13441 535 13539 633 ne
rect 13539 535 13893 633
tri 13893 535 13991 633 sw
tri 13991 535 14089 633 ne
rect 14089 535 14443 633
tri 14443 535 14541 633 sw
tri 14541 535 14639 633 ne
rect 14639 535 14993 633
tri 14993 535 15091 633 sw
tri 15091 535 15189 633 ne
rect 15189 535 15543 633
tri 15543 535 15641 633 sw
tri 15641 535 15739 633 ne
rect 15739 535 16093 633
tri 16093 535 16191 633 sw
tri 16191 535 16289 633 ne
rect 16289 535 16643 633
tri 16643 535 16741 633 sw
tri 16741 535 16839 633 ne
rect 16839 535 17193 633
tri 17193 535 17291 633 sw
tri 17291 535 17389 633 ne
rect 17389 535 17743 633
tri 17743 535 17841 633 sw
tri 17841 535 17939 633 ne
rect 17939 535 18293 633
tri 18293 535 18391 633 sw
tri 18391 535 18489 633 ne
rect 18489 535 18843 633
tri 18843 535 18941 633 sw
tri 18941 535 19039 633 ne
rect 19039 535 19393 633
tri 19393 535 19491 633 sw
tri 19491 535 19589 633 ne
rect 19589 613 20100 633
rect 20200 613 21800 713
rect 19589 535 21800 613
rect -500 487 241 535
rect -500 387 -400 487
rect -300 437 241 487
tri 241 437 339 535 sw
tri 339 437 437 535 ne
rect 437 437 791 535
tri 791 437 889 535 sw
tri 889 437 987 535 ne
rect 987 437 1341 535
tri 1341 437 1439 535 sw
tri 1439 437 1537 535 ne
rect 1537 437 1891 535
tri 1891 437 1989 535 sw
tri 1989 437 2087 535 ne
rect 2087 437 2441 535
tri 2441 437 2539 535 sw
tri 2539 437 2637 535 ne
rect 2637 437 2991 535
tri 2991 437 3089 535 sw
tri 3089 437 3187 535 ne
rect 3187 437 3541 535
tri 3541 437 3639 535 sw
tri 3639 437 3737 535 ne
rect 3737 437 4091 535
tri 4091 437 4189 535 sw
tri 4189 437 4287 535 ne
rect 4287 437 4641 535
tri 4641 437 4739 535 sw
tri 4739 437 4837 535 ne
rect 4837 437 5191 535
tri 5191 437 5289 535 sw
tri 5289 437 5387 535 ne
rect 5387 437 5741 535
tri 5741 437 5839 535 sw
tri 5839 437 5937 535 ne
rect 5937 437 6291 535
tri 6291 437 6389 535 sw
tri 6389 437 6487 535 ne
rect 6487 437 6841 535
tri 6841 437 6939 535 sw
tri 6939 437 7037 535 ne
rect 7037 437 7391 535
tri 7391 437 7489 535 sw
tri 7489 437 7587 535 ne
rect 7587 437 7941 535
tri 7941 437 8039 535 sw
tri 8039 437 8137 535 ne
rect 8137 437 8491 535
tri 8491 437 8589 535 sw
tri 8589 437 8687 535 ne
rect 8687 437 9041 535
tri 9041 437 9139 535 sw
tri 9139 437 9237 535 ne
rect 9237 437 9591 535
tri 9591 437 9689 535 sw
tri 9689 437 9787 535 ne
rect 9787 437 10141 535
tri 10141 437 10239 535 sw
tri 10239 437 10337 535 ne
rect 10337 437 10691 535
tri 10691 437 10789 535 sw
tri 10789 437 10887 535 ne
rect 10887 437 11241 535
tri 11241 437 11339 535 sw
tri 11339 437 11437 535 ne
rect 11437 437 11791 535
tri 11791 437 11889 535 sw
tri 11889 437 11987 535 ne
rect 11987 437 12341 535
tri 12341 437 12439 535 sw
tri 12439 437 12537 535 ne
rect 12537 437 12891 535
tri 12891 437 12989 535 sw
tri 12989 437 13087 535 ne
rect 13087 437 13441 535
tri 13441 437 13539 535 sw
tri 13539 437 13637 535 ne
rect 13637 437 13991 535
tri 13991 437 14089 535 sw
tri 14089 437 14187 535 ne
rect 14187 437 14541 535
tri 14541 437 14639 535 sw
tri 14639 437 14737 535 ne
rect 14737 437 15091 535
tri 15091 437 15189 535 sw
tri 15189 437 15287 535 ne
rect 15287 437 15641 535
tri 15641 437 15739 535 sw
tri 15739 437 15837 535 ne
rect 15837 437 16191 535
tri 16191 437 16289 535 sw
tri 16289 437 16387 535 ne
rect 16387 437 16741 535
tri 16741 437 16839 535 sw
tri 16839 437 16937 535 ne
rect 16937 437 17291 535
tri 17291 437 17389 535 sw
tri 17389 437 17487 535 ne
rect 17487 437 17841 535
tri 17841 437 17939 535 sw
tri 17939 437 18037 535 ne
rect 18037 437 18391 535
tri 18391 437 18489 535 sw
tri 18489 437 18587 535 ne
rect 18587 437 18941 535
tri 18941 437 19039 535 sw
tri 19039 437 19137 535 ne
rect 19137 437 19491 535
tri 19491 437 19589 535 sw
tri 19589 437 19687 535 ne
rect 19687 437 21800 535
rect -300 387 339 437
rect -500 339 339 387
tri 339 339 437 437 sw
tri 437 339 535 437 ne
rect 535 339 889 437
tri 889 339 987 437 sw
tri 987 339 1085 437 ne
rect 1085 339 1439 437
tri 1439 339 1537 437 sw
tri 1537 339 1635 437 ne
rect 1635 339 1989 437
tri 1989 339 2087 437 sw
tri 2087 339 2185 437 ne
rect 2185 339 2539 437
tri 2539 339 2637 437 sw
tri 2637 339 2735 437 ne
rect 2735 339 3089 437
tri 3089 339 3187 437 sw
tri 3187 339 3285 437 ne
rect 3285 339 3639 437
tri 3639 339 3737 437 sw
tri 3737 339 3835 437 ne
rect 3835 339 4189 437
tri 4189 339 4287 437 sw
tri 4287 339 4385 437 ne
rect 4385 339 4739 437
tri 4739 339 4837 437 sw
tri 4837 339 4935 437 ne
rect 4935 339 5289 437
tri 5289 339 5387 437 sw
tri 5387 339 5485 437 ne
rect 5485 339 5839 437
tri 5839 339 5937 437 sw
tri 5937 339 6035 437 ne
rect 6035 339 6389 437
tri 6389 339 6487 437 sw
tri 6487 339 6585 437 ne
rect 6585 339 6939 437
tri 6939 339 7037 437 sw
tri 7037 339 7135 437 ne
rect 7135 339 7489 437
tri 7489 339 7587 437 sw
tri 7587 339 7685 437 ne
rect 7685 339 8039 437
tri 8039 339 8137 437 sw
tri 8137 339 8235 437 ne
rect 8235 339 8589 437
tri 8589 339 8687 437 sw
tri 8687 339 8785 437 ne
rect 8785 339 9139 437
tri 9139 339 9237 437 sw
tri 9237 339 9335 437 ne
rect 9335 339 9689 437
tri 9689 339 9787 437 sw
tri 9787 339 9885 437 ne
rect 9885 339 10239 437
tri 10239 339 10337 437 sw
tri 10337 339 10435 437 ne
rect 10435 339 10789 437
tri 10789 339 10887 437 sw
tri 10887 339 10985 437 ne
rect 10985 339 11339 437
tri 11339 339 11437 437 sw
tri 11437 339 11535 437 ne
rect 11535 339 11889 437
tri 11889 339 11987 437 sw
tri 11987 339 12085 437 ne
rect 12085 339 12439 437
tri 12439 339 12537 437 sw
tri 12537 339 12635 437 ne
rect 12635 339 12989 437
tri 12989 339 13087 437 sw
tri 13087 339 13185 437 ne
rect 13185 339 13539 437
tri 13539 339 13637 437 sw
tri 13637 339 13735 437 ne
rect 13735 339 14089 437
tri 14089 339 14187 437 sw
tri 14187 339 14285 437 ne
rect 14285 339 14639 437
tri 14639 339 14737 437 sw
tri 14737 339 14835 437 ne
rect 14835 339 15189 437
tri 15189 339 15287 437 sw
tri 15287 339 15385 437 ne
rect 15385 339 15739 437
tri 15739 339 15837 437 sw
tri 15837 339 15935 437 ne
rect 15935 339 16289 437
tri 16289 339 16387 437 sw
tri 16387 339 16485 437 ne
rect 16485 339 16839 437
tri 16839 339 16937 437 sw
tri 16937 339 17035 437 ne
rect 17035 339 17389 437
tri 17389 339 17487 437 sw
tri 17487 339 17585 437 ne
rect 17585 339 17939 437
tri 17939 339 18037 437 sw
tri 18037 339 18135 437 ne
rect 18135 339 18489 437
tri 18489 339 18587 437 sw
tri 18587 339 18685 437 ne
rect 18685 339 19039 437
tri 19039 339 19137 437 sw
tri 19137 339 19235 437 ne
rect 19235 339 19589 437
tri 19589 339 19687 437 sw
rect -500 335 437 339
rect -500 215 215 335
rect 335 241 437 335
tri 437 241 535 339 sw
tri 535 241 633 339 ne
rect 633 335 987 339
rect 633 241 765 335
rect 335 215 535 241
rect -500 211 535 215
tri 535 211 565 241 sw
tri 633 211 663 241 ne
rect 663 215 765 241
rect 885 241 987 335
tri 987 241 1085 339 sw
tri 1085 241 1183 339 ne
rect 1183 335 1537 339
rect 1183 241 1315 335
rect 885 215 1085 241
rect 663 211 1085 215
tri 1085 211 1115 241 sw
tri 1183 211 1213 241 ne
rect 1213 215 1315 241
rect 1435 241 1537 335
tri 1537 241 1635 339 sw
tri 1635 241 1733 339 ne
rect 1733 335 2087 339
rect 1733 241 1865 335
rect 1435 215 1635 241
rect 1213 211 1635 215
tri 1635 211 1665 241 sw
tri 1733 211 1763 241 ne
rect 1763 215 1865 241
rect 1985 241 2087 335
tri 2087 241 2185 339 sw
tri 2185 241 2283 339 ne
rect 2283 335 2637 339
rect 2283 241 2415 335
rect 1985 215 2185 241
rect 1763 211 2185 215
tri 2185 211 2215 241 sw
tri 2283 211 2313 241 ne
rect 2313 215 2415 241
rect 2535 241 2637 335
tri 2637 241 2735 339 sw
tri 2735 241 2833 339 ne
rect 2833 335 3187 339
rect 2833 241 2965 335
rect 2535 215 2735 241
rect 2313 211 2735 215
tri 2735 211 2765 241 sw
tri 2833 211 2863 241 ne
rect 2863 215 2965 241
rect 3085 241 3187 335
tri 3187 241 3285 339 sw
tri 3285 241 3383 339 ne
rect 3383 335 3737 339
rect 3383 241 3515 335
rect 3085 215 3285 241
rect 2863 211 3285 215
tri 3285 211 3315 241 sw
tri 3383 211 3413 241 ne
rect 3413 215 3515 241
rect 3635 241 3737 335
tri 3737 241 3835 339 sw
tri 3835 241 3933 339 ne
rect 3933 335 4287 339
rect 3933 241 4065 335
rect 3635 215 3835 241
rect 3413 211 3835 215
tri 3835 211 3865 241 sw
tri 3933 211 3963 241 ne
rect 3963 215 4065 241
rect 4185 241 4287 335
tri 4287 241 4385 339 sw
tri 4385 241 4483 339 ne
rect 4483 335 4837 339
rect 4483 241 4615 335
rect 4185 215 4385 241
rect 3963 211 4385 215
tri 4385 211 4415 241 sw
tri 4483 211 4513 241 ne
rect 4513 215 4615 241
rect 4735 241 4837 335
tri 4837 241 4935 339 sw
tri 4935 241 5033 339 ne
rect 5033 335 5387 339
rect 5033 241 5165 335
rect 4735 215 4935 241
rect 4513 211 4935 215
tri 4935 211 4965 241 sw
tri 5033 211 5063 241 ne
rect 5063 215 5165 241
rect 5285 241 5387 335
tri 5387 241 5485 339 sw
tri 5485 241 5583 339 ne
rect 5583 335 5937 339
rect 5583 241 5715 335
rect 5285 215 5485 241
rect 5063 211 5485 215
tri 5485 211 5515 241 sw
tri 5583 211 5613 241 ne
rect 5613 215 5715 241
rect 5835 241 5937 335
tri 5937 241 6035 339 sw
tri 6035 241 6133 339 ne
rect 6133 335 6487 339
rect 6133 241 6265 335
rect 5835 215 6035 241
rect 5613 211 6035 215
tri 6035 211 6065 241 sw
tri 6133 211 6163 241 ne
rect 6163 215 6265 241
rect 6385 241 6487 335
tri 6487 241 6585 339 sw
tri 6585 241 6683 339 ne
rect 6683 335 7037 339
rect 6683 241 6815 335
rect 6385 215 6585 241
rect 6163 211 6585 215
tri 6585 211 6615 241 sw
tri 6683 211 6713 241 ne
rect 6713 215 6815 241
rect 6935 241 7037 335
tri 7037 241 7135 339 sw
tri 7135 241 7233 339 ne
rect 7233 335 7587 339
rect 7233 241 7365 335
rect 6935 215 7135 241
rect 6713 211 7135 215
tri 7135 211 7165 241 sw
tri 7233 211 7263 241 ne
rect 7263 215 7365 241
rect 7485 241 7587 335
tri 7587 241 7685 339 sw
tri 7685 241 7783 339 ne
rect 7783 335 8137 339
rect 7783 241 7915 335
rect 7485 215 7685 241
rect 7263 211 7685 215
tri 7685 211 7715 241 sw
tri 7783 211 7813 241 ne
rect 7813 215 7915 241
rect 8035 241 8137 335
tri 8137 241 8235 339 sw
tri 8235 241 8333 339 ne
rect 8333 335 8687 339
rect 8333 241 8465 335
rect 8035 215 8235 241
rect 7813 211 8235 215
tri 8235 211 8265 241 sw
tri 8333 211 8363 241 ne
rect 8363 215 8465 241
rect 8585 241 8687 335
tri 8687 241 8785 339 sw
tri 8785 241 8883 339 ne
rect 8883 335 9237 339
rect 8883 241 9015 335
rect 8585 215 8785 241
rect 8363 211 8785 215
tri 8785 211 8815 241 sw
tri 8883 211 8913 241 ne
rect 8913 215 9015 241
rect 9135 241 9237 335
tri 9237 241 9335 339 sw
tri 9335 241 9433 339 ne
rect 9433 335 9787 339
rect 9433 241 9565 335
rect 9135 215 9335 241
rect 8913 211 9335 215
tri 9335 211 9365 241 sw
tri 9433 211 9463 241 ne
rect 9463 215 9565 241
rect 9685 241 9787 335
tri 9787 241 9885 339 sw
tri 9885 241 9983 339 ne
rect 9983 335 10337 339
rect 9983 241 10115 335
rect 9685 215 9885 241
rect 9463 211 9885 215
tri 9885 211 9915 241 sw
tri 9983 211 10013 241 ne
rect 10013 215 10115 241
rect 10235 241 10337 335
tri 10337 241 10435 339 sw
tri 10435 241 10533 339 ne
rect 10533 335 10887 339
rect 10533 241 10665 335
rect 10235 215 10435 241
rect 10013 211 10435 215
tri 10435 211 10465 241 sw
tri 10533 211 10563 241 ne
rect 10563 215 10665 241
rect 10785 241 10887 335
tri 10887 241 10985 339 sw
tri 10985 241 11083 339 ne
rect 11083 335 11437 339
rect 11083 241 11215 335
rect 10785 215 10985 241
rect 10563 211 10985 215
tri 10985 211 11015 241 sw
tri 11083 211 11113 241 ne
rect 11113 215 11215 241
rect 11335 241 11437 335
tri 11437 241 11535 339 sw
tri 11535 241 11633 339 ne
rect 11633 335 11987 339
rect 11633 241 11765 335
rect 11335 215 11535 241
rect 11113 211 11535 215
tri 11535 211 11565 241 sw
tri 11633 211 11663 241 ne
rect 11663 215 11765 241
rect 11885 241 11987 335
tri 11987 241 12085 339 sw
tri 12085 241 12183 339 ne
rect 12183 335 12537 339
rect 12183 241 12315 335
rect 11885 215 12085 241
rect 11663 211 12085 215
tri 12085 211 12115 241 sw
tri 12183 211 12213 241 ne
rect 12213 215 12315 241
rect 12435 241 12537 335
tri 12537 241 12635 339 sw
tri 12635 241 12733 339 ne
rect 12733 335 13087 339
rect 12733 241 12865 335
rect 12435 215 12635 241
rect 12213 211 12635 215
tri 12635 211 12665 241 sw
tri 12733 211 12763 241 ne
rect 12763 215 12865 241
rect 12985 241 13087 335
tri 13087 241 13185 339 sw
tri 13185 241 13283 339 ne
rect 13283 335 13637 339
rect 13283 241 13415 335
rect 12985 215 13185 241
rect 12763 211 13185 215
tri 13185 211 13215 241 sw
tri 13283 211 13313 241 ne
rect 13313 215 13415 241
rect 13535 241 13637 335
tri 13637 241 13735 339 sw
tri 13735 241 13833 339 ne
rect 13833 335 14187 339
rect 13833 241 13965 335
rect 13535 215 13735 241
rect 13313 211 13735 215
tri 13735 211 13765 241 sw
tri 13833 211 13863 241 ne
rect 13863 215 13965 241
rect 14085 241 14187 335
tri 14187 241 14285 339 sw
tri 14285 241 14383 339 ne
rect 14383 335 14737 339
rect 14383 241 14515 335
rect 14085 215 14285 241
rect 13863 211 14285 215
tri 14285 211 14315 241 sw
tri 14383 211 14413 241 ne
rect 14413 215 14515 241
rect 14635 241 14737 335
tri 14737 241 14835 339 sw
tri 14835 241 14933 339 ne
rect 14933 335 15287 339
rect 14933 241 15065 335
rect 14635 215 14835 241
rect 14413 211 14835 215
tri 14835 211 14865 241 sw
tri 14933 211 14963 241 ne
rect 14963 215 15065 241
rect 15185 241 15287 335
tri 15287 241 15385 339 sw
tri 15385 241 15483 339 ne
rect 15483 335 15837 339
rect 15483 241 15615 335
rect 15185 215 15385 241
rect 14963 211 15385 215
tri 15385 211 15415 241 sw
tri 15483 211 15513 241 ne
rect 15513 215 15615 241
rect 15735 241 15837 335
tri 15837 241 15935 339 sw
tri 15935 241 16033 339 ne
rect 16033 335 16387 339
rect 16033 241 16165 335
rect 15735 215 15935 241
rect 15513 211 15935 215
tri 15935 211 15965 241 sw
tri 16033 211 16063 241 ne
rect 16063 215 16165 241
rect 16285 241 16387 335
tri 16387 241 16485 339 sw
tri 16485 241 16583 339 ne
rect 16583 335 16937 339
rect 16583 241 16715 335
rect 16285 215 16485 241
rect 16063 211 16485 215
tri 16485 211 16515 241 sw
tri 16583 211 16613 241 ne
rect 16613 215 16715 241
rect 16835 241 16937 335
tri 16937 241 17035 339 sw
tri 17035 241 17133 339 ne
rect 17133 335 17487 339
rect 17133 241 17265 335
rect 16835 215 17035 241
rect 16613 211 17035 215
tri 17035 211 17065 241 sw
tri 17133 211 17163 241 ne
rect 17163 215 17265 241
rect 17385 241 17487 335
tri 17487 241 17585 339 sw
tri 17585 241 17683 339 ne
rect 17683 335 18037 339
rect 17683 241 17815 335
rect 17385 215 17585 241
rect 17163 211 17585 215
tri 17585 211 17615 241 sw
tri 17683 211 17713 241 ne
rect 17713 215 17815 241
rect 17935 241 18037 335
tri 18037 241 18135 339 sw
tri 18135 241 18233 339 ne
rect 18233 335 18587 339
rect 18233 241 18365 335
rect 17935 215 18135 241
rect 17713 211 18135 215
tri 18135 211 18165 241 sw
tri 18233 211 18263 241 ne
rect 18263 215 18365 241
rect 18485 241 18587 335
tri 18587 241 18685 339 sw
tri 18685 241 18783 339 ne
rect 18783 335 19137 339
rect 18783 241 18915 335
rect 18485 215 18685 241
rect 18263 211 18685 215
tri 18685 211 18715 241 sw
tri 18783 211 18813 241 ne
rect 18813 215 18915 241
rect 19035 241 19137 335
tri 19137 241 19235 339 sw
tri 19235 241 19333 339 ne
rect 19333 335 20300 339
rect 19333 241 19465 335
rect 19035 215 19235 241
rect 18813 211 19235 215
tri 19235 211 19265 241 sw
tri 19333 211 19363 241 ne
rect 19363 215 19465 241
rect 19585 215 20300 335
rect 19363 211 20300 215
tri 113 113 211 211 ne
rect 211 113 565 211
tri 565 113 663 211 sw
tri 663 113 761 211 ne
rect 761 113 1115 211
tri 1115 113 1213 211 sw
tri 1213 113 1311 211 ne
rect 1311 113 1665 211
tri 1665 113 1763 211 sw
tri 1763 113 1861 211 ne
rect 1861 113 2215 211
tri 2215 113 2313 211 sw
tri 2313 113 2411 211 ne
rect 2411 113 2765 211
tri 2765 113 2863 211 sw
tri 2863 113 2961 211 ne
rect 2961 113 3315 211
tri 3315 113 3413 211 sw
tri 3413 113 3511 211 ne
rect 3511 113 3865 211
tri 3865 113 3963 211 sw
tri 3963 113 4061 211 ne
rect 4061 113 4415 211
tri 4415 113 4513 211 sw
tri 4513 113 4611 211 ne
rect 4611 113 4965 211
tri 4965 113 5063 211 sw
tri 5063 113 5161 211 ne
rect 5161 113 5515 211
tri 5515 113 5613 211 sw
tri 5613 113 5711 211 ne
rect 5711 113 6065 211
tri 6065 113 6163 211 sw
tri 6163 113 6261 211 ne
rect 6261 113 6615 211
tri 6615 113 6713 211 sw
tri 6713 113 6811 211 ne
rect 6811 113 7165 211
tri 7165 113 7263 211 sw
tri 7263 113 7361 211 ne
rect 7361 113 7715 211
tri 7715 113 7813 211 sw
tri 7813 113 7911 211 ne
rect 7911 113 8265 211
tri 8265 113 8363 211 sw
tri 8363 113 8461 211 ne
rect 8461 113 8815 211
tri 8815 113 8913 211 sw
tri 8913 113 9011 211 ne
rect 9011 113 9365 211
tri 9365 113 9463 211 sw
tri 9463 113 9561 211 ne
rect 9561 113 9915 211
tri 9915 113 10013 211 sw
tri 10013 113 10111 211 ne
rect 10111 113 10465 211
tri 10465 113 10563 211 sw
tri 10563 113 10661 211 ne
rect 10661 113 11015 211
tri 11015 113 11113 211 sw
tri 11113 113 11211 211 ne
rect 11211 113 11565 211
tri 11565 113 11663 211 sw
tri 11663 113 11761 211 ne
rect 11761 113 12115 211
tri 12115 113 12213 211 sw
tri 12213 113 12311 211 ne
rect 12311 113 12665 211
tri 12665 113 12763 211 sw
tri 12763 113 12861 211 ne
rect 12861 113 13215 211
tri 13215 113 13313 211 sw
tri 13313 113 13411 211 ne
rect 13411 113 13765 211
tri 13765 113 13863 211 sw
tri 13863 113 13961 211 ne
rect 13961 113 14315 211
tri 14315 113 14413 211 sw
tri 14413 113 14511 211 ne
rect 14511 113 14865 211
tri 14865 113 14963 211 sw
tri 14963 113 15061 211 ne
rect 15061 113 15415 211
tri 15415 113 15513 211 sw
tri 15513 113 15611 211 ne
rect 15611 113 15965 211
tri 15965 113 16063 211 sw
tri 16063 113 16161 211 ne
rect 16161 113 16515 211
tri 16515 113 16613 211 sw
tri 16613 113 16711 211 ne
rect 16711 113 17065 211
tri 17065 113 17163 211 sw
tri 17163 113 17261 211 ne
rect 17261 113 17615 211
tri 17615 113 17713 211 sw
tri 17713 113 17811 211 ne
rect 17811 113 18165 211
tri 18165 113 18263 211 sw
tri 18263 113 18361 211 ne
rect 18361 113 18715 211
tri 18715 113 18813 211 sw
tri 18813 113 18911 211 ne
rect 18911 113 19265 211
tri 19265 113 19363 211 sw
tri 19363 113 19461 211 ne
rect 211 -300 663 113
rect 211 -400 387 -300
rect 487 -400 663 -300
rect 211 -1000 663 -400
rect 761 -500 1213 113
rect 1311 -300 1763 113
rect 1311 -400 1487 -300
rect 1587 -400 1763 -300
rect 1311 -1000 1763 -400
rect 1861 -500 2313 113
rect 2411 -300 2863 113
rect 2411 -400 2587 -300
rect 2687 -400 2863 -300
rect 2411 -1000 2863 -400
rect 2961 -500 3413 113
rect 3511 -300 3963 113
rect 3511 -400 3687 -300
rect 3787 -400 3963 -300
rect 3511 -1000 3963 -400
rect 4061 -500 4513 113
rect 4611 -300 5063 113
rect 4611 -400 4787 -300
rect 4887 -400 5063 -300
rect 4611 -1000 5063 -400
rect 5161 -500 5613 113
rect 5711 -300 6163 113
rect 5711 -400 5887 -300
rect 5987 -400 6163 -300
rect 5711 -1000 6163 -400
rect 6261 -500 6713 113
rect 6811 -300 7263 113
rect 6811 -400 6987 -300
rect 7087 -400 7263 -300
rect 6811 -1000 7263 -400
rect 7361 -500 7813 113
rect 7911 -300 8363 113
rect 7911 -400 8087 -300
rect 8187 -400 8363 -300
rect 7911 -1000 8363 -400
rect 8461 -500 8913 113
rect 9011 -300 9463 113
rect 9011 -400 9187 -300
rect 9287 -400 9463 -300
rect 9011 -1000 9463 -400
rect 9561 -500 10013 113
rect 10111 -300 10563 113
rect 10111 -400 10287 -300
rect 10387 -400 10563 -300
rect 10111 -1000 10563 -400
rect 10661 -500 11113 113
rect 11211 -300 11663 113
rect 11211 -400 11387 -300
rect 11487 -400 11663 -300
rect 11211 -1000 11663 -400
rect 11761 -500 12213 113
rect 12311 -300 12763 113
rect 12311 -400 12487 -300
rect 12587 -400 12763 -300
rect 12311 -1000 12763 -400
rect 12861 -500 13313 113
rect 13411 -300 13863 113
rect 13411 -400 13587 -300
rect 13687 -400 13863 -300
rect 13411 -1000 13863 -400
rect 13961 -500 14413 113
rect 14511 -300 14963 113
rect 14511 -400 14687 -300
rect 14787 -400 14963 -300
rect 14511 -1000 14963 -400
rect 15061 -500 15513 113
rect 15611 -300 16063 113
rect 15611 -400 15787 -300
rect 15887 -400 16063 -300
rect 15611 -1000 16063 -400
rect 16161 -500 16613 113
rect 16711 -300 17163 113
rect 16711 -400 16887 -300
rect 16987 -400 17163 -300
rect 16711 -1000 17163 -400
rect 17261 -500 17713 113
rect 17811 -300 18263 113
rect 17811 -400 17987 -300
rect 18087 -400 18263 -300
rect 17811 -1000 18263 -400
rect 18361 -500 18813 113
rect 18911 -300 19363 113
rect 18911 -400 19087 -300
rect 19187 -400 19363 -300
rect 18911 -1000 19363 -400
rect 19461 -113 20300 211
rect 19461 -500 19913 -113
rect 20800 -1000 21800 437
rect 0 -2000 21800 -1000
<< via4 >>
rect 215 19465 335 19585
rect 765 19465 885 19585
rect 1315 19465 1435 19585
rect 1865 19465 1985 19585
rect 2415 19465 2535 19585
rect 2965 19465 3085 19585
rect 3515 19465 3635 19585
rect 4065 19465 4185 19585
rect 4615 19465 4735 19585
rect 5165 19465 5285 19585
rect 5715 19465 5835 19585
rect 6265 19465 6385 19585
rect 6815 19465 6935 19585
rect 7365 19465 7485 19585
rect 7915 19465 8035 19585
rect 8465 19465 8585 19585
rect 9015 19465 9135 19585
rect 9565 19465 9685 19585
rect 10115 19465 10235 19585
rect 10665 19465 10785 19585
rect 11215 19465 11335 19585
rect 11765 19465 11885 19585
rect 12315 19465 12435 19585
rect 12865 19465 12985 19585
rect 13415 19465 13535 19585
rect 13965 19465 14085 19585
rect 14515 19465 14635 19585
rect 15065 19465 15185 19585
rect 15615 19465 15735 19585
rect 16165 19465 16285 19585
rect 16715 19465 16835 19585
rect 17265 19465 17385 19585
rect 17815 19465 17935 19585
rect 18365 19465 18485 19585
rect 18915 19465 19035 19585
rect 19465 19465 19585 19585
rect 215 18915 335 19035
rect 19465 18915 19585 19035
rect 215 18365 335 18485
rect 19465 18365 19585 18485
rect 215 17815 335 17935
rect 19465 17815 19585 17935
rect 215 17265 335 17385
rect 19465 17265 19585 17385
rect 215 16715 335 16835
rect 19465 16715 19585 16835
rect 215 16165 335 16285
rect 19465 16165 19585 16285
rect 215 15615 335 15735
rect 19465 15615 19585 15735
rect 215 15065 335 15185
rect 19465 15065 19585 15185
rect 215 14515 335 14635
rect 19465 14515 19585 14635
rect 215 13965 335 14085
rect 19465 13965 19585 14085
rect 215 13415 335 13535
rect 19465 13415 19585 13535
rect 215 12865 335 12985
rect 19465 12865 19585 12985
rect 215 12315 335 12435
rect 19465 12315 19585 12435
rect 215 11765 335 11885
rect 19465 11765 19585 11885
rect 215 11215 335 11335
rect 19465 11215 19585 11335
rect 215 10665 335 10785
rect 19465 10665 19585 10785
rect 215 10115 335 10235
rect 19465 10115 19585 10235
rect 215 9565 335 9685
rect 19465 9565 19585 9685
rect 215 9015 335 9135
rect 19465 9015 19585 9135
rect 215 8465 335 8585
rect 19465 8465 19585 8585
rect 215 7915 335 8035
rect 19465 7915 19585 8035
rect 215 7365 335 7485
rect 19465 7365 19585 7485
rect 215 6815 335 6935
rect 19465 6815 19585 6935
rect 215 6265 335 6385
rect 19465 6265 19585 6385
rect 215 5715 335 5835
rect 19465 5715 19585 5835
rect 215 5165 335 5285
rect 19465 5165 19585 5285
rect 215 4615 335 4735
rect 19465 4615 19585 4735
rect 215 4065 335 4185
rect 19465 4065 19585 4185
rect 215 3515 335 3635
rect 19465 3515 19585 3635
rect 215 2965 335 3085
rect 19465 2965 19585 3085
rect 215 2415 335 2535
rect 19465 2415 19585 2535
rect 215 1865 335 1985
rect 19465 1865 19585 1985
rect 215 1315 335 1435
rect 19465 1315 19585 1435
rect 215 765 335 885
rect 19465 765 19585 885
rect 215 215 335 335
rect 765 215 885 335
rect 1315 215 1435 335
rect 1865 215 1985 335
rect 2415 215 2535 335
rect 2965 215 3085 335
rect 3515 215 3635 335
rect 4065 215 4185 335
rect 4615 215 4735 335
rect 5165 215 5285 335
rect 5715 215 5835 335
rect 6265 215 6385 335
rect 6815 215 6935 335
rect 7365 215 7485 335
rect 7915 215 8035 335
rect 8465 215 8585 335
rect 9015 215 9135 335
rect 9565 215 9685 335
rect 10115 215 10235 335
rect 10665 215 10785 335
rect 11215 215 11335 335
rect 11765 215 11885 335
rect 12315 215 12435 335
rect 12865 215 12985 335
rect 13415 215 13535 335
rect 13965 215 14085 335
rect 14515 215 14635 335
rect 15065 215 15185 335
rect 15615 215 15735 335
rect 16165 215 16285 335
rect 16715 215 16835 335
rect 17265 215 17385 335
rect 17815 215 17935 335
rect 18365 215 18485 335
rect 18915 215 19035 335
rect 19465 215 19585 335
<< metal5 >>
rect -2000 20800 19800 21800
rect -2000 19878 -1000 20800
rect -78 19878 233 20800
rect -2000 19585 233 19878
tri 233 19585 371 19723 sw
rect 472 19722 783 20300
tri 472 19585 609 19722 ne
rect 609 19585 783 19722
tri 783 19585 921 19723 sw
rect 1022 19722 1333 20800
tri 1022 19585 1159 19722 ne
rect 1159 19585 1333 19722
tri 1333 19585 1471 19723 sw
rect 1572 19722 1883 20300
tri 1572 19585 1709 19722 ne
rect 1709 19585 1883 19722
tri 1883 19585 2021 19723 sw
rect 2122 19722 2433 20800
tri 2122 19585 2259 19722 ne
rect 2259 19585 2433 19722
tri 2433 19585 2571 19723 sw
rect 2672 19722 2983 20300
tri 2672 19585 2809 19722 ne
rect 2809 19585 2983 19722
tri 2983 19585 3121 19723 sw
rect 3222 19722 3533 20800
tri 3222 19585 3359 19722 ne
rect 3359 19585 3533 19722
tri 3533 19585 3671 19723 sw
rect 3772 19722 4083 20300
tri 3772 19585 3909 19722 ne
rect 3909 19585 4083 19722
tri 4083 19585 4221 19723 sw
rect 4322 19722 4633 20800
tri 4322 19585 4459 19722 ne
rect 4459 19585 4633 19722
tri 4633 19585 4771 19723 sw
rect 4872 19722 5183 20300
tri 4872 19585 5009 19722 ne
rect 5009 19585 5183 19722
tri 5183 19585 5321 19723 sw
rect 5422 19722 5733 20800
tri 5422 19585 5559 19722 ne
rect 5559 19585 5733 19722
tri 5733 19585 5871 19723 sw
rect 5972 19722 6283 20300
tri 5972 19585 6109 19722 ne
rect 6109 19585 6283 19722
tri 6283 19585 6421 19723 sw
rect 6522 19722 6833 20800
tri 6522 19585 6659 19722 ne
rect 6659 19585 6833 19722
tri 6833 19585 6971 19723 sw
rect 7072 19722 7383 20300
tri 7072 19585 7209 19722 ne
rect 7209 19585 7383 19722
tri 7383 19585 7521 19723 sw
rect 7622 19722 7933 20800
tri 7622 19585 7759 19722 ne
rect 7759 19585 7933 19722
tri 7933 19585 8071 19723 sw
rect 8172 19722 8483 20300
tri 8172 19585 8309 19722 ne
rect 8309 19585 8483 19722
tri 8483 19585 8621 19723 sw
rect 8722 19722 9033 20800
tri 8722 19585 8859 19722 ne
rect 8859 19585 9033 19722
tri 9033 19585 9171 19723 sw
rect 9272 19722 9583 20300
tri 9272 19585 9409 19722 ne
rect 9409 19585 9583 19722
tri 9583 19585 9721 19723 sw
rect 9822 19722 10133 20800
tri 9822 19585 9959 19722 ne
rect 9959 19585 10133 19722
tri 10133 19585 10271 19723 sw
rect 10372 19722 10683 20300
tri 10372 19585 10509 19722 ne
rect 10509 19585 10683 19722
tri 10683 19585 10821 19723 sw
rect 10922 19722 11233 20800
tri 10922 19585 11059 19722 ne
rect 11059 19585 11233 19722
tri 11233 19585 11371 19723 sw
rect 11472 19722 11783 20300
tri 11472 19585 11609 19722 ne
rect 11609 19585 11783 19722
tri 11783 19585 11921 19723 sw
rect 12022 19722 12333 20800
tri 12022 19585 12159 19722 ne
rect 12159 19585 12333 19722
tri 12333 19585 12471 19723 sw
rect 12572 19722 12883 20300
tri 12572 19585 12709 19722 ne
rect 12709 19585 12883 19722
tri 12883 19585 13021 19723 sw
rect 13122 19722 13433 20800
tri 13122 19585 13259 19722 ne
rect 13259 19585 13433 19722
tri 13433 19585 13571 19723 sw
rect 13672 19722 13983 20300
tri 13672 19585 13809 19722 ne
rect 13809 19585 13983 19722
tri 13983 19585 14121 19723 sw
rect 14222 19722 14533 20800
tri 14222 19585 14359 19722 ne
rect 14359 19585 14533 19722
tri 14533 19585 14671 19723 sw
rect 14772 19722 15083 20300
tri 14772 19585 14909 19722 ne
rect 14909 19585 15083 19722
tri 15083 19585 15221 19723 sw
rect 15322 19722 15633 20800
tri 15322 19585 15459 19722 ne
rect 15459 19585 15633 19722
tri 15633 19585 15771 19723 sw
rect 15872 19722 16183 20300
tri 15872 19585 16009 19722 ne
rect 16009 19585 16183 19722
tri 16183 19585 16321 19723 sw
rect 16422 19722 16733 20800
tri 16422 19585 16559 19722 ne
rect 16559 19585 16733 19722
tri 16733 19585 16871 19723 sw
rect 16972 19722 17283 20300
tri 16972 19585 17109 19722 ne
rect 17109 19585 17283 19722
tri 17283 19585 17421 19723 sw
rect 17522 19722 17833 20800
tri 17522 19585 17659 19722 ne
rect 17659 19585 17833 19722
tri 17833 19585 17971 19723 sw
rect 18072 19722 18383 20300
tri 18072 19585 18209 19722 ne
rect 18209 19585 18383 19722
tri 18383 19585 18521 19723 sw
rect 18622 19722 18933 20800
tri 18622 19585 18759 19722 ne
rect 18759 19585 18933 19722
tri 18933 19585 19071 19723 sw
rect 19172 19722 19483 20300
tri 19172 19585 19309 19722 ne
rect 19309 19585 19483 19722
tri 19483 19585 19621 19723 sw
rect -2000 19567 215 19585
rect -2000 18778 -1000 19567
tri 77 19465 179 19567 ne
rect 179 19465 215 19567
rect 335 19465 371 19585
tri 179 19328 316 19465 ne
rect 316 19410 371 19465
tri 371 19410 546 19585 sw
tri 609 19465 729 19585 ne
rect 729 19465 765 19585
rect 885 19465 921 19585
rect 316 19328 546 19410
tri 546 19328 628 19410 sw
tri 729 19328 866 19465 ne
rect 866 19410 921 19465
tri 921 19410 1096 19585 sw
tri 1159 19465 1279 19585 ne
rect 1279 19465 1315 19585
rect 1435 19465 1471 19585
rect 866 19328 1096 19410
tri 1096 19328 1178 19410 sw
tri 1279 19328 1416 19465 ne
rect 1416 19410 1471 19465
tri 1471 19410 1646 19585 sw
tri 1709 19465 1829 19585 ne
rect 1829 19465 1865 19585
rect 1985 19465 2021 19585
rect 1416 19328 1646 19410
tri 1646 19328 1728 19410 sw
tri 1829 19328 1966 19465 ne
rect 1966 19410 2021 19465
tri 2021 19410 2196 19585 sw
tri 2259 19465 2379 19585 ne
rect 2379 19465 2415 19585
rect 2535 19465 2571 19585
rect 1966 19328 2196 19410
tri 2196 19328 2278 19410 sw
tri 2379 19328 2516 19465 ne
rect 2516 19410 2571 19465
tri 2571 19410 2746 19585 sw
tri 2809 19465 2929 19585 ne
rect 2929 19465 2965 19585
rect 3085 19465 3121 19585
rect 2516 19328 2746 19410
tri 2746 19328 2828 19410 sw
tri 2929 19328 3066 19465 ne
rect 3066 19410 3121 19465
tri 3121 19410 3296 19585 sw
tri 3359 19465 3479 19585 ne
rect 3479 19465 3515 19585
rect 3635 19465 3671 19585
rect 3066 19328 3296 19410
tri 3296 19328 3378 19410 sw
tri 3479 19328 3616 19465 ne
rect 3616 19410 3671 19465
tri 3671 19410 3846 19585 sw
tri 3909 19465 4029 19585 ne
rect 4029 19465 4065 19585
rect 4185 19465 4221 19585
rect 3616 19328 3846 19410
tri 3846 19328 3928 19410 sw
tri 4029 19328 4166 19465 ne
rect 4166 19410 4221 19465
tri 4221 19410 4396 19585 sw
tri 4459 19465 4579 19585 ne
rect 4579 19465 4615 19585
rect 4735 19465 4771 19585
rect 4166 19328 4396 19410
tri 4396 19328 4478 19410 sw
tri 4579 19328 4716 19465 ne
rect 4716 19410 4771 19465
tri 4771 19410 4946 19585 sw
tri 5009 19465 5129 19585 ne
rect 5129 19465 5165 19585
rect 5285 19465 5321 19585
rect 4716 19328 4946 19410
tri 4946 19328 5028 19410 sw
tri 5129 19328 5266 19465 ne
rect 5266 19410 5321 19465
tri 5321 19410 5496 19585 sw
tri 5559 19465 5679 19585 ne
rect 5679 19465 5715 19585
rect 5835 19465 5871 19585
rect 5266 19328 5496 19410
tri 5496 19328 5578 19410 sw
tri 5679 19328 5816 19465 ne
rect 5816 19410 5871 19465
tri 5871 19410 6046 19585 sw
tri 6109 19465 6229 19585 ne
rect 6229 19465 6265 19585
rect 6385 19465 6421 19585
rect 5816 19328 6046 19410
tri 6046 19328 6128 19410 sw
tri 6229 19328 6366 19465 ne
rect 6366 19410 6421 19465
tri 6421 19410 6596 19585 sw
tri 6659 19465 6779 19585 ne
rect 6779 19465 6815 19585
rect 6935 19465 6971 19585
rect 6366 19328 6596 19410
tri 6596 19328 6678 19410 sw
tri 6779 19328 6916 19465 ne
rect 6916 19410 6971 19465
tri 6971 19410 7146 19585 sw
tri 7209 19465 7329 19585 ne
rect 7329 19465 7365 19585
rect 7485 19465 7521 19585
rect 6916 19328 7146 19410
tri 7146 19328 7228 19410 sw
tri 7329 19328 7466 19465 ne
rect 7466 19410 7521 19465
tri 7521 19410 7696 19585 sw
tri 7759 19465 7879 19585 ne
rect 7879 19465 7915 19585
rect 8035 19465 8071 19585
rect 7466 19328 7696 19410
tri 7696 19328 7778 19410 sw
tri 7879 19328 8016 19465 ne
rect 8016 19410 8071 19465
tri 8071 19410 8246 19585 sw
tri 8309 19465 8429 19585 ne
rect 8429 19465 8465 19585
rect 8585 19465 8621 19585
rect 8016 19328 8246 19410
tri 8246 19328 8328 19410 sw
tri 8429 19328 8566 19465 ne
rect 8566 19410 8621 19465
tri 8621 19410 8796 19585 sw
tri 8859 19465 8979 19585 ne
rect 8979 19465 9015 19585
rect 9135 19465 9171 19585
rect 8566 19328 8796 19410
tri 8796 19328 8878 19410 sw
tri 8979 19328 9116 19465 ne
rect 9116 19410 9171 19465
tri 9171 19410 9346 19585 sw
tri 9409 19465 9529 19585 ne
rect 9529 19465 9565 19585
rect 9685 19465 9721 19585
rect 9116 19328 9346 19410
tri 9346 19328 9428 19410 sw
tri 9529 19328 9666 19465 ne
rect 9666 19410 9721 19465
tri 9721 19410 9896 19585 sw
tri 9959 19465 10079 19585 ne
rect 10079 19465 10115 19585
rect 10235 19465 10271 19585
rect 9666 19328 9896 19410
tri 9896 19328 9978 19410 sw
tri 10079 19328 10216 19465 ne
rect 10216 19410 10271 19465
tri 10271 19410 10446 19585 sw
tri 10509 19465 10629 19585 ne
rect 10629 19465 10665 19585
rect 10785 19465 10821 19585
rect 10216 19328 10446 19410
tri 10446 19328 10528 19410 sw
tri 10629 19328 10766 19465 ne
rect 10766 19410 10821 19465
tri 10821 19410 10996 19585 sw
tri 11059 19465 11179 19585 ne
rect 11179 19465 11215 19585
rect 11335 19465 11371 19585
rect 10766 19328 10996 19410
tri 10996 19328 11078 19410 sw
tri 11179 19328 11316 19465 ne
rect 11316 19410 11371 19465
tri 11371 19410 11546 19585 sw
tri 11609 19465 11729 19585 ne
rect 11729 19465 11765 19585
rect 11885 19465 11921 19585
rect 11316 19328 11546 19410
tri 11546 19328 11628 19410 sw
tri 11729 19328 11866 19465 ne
rect 11866 19410 11921 19465
tri 11921 19410 12096 19585 sw
tri 12159 19465 12279 19585 ne
rect 12279 19465 12315 19585
rect 12435 19465 12471 19585
rect 11866 19328 12096 19410
tri 12096 19328 12178 19410 sw
tri 12279 19328 12416 19465 ne
rect 12416 19410 12471 19465
tri 12471 19410 12646 19585 sw
tri 12709 19465 12829 19585 ne
rect 12829 19465 12865 19585
rect 12985 19465 13021 19585
rect 12416 19328 12646 19410
tri 12646 19328 12728 19410 sw
tri 12829 19328 12966 19465 ne
rect 12966 19410 13021 19465
tri 13021 19410 13196 19585 sw
tri 13259 19465 13379 19585 ne
rect 13379 19465 13415 19585
rect 13535 19465 13571 19585
rect 12966 19328 13196 19410
tri 13196 19328 13278 19410 sw
tri 13379 19328 13516 19465 ne
rect 13516 19410 13571 19465
tri 13571 19410 13746 19585 sw
tri 13809 19465 13929 19585 ne
rect 13929 19465 13965 19585
rect 14085 19465 14121 19585
rect 13516 19328 13746 19410
tri 13746 19328 13828 19410 sw
tri 13929 19328 14066 19465 ne
rect 14066 19410 14121 19465
tri 14121 19410 14296 19585 sw
tri 14359 19465 14479 19585 ne
rect 14479 19465 14515 19585
rect 14635 19465 14671 19585
rect 14066 19328 14296 19410
tri 14296 19328 14378 19410 sw
tri 14479 19328 14616 19465 ne
rect 14616 19410 14671 19465
tri 14671 19410 14846 19585 sw
tri 14909 19465 15029 19585 ne
rect 15029 19465 15065 19585
rect 15185 19465 15221 19585
rect 14616 19328 14846 19410
tri 14846 19328 14928 19410 sw
tri 15029 19328 15166 19465 ne
rect 15166 19410 15221 19465
tri 15221 19410 15396 19585 sw
tri 15459 19465 15579 19585 ne
rect 15579 19465 15615 19585
rect 15735 19465 15771 19585
rect 15166 19328 15396 19410
tri 15396 19328 15478 19410 sw
tri 15579 19328 15716 19465 ne
rect 15716 19410 15771 19465
tri 15771 19410 15946 19585 sw
tri 16009 19465 16129 19585 ne
rect 16129 19465 16165 19585
rect 16285 19465 16321 19585
rect 15716 19328 15946 19410
tri 15946 19328 16028 19410 sw
tri 16129 19328 16266 19465 ne
rect 16266 19410 16321 19465
tri 16321 19410 16496 19585 sw
tri 16559 19465 16679 19585 ne
rect 16679 19465 16715 19585
rect 16835 19465 16871 19585
rect 16266 19328 16496 19410
tri 16496 19328 16578 19410 sw
tri 16679 19328 16816 19465 ne
rect 16816 19410 16871 19465
tri 16871 19410 17046 19585 sw
tri 17109 19465 17229 19585 ne
rect 17229 19465 17265 19585
rect 17385 19465 17421 19585
rect 16816 19328 17046 19410
tri 17046 19328 17128 19410 sw
tri 17229 19328 17366 19465 ne
rect 17366 19410 17421 19465
tri 17421 19410 17596 19585 sw
tri 17659 19465 17779 19585 ne
rect 17779 19465 17815 19585
rect 17935 19465 17971 19585
rect 17366 19328 17596 19410
tri 17596 19328 17678 19410 sw
tri 17779 19328 17916 19465 ne
rect 17916 19410 17971 19465
tri 17971 19410 18146 19585 sw
tri 18209 19465 18329 19585 ne
rect 18329 19465 18365 19585
rect 18485 19465 18521 19585
rect 17916 19328 18146 19410
tri 18146 19328 18228 19410 sw
tri 18329 19328 18466 19465 ne
rect 18466 19410 18521 19465
tri 18521 19410 18696 19585 sw
tri 18759 19465 18879 19585 ne
rect 18879 19465 18915 19585
rect 19035 19465 19071 19585
rect 18466 19328 18696 19410
tri 18696 19328 18778 19410 sw
tri 18879 19328 19016 19465 ne
rect 19016 19410 19071 19465
tri 19071 19410 19246 19585 sw
tri 19309 19465 19429 19585 ne
rect 19429 19465 19465 19585
rect 19585 19483 19621 19585
tri 19621 19483 19723 19585 sw
rect 20800 19483 21800 19800
rect 19585 19465 21800 19483
rect 19016 19328 19246 19410
tri 19246 19328 19328 19410 sw
tri 19429 19328 19566 19465 ne
rect 19566 19328 21800 19465
rect -500 19172 78 19328
tri 78 19172 234 19328 sw
tri 316 19172 472 19328 ne
rect 472 19172 628 19328
tri 628 19172 784 19328 sw
tri 866 19172 1022 19328 ne
rect 1022 19172 1178 19328
tri 1178 19172 1334 19328 sw
tri 1416 19172 1572 19328 ne
rect 1572 19172 1728 19328
tri 1728 19172 1884 19328 sw
tri 1966 19172 2122 19328 ne
rect 2122 19172 2278 19328
tri 2278 19172 2434 19328 sw
tri 2516 19172 2672 19328 ne
rect 2672 19172 2828 19328
tri 2828 19172 2984 19328 sw
tri 3066 19172 3222 19328 ne
rect 3222 19172 3378 19328
tri 3378 19172 3534 19328 sw
tri 3616 19172 3772 19328 ne
rect 3772 19172 3928 19328
tri 3928 19172 4084 19328 sw
tri 4166 19172 4322 19328 ne
rect 4322 19172 4478 19328
tri 4478 19172 4634 19328 sw
tri 4716 19172 4872 19328 ne
rect 4872 19172 5028 19328
tri 5028 19172 5184 19328 sw
tri 5266 19172 5422 19328 ne
rect 5422 19172 5578 19328
tri 5578 19172 5734 19328 sw
tri 5816 19172 5972 19328 ne
rect 5972 19172 6128 19328
tri 6128 19172 6284 19328 sw
tri 6366 19172 6522 19328 ne
rect 6522 19172 6678 19328
tri 6678 19172 6834 19328 sw
tri 6916 19172 7072 19328 ne
rect 7072 19172 7228 19328
tri 7228 19172 7384 19328 sw
tri 7466 19172 7622 19328 ne
rect 7622 19172 7778 19328
tri 7778 19172 7934 19328 sw
tri 8016 19172 8172 19328 ne
rect 8172 19172 8328 19328
tri 8328 19172 8484 19328 sw
tri 8566 19172 8722 19328 ne
rect 8722 19172 8878 19328
tri 8878 19172 9034 19328 sw
tri 9116 19172 9272 19328 ne
rect 9272 19172 9428 19328
tri 9428 19172 9584 19328 sw
tri 9666 19172 9822 19328 ne
rect 9822 19172 9978 19328
tri 9978 19172 10134 19328 sw
tri 10216 19172 10372 19328 ne
rect 10372 19172 10528 19328
tri 10528 19172 10684 19328 sw
tri 10766 19172 10922 19328 ne
rect 10922 19172 11078 19328
tri 11078 19172 11234 19328 sw
tri 11316 19172 11472 19328 ne
rect 11472 19172 11628 19328
tri 11628 19172 11784 19328 sw
tri 11866 19172 12022 19328 ne
rect 12022 19172 12178 19328
tri 12178 19172 12334 19328 sw
tri 12416 19172 12572 19328 ne
rect 12572 19172 12728 19328
tri 12728 19172 12884 19328 sw
tri 12966 19172 13122 19328 ne
rect 13122 19172 13278 19328
tri 13278 19172 13434 19328 sw
tri 13516 19172 13672 19328 ne
rect 13672 19172 13828 19328
tri 13828 19172 13984 19328 sw
tri 14066 19172 14222 19328 ne
rect 14222 19172 14378 19328
tri 14378 19172 14534 19328 sw
tri 14616 19172 14772 19328 ne
rect 14772 19172 14928 19328
tri 14928 19172 15084 19328 sw
tri 15166 19172 15322 19328 ne
rect 15322 19172 15478 19328
tri 15478 19172 15634 19328 sw
tri 15716 19172 15872 19328 ne
rect 15872 19172 16028 19328
tri 16028 19172 16184 19328 sw
tri 16266 19172 16422 19328 ne
rect 16422 19172 16578 19328
tri 16578 19172 16734 19328 sw
tri 16816 19172 16972 19328 ne
rect 16972 19172 17128 19328
tri 17128 19172 17284 19328 sw
tri 17366 19172 17522 19328 ne
rect 17522 19172 17678 19328
tri 17678 19172 17834 19328 sw
tri 17916 19172 18072 19328 ne
rect 18072 19172 18228 19328
tri 18228 19172 18384 19328 sw
tri 18466 19172 18622 19328 ne
rect 18622 19172 18778 19328
tri 18778 19172 18934 19328 sw
tri 19016 19172 19172 19328 ne
rect 19172 19172 19328 19328
tri 19328 19172 19484 19328 sw
tri 19566 19172 19722 19328 ne
rect 19722 19172 21800 19328
rect -500 19035 234 19172
tri 234 19035 371 19172 sw
tri 472 19035 609 19172 ne
rect 609 19035 784 19172
tri 784 19035 921 19172 sw
tri 1022 19035 1159 19172 ne
rect 1159 19035 1334 19172
tri 1334 19035 1471 19172 sw
tri 1572 19035 1709 19172 ne
rect 1709 19035 1884 19172
tri 1884 19035 2021 19172 sw
tri 2122 19035 2259 19172 ne
rect 2259 19035 2434 19172
tri 2434 19035 2571 19172 sw
tri 2672 19035 2809 19172 ne
rect 2809 19035 2984 19172
tri 2984 19035 3121 19172 sw
tri 3222 19035 3359 19172 ne
rect 3359 19035 3534 19172
tri 3534 19035 3671 19172 sw
tri 3772 19035 3909 19172 ne
rect 3909 19035 4084 19172
tri 4084 19035 4221 19172 sw
tri 4322 19035 4459 19172 ne
rect 4459 19035 4634 19172
tri 4634 19035 4771 19172 sw
tri 4872 19035 5009 19172 ne
rect 5009 19035 5184 19172
tri 5184 19035 5321 19172 sw
tri 5422 19035 5559 19172 ne
rect 5559 19035 5734 19172
tri 5734 19035 5871 19172 sw
tri 5972 19035 6109 19172 ne
rect 6109 19035 6284 19172
tri 6284 19035 6421 19172 sw
tri 6522 19035 6659 19172 ne
rect 6659 19035 6834 19172
tri 6834 19035 6971 19172 sw
tri 7072 19035 7209 19172 ne
rect 7209 19035 7384 19172
tri 7384 19035 7521 19172 sw
tri 7622 19035 7759 19172 ne
rect 7759 19035 7934 19172
tri 7934 19035 8071 19172 sw
tri 8172 19035 8309 19172 ne
rect 8309 19035 8484 19172
tri 8484 19035 8621 19172 sw
tri 8722 19035 8859 19172 ne
rect 8859 19035 9034 19172
tri 9034 19035 9171 19172 sw
tri 9272 19035 9409 19172 ne
rect 9409 19035 9584 19172
tri 9584 19035 9721 19172 sw
tri 9822 19035 9959 19172 ne
rect 9959 19035 10134 19172
tri 10134 19035 10271 19172 sw
tri 10372 19035 10509 19172 ne
rect 10509 19035 10684 19172
tri 10684 19035 10821 19172 sw
tri 10922 19035 11059 19172 ne
rect 11059 19035 11234 19172
tri 11234 19035 11371 19172 sw
tri 11472 19035 11609 19172 ne
rect 11609 19035 11784 19172
tri 11784 19035 11921 19172 sw
tri 12022 19035 12159 19172 ne
rect 12159 19035 12334 19172
tri 12334 19035 12471 19172 sw
tri 12572 19035 12709 19172 ne
rect 12709 19035 12884 19172
tri 12884 19035 13021 19172 sw
tri 13122 19035 13259 19172 ne
rect 13259 19035 13434 19172
tri 13434 19035 13571 19172 sw
tri 13672 19035 13809 19172 ne
rect 13809 19035 13984 19172
tri 13984 19035 14121 19172 sw
tri 14222 19035 14359 19172 ne
rect 14359 19035 14534 19172
tri 14534 19035 14671 19172 sw
tri 14772 19035 14909 19172 ne
rect 14909 19035 15084 19172
tri 15084 19035 15221 19172 sw
tri 15322 19035 15459 19172 ne
rect 15459 19035 15634 19172
tri 15634 19035 15771 19172 sw
tri 15872 19035 16009 19172 ne
rect 16009 19035 16184 19172
tri 16184 19035 16321 19172 sw
tri 16422 19035 16559 19172 ne
rect 16559 19035 16734 19172
tri 16734 19035 16871 19172 sw
tri 16972 19035 17109 19172 ne
rect 17109 19035 17284 19172
tri 17284 19035 17421 19172 sw
tri 17522 19035 17659 19172 ne
rect 17659 19035 17834 19172
tri 17834 19035 17971 19172 sw
tri 18072 19035 18209 19172 ne
rect 18209 19035 18384 19172
tri 18384 19035 18521 19172 sw
tri 18622 19035 18759 19172 ne
rect 18759 19035 18934 19172
tri 18934 19035 19071 19172 sw
tri 19172 19035 19309 19172 ne
rect 19309 19035 19484 19172
tri 19484 19035 19621 19172 sw
rect -500 19017 215 19035
tri 77 18915 179 19017 ne
rect 179 18915 215 19017
rect 335 18915 371 19035
tri 179 18778 316 18915 ne
rect 316 18860 371 18915
tri 371 18860 546 19035 sw
tri 609 18915 729 19035 ne
rect 729 18915 765 19035
rect 885 18915 921 19035
rect 316 18778 546 18860
tri 546 18778 628 18860 sw
tri 729 18778 866 18915 ne
rect 866 18860 921 18915
tri 921 18860 1096 19035 sw
tri 1159 18915 1279 19035 ne
rect 1279 18915 1315 19035
rect 1435 18915 1471 19035
rect 866 18778 1096 18860
tri 1096 18778 1178 18860 sw
tri 1279 18778 1416 18915 ne
rect 1416 18860 1471 18915
tri 1471 18860 1646 19035 sw
tri 1709 18915 1829 19035 ne
rect 1829 18915 1865 19035
rect 1985 18915 2021 19035
rect 1416 18778 1646 18860
tri 1646 18778 1728 18860 sw
tri 1829 18778 1966 18915 ne
rect 1966 18860 2021 18915
tri 2021 18860 2196 19035 sw
tri 2259 18915 2379 19035 ne
rect 2379 18915 2415 19035
rect 2535 18915 2571 19035
rect 1966 18778 2196 18860
tri 2196 18778 2278 18860 sw
tri 2379 18778 2516 18915 ne
rect 2516 18860 2571 18915
tri 2571 18860 2746 19035 sw
tri 2809 18915 2929 19035 ne
rect 2929 18915 2965 19035
rect 3085 18915 3121 19035
rect 2516 18778 2746 18860
tri 2746 18778 2828 18860 sw
tri 2929 18778 3066 18915 ne
rect 3066 18860 3121 18915
tri 3121 18860 3296 19035 sw
tri 3359 18915 3479 19035 ne
rect 3479 18915 3515 19035
rect 3635 18915 3671 19035
rect 3066 18778 3296 18860
tri 3296 18778 3378 18860 sw
tri 3479 18778 3616 18915 ne
rect 3616 18860 3671 18915
tri 3671 18860 3846 19035 sw
tri 3909 18915 4029 19035 ne
rect 4029 18915 4065 19035
rect 4185 18915 4221 19035
rect 3616 18778 3846 18860
tri 3846 18778 3928 18860 sw
tri 4029 18778 4166 18915 ne
rect 4166 18860 4221 18915
tri 4221 18860 4396 19035 sw
tri 4459 18915 4579 19035 ne
rect 4579 18915 4615 19035
rect 4735 18915 4771 19035
rect 4166 18778 4396 18860
tri 4396 18778 4478 18860 sw
tri 4579 18778 4716 18915 ne
rect 4716 18860 4771 18915
tri 4771 18860 4946 19035 sw
tri 5009 18915 5129 19035 ne
rect 5129 18915 5165 19035
rect 5285 18915 5321 19035
rect 4716 18778 4946 18860
tri 4946 18778 5028 18860 sw
tri 5129 18778 5266 18915 ne
rect 5266 18860 5321 18915
tri 5321 18860 5496 19035 sw
tri 5559 18915 5679 19035 ne
rect 5679 18915 5715 19035
rect 5835 18915 5871 19035
rect 5266 18778 5496 18860
tri 5496 18778 5578 18860 sw
tri 5679 18778 5816 18915 ne
rect 5816 18860 5871 18915
tri 5871 18860 6046 19035 sw
tri 6109 18915 6229 19035 ne
rect 6229 18915 6265 19035
rect 6385 18915 6421 19035
rect 5816 18778 6046 18860
tri 6046 18778 6128 18860 sw
tri 6229 18778 6366 18915 ne
rect 6366 18860 6421 18915
tri 6421 18860 6596 19035 sw
tri 6659 18915 6779 19035 ne
rect 6779 18915 6815 19035
rect 6935 18915 6971 19035
rect 6366 18778 6596 18860
tri 6596 18778 6678 18860 sw
tri 6779 18778 6916 18915 ne
rect 6916 18860 6971 18915
tri 6971 18860 7146 19035 sw
tri 7209 18915 7329 19035 ne
rect 7329 18915 7365 19035
rect 7485 18915 7521 19035
rect 6916 18778 7146 18860
tri 7146 18778 7228 18860 sw
tri 7329 18778 7466 18915 ne
rect 7466 18860 7521 18915
tri 7521 18860 7696 19035 sw
tri 7759 18915 7879 19035 ne
rect 7879 18915 7915 19035
rect 8035 18915 8071 19035
rect 7466 18778 7696 18860
tri 7696 18778 7778 18860 sw
tri 7879 18778 8016 18915 ne
rect 8016 18860 8071 18915
tri 8071 18860 8246 19035 sw
tri 8309 18915 8429 19035 ne
rect 8429 18915 8465 19035
rect 8585 18915 8621 19035
rect 8016 18778 8246 18860
tri 8246 18778 8328 18860 sw
tri 8429 18778 8566 18915 ne
rect 8566 18860 8621 18915
tri 8621 18860 8796 19035 sw
tri 8859 18915 8979 19035 ne
rect 8979 18915 9015 19035
rect 9135 18915 9171 19035
rect 8566 18778 8796 18860
tri 8796 18778 8878 18860 sw
tri 8979 18778 9116 18915 ne
rect 9116 18860 9171 18915
tri 9171 18860 9346 19035 sw
tri 9409 18915 9529 19035 ne
rect 9529 18915 9565 19035
rect 9685 18915 9721 19035
rect 9116 18778 9346 18860
tri 9346 18778 9428 18860 sw
tri 9529 18778 9666 18915 ne
rect 9666 18860 9721 18915
tri 9721 18860 9896 19035 sw
tri 9959 18915 10079 19035 ne
rect 10079 18915 10115 19035
rect 10235 18915 10271 19035
rect 9666 18778 9896 18860
tri 9896 18778 9978 18860 sw
tri 10079 18778 10216 18915 ne
rect 10216 18860 10271 18915
tri 10271 18860 10446 19035 sw
tri 10509 18915 10629 19035 ne
rect 10629 18915 10665 19035
rect 10785 18915 10821 19035
rect 10216 18778 10446 18860
tri 10446 18778 10528 18860 sw
tri 10629 18778 10766 18915 ne
rect 10766 18860 10821 18915
tri 10821 18860 10996 19035 sw
tri 11059 18915 11179 19035 ne
rect 11179 18915 11215 19035
rect 11335 18915 11371 19035
rect 10766 18778 10996 18860
tri 10996 18778 11078 18860 sw
tri 11179 18778 11316 18915 ne
rect 11316 18860 11371 18915
tri 11371 18860 11546 19035 sw
tri 11609 18915 11729 19035 ne
rect 11729 18915 11765 19035
rect 11885 18915 11921 19035
rect 11316 18778 11546 18860
tri 11546 18778 11628 18860 sw
tri 11729 18778 11866 18915 ne
rect 11866 18860 11921 18915
tri 11921 18860 12096 19035 sw
tri 12159 18915 12279 19035 ne
rect 12279 18915 12315 19035
rect 12435 18915 12471 19035
rect 11866 18778 12096 18860
tri 12096 18778 12178 18860 sw
tri 12279 18778 12416 18915 ne
rect 12416 18860 12471 18915
tri 12471 18860 12646 19035 sw
tri 12709 18915 12829 19035 ne
rect 12829 18915 12865 19035
rect 12985 18915 13021 19035
rect 12416 18778 12646 18860
tri 12646 18778 12728 18860 sw
tri 12829 18778 12966 18915 ne
rect 12966 18860 13021 18915
tri 13021 18860 13196 19035 sw
tri 13259 18915 13379 19035 ne
rect 13379 18915 13415 19035
rect 13535 18915 13571 19035
rect 12966 18778 13196 18860
tri 13196 18778 13278 18860 sw
tri 13379 18778 13516 18915 ne
rect 13516 18860 13571 18915
tri 13571 18860 13746 19035 sw
tri 13809 18915 13929 19035 ne
rect 13929 18915 13965 19035
rect 14085 18915 14121 19035
rect 13516 18778 13746 18860
tri 13746 18778 13828 18860 sw
tri 13929 18778 14066 18915 ne
rect 14066 18860 14121 18915
tri 14121 18860 14296 19035 sw
tri 14359 18915 14479 19035 ne
rect 14479 18915 14515 19035
rect 14635 18915 14671 19035
rect 14066 18778 14296 18860
tri 14296 18778 14378 18860 sw
tri 14479 18778 14616 18915 ne
rect 14616 18860 14671 18915
tri 14671 18860 14846 19035 sw
tri 14909 18915 15029 19035 ne
rect 15029 18915 15065 19035
rect 15185 18915 15221 19035
rect 14616 18778 14846 18860
tri 14846 18778 14928 18860 sw
tri 15029 18778 15166 18915 ne
rect 15166 18860 15221 18915
tri 15221 18860 15396 19035 sw
tri 15459 18915 15579 19035 ne
rect 15579 18915 15615 19035
rect 15735 18915 15771 19035
rect 15166 18778 15396 18860
tri 15396 18778 15478 18860 sw
tri 15579 18778 15716 18915 ne
rect 15716 18860 15771 18915
tri 15771 18860 15946 19035 sw
tri 16009 18915 16129 19035 ne
rect 16129 18915 16165 19035
rect 16285 18915 16321 19035
rect 15716 18778 15946 18860
tri 15946 18778 16028 18860 sw
tri 16129 18778 16266 18915 ne
rect 16266 18860 16321 18915
tri 16321 18860 16496 19035 sw
tri 16559 18915 16679 19035 ne
rect 16679 18915 16715 19035
rect 16835 18915 16871 19035
rect 16266 18778 16496 18860
tri 16496 18778 16578 18860 sw
tri 16679 18778 16816 18915 ne
rect 16816 18860 16871 18915
tri 16871 18860 17046 19035 sw
tri 17109 18915 17229 19035 ne
rect 17229 18915 17265 19035
rect 17385 18915 17421 19035
rect 16816 18778 17046 18860
tri 17046 18778 17128 18860 sw
tri 17229 18778 17366 18915 ne
rect 17366 18860 17421 18915
tri 17421 18860 17596 19035 sw
tri 17659 18915 17779 19035 ne
rect 17779 18915 17815 19035
rect 17935 18915 17971 19035
rect 17366 18778 17596 18860
tri 17596 18778 17678 18860 sw
tri 17779 18778 17916 18915 ne
rect 17916 18860 17971 18915
tri 17971 18860 18146 19035 sw
tri 18209 18915 18329 19035 ne
rect 18329 18915 18365 19035
rect 18485 18915 18521 19035
rect 17916 18778 18146 18860
tri 18146 18778 18228 18860 sw
tri 18329 18778 18466 18915 ne
rect 18466 18860 18521 18915
tri 18521 18860 18696 19035 sw
tri 18759 18915 18879 19035 ne
rect 18879 18915 18915 19035
rect 19035 18915 19071 19035
rect 18466 18778 18696 18860
tri 18696 18778 18778 18860 sw
tri 18879 18778 19016 18915 ne
rect 19016 18860 19071 18915
tri 19071 18860 19246 19035 sw
tri 19309 18915 19429 19035 ne
rect 19429 18915 19465 19035
rect 19585 18933 19621 19035
tri 19621 18933 19723 19035 sw
rect 19585 18915 20300 18933
rect 19016 18778 19246 18860
tri 19246 18778 19328 18860 sw
tri 19429 18778 19566 18915 ne
rect 19566 18778 20300 18915
rect -2000 18622 78 18778
tri 78 18622 234 18778 sw
tri 316 18622 472 18778 ne
rect 472 18622 628 18778
tri 628 18622 784 18778 sw
tri 866 18622 1022 18778 ne
rect 1022 18622 1178 18778
tri 1178 18622 1334 18778 sw
tri 1416 18622 1572 18778 ne
rect 1572 18622 1728 18778
tri 1728 18622 1884 18778 sw
tri 1966 18622 2122 18778 ne
rect 2122 18622 2278 18778
tri 2278 18622 2434 18778 sw
tri 2516 18622 2672 18778 ne
rect 2672 18622 2828 18778
tri 2828 18622 2984 18778 sw
tri 3066 18622 3222 18778 ne
rect 3222 18622 3378 18778
tri 3378 18622 3534 18778 sw
tri 3616 18622 3772 18778 ne
rect 3772 18622 3928 18778
tri 3928 18622 4084 18778 sw
tri 4166 18622 4322 18778 ne
rect 4322 18622 4478 18778
tri 4478 18622 4634 18778 sw
tri 4716 18622 4872 18778 ne
rect 4872 18622 5028 18778
tri 5028 18622 5184 18778 sw
tri 5266 18622 5422 18778 ne
rect 5422 18622 5578 18778
tri 5578 18622 5734 18778 sw
tri 5816 18622 5972 18778 ne
rect 5972 18622 6128 18778
tri 6128 18622 6284 18778 sw
tri 6366 18622 6522 18778 ne
rect 6522 18622 6678 18778
tri 6678 18622 6834 18778 sw
tri 6916 18622 7072 18778 ne
rect 7072 18622 7228 18778
tri 7228 18622 7384 18778 sw
tri 7466 18622 7622 18778 ne
rect 7622 18622 7778 18778
tri 7778 18622 7934 18778 sw
tri 8016 18622 8172 18778 ne
rect 8172 18622 8328 18778
tri 8328 18622 8484 18778 sw
tri 8566 18622 8722 18778 ne
rect 8722 18622 8878 18778
tri 8878 18622 9034 18778 sw
tri 9116 18622 9272 18778 ne
rect 9272 18622 9428 18778
tri 9428 18622 9584 18778 sw
tri 9666 18622 9822 18778 ne
rect 9822 18622 9978 18778
tri 9978 18622 10134 18778 sw
tri 10216 18622 10372 18778 ne
rect 10372 18622 10528 18778
tri 10528 18622 10684 18778 sw
tri 10766 18622 10922 18778 ne
rect 10922 18622 11078 18778
tri 11078 18622 11234 18778 sw
tri 11316 18622 11472 18778 ne
rect 11472 18622 11628 18778
tri 11628 18622 11784 18778 sw
tri 11866 18622 12022 18778 ne
rect 12022 18622 12178 18778
tri 12178 18622 12334 18778 sw
tri 12416 18622 12572 18778 ne
rect 12572 18622 12728 18778
tri 12728 18622 12884 18778 sw
tri 12966 18622 13122 18778 ne
rect 13122 18622 13278 18778
tri 13278 18622 13434 18778 sw
tri 13516 18622 13672 18778 ne
rect 13672 18622 13828 18778
tri 13828 18622 13984 18778 sw
tri 14066 18622 14222 18778 ne
rect 14222 18622 14378 18778
tri 14378 18622 14534 18778 sw
tri 14616 18622 14772 18778 ne
rect 14772 18622 14928 18778
tri 14928 18622 15084 18778 sw
tri 15166 18622 15322 18778 ne
rect 15322 18622 15478 18778
tri 15478 18622 15634 18778 sw
tri 15716 18622 15872 18778 ne
rect 15872 18622 16028 18778
tri 16028 18622 16184 18778 sw
tri 16266 18622 16422 18778 ne
rect 16422 18622 16578 18778
tri 16578 18622 16734 18778 sw
tri 16816 18622 16972 18778 ne
rect 16972 18622 17128 18778
tri 17128 18622 17284 18778 sw
tri 17366 18622 17522 18778 ne
rect 17522 18622 17678 18778
tri 17678 18622 17834 18778 sw
tri 17916 18622 18072 18778 ne
rect 18072 18622 18228 18778
tri 18228 18622 18384 18778 sw
tri 18466 18622 18622 18778 ne
rect 18622 18622 18778 18778
tri 18778 18622 18934 18778 sw
tri 19016 18622 19172 18778 ne
rect 19172 18622 19328 18778
tri 19328 18622 19484 18778 sw
tri 19566 18622 19722 18778 ne
rect 19722 18622 20300 18778
rect -2000 18485 234 18622
tri 234 18485 371 18622 sw
tri 472 18485 609 18622 ne
rect 609 18485 784 18622
tri 784 18485 921 18622 sw
tri 1022 18485 1159 18622 ne
rect 1159 18485 1334 18622
tri 1334 18485 1471 18622 sw
tri 1572 18485 1709 18622 ne
rect 1709 18485 1884 18622
tri 1884 18485 2021 18622 sw
tri 2122 18485 2259 18622 ne
rect 2259 18485 2434 18622
tri 2434 18485 2571 18622 sw
tri 2672 18485 2809 18622 ne
rect 2809 18485 2984 18622
tri 2984 18485 3121 18622 sw
tri 3222 18485 3359 18622 ne
rect 3359 18485 3534 18622
tri 3534 18485 3671 18622 sw
tri 3772 18485 3909 18622 ne
rect 3909 18485 4084 18622
tri 4084 18485 4221 18622 sw
tri 4322 18485 4459 18622 ne
rect 4459 18485 4634 18622
tri 4634 18485 4771 18622 sw
tri 4872 18485 5009 18622 ne
rect 5009 18485 5184 18622
tri 5184 18485 5321 18622 sw
tri 5422 18485 5559 18622 ne
rect 5559 18485 5734 18622
tri 5734 18485 5871 18622 sw
tri 5972 18485 6109 18622 ne
rect 6109 18485 6284 18622
tri 6284 18485 6421 18622 sw
tri 6522 18485 6659 18622 ne
rect 6659 18485 6834 18622
tri 6834 18485 6971 18622 sw
tri 7072 18485 7209 18622 ne
rect 7209 18485 7384 18622
tri 7384 18485 7521 18622 sw
tri 7622 18485 7759 18622 ne
rect 7759 18485 7934 18622
tri 7934 18485 8071 18622 sw
tri 8172 18485 8309 18622 ne
rect 8309 18485 8484 18622
tri 8484 18485 8621 18622 sw
tri 8722 18485 8859 18622 ne
rect 8859 18485 9034 18622
tri 9034 18485 9171 18622 sw
tri 9272 18485 9409 18622 ne
rect 9409 18485 9584 18622
tri 9584 18485 9721 18622 sw
tri 9822 18485 9959 18622 ne
rect 9959 18485 10134 18622
tri 10134 18485 10271 18622 sw
tri 10372 18485 10509 18622 ne
rect 10509 18485 10684 18622
tri 10684 18485 10821 18622 sw
tri 10922 18485 11059 18622 ne
rect 11059 18485 11234 18622
tri 11234 18485 11371 18622 sw
tri 11472 18485 11609 18622 ne
rect 11609 18485 11784 18622
tri 11784 18485 11921 18622 sw
tri 12022 18485 12159 18622 ne
rect 12159 18485 12334 18622
tri 12334 18485 12471 18622 sw
tri 12572 18485 12709 18622 ne
rect 12709 18485 12884 18622
tri 12884 18485 13021 18622 sw
tri 13122 18485 13259 18622 ne
rect 13259 18485 13434 18622
tri 13434 18485 13571 18622 sw
tri 13672 18485 13809 18622 ne
rect 13809 18485 13984 18622
tri 13984 18485 14121 18622 sw
tri 14222 18485 14359 18622 ne
rect 14359 18485 14534 18622
tri 14534 18485 14671 18622 sw
tri 14772 18485 14909 18622 ne
rect 14909 18485 15084 18622
tri 15084 18485 15221 18622 sw
tri 15322 18485 15459 18622 ne
rect 15459 18485 15634 18622
tri 15634 18485 15771 18622 sw
tri 15872 18485 16009 18622 ne
rect 16009 18485 16184 18622
tri 16184 18485 16321 18622 sw
tri 16422 18485 16559 18622 ne
rect 16559 18485 16734 18622
tri 16734 18485 16871 18622 sw
tri 16972 18485 17109 18622 ne
rect 17109 18485 17284 18622
tri 17284 18485 17421 18622 sw
tri 17522 18485 17659 18622 ne
rect 17659 18485 17834 18622
tri 17834 18485 17971 18622 sw
tri 18072 18485 18209 18622 ne
rect 18209 18485 18384 18622
tri 18384 18485 18521 18622 sw
tri 18622 18485 18759 18622 ne
rect 18759 18485 18934 18622
tri 18934 18485 19071 18622 sw
tri 19172 18485 19309 18622 ne
rect 19309 18485 19484 18622
tri 19484 18485 19621 18622 sw
rect -2000 18467 215 18485
rect -2000 17678 -1000 18467
tri 77 18365 179 18467 ne
rect 179 18365 215 18467
rect 335 18365 371 18485
tri 179 18228 316 18365 ne
rect 316 18310 371 18365
tri 371 18310 546 18485 sw
tri 609 18365 729 18485 ne
rect 729 18365 765 18485
rect 885 18365 921 18485
rect 316 18228 546 18310
tri 546 18228 628 18310 sw
tri 729 18228 866 18365 ne
rect 866 18310 921 18365
tri 921 18310 1096 18485 sw
tri 1159 18365 1279 18485 ne
rect 1279 18365 1315 18485
rect 1435 18365 1471 18485
rect 866 18228 1096 18310
tri 1096 18228 1178 18310 sw
tri 1279 18228 1416 18365 ne
rect 1416 18310 1471 18365
tri 1471 18310 1646 18485 sw
tri 1709 18365 1829 18485 ne
rect 1829 18365 1865 18485
rect 1985 18365 2021 18485
rect 1416 18228 1646 18310
tri 1646 18228 1728 18310 sw
tri 1829 18228 1966 18365 ne
rect 1966 18310 2021 18365
tri 2021 18310 2196 18485 sw
tri 2259 18365 2379 18485 ne
rect 2379 18365 2415 18485
rect 2535 18365 2571 18485
rect 1966 18228 2196 18310
tri 2196 18228 2278 18310 sw
tri 2379 18228 2516 18365 ne
rect 2516 18310 2571 18365
tri 2571 18310 2746 18485 sw
tri 2809 18365 2929 18485 ne
rect 2929 18365 2965 18485
rect 3085 18365 3121 18485
rect 2516 18228 2746 18310
tri 2746 18228 2828 18310 sw
tri 2929 18228 3066 18365 ne
rect 3066 18310 3121 18365
tri 3121 18310 3296 18485 sw
tri 3359 18365 3479 18485 ne
rect 3479 18365 3515 18485
rect 3635 18365 3671 18485
rect 3066 18228 3296 18310
tri 3296 18228 3378 18310 sw
tri 3479 18228 3616 18365 ne
rect 3616 18310 3671 18365
tri 3671 18310 3846 18485 sw
tri 3909 18365 4029 18485 ne
rect 4029 18365 4065 18485
rect 4185 18365 4221 18485
rect 3616 18228 3846 18310
tri 3846 18228 3928 18310 sw
tri 4029 18228 4166 18365 ne
rect 4166 18310 4221 18365
tri 4221 18310 4396 18485 sw
tri 4459 18365 4579 18485 ne
rect 4579 18365 4615 18485
rect 4735 18365 4771 18485
rect 4166 18228 4396 18310
tri 4396 18228 4478 18310 sw
tri 4579 18228 4716 18365 ne
rect 4716 18310 4771 18365
tri 4771 18310 4946 18485 sw
tri 5009 18365 5129 18485 ne
rect 5129 18365 5165 18485
rect 5285 18365 5321 18485
rect 4716 18228 4946 18310
tri 4946 18228 5028 18310 sw
tri 5129 18228 5266 18365 ne
rect 5266 18310 5321 18365
tri 5321 18310 5496 18485 sw
tri 5559 18365 5679 18485 ne
rect 5679 18365 5715 18485
rect 5835 18365 5871 18485
rect 5266 18228 5496 18310
tri 5496 18228 5578 18310 sw
tri 5679 18228 5816 18365 ne
rect 5816 18310 5871 18365
tri 5871 18310 6046 18485 sw
tri 6109 18365 6229 18485 ne
rect 6229 18365 6265 18485
rect 6385 18365 6421 18485
rect 5816 18228 6046 18310
tri 6046 18228 6128 18310 sw
tri 6229 18228 6366 18365 ne
rect 6366 18310 6421 18365
tri 6421 18310 6596 18485 sw
tri 6659 18365 6779 18485 ne
rect 6779 18365 6815 18485
rect 6935 18365 6971 18485
rect 6366 18228 6596 18310
tri 6596 18228 6678 18310 sw
tri 6779 18228 6916 18365 ne
rect 6916 18310 6971 18365
tri 6971 18310 7146 18485 sw
tri 7209 18365 7329 18485 ne
rect 7329 18365 7365 18485
rect 7485 18365 7521 18485
rect 6916 18228 7146 18310
tri 7146 18228 7228 18310 sw
tri 7329 18228 7466 18365 ne
rect 7466 18310 7521 18365
tri 7521 18310 7696 18485 sw
tri 7759 18365 7879 18485 ne
rect 7879 18365 7915 18485
rect 8035 18365 8071 18485
rect 7466 18228 7696 18310
tri 7696 18228 7778 18310 sw
tri 7879 18228 8016 18365 ne
rect 8016 18310 8071 18365
tri 8071 18310 8246 18485 sw
tri 8309 18365 8429 18485 ne
rect 8429 18365 8465 18485
rect 8585 18365 8621 18485
rect 8016 18228 8246 18310
tri 8246 18228 8328 18310 sw
tri 8429 18228 8566 18365 ne
rect 8566 18310 8621 18365
tri 8621 18310 8796 18485 sw
tri 8859 18365 8979 18485 ne
rect 8979 18365 9015 18485
rect 9135 18365 9171 18485
rect 8566 18228 8796 18310
tri 8796 18228 8878 18310 sw
tri 8979 18228 9116 18365 ne
rect 9116 18310 9171 18365
tri 9171 18310 9346 18485 sw
tri 9409 18365 9529 18485 ne
rect 9529 18365 9565 18485
rect 9685 18365 9721 18485
rect 9116 18228 9346 18310
tri 9346 18228 9428 18310 sw
tri 9529 18228 9666 18365 ne
rect 9666 18310 9721 18365
tri 9721 18310 9896 18485 sw
tri 9959 18365 10079 18485 ne
rect 10079 18365 10115 18485
rect 10235 18365 10271 18485
rect 9666 18228 9896 18310
tri 9896 18228 9978 18310 sw
tri 10079 18228 10216 18365 ne
rect 10216 18310 10271 18365
tri 10271 18310 10446 18485 sw
tri 10509 18365 10629 18485 ne
rect 10629 18365 10665 18485
rect 10785 18365 10821 18485
rect 10216 18228 10446 18310
tri 10446 18228 10528 18310 sw
tri 10629 18228 10766 18365 ne
rect 10766 18310 10821 18365
tri 10821 18310 10996 18485 sw
tri 11059 18365 11179 18485 ne
rect 11179 18365 11215 18485
rect 11335 18365 11371 18485
rect 10766 18228 10996 18310
tri 10996 18228 11078 18310 sw
tri 11179 18228 11316 18365 ne
rect 11316 18310 11371 18365
tri 11371 18310 11546 18485 sw
tri 11609 18365 11729 18485 ne
rect 11729 18365 11765 18485
rect 11885 18365 11921 18485
rect 11316 18228 11546 18310
tri 11546 18228 11628 18310 sw
tri 11729 18228 11866 18365 ne
rect 11866 18310 11921 18365
tri 11921 18310 12096 18485 sw
tri 12159 18365 12279 18485 ne
rect 12279 18365 12315 18485
rect 12435 18365 12471 18485
rect 11866 18228 12096 18310
tri 12096 18228 12178 18310 sw
tri 12279 18228 12416 18365 ne
rect 12416 18310 12471 18365
tri 12471 18310 12646 18485 sw
tri 12709 18365 12829 18485 ne
rect 12829 18365 12865 18485
rect 12985 18365 13021 18485
rect 12416 18228 12646 18310
tri 12646 18228 12728 18310 sw
tri 12829 18228 12966 18365 ne
rect 12966 18310 13021 18365
tri 13021 18310 13196 18485 sw
tri 13259 18365 13379 18485 ne
rect 13379 18365 13415 18485
rect 13535 18365 13571 18485
rect 12966 18228 13196 18310
tri 13196 18228 13278 18310 sw
tri 13379 18228 13516 18365 ne
rect 13516 18310 13571 18365
tri 13571 18310 13746 18485 sw
tri 13809 18365 13929 18485 ne
rect 13929 18365 13965 18485
rect 14085 18365 14121 18485
rect 13516 18228 13746 18310
tri 13746 18228 13828 18310 sw
tri 13929 18228 14066 18365 ne
rect 14066 18310 14121 18365
tri 14121 18310 14296 18485 sw
tri 14359 18365 14479 18485 ne
rect 14479 18365 14515 18485
rect 14635 18365 14671 18485
rect 14066 18228 14296 18310
tri 14296 18228 14378 18310 sw
tri 14479 18228 14616 18365 ne
rect 14616 18310 14671 18365
tri 14671 18310 14846 18485 sw
tri 14909 18365 15029 18485 ne
rect 15029 18365 15065 18485
rect 15185 18365 15221 18485
rect 14616 18228 14846 18310
tri 14846 18228 14928 18310 sw
tri 15029 18228 15166 18365 ne
rect 15166 18310 15221 18365
tri 15221 18310 15396 18485 sw
tri 15459 18365 15579 18485 ne
rect 15579 18365 15615 18485
rect 15735 18365 15771 18485
rect 15166 18228 15396 18310
tri 15396 18228 15478 18310 sw
tri 15579 18228 15716 18365 ne
rect 15716 18310 15771 18365
tri 15771 18310 15946 18485 sw
tri 16009 18365 16129 18485 ne
rect 16129 18365 16165 18485
rect 16285 18365 16321 18485
rect 15716 18228 15946 18310
tri 15946 18228 16028 18310 sw
tri 16129 18228 16266 18365 ne
rect 16266 18310 16321 18365
tri 16321 18310 16496 18485 sw
tri 16559 18365 16679 18485 ne
rect 16679 18365 16715 18485
rect 16835 18365 16871 18485
rect 16266 18228 16496 18310
tri 16496 18228 16578 18310 sw
tri 16679 18228 16816 18365 ne
rect 16816 18310 16871 18365
tri 16871 18310 17046 18485 sw
tri 17109 18365 17229 18485 ne
rect 17229 18365 17265 18485
rect 17385 18365 17421 18485
rect 16816 18228 17046 18310
tri 17046 18228 17128 18310 sw
tri 17229 18228 17366 18365 ne
rect 17366 18310 17421 18365
tri 17421 18310 17596 18485 sw
tri 17659 18365 17779 18485 ne
rect 17779 18365 17815 18485
rect 17935 18365 17971 18485
rect 17366 18228 17596 18310
tri 17596 18228 17678 18310 sw
tri 17779 18228 17916 18365 ne
rect 17916 18310 17971 18365
tri 17971 18310 18146 18485 sw
tri 18209 18365 18329 18485 ne
rect 18329 18365 18365 18485
rect 18485 18365 18521 18485
rect 17916 18228 18146 18310
tri 18146 18228 18228 18310 sw
tri 18329 18228 18466 18365 ne
rect 18466 18310 18521 18365
tri 18521 18310 18696 18485 sw
tri 18759 18365 18879 18485 ne
rect 18879 18365 18915 18485
rect 19035 18365 19071 18485
rect 18466 18228 18696 18310
tri 18696 18228 18778 18310 sw
tri 18879 18228 19016 18365 ne
rect 19016 18310 19071 18365
tri 19071 18310 19246 18485 sw
tri 19309 18365 19429 18485 ne
rect 19429 18365 19465 18485
rect 19585 18383 19621 18485
tri 19621 18383 19723 18485 sw
rect 20800 18383 21800 19172
rect 19585 18365 21800 18383
rect 19016 18228 19246 18310
tri 19246 18228 19328 18310 sw
tri 19429 18228 19566 18365 ne
rect 19566 18228 21800 18365
rect -500 18072 78 18228
tri 78 18072 234 18228 sw
tri 316 18072 472 18228 ne
rect 472 18072 628 18228
tri 628 18072 784 18228 sw
tri 866 18072 1022 18228 ne
rect 1022 18072 1178 18228
tri 1178 18072 1334 18228 sw
tri 1416 18072 1572 18228 ne
rect 1572 18072 1728 18228
tri 1728 18072 1884 18228 sw
tri 1966 18072 2122 18228 ne
rect 2122 18072 2278 18228
tri 2278 18072 2434 18228 sw
tri 2516 18072 2672 18228 ne
rect 2672 18072 2828 18228
tri 2828 18072 2984 18228 sw
tri 3066 18072 3222 18228 ne
rect 3222 18072 3378 18228
tri 3378 18072 3534 18228 sw
tri 3616 18072 3772 18228 ne
rect 3772 18072 3928 18228
tri 3928 18072 4084 18228 sw
tri 4166 18072 4322 18228 ne
rect 4322 18072 4478 18228
tri 4478 18072 4634 18228 sw
tri 4716 18072 4872 18228 ne
rect 4872 18072 5028 18228
tri 5028 18072 5184 18228 sw
tri 5266 18072 5422 18228 ne
rect 5422 18072 5578 18228
tri 5578 18072 5734 18228 sw
tri 5816 18072 5972 18228 ne
rect 5972 18072 6128 18228
tri 6128 18072 6284 18228 sw
tri 6366 18072 6522 18228 ne
rect 6522 18072 6678 18228
tri 6678 18072 6834 18228 sw
tri 6916 18072 7072 18228 ne
rect 7072 18072 7228 18228
tri 7228 18072 7384 18228 sw
tri 7466 18072 7622 18228 ne
rect 7622 18072 7778 18228
tri 7778 18072 7934 18228 sw
tri 8016 18072 8172 18228 ne
rect 8172 18072 8328 18228
tri 8328 18072 8484 18228 sw
tri 8566 18072 8722 18228 ne
rect 8722 18072 8878 18228
tri 8878 18072 9034 18228 sw
tri 9116 18072 9272 18228 ne
rect 9272 18072 9428 18228
tri 9428 18072 9584 18228 sw
tri 9666 18072 9822 18228 ne
rect 9822 18072 9978 18228
tri 9978 18072 10134 18228 sw
tri 10216 18072 10372 18228 ne
rect 10372 18072 10528 18228
tri 10528 18072 10684 18228 sw
tri 10766 18072 10922 18228 ne
rect 10922 18072 11078 18228
tri 11078 18072 11234 18228 sw
tri 11316 18072 11472 18228 ne
rect 11472 18072 11628 18228
tri 11628 18072 11784 18228 sw
tri 11866 18072 12022 18228 ne
rect 12022 18072 12178 18228
tri 12178 18072 12334 18228 sw
tri 12416 18072 12572 18228 ne
rect 12572 18072 12728 18228
tri 12728 18072 12884 18228 sw
tri 12966 18072 13122 18228 ne
rect 13122 18072 13278 18228
tri 13278 18072 13434 18228 sw
tri 13516 18072 13672 18228 ne
rect 13672 18072 13828 18228
tri 13828 18072 13984 18228 sw
tri 14066 18072 14222 18228 ne
rect 14222 18072 14378 18228
tri 14378 18072 14534 18228 sw
tri 14616 18072 14772 18228 ne
rect 14772 18072 14928 18228
tri 14928 18072 15084 18228 sw
tri 15166 18072 15322 18228 ne
rect 15322 18072 15478 18228
tri 15478 18072 15634 18228 sw
tri 15716 18072 15872 18228 ne
rect 15872 18072 16028 18228
tri 16028 18072 16184 18228 sw
tri 16266 18072 16422 18228 ne
rect 16422 18072 16578 18228
tri 16578 18072 16734 18228 sw
tri 16816 18072 16972 18228 ne
rect 16972 18072 17128 18228
tri 17128 18072 17284 18228 sw
tri 17366 18072 17522 18228 ne
rect 17522 18072 17678 18228
tri 17678 18072 17834 18228 sw
tri 17916 18072 18072 18228 ne
rect 18072 18072 18228 18228
tri 18228 18072 18384 18228 sw
tri 18466 18072 18622 18228 ne
rect 18622 18072 18778 18228
tri 18778 18072 18934 18228 sw
tri 19016 18072 19172 18228 ne
rect 19172 18072 19328 18228
tri 19328 18072 19484 18228 sw
tri 19566 18072 19722 18228 ne
rect 19722 18072 21800 18228
rect -500 17935 234 18072
tri 234 17935 371 18072 sw
tri 472 17935 609 18072 ne
rect 609 17935 784 18072
tri 784 17935 921 18072 sw
tri 1022 17935 1159 18072 ne
rect 1159 17935 1334 18072
tri 1334 17935 1471 18072 sw
tri 1572 17935 1709 18072 ne
rect 1709 17935 1884 18072
tri 1884 17935 2021 18072 sw
tri 2122 17935 2259 18072 ne
rect 2259 17935 2434 18072
tri 2434 17935 2571 18072 sw
tri 2672 17935 2809 18072 ne
rect 2809 17935 2984 18072
tri 2984 17935 3121 18072 sw
tri 3222 17935 3359 18072 ne
rect 3359 17935 3534 18072
tri 3534 17935 3671 18072 sw
tri 3772 17935 3909 18072 ne
rect 3909 17935 4084 18072
tri 4084 17935 4221 18072 sw
tri 4322 17935 4459 18072 ne
rect 4459 17935 4634 18072
tri 4634 17935 4771 18072 sw
tri 4872 17935 5009 18072 ne
rect 5009 17935 5184 18072
tri 5184 17935 5321 18072 sw
tri 5422 17935 5559 18072 ne
rect 5559 17935 5734 18072
tri 5734 17935 5871 18072 sw
tri 5972 17935 6109 18072 ne
rect 6109 17935 6284 18072
tri 6284 17935 6421 18072 sw
tri 6522 17935 6659 18072 ne
rect 6659 17935 6834 18072
tri 6834 17935 6971 18072 sw
tri 7072 17935 7209 18072 ne
rect 7209 17935 7384 18072
tri 7384 17935 7521 18072 sw
tri 7622 17935 7759 18072 ne
rect 7759 17935 7934 18072
tri 7934 17935 8071 18072 sw
tri 8172 17935 8309 18072 ne
rect 8309 17935 8484 18072
tri 8484 17935 8621 18072 sw
tri 8722 17935 8859 18072 ne
rect 8859 17935 9034 18072
tri 9034 17935 9171 18072 sw
tri 9272 17935 9409 18072 ne
rect 9409 17935 9584 18072
tri 9584 17935 9721 18072 sw
tri 9822 17935 9959 18072 ne
rect 9959 17935 10134 18072
tri 10134 17935 10271 18072 sw
tri 10372 17935 10509 18072 ne
rect 10509 17935 10684 18072
tri 10684 17935 10821 18072 sw
tri 10922 17935 11059 18072 ne
rect 11059 17935 11234 18072
tri 11234 17935 11371 18072 sw
tri 11472 17935 11609 18072 ne
rect 11609 17935 11784 18072
tri 11784 17935 11921 18072 sw
tri 12022 17935 12159 18072 ne
rect 12159 17935 12334 18072
tri 12334 17935 12471 18072 sw
tri 12572 17935 12709 18072 ne
rect 12709 17935 12884 18072
tri 12884 17935 13021 18072 sw
tri 13122 17935 13259 18072 ne
rect 13259 17935 13434 18072
tri 13434 17935 13571 18072 sw
tri 13672 17935 13809 18072 ne
rect 13809 17935 13984 18072
tri 13984 17935 14121 18072 sw
tri 14222 17935 14359 18072 ne
rect 14359 17935 14534 18072
tri 14534 17935 14671 18072 sw
tri 14772 17935 14909 18072 ne
rect 14909 17935 15084 18072
tri 15084 17935 15221 18072 sw
tri 15322 17935 15459 18072 ne
rect 15459 17935 15634 18072
tri 15634 17935 15771 18072 sw
tri 15872 17935 16009 18072 ne
rect 16009 17935 16184 18072
tri 16184 17935 16321 18072 sw
tri 16422 17935 16559 18072 ne
rect 16559 17935 16734 18072
tri 16734 17935 16871 18072 sw
tri 16972 17935 17109 18072 ne
rect 17109 17935 17284 18072
tri 17284 17935 17421 18072 sw
tri 17522 17935 17659 18072 ne
rect 17659 17935 17834 18072
tri 17834 17935 17971 18072 sw
tri 18072 17935 18209 18072 ne
rect 18209 17935 18384 18072
tri 18384 17935 18521 18072 sw
tri 18622 17935 18759 18072 ne
rect 18759 17935 18934 18072
tri 18934 17935 19071 18072 sw
tri 19172 17935 19309 18072 ne
rect 19309 17935 19484 18072
tri 19484 17935 19621 18072 sw
rect -500 17917 215 17935
tri 77 17815 179 17917 ne
rect 179 17815 215 17917
rect 335 17815 371 17935
tri 179 17678 316 17815 ne
rect 316 17760 371 17815
tri 371 17760 546 17935 sw
tri 609 17815 729 17935 ne
rect 729 17815 765 17935
rect 885 17815 921 17935
rect 316 17678 546 17760
tri 546 17678 628 17760 sw
tri 729 17678 866 17815 ne
rect 866 17760 921 17815
tri 921 17760 1096 17935 sw
tri 1159 17815 1279 17935 ne
rect 1279 17815 1315 17935
rect 1435 17815 1471 17935
rect 866 17678 1096 17760
tri 1096 17678 1178 17760 sw
tri 1279 17678 1416 17815 ne
rect 1416 17760 1471 17815
tri 1471 17760 1646 17935 sw
tri 1709 17815 1829 17935 ne
rect 1829 17815 1865 17935
rect 1985 17815 2021 17935
rect 1416 17678 1646 17760
tri 1646 17678 1728 17760 sw
tri 1829 17678 1966 17815 ne
rect 1966 17760 2021 17815
tri 2021 17760 2196 17935 sw
tri 2259 17815 2379 17935 ne
rect 2379 17815 2415 17935
rect 2535 17815 2571 17935
rect 1966 17678 2196 17760
tri 2196 17678 2278 17760 sw
tri 2379 17678 2516 17815 ne
rect 2516 17760 2571 17815
tri 2571 17760 2746 17935 sw
tri 2809 17815 2929 17935 ne
rect 2929 17815 2965 17935
rect 3085 17815 3121 17935
rect 2516 17678 2746 17760
tri 2746 17678 2828 17760 sw
tri 2929 17678 3066 17815 ne
rect 3066 17760 3121 17815
tri 3121 17760 3296 17935 sw
tri 3359 17815 3479 17935 ne
rect 3479 17815 3515 17935
rect 3635 17815 3671 17935
rect 3066 17678 3296 17760
tri 3296 17678 3378 17760 sw
tri 3479 17678 3616 17815 ne
rect 3616 17760 3671 17815
tri 3671 17760 3846 17935 sw
tri 3909 17815 4029 17935 ne
rect 4029 17815 4065 17935
rect 4185 17815 4221 17935
rect 3616 17678 3846 17760
tri 3846 17678 3928 17760 sw
tri 4029 17678 4166 17815 ne
rect 4166 17760 4221 17815
tri 4221 17760 4396 17935 sw
tri 4459 17815 4579 17935 ne
rect 4579 17815 4615 17935
rect 4735 17815 4771 17935
rect 4166 17678 4396 17760
tri 4396 17678 4478 17760 sw
tri 4579 17678 4716 17815 ne
rect 4716 17760 4771 17815
tri 4771 17760 4946 17935 sw
tri 5009 17815 5129 17935 ne
rect 5129 17815 5165 17935
rect 5285 17815 5321 17935
rect 4716 17678 4946 17760
tri 4946 17678 5028 17760 sw
tri 5129 17678 5266 17815 ne
rect 5266 17760 5321 17815
tri 5321 17760 5496 17935 sw
tri 5559 17815 5679 17935 ne
rect 5679 17815 5715 17935
rect 5835 17815 5871 17935
rect 5266 17678 5496 17760
tri 5496 17678 5578 17760 sw
tri 5679 17678 5816 17815 ne
rect 5816 17760 5871 17815
tri 5871 17760 6046 17935 sw
tri 6109 17815 6229 17935 ne
rect 6229 17815 6265 17935
rect 6385 17815 6421 17935
rect 5816 17678 6046 17760
tri 6046 17678 6128 17760 sw
tri 6229 17678 6366 17815 ne
rect 6366 17760 6421 17815
tri 6421 17760 6596 17935 sw
tri 6659 17815 6779 17935 ne
rect 6779 17815 6815 17935
rect 6935 17815 6971 17935
rect 6366 17678 6596 17760
tri 6596 17678 6678 17760 sw
tri 6779 17678 6916 17815 ne
rect 6916 17760 6971 17815
tri 6971 17760 7146 17935 sw
tri 7209 17815 7329 17935 ne
rect 7329 17815 7365 17935
rect 7485 17815 7521 17935
rect 6916 17678 7146 17760
tri 7146 17678 7228 17760 sw
tri 7329 17678 7466 17815 ne
rect 7466 17760 7521 17815
tri 7521 17760 7696 17935 sw
tri 7759 17815 7879 17935 ne
rect 7879 17815 7915 17935
rect 8035 17815 8071 17935
rect 7466 17678 7696 17760
tri 7696 17678 7778 17760 sw
tri 7879 17678 8016 17815 ne
rect 8016 17760 8071 17815
tri 8071 17760 8246 17935 sw
tri 8309 17815 8429 17935 ne
rect 8429 17815 8465 17935
rect 8585 17815 8621 17935
rect 8016 17678 8246 17760
tri 8246 17678 8328 17760 sw
tri 8429 17678 8566 17815 ne
rect 8566 17760 8621 17815
tri 8621 17760 8796 17935 sw
tri 8859 17815 8979 17935 ne
rect 8979 17815 9015 17935
rect 9135 17815 9171 17935
rect 8566 17678 8796 17760
tri 8796 17678 8878 17760 sw
tri 8979 17678 9116 17815 ne
rect 9116 17760 9171 17815
tri 9171 17760 9346 17935 sw
tri 9409 17815 9529 17935 ne
rect 9529 17815 9565 17935
rect 9685 17815 9721 17935
rect 9116 17678 9346 17760
tri 9346 17678 9428 17760 sw
tri 9529 17678 9666 17815 ne
rect 9666 17760 9721 17815
tri 9721 17760 9896 17935 sw
tri 9959 17815 10079 17935 ne
rect 10079 17815 10115 17935
rect 10235 17815 10271 17935
rect 9666 17678 9896 17760
tri 9896 17678 9978 17760 sw
tri 10079 17678 10216 17815 ne
rect 10216 17760 10271 17815
tri 10271 17760 10446 17935 sw
tri 10509 17815 10629 17935 ne
rect 10629 17815 10665 17935
rect 10785 17815 10821 17935
rect 10216 17678 10446 17760
tri 10446 17678 10528 17760 sw
tri 10629 17678 10766 17815 ne
rect 10766 17760 10821 17815
tri 10821 17760 10996 17935 sw
tri 11059 17815 11179 17935 ne
rect 11179 17815 11215 17935
rect 11335 17815 11371 17935
rect 10766 17678 10996 17760
tri 10996 17678 11078 17760 sw
tri 11179 17678 11316 17815 ne
rect 11316 17760 11371 17815
tri 11371 17760 11546 17935 sw
tri 11609 17815 11729 17935 ne
rect 11729 17815 11765 17935
rect 11885 17815 11921 17935
rect 11316 17678 11546 17760
tri 11546 17678 11628 17760 sw
tri 11729 17678 11866 17815 ne
rect 11866 17760 11921 17815
tri 11921 17760 12096 17935 sw
tri 12159 17815 12279 17935 ne
rect 12279 17815 12315 17935
rect 12435 17815 12471 17935
rect 11866 17678 12096 17760
tri 12096 17678 12178 17760 sw
tri 12279 17678 12416 17815 ne
rect 12416 17760 12471 17815
tri 12471 17760 12646 17935 sw
tri 12709 17815 12829 17935 ne
rect 12829 17815 12865 17935
rect 12985 17815 13021 17935
rect 12416 17678 12646 17760
tri 12646 17678 12728 17760 sw
tri 12829 17678 12966 17815 ne
rect 12966 17760 13021 17815
tri 13021 17760 13196 17935 sw
tri 13259 17815 13379 17935 ne
rect 13379 17815 13415 17935
rect 13535 17815 13571 17935
rect 12966 17678 13196 17760
tri 13196 17678 13278 17760 sw
tri 13379 17678 13516 17815 ne
rect 13516 17760 13571 17815
tri 13571 17760 13746 17935 sw
tri 13809 17815 13929 17935 ne
rect 13929 17815 13965 17935
rect 14085 17815 14121 17935
rect 13516 17678 13746 17760
tri 13746 17678 13828 17760 sw
tri 13929 17678 14066 17815 ne
rect 14066 17760 14121 17815
tri 14121 17760 14296 17935 sw
tri 14359 17815 14479 17935 ne
rect 14479 17815 14515 17935
rect 14635 17815 14671 17935
rect 14066 17678 14296 17760
tri 14296 17678 14378 17760 sw
tri 14479 17678 14616 17815 ne
rect 14616 17760 14671 17815
tri 14671 17760 14846 17935 sw
tri 14909 17815 15029 17935 ne
rect 15029 17815 15065 17935
rect 15185 17815 15221 17935
rect 14616 17678 14846 17760
tri 14846 17678 14928 17760 sw
tri 15029 17678 15166 17815 ne
rect 15166 17760 15221 17815
tri 15221 17760 15396 17935 sw
tri 15459 17815 15579 17935 ne
rect 15579 17815 15615 17935
rect 15735 17815 15771 17935
rect 15166 17678 15396 17760
tri 15396 17678 15478 17760 sw
tri 15579 17678 15716 17815 ne
rect 15716 17760 15771 17815
tri 15771 17760 15946 17935 sw
tri 16009 17815 16129 17935 ne
rect 16129 17815 16165 17935
rect 16285 17815 16321 17935
rect 15716 17678 15946 17760
tri 15946 17678 16028 17760 sw
tri 16129 17678 16266 17815 ne
rect 16266 17760 16321 17815
tri 16321 17760 16496 17935 sw
tri 16559 17815 16679 17935 ne
rect 16679 17815 16715 17935
rect 16835 17815 16871 17935
rect 16266 17678 16496 17760
tri 16496 17678 16578 17760 sw
tri 16679 17678 16816 17815 ne
rect 16816 17760 16871 17815
tri 16871 17760 17046 17935 sw
tri 17109 17815 17229 17935 ne
rect 17229 17815 17265 17935
rect 17385 17815 17421 17935
rect 16816 17678 17046 17760
tri 17046 17678 17128 17760 sw
tri 17229 17678 17366 17815 ne
rect 17366 17760 17421 17815
tri 17421 17760 17596 17935 sw
tri 17659 17815 17779 17935 ne
rect 17779 17815 17815 17935
rect 17935 17815 17971 17935
rect 17366 17678 17596 17760
tri 17596 17678 17678 17760 sw
tri 17779 17678 17916 17815 ne
rect 17916 17760 17971 17815
tri 17971 17760 18146 17935 sw
tri 18209 17815 18329 17935 ne
rect 18329 17815 18365 17935
rect 18485 17815 18521 17935
rect 17916 17678 18146 17760
tri 18146 17678 18228 17760 sw
tri 18329 17678 18466 17815 ne
rect 18466 17760 18521 17815
tri 18521 17760 18696 17935 sw
tri 18759 17815 18879 17935 ne
rect 18879 17815 18915 17935
rect 19035 17815 19071 17935
rect 18466 17678 18696 17760
tri 18696 17678 18778 17760 sw
tri 18879 17678 19016 17815 ne
rect 19016 17760 19071 17815
tri 19071 17760 19246 17935 sw
tri 19309 17815 19429 17935 ne
rect 19429 17815 19465 17935
rect 19585 17833 19621 17935
tri 19621 17833 19723 17935 sw
rect 19585 17815 20300 17833
rect 19016 17678 19246 17760
tri 19246 17678 19328 17760 sw
tri 19429 17678 19566 17815 ne
rect 19566 17678 20300 17815
rect -2000 17522 78 17678
tri 78 17522 234 17678 sw
tri 316 17522 472 17678 ne
rect 472 17522 628 17678
tri 628 17522 784 17678 sw
tri 866 17522 1022 17678 ne
rect 1022 17522 1178 17678
tri 1178 17522 1334 17678 sw
tri 1416 17522 1572 17678 ne
rect 1572 17522 1728 17678
tri 1728 17522 1884 17678 sw
tri 1966 17522 2122 17678 ne
rect 2122 17522 2278 17678
tri 2278 17522 2434 17678 sw
tri 2516 17522 2672 17678 ne
rect 2672 17522 2828 17678
tri 2828 17522 2984 17678 sw
tri 3066 17522 3222 17678 ne
rect 3222 17522 3378 17678
tri 3378 17522 3534 17678 sw
tri 3616 17522 3772 17678 ne
rect 3772 17522 3928 17678
tri 3928 17522 4084 17678 sw
tri 4166 17522 4322 17678 ne
rect 4322 17522 4478 17678
tri 4478 17522 4634 17678 sw
tri 4716 17522 4872 17678 ne
rect 4872 17522 5028 17678
tri 5028 17522 5184 17678 sw
tri 5266 17522 5422 17678 ne
rect 5422 17522 5578 17678
tri 5578 17522 5734 17678 sw
tri 5816 17522 5972 17678 ne
rect 5972 17522 6128 17678
tri 6128 17522 6284 17678 sw
tri 6366 17522 6522 17678 ne
rect 6522 17522 6678 17678
tri 6678 17522 6834 17678 sw
tri 6916 17522 7072 17678 ne
rect 7072 17522 7228 17678
tri 7228 17522 7384 17678 sw
tri 7466 17522 7622 17678 ne
rect 7622 17522 7778 17678
tri 7778 17522 7934 17678 sw
tri 8016 17522 8172 17678 ne
rect 8172 17522 8328 17678
tri 8328 17522 8484 17678 sw
tri 8566 17522 8722 17678 ne
rect 8722 17522 8878 17678
tri 8878 17522 9034 17678 sw
tri 9116 17522 9272 17678 ne
rect 9272 17522 9428 17678
tri 9428 17522 9584 17678 sw
tri 9666 17522 9822 17678 ne
rect 9822 17522 9978 17678
tri 9978 17522 10134 17678 sw
tri 10216 17522 10372 17678 ne
rect 10372 17522 10528 17678
tri 10528 17522 10684 17678 sw
tri 10766 17522 10922 17678 ne
rect 10922 17522 11078 17678
tri 11078 17522 11234 17678 sw
tri 11316 17522 11472 17678 ne
rect 11472 17522 11628 17678
tri 11628 17522 11784 17678 sw
tri 11866 17522 12022 17678 ne
rect 12022 17522 12178 17678
tri 12178 17522 12334 17678 sw
tri 12416 17522 12572 17678 ne
rect 12572 17522 12728 17678
tri 12728 17522 12884 17678 sw
tri 12966 17522 13122 17678 ne
rect 13122 17522 13278 17678
tri 13278 17522 13434 17678 sw
tri 13516 17522 13672 17678 ne
rect 13672 17522 13828 17678
tri 13828 17522 13984 17678 sw
tri 14066 17522 14222 17678 ne
rect 14222 17522 14378 17678
tri 14378 17522 14534 17678 sw
tri 14616 17522 14772 17678 ne
rect 14772 17522 14928 17678
tri 14928 17522 15084 17678 sw
tri 15166 17522 15322 17678 ne
rect 15322 17522 15478 17678
tri 15478 17522 15634 17678 sw
tri 15716 17522 15872 17678 ne
rect 15872 17522 16028 17678
tri 16028 17522 16184 17678 sw
tri 16266 17522 16422 17678 ne
rect 16422 17522 16578 17678
tri 16578 17522 16734 17678 sw
tri 16816 17522 16972 17678 ne
rect 16972 17522 17128 17678
tri 17128 17522 17284 17678 sw
tri 17366 17522 17522 17678 ne
rect 17522 17522 17678 17678
tri 17678 17522 17834 17678 sw
tri 17916 17522 18072 17678 ne
rect 18072 17522 18228 17678
tri 18228 17522 18384 17678 sw
tri 18466 17522 18622 17678 ne
rect 18622 17522 18778 17678
tri 18778 17522 18934 17678 sw
tri 19016 17522 19172 17678 ne
rect 19172 17522 19328 17678
tri 19328 17522 19484 17678 sw
tri 19566 17522 19722 17678 ne
rect 19722 17522 20300 17678
rect -2000 17385 234 17522
tri 234 17385 371 17522 sw
tri 472 17385 609 17522 ne
rect 609 17385 784 17522
tri 784 17385 921 17522 sw
tri 1022 17385 1159 17522 ne
rect 1159 17385 1334 17522
tri 1334 17385 1471 17522 sw
tri 1572 17385 1709 17522 ne
rect 1709 17385 1884 17522
tri 1884 17385 2021 17522 sw
tri 2122 17385 2259 17522 ne
rect 2259 17385 2434 17522
tri 2434 17385 2571 17522 sw
tri 2672 17385 2809 17522 ne
rect 2809 17385 2984 17522
tri 2984 17385 3121 17522 sw
tri 3222 17385 3359 17522 ne
rect 3359 17385 3534 17522
tri 3534 17385 3671 17522 sw
tri 3772 17385 3909 17522 ne
rect 3909 17385 4084 17522
tri 4084 17385 4221 17522 sw
tri 4322 17385 4459 17522 ne
rect 4459 17385 4634 17522
tri 4634 17385 4771 17522 sw
tri 4872 17385 5009 17522 ne
rect 5009 17385 5184 17522
tri 5184 17385 5321 17522 sw
tri 5422 17385 5559 17522 ne
rect 5559 17385 5734 17522
tri 5734 17385 5871 17522 sw
tri 5972 17385 6109 17522 ne
rect 6109 17385 6284 17522
tri 6284 17385 6421 17522 sw
tri 6522 17385 6659 17522 ne
rect 6659 17385 6834 17522
tri 6834 17385 6971 17522 sw
tri 7072 17385 7209 17522 ne
rect 7209 17385 7384 17522
tri 7384 17385 7521 17522 sw
tri 7622 17385 7759 17522 ne
rect 7759 17385 7934 17522
tri 7934 17385 8071 17522 sw
tri 8172 17385 8309 17522 ne
rect 8309 17385 8484 17522
tri 8484 17385 8621 17522 sw
tri 8722 17385 8859 17522 ne
rect 8859 17385 9034 17522
tri 9034 17385 9171 17522 sw
tri 9272 17385 9409 17522 ne
rect 9409 17385 9584 17522
tri 9584 17385 9721 17522 sw
tri 9822 17385 9959 17522 ne
rect 9959 17385 10134 17522
tri 10134 17385 10271 17522 sw
tri 10372 17385 10509 17522 ne
rect 10509 17385 10684 17522
tri 10684 17385 10821 17522 sw
tri 10922 17385 11059 17522 ne
rect 11059 17385 11234 17522
tri 11234 17385 11371 17522 sw
tri 11472 17385 11609 17522 ne
rect 11609 17385 11784 17522
tri 11784 17385 11921 17522 sw
tri 12022 17385 12159 17522 ne
rect 12159 17385 12334 17522
tri 12334 17385 12471 17522 sw
tri 12572 17385 12709 17522 ne
rect 12709 17385 12884 17522
tri 12884 17385 13021 17522 sw
tri 13122 17385 13259 17522 ne
rect 13259 17385 13434 17522
tri 13434 17385 13571 17522 sw
tri 13672 17385 13809 17522 ne
rect 13809 17385 13984 17522
tri 13984 17385 14121 17522 sw
tri 14222 17385 14359 17522 ne
rect 14359 17385 14534 17522
tri 14534 17385 14671 17522 sw
tri 14772 17385 14909 17522 ne
rect 14909 17385 15084 17522
tri 15084 17385 15221 17522 sw
tri 15322 17385 15459 17522 ne
rect 15459 17385 15634 17522
tri 15634 17385 15771 17522 sw
tri 15872 17385 16009 17522 ne
rect 16009 17385 16184 17522
tri 16184 17385 16321 17522 sw
tri 16422 17385 16559 17522 ne
rect 16559 17385 16734 17522
tri 16734 17385 16871 17522 sw
tri 16972 17385 17109 17522 ne
rect 17109 17385 17284 17522
tri 17284 17385 17421 17522 sw
tri 17522 17385 17659 17522 ne
rect 17659 17385 17834 17522
tri 17834 17385 17971 17522 sw
tri 18072 17385 18209 17522 ne
rect 18209 17385 18384 17522
tri 18384 17385 18521 17522 sw
tri 18622 17385 18759 17522 ne
rect 18759 17385 18934 17522
tri 18934 17385 19071 17522 sw
tri 19172 17385 19309 17522 ne
rect 19309 17385 19484 17522
tri 19484 17385 19621 17522 sw
rect -2000 17367 215 17385
rect -2000 16578 -1000 17367
tri 77 17265 179 17367 ne
rect 179 17265 215 17367
rect 335 17265 371 17385
tri 179 17128 316 17265 ne
rect 316 17210 371 17265
tri 371 17210 546 17385 sw
tri 609 17265 729 17385 ne
rect 729 17265 765 17385
rect 885 17265 921 17385
rect 316 17128 546 17210
tri 546 17128 628 17210 sw
tri 729 17128 866 17265 ne
rect 866 17210 921 17265
tri 921 17210 1096 17385 sw
tri 1159 17265 1279 17385 ne
rect 1279 17265 1315 17385
rect 1435 17265 1471 17385
rect 866 17128 1096 17210
tri 1096 17128 1178 17210 sw
tri 1279 17128 1416 17265 ne
rect 1416 17210 1471 17265
tri 1471 17210 1646 17385 sw
tri 1709 17265 1829 17385 ne
rect 1829 17265 1865 17385
rect 1985 17265 2021 17385
rect 1416 17128 1646 17210
tri 1646 17128 1728 17210 sw
tri 1829 17128 1966 17265 ne
rect 1966 17210 2021 17265
tri 2021 17210 2196 17385 sw
tri 2259 17265 2379 17385 ne
rect 2379 17265 2415 17385
rect 2535 17265 2571 17385
rect 1966 17128 2196 17210
tri 2196 17128 2278 17210 sw
tri 2379 17128 2516 17265 ne
rect 2516 17210 2571 17265
tri 2571 17210 2746 17385 sw
tri 2809 17265 2929 17385 ne
rect 2929 17265 2965 17385
rect 3085 17265 3121 17385
rect 2516 17128 2746 17210
tri 2746 17128 2828 17210 sw
tri 2929 17128 3066 17265 ne
rect 3066 17210 3121 17265
tri 3121 17210 3296 17385 sw
tri 3359 17265 3479 17385 ne
rect 3479 17265 3515 17385
rect 3635 17265 3671 17385
rect 3066 17128 3296 17210
tri 3296 17128 3378 17210 sw
tri 3479 17128 3616 17265 ne
rect 3616 17210 3671 17265
tri 3671 17210 3846 17385 sw
tri 3909 17265 4029 17385 ne
rect 4029 17265 4065 17385
rect 4185 17265 4221 17385
rect 3616 17128 3846 17210
tri 3846 17128 3928 17210 sw
tri 4029 17128 4166 17265 ne
rect 4166 17210 4221 17265
tri 4221 17210 4396 17385 sw
tri 4459 17265 4579 17385 ne
rect 4579 17265 4615 17385
rect 4735 17265 4771 17385
rect 4166 17128 4396 17210
tri 4396 17128 4478 17210 sw
tri 4579 17128 4716 17265 ne
rect 4716 17210 4771 17265
tri 4771 17210 4946 17385 sw
tri 5009 17265 5129 17385 ne
rect 5129 17265 5165 17385
rect 5285 17265 5321 17385
rect 4716 17128 4946 17210
tri 4946 17128 5028 17210 sw
tri 5129 17128 5266 17265 ne
rect 5266 17210 5321 17265
tri 5321 17210 5496 17385 sw
tri 5559 17265 5679 17385 ne
rect 5679 17265 5715 17385
rect 5835 17265 5871 17385
rect 5266 17128 5496 17210
tri 5496 17128 5578 17210 sw
tri 5679 17128 5816 17265 ne
rect 5816 17210 5871 17265
tri 5871 17210 6046 17385 sw
tri 6109 17265 6229 17385 ne
rect 6229 17265 6265 17385
rect 6385 17265 6421 17385
rect 5816 17128 6046 17210
tri 6046 17128 6128 17210 sw
tri 6229 17128 6366 17265 ne
rect 6366 17210 6421 17265
tri 6421 17210 6596 17385 sw
tri 6659 17265 6779 17385 ne
rect 6779 17265 6815 17385
rect 6935 17265 6971 17385
rect 6366 17128 6596 17210
tri 6596 17128 6678 17210 sw
tri 6779 17128 6916 17265 ne
rect 6916 17210 6971 17265
tri 6971 17210 7146 17385 sw
tri 7209 17265 7329 17385 ne
rect 7329 17265 7365 17385
rect 7485 17265 7521 17385
rect 6916 17128 7146 17210
tri 7146 17128 7228 17210 sw
tri 7329 17128 7466 17265 ne
rect 7466 17210 7521 17265
tri 7521 17210 7696 17385 sw
tri 7759 17265 7879 17385 ne
rect 7879 17265 7915 17385
rect 8035 17265 8071 17385
rect 7466 17128 7696 17210
tri 7696 17128 7778 17210 sw
tri 7879 17128 8016 17265 ne
rect 8016 17210 8071 17265
tri 8071 17210 8246 17385 sw
tri 8309 17265 8429 17385 ne
rect 8429 17265 8465 17385
rect 8585 17265 8621 17385
rect 8016 17128 8246 17210
tri 8246 17128 8328 17210 sw
tri 8429 17128 8566 17265 ne
rect 8566 17210 8621 17265
tri 8621 17210 8796 17385 sw
tri 8859 17265 8979 17385 ne
rect 8979 17265 9015 17385
rect 9135 17265 9171 17385
rect 8566 17128 8796 17210
tri 8796 17128 8878 17210 sw
tri 8979 17128 9116 17265 ne
rect 9116 17210 9171 17265
tri 9171 17210 9346 17385 sw
tri 9409 17265 9529 17385 ne
rect 9529 17265 9565 17385
rect 9685 17265 9721 17385
rect 9116 17128 9346 17210
tri 9346 17128 9428 17210 sw
tri 9529 17128 9666 17265 ne
rect 9666 17210 9721 17265
tri 9721 17210 9896 17385 sw
tri 9959 17265 10079 17385 ne
rect 10079 17265 10115 17385
rect 10235 17265 10271 17385
rect 9666 17128 9896 17210
tri 9896 17128 9978 17210 sw
tri 10079 17128 10216 17265 ne
rect 10216 17210 10271 17265
tri 10271 17210 10446 17385 sw
tri 10509 17265 10629 17385 ne
rect 10629 17265 10665 17385
rect 10785 17265 10821 17385
rect 10216 17128 10446 17210
tri 10446 17128 10528 17210 sw
tri 10629 17128 10766 17265 ne
rect 10766 17210 10821 17265
tri 10821 17210 10996 17385 sw
tri 11059 17265 11179 17385 ne
rect 11179 17265 11215 17385
rect 11335 17265 11371 17385
rect 10766 17128 10996 17210
tri 10996 17128 11078 17210 sw
tri 11179 17128 11316 17265 ne
rect 11316 17210 11371 17265
tri 11371 17210 11546 17385 sw
tri 11609 17265 11729 17385 ne
rect 11729 17265 11765 17385
rect 11885 17265 11921 17385
rect 11316 17128 11546 17210
tri 11546 17128 11628 17210 sw
tri 11729 17128 11866 17265 ne
rect 11866 17210 11921 17265
tri 11921 17210 12096 17385 sw
tri 12159 17265 12279 17385 ne
rect 12279 17265 12315 17385
rect 12435 17265 12471 17385
rect 11866 17128 12096 17210
tri 12096 17128 12178 17210 sw
tri 12279 17128 12416 17265 ne
rect 12416 17210 12471 17265
tri 12471 17210 12646 17385 sw
tri 12709 17265 12829 17385 ne
rect 12829 17265 12865 17385
rect 12985 17265 13021 17385
rect 12416 17128 12646 17210
tri 12646 17128 12728 17210 sw
tri 12829 17128 12966 17265 ne
rect 12966 17210 13021 17265
tri 13021 17210 13196 17385 sw
tri 13259 17265 13379 17385 ne
rect 13379 17265 13415 17385
rect 13535 17265 13571 17385
rect 12966 17128 13196 17210
tri 13196 17128 13278 17210 sw
tri 13379 17128 13516 17265 ne
rect 13516 17210 13571 17265
tri 13571 17210 13746 17385 sw
tri 13809 17265 13929 17385 ne
rect 13929 17265 13965 17385
rect 14085 17265 14121 17385
rect 13516 17128 13746 17210
tri 13746 17128 13828 17210 sw
tri 13929 17128 14066 17265 ne
rect 14066 17210 14121 17265
tri 14121 17210 14296 17385 sw
tri 14359 17265 14479 17385 ne
rect 14479 17265 14515 17385
rect 14635 17265 14671 17385
rect 14066 17128 14296 17210
tri 14296 17128 14378 17210 sw
tri 14479 17128 14616 17265 ne
rect 14616 17210 14671 17265
tri 14671 17210 14846 17385 sw
tri 14909 17265 15029 17385 ne
rect 15029 17265 15065 17385
rect 15185 17265 15221 17385
rect 14616 17128 14846 17210
tri 14846 17128 14928 17210 sw
tri 15029 17128 15166 17265 ne
rect 15166 17210 15221 17265
tri 15221 17210 15396 17385 sw
tri 15459 17265 15579 17385 ne
rect 15579 17265 15615 17385
rect 15735 17265 15771 17385
rect 15166 17128 15396 17210
tri 15396 17128 15478 17210 sw
tri 15579 17128 15716 17265 ne
rect 15716 17210 15771 17265
tri 15771 17210 15946 17385 sw
tri 16009 17265 16129 17385 ne
rect 16129 17265 16165 17385
rect 16285 17265 16321 17385
rect 15716 17128 15946 17210
tri 15946 17128 16028 17210 sw
tri 16129 17128 16266 17265 ne
rect 16266 17210 16321 17265
tri 16321 17210 16496 17385 sw
tri 16559 17265 16679 17385 ne
rect 16679 17265 16715 17385
rect 16835 17265 16871 17385
rect 16266 17128 16496 17210
tri 16496 17128 16578 17210 sw
tri 16679 17128 16816 17265 ne
rect 16816 17210 16871 17265
tri 16871 17210 17046 17385 sw
tri 17109 17265 17229 17385 ne
rect 17229 17265 17265 17385
rect 17385 17265 17421 17385
rect 16816 17128 17046 17210
tri 17046 17128 17128 17210 sw
tri 17229 17128 17366 17265 ne
rect 17366 17210 17421 17265
tri 17421 17210 17596 17385 sw
tri 17659 17265 17779 17385 ne
rect 17779 17265 17815 17385
rect 17935 17265 17971 17385
rect 17366 17128 17596 17210
tri 17596 17128 17678 17210 sw
tri 17779 17128 17916 17265 ne
rect 17916 17210 17971 17265
tri 17971 17210 18146 17385 sw
tri 18209 17265 18329 17385 ne
rect 18329 17265 18365 17385
rect 18485 17265 18521 17385
rect 17916 17128 18146 17210
tri 18146 17128 18228 17210 sw
tri 18329 17128 18466 17265 ne
rect 18466 17210 18521 17265
tri 18521 17210 18696 17385 sw
tri 18759 17265 18879 17385 ne
rect 18879 17265 18915 17385
rect 19035 17265 19071 17385
rect 18466 17128 18696 17210
tri 18696 17128 18778 17210 sw
tri 18879 17128 19016 17265 ne
rect 19016 17210 19071 17265
tri 19071 17210 19246 17385 sw
tri 19309 17265 19429 17385 ne
rect 19429 17265 19465 17385
rect 19585 17283 19621 17385
tri 19621 17283 19723 17385 sw
rect 20800 17283 21800 18072
rect 19585 17265 21800 17283
rect 19016 17128 19246 17210
tri 19246 17128 19328 17210 sw
tri 19429 17128 19566 17265 ne
rect 19566 17128 21800 17265
rect -500 16972 78 17128
tri 78 16972 234 17128 sw
tri 316 16972 472 17128 ne
rect 472 16972 628 17128
tri 628 16972 784 17128 sw
tri 866 16972 1022 17128 ne
rect 1022 16972 1178 17128
tri 1178 16972 1334 17128 sw
tri 1416 16972 1572 17128 ne
rect 1572 16972 1728 17128
tri 1728 16972 1884 17128 sw
tri 1966 16972 2122 17128 ne
rect 2122 16972 2278 17128
tri 2278 16972 2434 17128 sw
tri 2516 16972 2672 17128 ne
rect 2672 16972 2828 17128
tri 2828 16972 2984 17128 sw
tri 3066 16972 3222 17128 ne
rect 3222 16972 3378 17128
tri 3378 16972 3534 17128 sw
tri 3616 16972 3772 17128 ne
rect 3772 16972 3928 17128
tri 3928 16972 4084 17128 sw
tri 4166 16972 4322 17128 ne
rect 4322 16972 4478 17128
tri 4478 16972 4634 17128 sw
tri 4716 16972 4872 17128 ne
rect 4872 16972 5028 17128
tri 5028 16972 5184 17128 sw
tri 5266 16972 5422 17128 ne
rect 5422 16972 5578 17128
tri 5578 16972 5734 17128 sw
tri 5816 16972 5972 17128 ne
rect 5972 16972 6128 17128
tri 6128 16972 6284 17128 sw
tri 6366 16972 6522 17128 ne
rect 6522 16972 6678 17128
tri 6678 16972 6834 17128 sw
tri 6916 16972 7072 17128 ne
rect 7072 16972 7228 17128
tri 7228 16972 7384 17128 sw
tri 7466 16972 7622 17128 ne
rect 7622 16972 7778 17128
tri 7778 16972 7934 17128 sw
tri 8016 16972 8172 17128 ne
rect 8172 16972 8328 17128
tri 8328 16972 8484 17128 sw
tri 8566 16972 8722 17128 ne
rect 8722 16972 8878 17128
tri 8878 16972 9034 17128 sw
tri 9116 16972 9272 17128 ne
rect 9272 16972 9428 17128
tri 9428 16972 9584 17128 sw
tri 9666 16972 9822 17128 ne
rect 9822 16972 9978 17128
tri 9978 16972 10134 17128 sw
tri 10216 16972 10372 17128 ne
rect 10372 16972 10528 17128
tri 10528 16972 10684 17128 sw
tri 10766 16972 10922 17128 ne
rect 10922 16972 11078 17128
tri 11078 16972 11234 17128 sw
tri 11316 16972 11472 17128 ne
rect 11472 16972 11628 17128
tri 11628 16972 11784 17128 sw
tri 11866 16972 12022 17128 ne
rect 12022 16972 12178 17128
tri 12178 16972 12334 17128 sw
tri 12416 16972 12572 17128 ne
rect 12572 16972 12728 17128
tri 12728 16972 12884 17128 sw
tri 12966 16972 13122 17128 ne
rect 13122 16972 13278 17128
tri 13278 16972 13434 17128 sw
tri 13516 16972 13672 17128 ne
rect 13672 16972 13828 17128
tri 13828 16972 13984 17128 sw
tri 14066 16972 14222 17128 ne
rect 14222 16972 14378 17128
tri 14378 16972 14534 17128 sw
tri 14616 16972 14772 17128 ne
rect 14772 16972 14928 17128
tri 14928 16972 15084 17128 sw
tri 15166 16972 15322 17128 ne
rect 15322 16972 15478 17128
tri 15478 16972 15634 17128 sw
tri 15716 16972 15872 17128 ne
rect 15872 16972 16028 17128
tri 16028 16972 16184 17128 sw
tri 16266 16972 16422 17128 ne
rect 16422 16972 16578 17128
tri 16578 16972 16734 17128 sw
tri 16816 16972 16972 17128 ne
rect 16972 16972 17128 17128
tri 17128 16972 17284 17128 sw
tri 17366 16972 17522 17128 ne
rect 17522 16972 17678 17128
tri 17678 16972 17834 17128 sw
tri 17916 16972 18072 17128 ne
rect 18072 16972 18228 17128
tri 18228 16972 18384 17128 sw
tri 18466 16972 18622 17128 ne
rect 18622 16972 18778 17128
tri 18778 16972 18934 17128 sw
tri 19016 16972 19172 17128 ne
rect 19172 16972 19328 17128
tri 19328 16972 19484 17128 sw
tri 19566 16972 19722 17128 ne
rect 19722 16972 21800 17128
rect -500 16835 234 16972
tri 234 16835 371 16972 sw
tri 472 16835 609 16972 ne
rect 609 16835 784 16972
tri 784 16835 921 16972 sw
tri 1022 16835 1159 16972 ne
rect 1159 16835 1334 16972
tri 1334 16835 1471 16972 sw
tri 1572 16835 1709 16972 ne
rect 1709 16835 1884 16972
tri 1884 16835 2021 16972 sw
tri 2122 16835 2259 16972 ne
rect 2259 16835 2434 16972
tri 2434 16835 2571 16972 sw
tri 2672 16835 2809 16972 ne
rect 2809 16835 2984 16972
tri 2984 16835 3121 16972 sw
tri 3222 16835 3359 16972 ne
rect 3359 16835 3534 16972
tri 3534 16835 3671 16972 sw
tri 3772 16835 3909 16972 ne
rect 3909 16835 4084 16972
tri 4084 16835 4221 16972 sw
tri 4322 16835 4459 16972 ne
rect 4459 16835 4634 16972
tri 4634 16835 4771 16972 sw
tri 4872 16835 5009 16972 ne
rect 5009 16835 5184 16972
tri 5184 16835 5321 16972 sw
tri 5422 16835 5559 16972 ne
rect 5559 16835 5734 16972
tri 5734 16835 5871 16972 sw
tri 5972 16835 6109 16972 ne
rect 6109 16835 6284 16972
tri 6284 16835 6421 16972 sw
tri 6522 16835 6659 16972 ne
rect 6659 16835 6834 16972
tri 6834 16835 6971 16972 sw
tri 7072 16835 7209 16972 ne
rect 7209 16835 7384 16972
tri 7384 16835 7521 16972 sw
tri 7622 16835 7759 16972 ne
rect 7759 16835 7934 16972
tri 7934 16835 8071 16972 sw
tri 8172 16835 8309 16972 ne
rect 8309 16835 8484 16972
tri 8484 16835 8621 16972 sw
tri 8722 16835 8859 16972 ne
rect 8859 16835 9034 16972
tri 9034 16835 9171 16972 sw
tri 9272 16835 9409 16972 ne
rect 9409 16835 9584 16972
tri 9584 16835 9721 16972 sw
tri 9822 16835 9959 16972 ne
rect 9959 16835 10134 16972
tri 10134 16835 10271 16972 sw
tri 10372 16835 10509 16972 ne
rect 10509 16835 10684 16972
tri 10684 16835 10821 16972 sw
tri 10922 16835 11059 16972 ne
rect 11059 16835 11234 16972
tri 11234 16835 11371 16972 sw
tri 11472 16835 11609 16972 ne
rect 11609 16835 11784 16972
tri 11784 16835 11921 16972 sw
tri 12022 16835 12159 16972 ne
rect 12159 16835 12334 16972
tri 12334 16835 12471 16972 sw
tri 12572 16835 12709 16972 ne
rect 12709 16835 12884 16972
tri 12884 16835 13021 16972 sw
tri 13122 16835 13259 16972 ne
rect 13259 16835 13434 16972
tri 13434 16835 13571 16972 sw
tri 13672 16835 13809 16972 ne
rect 13809 16835 13984 16972
tri 13984 16835 14121 16972 sw
tri 14222 16835 14359 16972 ne
rect 14359 16835 14534 16972
tri 14534 16835 14671 16972 sw
tri 14772 16835 14909 16972 ne
rect 14909 16835 15084 16972
tri 15084 16835 15221 16972 sw
tri 15322 16835 15459 16972 ne
rect 15459 16835 15634 16972
tri 15634 16835 15771 16972 sw
tri 15872 16835 16009 16972 ne
rect 16009 16835 16184 16972
tri 16184 16835 16321 16972 sw
tri 16422 16835 16559 16972 ne
rect 16559 16835 16734 16972
tri 16734 16835 16871 16972 sw
tri 16972 16835 17109 16972 ne
rect 17109 16835 17284 16972
tri 17284 16835 17421 16972 sw
tri 17522 16835 17659 16972 ne
rect 17659 16835 17834 16972
tri 17834 16835 17971 16972 sw
tri 18072 16835 18209 16972 ne
rect 18209 16835 18384 16972
tri 18384 16835 18521 16972 sw
tri 18622 16835 18759 16972 ne
rect 18759 16835 18934 16972
tri 18934 16835 19071 16972 sw
tri 19172 16835 19309 16972 ne
rect 19309 16835 19484 16972
tri 19484 16835 19621 16972 sw
rect -500 16817 215 16835
tri 77 16715 179 16817 ne
rect 179 16715 215 16817
rect 335 16715 371 16835
tri 179 16578 316 16715 ne
rect 316 16660 371 16715
tri 371 16660 546 16835 sw
tri 609 16715 729 16835 ne
rect 729 16715 765 16835
rect 885 16715 921 16835
rect 316 16578 546 16660
tri 546 16578 628 16660 sw
tri 729 16578 866 16715 ne
rect 866 16660 921 16715
tri 921 16660 1096 16835 sw
tri 1159 16715 1279 16835 ne
rect 1279 16715 1315 16835
rect 1435 16715 1471 16835
rect 866 16578 1096 16660
tri 1096 16578 1178 16660 sw
tri 1279 16578 1416 16715 ne
rect 1416 16660 1471 16715
tri 1471 16660 1646 16835 sw
tri 1709 16715 1829 16835 ne
rect 1829 16715 1865 16835
rect 1985 16715 2021 16835
rect 1416 16578 1646 16660
tri 1646 16578 1728 16660 sw
tri 1829 16578 1966 16715 ne
rect 1966 16660 2021 16715
tri 2021 16660 2196 16835 sw
tri 2259 16715 2379 16835 ne
rect 2379 16715 2415 16835
rect 2535 16715 2571 16835
rect 1966 16578 2196 16660
tri 2196 16578 2278 16660 sw
tri 2379 16578 2516 16715 ne
rect 2516 16660 2571 16715
tri 2571 16660 2746 16835 sw
tri 2809 16715 2929 16835 ne
rect 2929 16715 2965 16835
rect 3085 16715 3121 16835
rect 2516 16578 2746 16660
tri 2746 16578 2828 16660 sw
tri 2929 16578 3066 16715 ne
rect 3066 16660 3121 16715
tri 3121 16660 3296 16835 sw
tri 3359 16715 3479 16835 ne
rect 3479 16715 3515 16835
rect 3635 16715 3671 16835
rect 3066 16578 3296 16660
tri 3296 16578 3378 16660 sw
tri 3479 16578 3616 16715 ne
rect 3616 16660 3671 16715
tri 3671 16660 3846 16835 sw
tri 3909 16715 4029 16835 ne
rect 4029 16715 4065 16835
rect 4185 16715 4221 16835
rect 3616 16578 3846 16660
tri 3846 16578 3928 16660 sw
tri 4029 16578 4166 16715 ne
rect 4166 16660 4221 16715
tri 4221 16660 4396 16835 sw
tri 4459 16715 4579 16835 ne
rect 4579 16715 4615 16835
rect 4735 16715 4771 16835
rect 4166 16578 4396 16660
tri 4396 16578 4478 16660 sw
tri 4579 16578 4716 16715 ne
rect 4716 16660 4771 16715
tri 4771 16660 4946 16835 sw
tri 5009 16715 5129 16835 ne
rect 5129 16715 5165 16835
rect 5285 16715 5321 16835
rect 4716 16578 4946 16660
tri 4946 16578 5028 16660 sw
tri 5129 16578 5266 16715 ne
rect 5266 16660 5321 16715
tri 5321 16660 5496 16835 sw
tri 5559 16715 5679 16835 ne
rect 5679 16715 5715 16835
rect 5835 16715 5871 16835
rect 5266 16578 5496 16660
tri 5496 16578 5578 16660 sw
tri 5679 16578 5816 16715 ne
rect 5816 16660 5871 16715
tri 5871 16660 6046 16835 sw
tri 6109 16715 6229 16835 ne
rect 6229 16715 6265 16835
rect 6385 16715 6421 16835
rect 5816 16578 6046 16660
tri 6046 16578 6128 16660 sw
tri 6229 16578 6366 16715 ne
rect 6366 16660 6421 16715
tri 6421 16660 6596 16835 sw
tri 6659 16715 6779 16835 ne
rect 6779 16715 6815 16835
rect 6935 16715 6971 16835
rect 6366 16578 6596 16660
tri 6596 16578 6678 16660 sw
tri 6779 16578 6916 16715 ne
rect 6916 16660 6971 16715
tri 6971 16660 7146 16835 sw
tri 7209 16715 7329 16835 ne
rect 7329 16715 7365 16835
rect 7485 16715 7521 16835
rect 6916 16578 7146 16660
tri 7146 16578 7228 16660 sw
tri 7329 16578 7466 16715 ne
rect 7466 16660 7521 16715
tri 7521 16660 7696 16835 sw
tri 7759 16715 7879 16835 ne
rect 7879 16715 7915 16835
rect 8035 16715 8071 16835
rect 7466 16578 7696 16660
tri 7696 16578 7778 16660 sw
tri 7879 16578 8016 16715 ne
rect 8016 16660 8071 16715
tri 8071 16660 8246 16835 sw
tri 8309 16715 8429 16835 ne
rect 8429 16715 8465 16835
rect 8585 16715 8621 16835
rect 8016 16578 8246 16660
tri 8246 16578 8328 16660 sw
tri 8429 16578 8566 16715 ne
rect 8566 16660 8621 16715
tri 8621 16660 8796 16835 sw
tri 8859 16715 8979 16835 ne
rect 8979 16715 9015 16835
rect 9135 16715 9171 16835
rect 8566 16578 8796 16660
tri 8796 16578 8878 16660 sw
tri 8979 16578 9116 16715 ne
rect 9116 16660 9171 16715
tri 9171 16660 9346 16835 sw
tri 9409 16715 9529 16835 ne
rect 9529 16715 9565 16835
rect 9685 16715 9721 16835
rect 9116 16578 9346 16660
tri 9346 16578 9428 16660 sw
tri 9529 16578 9666 16715 ne
rect 9666 16660 9721 16715
tri 9721 16660 9896 16835 sw
tri 9959 16715 10079 16835 ne
rect 10079 16715 10115 16835
rect 10235 16715 10271 16835
rect 9666 16578 9896 16660
tri 9896 16578 9978 16660 sw
tri 10079 16578 10216 16715 ne
rect 10216 16660 10271 16715
tri 10271 16660 10446 16835 sw
tri 10509 16715 10629 16835 ne
rect 10629 16715 10665 16835
rect 10785 16715 10821 16835
rect 10216 16578 10446 16660
tri 10446 16578 10528 16660 sw
tri 10629 16578 10766 16715 ne
rect 10766 16660 10821 16715
tri 10821 16660 10996 16835 sw
tri 11059 16715 11179 16835 ne
rect 11179 16715 11215 16835
rect 11335 16715 11371 16835
rect 10766 16578 10996 16660
tri 10996 16578 11078 16660 sw
tri 11179 16578 11316 16715 ne
rect 11316 16660 11371 16715
tri 11371 16660 11546 16835 sw
tri 11609 16715 11729 16835 ne
rect 11729 16715 11765 16835
rect 11885 16715 11921 16835
rect 11316 16578 11546 16660
tri 11546 16578 11628 16660 sw
tri 11729 16578 11866 16715 ne
rect 11866 16660 11921 16715
tri 11921 16660 12096 16835 sw
tri 12159 16715 12279 16835 ne
rect 12279 16715 12315 16835
rect 12435 16715 12471 16835
rect 11866 16578 12096 16660
tri 12096 16578 12178 16660 sw
tri 12279 16578 12416 16715 ne
rect 12416 16660 12471 16715
tri 12471 16660 12646 16835 sw
tri 12709 16715 12829 16835 ne
rect 12829 16715 12865 16835
rect 12985 16715 13021 16835
rect 12416 16578 12646 16660
tri 12646 16578 12728 16660 sw
tri 12829 16578 12966 16715 ne
rect 12966 16660 13021 16715
tri 13021 16660 13196 16835 sw
tri 13259 16715 13379 16835 ne
rect 13379 16715 13415 16835
rect 13535 16715 13571 16835
rect 12966 16578 13196 16660
tri 13196 16578 13278 16660 sw
tri 13379 16578 13516 16715 ne
rect 13516 16660 13571 16715
tri 13571 16660 13746 16835 sw
tri 13809 16715 13929 16835 ne
rect 13929 16715 13965 16835
rect 14085 16715 14121 16835
rect 13516 16578 13746 16660
tri 13746 16578 13828 16660 sw
tri 13929 16578 14066 16715 ne
rect 14066 16660 14121 16715
tri 14121 16660 14296 16835 sw
tri 14359 16715 14479 16835 ne
rect 14479 16715 14515 16835
rect 14635 16715 14671 16835
rect 14066 16578 14296 16660
tri 14296 16578 14378 16660 sw
tri 14479 16578 14616 16715 ne
rect 14616 16660 14671 16715
tri 14671 16660 14846 16835 sw
tri 14909 16715 15029 16835 ne
rect 15029 16715 15065 16835
rect 15185 16715 15221 16835
rect 14616 16578 14846 16660
tri 14846 16578 14928 16660 sw
tri 15029 16578 15166 16715 ne
rect 15166 16660 15221 16715
tri 15221 16660 15396 16835 sw
tri 15459 16715 15579 16835 ne
rect 15579 16715 15615 16835
rect 15735 16715 15771 16835
rect 15166 16578 15396 16660
tri 15396 16578 15478 16660 sw
tri 15579 16578 15716 16715 ne
rect 15716 16660 15771 16715
tri 15771 16660 15946 16835 sw
tri 16009 16715 16129 16835 ne
rect 16129 16715 16165 16835
rect 16285 16715 16321 16835
rect 15716 16578 15946 16660
tri 15946 16578 16028 16660 sw
tri 16129 16578 16266 16715 ne
rect 16266 16660 16321 16715
tri 16321 16660 16496 16835 sw
tri 16559 16715 16679 16835 ne
rect 16679 16715 16715 16835
rect 16835 16715 16871 16835
rect 16266 16578 16496 16660
tri 16496 16578 16578 16660 sw
tri 16679 16578 16816 16715 ne
rect 16816 16660 16871 16715
tri 16871 16660 17046 16835 sw
tri 17109 16715 17229 16835 ne
rect 17229 16715 17265 16835
rect 17385 16715 17421 16835
rect 16816 16578 17046 16660
tri 17046 16578 17128 16660 sw
tri 17229 16578 17366 16715 ne
rect 17366 16660 17421 16715
tri 17421 16660 17596 16835 sw
tri 17659 16715 17779 16835 ne
rect 17779 16715 17815 16835
rect 17935 16715 17971 16835
rect 17366 16578 17596 16660
tri 17596 16578 17678 16660 sw
tri 17779 16578 17916 16715 ne
rect 17916 16660 17971 16715
tri 17971 16660 18146 16835 sw
tri 18209 16715 18329 16835 ne
rect 18329 16715 18365 16835
rect 18485 16715 18521 16835
rect 17916 16578 18146 16660
tri 18146 16578 18228 16660 sw
tri 18329 16578 18466 16715 ne
rect 18466 16660 18521 16715
tri 18521 16660 18696 16835 sw
tri 18759 16715 18879 16835 ne
rect 18879 16715 18915 16835
rect 19035 16715 19071 16835
rect 18466 16578 18696 16660
tri 18696 16578 18778 16660 sw
tri 18879 16578 19016 16715 ne
rect 19016 16660 19071 16715
tri 19071 16660 19246 16835 sw
tri 19309 16715 19429 16835 ne
rect 19429 16715 19465 16835
rect 19585 16733 19621 16835
tri 19621 16733 19723 16835 sw
rect 19585 16715 20300 16733
rect 19016 16578 19246 16660
tri 19246 16578 19328 16660 sw
tri 19429 16578 19566 16715 ne
rect 19566 16578 20300 16715
rect -2000 16422 78 16578
tri 78 16422 234 16578 sw
tri 316 16422 472 16578 ne
rect 472 16422 628 16578
tri 628 16422 784 16578 sw
tri 866 16422 1022 16578 ne
rect 1022 16422 1178 16578
tri 1178 16422 1334 16578 sw
tri 1416 16422 1572 16578 ne
rect 1572 16422 1728 16578
tri 1728 16422 1884 16578 sw
tri 1966 16422 2122 16578 ne
rect 2122 16422 2278 16578
tri 2278 16422 2434 16578 sw
tri 2516 16422 2672 16578 ne
rect 2672 16422 2828 16578
tri 2828 16422 2984 16578 sw
tri 3066 16422 3222 16578 ne
rect 3222 16422 3378 16578
tri 3378 16422 3534 16578 sw
tri 3616 16422 3772 16578 ne
rect 3772 16422 3928 16578
tri 3928 16422 4084 16578 sw
tri 4166 16422 4322 16578 ne
rect 4322 16422 4478 16578
tri 4478 16422 4634 16578 sw
tri 4716 16422 4872 16578 ne
rect 4872 16422 5028 16578
tri 5028 16422 5184 16578 sw
tri 5266 16422 5422 16578 ne
rect 5422 16422 5578 16578
tri 5578 16422 5734 16578 sw
tri 5816 16422 5972 16578 ne
rect 5972 16422 6128 16578
tri 6128 16422 6284 16578 sw
tri 6366 16422 6522 16578 ne
rect 6522 16422 6678 16578
tri 6678 16422 6834 16578 sw
tri 6916 16422 7072 16578 ne
rect 7072 16422 7228 16578
tri 7228 16422 7384 16578 sw
tri 7466 16422 7622 16578 ne
rect 7622 16422 7778 16578
tri 7778 16422 7934 16578 sw
tri 8016 16422 8172 16578 ne
rect 8172 16422 8328 16578
tri 8328 16422 8484 16578 sw
tri 8566 16422 8722 16578 ne
rect 8722 16422 8878 16578
tri 8878 16422 9034 16578 sw
tri 9116 16422 9272 16578 ne
rect 9272 16422 9428 16578
tri 9428 16422 9584 16578 sw
tri 9666 16422 9822 16578 ne
rect 9822 16422 9978 16578
tri 9978 16422 10134 16578 sw
tri 10216 16422 10372 16578 ne
rect 10372 16422 10528 16578
tri 10528 16422 10684 16578 sw
tri 10766 16422 10922 16578 ne
rect 10922 16422 11078 16578
tri 11078 16422 11234 16578 sw
tri 11316 16422 11472 16578 ne
rect 11472 16422 11628 16578
tri 11628 16422 11784 16578 sw
tri 11866 16422 12022 16578 ne
rect 12022 16422 12178 16578
tri 12178 16422 12334 16578 sw
tri 12416 16422 12572 16578 ne
rect 12572 16422 12728 16578
tri 12728 16422 12884 16578 sw
tri 12966 16422 13122 16578 ne
rect 13122 16422 13278 16578
tri 13278 16422 13434 16578 sw
tri 13516 16422 13672 16578 ne
rect 13672 16422 13828 16578
tri 13828 16422 13984 16578 sw
tri 14066 16422 14222 16578 ne
rect 14222 16422 14378 16578
tri 14378 16422 14534 16578 sw
tri 14616 16422 14772 16578 ne
rect 14772 16422 14928 16578
tri 14928 16422 15084 16578 sw
tri 15166 16422 15322 16578 ne
rect 15322 16422 15478 16578
tri 15478 16422 15634 16578 sw
tri 15716 16422 15872 16578 ne
rect 15872 16422 16028 16578
tri 16028 16422 16184 16578 sw
tri 16266 16422 16422 16578 ne
rect 16422 16422 16578 16578
tri 16578 16422 16734 16578 sw
tri 16816 16422 16972 16578 ne
rect 16972 16422 17128 16578
tri 17128 16422 17284 16578 sw
tri 17366 16422 17522 16578 ne
rect 17522 16422 17678 16578
tri 17678 16422 17834 16578 sw
tri 17916 16422 18072 16578 ne
rect 18072 16422 18228 16578
tri 18228 16422 18384 16578 sw
tri 18466 16422 18622 16578 ne
rect 18622 16422 18778 16578
tri 18778 16422 18934 16578 sw
tri 19016 16422 19172 16578 ne
rect 19172 16422 19328 16578
tri 19328 16422 19484 16578 sw
tri 19566 16422 19722 16578 ne
rect 19722 16422 20300 16578
rect -2000 16285 234 16422
tri 234 16285 371 16422 sw
tri 472 16285 609 16422 ne
rect 609 16285 784 16422
tri 784 16285 921 16422 sw
tri 1022 16285 1159 16422 ne
rect 1159 16285 1334 16422
tri 1334 16285 1471 16422 sw
tri 1572 16285 1709 16422 ne
rect 1709 16285 1884 16422
tri 1884 16285 2021 16422 sw
tri 2122 16285 2259 16422 ne
rect 2259 16285 2434 16422
tri 2434 16285 2571 16422 sw
tri 2672 16285 2809 16422 ne
rect 2809 16285 2984 16422
tri 2984 16285 3121 16422 sw
tri 3222 16285 3359 16422 ne
rect 3359 16285 3534 16422
tri 3534 16285 3671 16422 sw
tri 3772 16285 3909 16422 ne
rect 3909 16285 4084 16422
tri 4084 16285 4221 16422 sw
tri 4322 16285 4459 16422 ne
rect 4459 16285 4634 16422
tri 4634 16285 4771 16422 sw
tri 4872 16285 5009 16422 ne
rect 5009 16285 5184 16422
tri 5184 16285 5321 16422 sw
tri 5422 16285 5559 16422 ne
rect 5559 16285 5734 16422
tri 5734 16285 5871 16422 sw
tri 5972 16285 6109 16422 ne
rect 6109 16285 6284 16422
tri 6284 16285 6421 16422 sw
tri 6522 16285 6659 16422 ne
rect 6659 16285 6834 16422
tri 6834 16285 6971 16422 sw
tri 7072 16285 7209 16422 ne
rect 7209 16285 7384 16422
tri 7384 16285 7521 16422 sw
tri 7622 16285 7759 16422 ne
rect 7759 16285 7934 16422
tri 7934 16285 8071 16422 sw
tri 8172 16285 8309 16422 ne
rect 8309 16285 8484 16422
tri 8484 16285 8621 16422 sw
tri 8722 16285 8859 16422 ne
rect 8859 16285 9034 16422
tri 9034 16285 9171 16422 sw
tri 9272 16285 9409 16422 ne
rect 9409 16285 9584 16422
tri 9584 16285 9721 16422 sw
tri 9822 16285 9959 16422 ne
rect 9959 16285 10134 16422
tri 10134 16285 10271 16422 sw
tri 10372 16285 10509 16422 ne
rect 10509 16285 10684 16422
tri 10684 16285 10821 16422 sw
tri 10922 16285 11059 16422 ne
rect 11059 16285 11234 16422
tri 11234 16285 11371 16422 sw
tri 11472 16285 11609 16422 ne
rect 11609 16285 11784 16422
tri 11784 16285 11921 16422 sw
tri 12022 16285 12159 16422 ne
rect 12159 16285 12334 16422
tri 12334 16285 12471 16422 sw
tri 12572 16285 12709 16422 ne
rect 12709 16285 12884 16422
tri 12884 16285 13021 16422 sw
tri 13122 16285 13259 16422 ne
rect 13259 16285 13434 16422
tri 13434 16285 13571 16422 sw
tri 13672 16285 13809 16422 ne
rect 13809 16285 13984 16422
tri 13984 16285 14121 16422 sw
tri 14222 16285 14359 16422 ne
rect 14359 16285 14534 16422
tri 14534 16285 14671 16422 sw
tri 14772 16285 14909 16422 ne
rect 14909 16285 15084 16422
tri 15084 16285 15221 16422 sw
tri 15322 16285 15459 16422 ne
rect 15459 16285 15634 16422
tri 15634 16285 15771 16422 sw
tri 15872 16285 16009 16422 ne
rect 16009 16285 16184 16422
tri 16184 16285 16321 16422 sw
tri 16422 16285 16559 16422 ne
rect 16559 16285 16734 16422
tri 16734 16285 16871 16422 sw
tri 16972 16285 17109 16422 ne
rect 17109 16285 17284 16422
tri 17284 16285 17421 16422 sw
tri 17522 16285 17659 16422 ne
rect 17659 16285 17834 16422
tri 17834 16285 17971 16422 sw
tri 18072 16285 18209 16422 ne
rect 18209 16285 18384 16422
tri 18384 16285 18521 16422 sw
tri 18622 16285 18759 16422 ne
rect 18759 16285 18934 16422
tri 18934 16285 19071 16422 sw
tri 19172 16285 19309 16422 ne
rect 19309 16285 19484 16422
tri 19484 16285 19621 16422 sw
rect -2000 16267 215 16285
rect -2000 15478 -1000 16267
tri 77 16165 179 16267 ne
rect 179 16165 215 16267
rect 335 16165 371 16285
tri 179 16028 316 16165 ne
rect 316 16110 371 16165
tri 371 16110 546 16285 sw
tri 609 16165 729 16285 ne
rect 729 16165 765 16285
rect 885 16165 921 16285
rect 316 16028 546 16110
tri 546 16028 628 16110 sw
tri 729 16028 866 16165 ne
rect 866 16110 921 16165
tri 921 16110 1096 16285 sw
tri 1159 16165 1279 16285 ne
rect 1279 16165 1315 16285
rect 1435 16165 1471 16285
rect 866 16028 1096 16110
tri 1096 16028 1178 16110 sw
tri 1279 16028 1416 16165 ne
rect 1416 16110 1471 16165
tri 1471 16110 1646 16285 sw
tri 1709 16165 1829 16285 ne
rect 1829 16165 1865 16285
rect 1985 16165 2021 16285
rect 1416 16028 1646 16110
tri 1646 16028 1728 16110 sw
tri 1829 16028 1966 16165 ne
rect 1966 16110 2021 16165
tri 2021 16110 2196 16285 sw
tri 2259 16165 2379 16285 ne
rect 2379 16165 2415 16285
rect 2535 16165 2571 16285
rect 1966 16028 2196 16110
tri 2196 16028 2278 16110 sw
tri 2379 16028 2516 16165 ne
rect 2516 16110 2571 16165
tri 2571 16110 2746 16285 sw
tri 2809 16165 2929 16285 ne
rect 2929 16165 2965 16285
rect 3085 16165 3121 16285
rect 2516 16028 2746 16110
tri 2746 16028 2828 16110 sw
tri 2929 16028 3066 16165 ne
rect 3066 16110 3121 16165
tri 3121 16110 3296 16285 sw
tri 3359 16165 3479 16285 ne
rect 3479 16165 3515 16285
rect 3635 16165 3671 16285
rect 3066 16028 3296 16110
tri 3296 16028 3378 16110 sw
tri 3479 16028 3616 16165 ne
rect 3616 16110 3671 16165
tri 3671 16110 3846 16285 sw
tri 3909 16165 4029 16285 ne
rect 4029 16165 4065 16285
rect 4185 16165 4221 16285
rect 3616 16028 3846 16110
tri 3846 16028 3928 16110 sw
tri 4029 16028 4166 16165 ne
rect 4166 16110 4221 16165
tri 4221 16110 4396 16285 sw
tri 4459 16165 4579 16285 ne
rect 4579 16165 4615 16285
rect 4735 16165 4771 16285
rect 4166 16028 4396 16110
tri 4396 16028 4478 16110 sw
tri 4579 16028 4716 16165 ne
rect 4716 16110 4771 16165
tri 4771 16110 4946 16285 sw
tri 5009 16165 5129 16285 ne
rect 5129 16165 5165 16285
rect 5285 16165 5321 16285
rect 4716 16028 4946 16110
tri 4946 16028 5028 16110 sw
tri 5129 16028 5266 16165 ne
rect 5266 16110 5321 16165
tri 5321 16110 5496 16285 sw
tri 5559 16165 5679 16285 ne
rect 5679 16165 5715 16285
rect 5835 16165 5871 16285
rect 5266 16028 5496 16110
tri 5496 16028 5578 16110 sw
tri 5679 16028 5816 16165 ne
rect 5816 16110 5871 16165
tri 5871 16110 6046 16285 sw
tri 6109 16165 6229 16285 ne
rect 6229 16165 6265 16285
rect 6385 16165 6421 16285
rect 5816 16028 6046 16110
tri 6046 16028 6128 16110 sw
tri 6229 16028 6366 16165 ne
rect 6366 16110 6421 16165
tri 6421 16110 6596 16285 sw
tri 6659 16165 6779 16285 ne
rect 6779 16165 6815 16285
rect 6935 16165 6971 16285
rect 6366 16028 6596 16110
tri 6596 16028 6678 16110 sw
tri 6779 16028 6916 16165 ne
rect 6916 16110 6971 16165
tri 6971 16110 7146 16285 sw
tri 7209 16165 7329 16285 ne
rect 7329 16165 7365 16285
rect 7485 16165 7521 16285
rect 6916 16028 7146 16110
tri 7146 16028 7228 16110 sw
tri 7329 16028 7466 16165 ne
rect 7466 16110 7521 16165
tri 7521 16110 7696 16285 sw
tri 7759 16165 7879 16285 ne
rect 7879 16165 7915 16285
rect 8035 16165 8071 16285
rect 7466 16028 7696 16110
tri 7696 16028 7778 16110 sw
tri 7879 16028 8016 16165 ne
rect 8016 16110 8071 16165
tri 8071 16110 8246 16285 sw
tri 8309 16165 8429 16285 ne
rect 8429 16165 8465 16285
rect 8585 16165 8621 16285
rect 8016 16028 8246 16110
tri 8246 16028 8328 16110 sw
tri 8429 16028 8566 16165 ne
rect 8566 16110 8621 16165
tri 8621 16110 8796 16285 sw
tri 8859 16165 8979 16285 ne
rect 8979 16165 9015 16285
rect 9135 16165 9171 16285
rect 8566 16028 8796 16110
tri 8796 16028 8878 16110 sw
tri 8979 16028 9116 16165 ne
rect 9116 16110 9171 16165
tri 9171 16110 9346 16285 sw
tri 9409 16165 9529 16285 ne
rect 9529 16165 9565 16285
rect 9685 16165 9721 16285
rect 9116 16028 9346 16110
tri 9346 16028 9428 16110 sw
tri 9529 16028 9666 16165 ne
rect 9666 16110 9721 16165
tri 9721 16110 9896 16285 sw
tri 9959 16165 10079 16285 ne
rect 10079 16165 10115 16285
rect 10235 16165 10271 16285
rect 9666 16028 9896 16110
tri 9896 16028 9978 16110 sw
tri 10079 16028 10216 16165 ne
rect 10216 16110 10271 16165
tri 10271 16110 10446 16285 sw
tri 10509 16165 10629 16285 ne
rect 10629 16165 10665 16285
rect 10785 16165 10821 16285
rect 10216 16028 10446 16110
tri 10446 16028 10528 16110 sw
tri 10629 16028 10766 16165 ne
rect 10766 16110 10821 16165
tri 10821 16110 10996 16285 sw
tri 11059 16165 11179 16285 ne
rect 11179 16165 11215 16285
rect 11335 16165 11371 16285
rect 10766 16028 10996 16110
tri 10996 16028 11078 16110 sw
tri 11179 16028 11316 16165 ne
rect 11316 16110 11371 16165
tri 11371 16110 11546 16285 sw
tri 11609 16165 11729 16285 ne
rect 11729 16165 11765 16285
rect 11885 16165 11921 16285
rect 11316 16028 11546 16110
tri 11546 16028 11628 16110 sw
tri 11729 16028 11866 16165 ne
rect 11866 16110 11921 16165
tri 11921 16110 12096 16285 sw
tri 12159 16165 12279 16285 ne
rect 12279 16165 12315 16285
rect 12435 16165 12471 16285
rect 11866 16028 12096 16110
tri 12096 16028 12178 16110 sw
tri 12279 16028 12416 16165 ne
rect 12416 16110 12471 16165
tri 12471 16110 12646 16285 sw
tri 12709 16165 12829 16285 ne
rect 12829 16165 12865 16285
rect 12985 16165 13021 16285
rect 12416 16028 12646 16110
tri 12646 16028 12728 16110 sw
tri 12829 16028 12966 16165 ne
rect 12966 16110 13021 16165
tri 13021 16110 13196 16285 sw
tri 13259 16165 13379 16285 ne
rect 13379 16165 13415 16285
rect 13535 16165 13571 16285
rect 12966 16028 13196 16110
tri 13196 16028 13278 16110 sw
tri 13379 16028 13516 16165 ne
rect 13516 16110 13571 16165
tri 13571 16110 13746 16285 sw
tri 13809 16165 13929 16285 ne
rect 13929 16165 13965 16285
rect 14085 16165 14121 16285
rect 13516 16028 13746 16110
tri 13746 16028 13828 16110 sw
tri 13929 16028 14066 16165 ne
rect 14066 16110 14121 16165
tri 14121 16110 14296 16285 sw
tri 14359 16165 14479 16285 ne
rect 14479 16165 14515 16285
rect 14635 16165 14671 16285
rect 14066 16028 14296 16110
tri 14296 16028 14378 16110 sw
tri 14479 16028 14616 16165 ne
rect 14616 16110 14671 16165
tri 14671 16110 14846 16285 sw
tri 14909 16165 15029 16285 ne
rect 15029 16165 15065 16285
rect 15185 16165 15221 16285
rect 14616 16028 14846 16110
tri 14846 16028 14928 16110 sw
tri 15029 16028 15166 16165 ne
rect 15166 16110 15221 16165
tri 15221 16110 15396 16285 sw
tri 15459 16165 15579 16285 ne
rect 15579 16165 15615 16285
rect 15735 16165 15771 16285
rect 15166 16028 15396 16110
tri 15396 16028 15478 16110 sw
tri 15579 16028 15716 16165 ne
rect 15716 16110 15771 16165
tri 15771 16110 15946 16285 sw
tri 16009 16165 16129 16285 ne
rect 16129 16165 16165 16285
rect 16285 16165 16321 16285
rect 15716 16028 15946 16110
tri 15946 16028 16028 16110 sw
tri 16129 16028 16266 16165 ne
rect 16266 16110 16321 16165
tri 16321 16110 16496 16285 sw
tri 16559 16165 16679 16285 ne
rect 16679 16165 16715 16285
rect 16835 16165 16871 16285
rect 16266 16028 16496 16110
tri 16496 16028 16578 16110 sw
tri 16679 16028 16816 16165 ne
rect 16816 16110 16871 16165
tri 16871 16110 17046 16285 sw
tri 17109 16165 17229 16285 ne
rect 17229 16165 17265 16285
rect 17385 16165 17421 16285
rect 16816 16028 17046 16110
tri 17046 16028 17128 16110 sw
tri 17229 16028 17366 16165 ne
rect 17366 16110 17421 16165
tri 17421 16110 17596 16285 sw
tri 17659 16165 17779 16285 ne
rect 17779 16165 17815 16285
rect 17935 16165 17971 16285
rect 17366 16028 17596 16110
tri 17596 16028 17678 16110 sw
tri 17779 16028 17916 16165 ne
rect 17916 16110 17971 16165
tri 17971 16110 18146 16285 sw
tri 18209 16165 18329 16285 ne
rect 18329 16165 18365 16285
rect 18485 16165 18521 16285
rect 17916 16028 18146 16110
tri 18146 16028 18228 16110 sw
tri 18329 16028 18466 16165 ne
rect 18466 16110 18521 16165
tri 18521 16110 18696 16285 sw
tri 18759 16165 18879 16285 ne
rect 18879 16165 18915 16285
rect 19035 16165 19071 16285
rect 18466 16028 18696 16110
tri 18696 16028 18778 16110 sw
tri 18879 16028 19016 16165 ne
rect 19016 16110 19071 16165
tri 19071 16110 19246 16285 sw
tri 19309 16165 19429 16285 ne
rect 19429 16165 19465 16285
rect 19585 16183 19621 16285
tri 19621 16183 19723 16285 sw
rect 20800 16183 21800 16972
rect 19585 16165 21800 16183
rect 19016 16028 19246 16110
tri 19246 16028 19328 16110 sw
tri 19429 16028 19566 16165 ne
rect 19566 16028 21800 16165
rect -500 15872 78 16028
tri 78 15872 234 16028 sw
tri 316 15872 472 16028 ne
rect 472 15872 628 16028
tri 628 15872 784 16028 sw
tri 866 15872 1022 16028 ne
rect 1022 15872 1178 16028
tri 1178 15872 1334 16028 sw
tri 1416 15872 1572 16028 ne
rect 1572 15872 1728 16028
tri 1728 15872 1884 16028 sw
tri 1966 15872 2122 16028 ne
rect 2122 15872 2278 16028
tri 2278 15872 2434 16028 sw
tri 2516 15872 2672 16028 ne
rect 2672 15872 2828 16028
tri 2828 15872 2984 16028 sw
tri 3066 15872 3222 16028 ne
rect 3222 15872 3378 16028
tri 3378 15872 3534 16028 sw
tri 3616 15872 3772 16028 ne
rect 3772 15872 3928 16028
tri 3928 15872 4084 16028 sw
tri 4166 15872 4322 16028 ne
rect 4322 15872 4478 16028
tri 4478 15872 4634 16028 sw
tri 4716 15872 4872 16028 ne
rect 4872 15872 5028 16028
tri 5028 15872 5184 16028 sw
tri 5266 15872 5422 16028 ne
rect 5422 15872 5578 16028
tri 5578 15872 5734 16028 sw
tri 5816 15872 5972 16028 ne
rect 5972 15872 6128 16028
tri 6128 15872 6284 16028 sw
tri 6366 15872 6522 16028 ne
rect 6522 15872 6678 16028
tri 6678 15872 6834 16028 sw
tri 6916 15872 7072 16028 ne
rect 7072 15872 7228 16028
tri 7228 15872 7384 16028 sw
tri 7466 15872 7622 16028 ne
rect 7622 15872 7778 16028
tri 7778 15872 7934 16028 sw
tri 8016 15872 8172 16028 ne
rect 8172 15872 8328 16028
tri 8328 15872 8484 16028 sw
tri 8566 15872 8722 16028 ne
rect 8722 15872 8878 16028
tri 8878 15872 9034 16028 sw
tri 9116 15872 9272 16028 ne
rect 9272 15872 9428 16028
tri 9428 15872 9584 16028 sw
tri 9666 15872 9822 16028 ne
rect 9822 15872 9978 16028
tri 9978 15872 10134 16028 sw
tri 10216 15872 10372 16028 ne
rect 10372 15872 10528 16028
tri 10528 15872 10684 16028 sw
tri 10766 15872 10922 16028 ne
rect 10922 15872 11078 16028
tri 11078 15872 11234 16028 sw
tri 11316 15872 11472 16028 ne
rect 11472 15872 11628 16028
tri 11628 15872 11784 16028 sw
tri 11866 15872 12022 16028 ne
rect 12022 15872 12178 16028
tri 12178 15872 12334 16028 sw
tri 12416 15872 12572 16028 ne
rect 12572 15872 12728 16028
tri 12728 15872 12884 16028 sw
tri 12966 15872 13122 16028 ne
rect 13122 15872 13278 16028
tri 13278 15872 13434 16028 sw
tri 13516 15872 13672 16028 ne
rect 13672 15872 13828 16028
tri 13828 15872 13984 16028 sw
tri 14066 15872 14222 16028 ne
rect 14222 15872 14378 16028
tri 14378 15872 14534 16028 sw
tri 14616 15872 14772 16028 ne
rect 14772 15872 14928 16028
tri 14928 15872 15084 16028 sw
tri 15166 15872 15322 16028 ne
rect 15322 15872 15478 16028
tri 15478 15872 15634 16028 sw
tri 15716 15872 15872 16028 ne
rect 15872 15872 16028 16028
tri 16028 15872 16184 16028 sw
tri 16266 15872 16422 16028 ne
rect 16422 15872 16578 16028
tri 16578 15872 16734 16028 sw
tri 16816 15872 16972 16028 ne
rect 16972 15872 17128 16028
tri 17128 15872 17284 16028 sw
tri 17366 15872 17522 16028 ne
rect 17522 15872 17678 16028
tri 17678 15872 17834 16028 sw
tri 17916 15872 18072 16028 ne
rect 18072 15872 18228 16028
tri 18228 15872 18384 16028 sw
tri 18466 15872 18622 16028 ne
rect 18622 15872 18778 16028
tri 18778 15872 18934 16028 sw
tri 19016 15872 19172 16028 ne
rect 19172 15872 19328 16028
tri 19328 15872 19484 16028 sw
tri 19566 15872 19722 16028 ne
rect 19722 15872 21800 16028
rect -500 15735 234 15872
tri 234 15735 371 15872 sw
tri 472 15735 609 15872 ne
rect 609 15735 784 15872
tri 784 15735 921 15872 sw
tri 1022 15735 1159 15872 ne
rect 1159 15735 1334 15872
tri 1334 15735 1471 15872 sw
tri 1572 15735 1709 15872 ne
rect 1709 15735 1884 15872
tri 1884 15735 2021 15872 sw
tri 2122 15735 2259 15872 ne
rect 2259 15735 2434 15872
tri 2434 15735 2571 15872 sw
tri 2672 15735 2809 15872 ne
rect 2809 15735 2984 15872
tri 2984 15735 3121 15872 sw
tri 3222 15735 3359 15872 ne
rect 3359 15735 3534 15872
tri 3534 15735 3671 15872 sw
tri 3772 15735 3909 15872 ne
rect 3909 15735 4084 15872
tri 4084 15735 4221 15872 sw
tri 4322 15735 4459 15872 ne
rect 4459 15735 4634 15872
tri 4634 15735 4771 15872 sw
tri 4872 15735 5009 15872 ne
rect 5009 15735 5184 15872
tri 5184 15735 5321 15872 sw
tri 5422 15735 5559 15872 ne
rect 5559 15735 5734 15872
tri 5734 15735 5871 15872 sw
tri 5972 15735 6109 15872 ne
rect 6109 15735 6284 15872
tri 6284 15735 6421 15872 sw
tri 6522 15735 6659 15872 ne
rect 6659 15735 6834 15872
tri 6834 15735 6971 15872 sw
tri 7072 15735 7209 15872 ne
rect 7209 15735 7384 15872
tri 7384 15735 7521 15872 sw
tri 7622 15735 7759 15872 ne
rect 7759 15735 7934 15872
tri 7934 15735 8071 15872 sw
tri 8172 15735 8309 15872 ne
rect 8309 15735 8484 15872
tri 8484 15735 8621 15872 sw
tri 8722 15735 8859 15872 ne
rect 8859 15735 9034 15872
tri 9034 15735 9171 15872 sw
tri 9272 15735 9409 15872 ne
rect 9409 15735 9584 15872
tri 9584 15735 9721 15872 sw
tri 9822 15735 9959 15872 ne
rect 9959 15735 10134 15872
tri 10134 15735 10271 15872 sw
tri 10372 15735 10509 15872 ne
rect 10509 15735 10684 15872
tri 10684 15735 10821 15872 sw
tri 10922 15735 11059 15872 ne
rect 11059 15735 11234 15872
tri 11234 15735 11371 15872 sw
tri 11472 15735 11609 15872 ne
rect 11609 15735 11784 15872
tri 11784 15735 11921 15872 sw
tri 12022 15735 12159 15872 ne
rect 12159 15735 12334 15872
tri 12334 15735 12471 15872 sw
tri 12572 15735 12709 15872 ne
rect 12709 15735 12884 15872
tri 12884 15735 13021 15872 sw
tri 13122 15735 13259 15872 ne
rect 13259 15735 13434 15872
tri 13434 15735 13571 15872 sw
tri 13672 15735 13809 15872 ne
rect 13809 15735 13984 15872
tri 13984 15735 14121 15872 sw
tri 14222 15735 14359 15872 ne
rect 14359 15735 14534 15872
tri 14534 15735 14671 15872 sw
tri 14772 15735 14909 15872 ne
rect 14909 15735 15084 15872
tri 15084 15735 15221 15872 sw
tri 15322 15735 15459 15872 ne
rect 15459 15735 15634 15872
tri 15634 15735 15771 15872 sw
tri 15872 15735 16009 15872 ne
rect 16009 15735 16184 15872
tri 16184 15735 16321 15872 sw
tri 16422 15735 16559 15872 ne
rect 16559 15735 16734 15872
tri 16734 15735 16871 15872 sw
tri 16972 15735 17109 15872 ne
rect 17109 15735 17284 15872
tri 17284 15735 17421 15872 sw
tri 17522 15735 17659 15872 ne
rect 17659 15735 17834 15872
tri 17834 15735 17971 15872 sw
tri 18072 15735 18209 15872 ne
rect 18209 15735 18384 15872
tri 18384 15735 18521 15872 sw
tri 18622 15735 18759 15872 ne
rect 18759 15735 18934 15872
tri 18934 15735 19071 15872 sw
tri 19172 15735 19309 15872 ne
rect 19309 15735 19484 15872
tri 19484 15735 19621 15872 sw
rect -500 15717 215 15735
tri 77 15615 179 15717 ne
rect 179 15615 215 15717
rect 335 15615 371 15735
tri 179 15478 316 15615 ne
rect 316 15560 371 15615
tri 371 15560 546 15735 sw
tri 609 15615 729 15735 ne
rect 729 15615 765 15735
rect 885 15615 921 15735
rect 316 15478 546 15560
tri 546 15478 628 15560 sw
tri 729 15478 866 15615 ne
rect 866 15560 921 15615
tri 921 15560 1096 15735 sw
tri 1159 15615 1279 15735 ne
rect 1279 15615 1315 15735
rect 1435 15615 1471 15735
rect 866 15478 1096 15560
tri 1096 15478 1178 15560 sw
tri 1279 15478 1416 15615 ne
rect 1416 15560 1471 15615
tri 1471 15560 1646 15735 sw
tri 1709 15615 1829 15735 ne
rect 1829 15615 1865 15735
rect 1985 15615 2021 15735
rect 1416 15478 1646 15560
tri 1646 15478 1728 15560 sw
tri 1829 15478 1966 15615 ne
rect 1966 15560 2021 15615
tri 2021 15560 2196 15735 sw
tri 2259 15615 2379 15735 ne
rect 2379 15615 2415 15735
rect 2535 15615 2571 15735
rect 1966 15478 2196 15560
tri 2196 15478 2278 15560 sw
tri 2379 15478 2516 15615 ne
rect 2516 15560 2571 15615
tri 2571 15560 2746 15735 sw
tri 2809 15615 2929 15735 ne
rect 2929 15615 2965 15735
rect 3085 15615 3121 15735
rect 2516 15478 2746 15560
tri 2746 15478 2828 15560 sw
tri 2929 15478 3066 15615 ne
rect 3066 15560 3121 15615
tri 3121 15560 3296 15735 sw
tri 3359 15615 3479 15735 ne
rect 3479 15615 3515 15735
rect 3635 15615 3671 15735
rect 3066 15478 3296 15560
tri 3296 15478 3378 15560 sw
tri 3479 15478 3616 15615 ne
rect 3616 15560 3671 15615
tri 3671 15560 3846 15735 sw
tri 3909 15615 4029 15735 ne
rect 4029 15615 4065 15735
rect 4185 15615 4221 15735
rect 3616 15478 3846 15560
tri 3846 15478 3928 15560 sw
tri 4029 15478 4166 15615 ne
rect 4166 15560 4221 15615
tri 4221 15560 4396 15735 sw
tri 4459 15615 4579 15735 ne
rect 4579 15615 4615 15735
rect 4735 15615 4771 15735
rect 4166 15478 4396 15560
tri 4396 15478 4478 15560 sw
tri 4579 15478 4716 15615 ne
rect 4716 15560 4771 15615
tri 4771 15560 4946 15735 sw
tri 5009 15615 5129 15735 ne
rect 5129 15615 5165 15735
rect 5285 15615 5321 15735
rect 4716 15478 4946 15560
tri 4946 15478 5028 15560 sw
tri 5129 15478 5266 15615 ne
rect 5266 15560 5321 15615
tri 5321 15560 5496 15735 sw
tri 5559 15615 5679 15735 ne
rect 5679 15615 5715 15735
rect 5835 15615 5871 15735
rect 5266 15478 5496 15560
tri 5496 15478 5578 15560 sw
tri 5679 15478 5816 15615 ne
rect 5816 15560 5871 15615
tri 5871 15560 6046 15735 sw
tri 6109 15615 6229 15735 ne
rect 6229 15615 6265 15735
rect 6385 15615 6421 15735
rect 5816 15478 6046 15560
tri 6046 15478 6128 15560 sw
tri 6229 15478 6366 15615 ne
rect 6366 15560 6421 15615
tri 6421 15560 6596 15735 sw
tri 6659 15615 6779 15735 ne
rect 6779 15615 6815 15735
rect 6935 15615 6971 15735
rect 6366 15478 6596 15560
tri 6596 15478 6678 15560 sw
tri 6779 15478 6916 15615 ne
rect 6916 15560 6971 15615
tri 6971 15560 7146 15735 sw
tri 7209 15615 7329 15735 ne
rect 7329 15615 7365 15735
rect 7485 15615 7521 15735
rect 6916 15478 7146 15560
tri 7146 15478 7228 15560 sw
tri 7329 15478 7466 15615 ne
rect 7466 15560 7521 15615
tri 7521 15560 7696 15735 sw
tri 7759 15615 7879 15735 ne
rect 7879 15615 7915 15735
rect 8035 15615 8071 15735
rect 7466 15478 7696 15560
tri 7696 15478 7778 15560 sw
tri 7879 15478 8016 15615 ne
rect 8016 15560 8071 15615
tri 8071 15560 8246 15735 sw
tri 8309 15615 8429 15735 ne
rect 8429 15615 8465 15735
rect 8585 15615 8621 15735
rect 8016 15478 8246 15560
tri 8246 15478 8328 15560 sw
tri 8429 15478 8566 15615 ne
rect 8566 15560 8621 15615
tri 8621 15560 8796 15735 sw
tri 8859 15615 8979 15735 ne
rect 8979 15615 9015 15735
rect 9135 15615 9171 15735
rect 8566 15478 8796 15560
tri 8796 15478 8878 15560 sw
tri 8979 15478 9116 15615 ne
rect 9116 15560 9171 15615
tri 9171 15560 9346 15735 sw
tri 9409 15615 9529 15735 ne
rect 9529 15615 9565 15735
rect 9685 15615 9721 15735
rect 9116 15478 9346 15560
tri 9346 15478 9428 15560 sw
tri 9529 15478 9666 15615 ne
rect 9666 15560 9721 15615
tri 9721 15560 9896 15735 sw
tri 9959 15615 10079 15735 ne
rect 10079 15615 10115 15735
rect 10235 15615 10271 15735
rect 9666 15478 9896 15560
tri 9896 15478 9978 15560 sw
tri 10079 15478 10216 15615 ne
rect 10216 15560 10271 15615
tri 10271 15560 10446 15735 sw
tri 10509 15615 10629 15735 ne
rect 10629 15615 10665 15735
rect 10785 15615 10821 15735
rect 10216 15478 10446 15560
tri 10446 15478 10528 15560 sw
tri 10629 15478 10766 15615 ne
rect 10766 15560 10821 15615
tri 10821 15560 10996 15735 sw
tri 11059 15615 11179 15735 ne
rect 11179 15615 11215 15735
rect 11335 15615 11371 15735
rect 10766 15478 10996 15560
tri 10996 15478 11078 15560 sw
tri 11179 15478 11316 15615 ne
rect 11316 15560 11371 15615
tri 11371 15560 11546 15735 sw
tri 11609 15615 11729 15735 ne
rect 11729 15615 11765 15735
rect 11885 15615 11921 15735
rect 11316 15478 11546 15560
tri 11546 15478 11628 15560 sw
tri 11729 15478 11866 15615 ne
rect 11866 15560 11921 15615
tri 11921 15560 12096 15735 sw
tri 12159 15615 12279 15735 ne
rect 12279 15615 12315 15735
rect 12435 15615 12471 15735
rect 11866 15478 12096 15560
tri 12096 15478 12178 15560 sw
tri 12279 15478 12416 15615 ne
rect 12416 15560 12471 15615
tri 12471 15560 12646 15735 sw
tri 12709 15615 12829 15735 ne
rect 12829 15615 12865 15735
rect 12985 15615 13021 15735
rect 12416 15478 12646 15560
tri 12646 15478 12728 15560 sw
tri 12829 15478 12966 15615 ne
rect 12966 15560 13021 15615
tri 13021 15560 13196 15735 sw
tri 13259 15615 13379 15735 ne
rect 13379 15615 13415 15735
rect 13535 15615 13571 15735
rect 12966 15478 13196 15560
tri 13196 15478 13278 15560 sw
tri 13379 15478 13516 15615 ne
rect 13516 15560 13571 15615
tri 13571 15560 13746 15735 sw
tri 13809 15615 13929 15735 ne
rect 13929 15615 13965 15735
rect 14085 15615 14121 15735
rect 13516 15478 13746 15560
tri 13746 15478 13828 15560 sw
tri 13929 15478 14066 15615 ne
rect 14066 15560 14121 15615
tri 14121 15560 14296 15735 sw
tri 14359 15615 14479 15735 ne
rect 14479 15615 14515 15735
rect 14635 15615 14671 15735
rect 14066 15478 14296 15560
tri 14296 15478 14378 15560 sw
tri 14479 15478 14616 15615 ne
rect 14616 15560 14671 15615
tri 14671 15560 14846 15735 sw
tri 14909 15615 15029 15735 ne
rect 15029 15615 15065 15735
rect 15185 15615 15221 15735
rect 14616 15478 14846 15560
tri 14846 15478 14928 15560 sw
tri 15029 15478 15166 15615 ne
rect 15166 15560 15221 15615
tri 15221 15560 15396 15735 sw
tri 15459 15615 15579 15735 ne
rect 15579 15615 15615 15735
rect 15735 15615 15771 15735
rect 15166 15478 15396 15560
tri 15396 15478 15478 15560 sw
tri 15579 15478 15716 15615 ne
rect 15716 15560 15771 15615
tri 15771 15560 15946 15735 sw
tri 16009 15615 16129 15735 ne
rect 16129 15615 16165 15735
rect 16285 15615 16321 15735
rect 15716 15478 15946 15560
tri 15946 15478 16028 15560 sw
tri 16129 15478 16266 15615 ne
rect 16266 15560 16321 15615
tri 16321 15560 16496 15735 sw
tri 16559 15615 16679 15735 ne
rect 16679 15615 16715 15735
rect 16835 15615 16871 15735
rect 16266 15478 16496 15560
tri 16496 15478 16578 15560 sw
tri 16679 15478 16816 15615 ne
rect 16816 15560 16871 15615
tri 16871 15560 17046 15735 sw
tri 17109 15615 17229 15735 ne
rect 17229 15615 17265 15735
rect 17385 15615 17421 15735
rect 16816 15478 17046 15560
tri 17046 15478 17128 15560 sw
tri 17229 15478 17366 15615 ne
rect 17366 15560 17421 15615
tri 17421 15560 17596 15735 sw
tri 17659 15615 17779 15735 ne
rect 17779 15615 17815 15735
rect 17935 15615 17971 15735
rect 17366 15478 17596 15560
tri 17596 15478 17678 15560 sw
tri 17779 15478 17916 15615 ne
rect 17916 15560 17971 15615
tri 17971 15560 18146 15735 sw
tri 18209 15615 18329 15735 ne
rect 18329 15615 18365 15735
rect 18485 15615 18521 15735
rect 17916 15478 18146 15560
tri 18146 15478 18228 15560 sw
tri 18329 15478 18466 15615 ne
rect 18466 15560 18521 15615
tri 18521 15560 18696 15735 sw
tri 18759 15615 18879 15735 ne
rect 18879 15615 18915 15735
rect 19035 15615 19071 15735
rect 18466 15478 18696 15560
tri 18696 15478 18778 15560 sw
tri 18879 15478 19016 15615 ne
rect 19016 15560 19071 15615
tri 19071 15560 19246 15735 sw
tri 19309 15615 19429 15735 ne
rect 19429 15615 19465 15735
rect 19585 15633 19621 15735
tri 19621 15633 19723 15735 sw
rect 19585 15615 20300 15633
rect 19016 15478 19246 15560
tri 19246 15478 19328 15560 sw
tri 19429 15478 19566 15615 ne
rect 19566 15478 20300 15615
rect -2000 15322 78 15478
tri 78 15322 234 15478 sw
tri 316 15322 472 15478 ne
rect 472 15322 628 15478
tri 628 15322 784 15478 sw
tri 866 15322 1022 15478 ne
rect 1022 15322 1178 15478
tri 1178 15322 1334 15478 sw
tri 1416 15322 1572 15478 ne
rect 1572 15322 1728 15478
tri 1728 15322 1884 15478 sw
tri 1966 15322 2122 15478 ne
rect 2122 15322 2278 15478
tri 2278 15322 2434 15478 sw
tri 2516 15322 2672 15478 ne
rect 2672 15322 2828 15478
tri 2828 15322 2984 15478 sw
tri 3066 15322 3222 15478 ne
rect 3222 15322 3378 15478
tri 3378 15322 3534 15478 sw
tri 3616 15322 3772 15478 ne
rect 3772 15322 3928 15478
tri 3928 15322 4084 15478 sw
tri 4166 15322 4322 15478 ne
rect 4322 15322 4478 15478
tri 4478 15322 4634 15478 sw
tri 4716 15322 4872 15478 ne
rect 4872 15322 5028 15478
tri 5028 15322 5184 15478 sw
tri 5266 15322 5422 15478 ne
rect 5422 15322 5578 15478
tri 5578 15322 5734 15478 sw
tri 5816 15322 5972 15478 ne
rect 5972 15322 6128 15478
tri 6128 15322 6284 15478 sw
tri 6366 15322 6522 15478 ne
rect 6522 15322 6678 15478
tri 6678 15322 6834 15478 sw
tri 6916 15322 7072 15478 ne
rect 7072 15322 7228 15478
tri 7228 15322 7384 15478 sw
tri 7466 15322 7622 15478 ne
rect 7622 15322 7778 15478
tri 7778 15322 7934 15478 sw
tri 8016 15322 8172 15478 ne
rect 8172 15322 8328 15478
tri 8328 15322 8484 15478 sw
tri 8566 15322 8722 15478 ne
rect 8722 15322 8878 15478
tri 8878 15322 9034 15478 sw
tri 9116 15322 9272 15478 ne
rect 9272 15322 9428 15478
tri 9428 15322 9584 15478 sw
tri 9666 15322 9822 15478 ne
rect 9822 15322 9978 15478
tri 9978 15322 10134 15478 sw
tri 10216 15322 10372 15478 ne
rect 10372 15322 10528 15478
tri 10528 15322 10684 15478 sw
tri 10766 15322 10922 15478 ne
rect 10922 15322 11078 15478
tri 11078 15322 11234 15478 sw
tri 11316 15322 11472 15478 ne
rect 11472 15322 11628 15478
tri 11628 15322 11784 15478 sw
tri 11866 15322 12022 15478 ne
rect 12022 15322 12178 15478
tri 12178 15322 12334 15478 sw
tri 12416 15322 12572 15478 ne
rect 12572 15322 12728 15478
tri 12728 15322 12884 15478 sw
tri 12966 15322 13122 15478 ne
rect 13122 15322 13278 15478
tri 13278 15322 13434 15478 sw
tri 13516 15322 13672 15478 ne
rect 13672 15322 13828 15478
tri 13828 15322 13984 15478 sw
tri 14066 15322 14222 15478 ne
rect 14222 15322 14378 15478
tri 14378 15322 14534 15478 sw
tri 14616 15322 14772 15478 ne
rect 14772 15322 14928 15478
tri 14928 15322 15084 15478 sw
tri 15166 15322 15322 15478 ne
rect 15322 15322 15478 15478
tri 15478 15322 15634 15478 sw
tri 15716 15322 15872 15478 ne
rect 15872 15322 16028 15478
tri 16028 15322 16184 15478 sw
tri 16266 15322 16422 15478 ne
rect 16422 15322 16578 15478
tri 16578 15322 16734 15478 sw
tri 16816 15322 16972 15478 ne
rect 16972 15322 17128 15478
tri 17128 15322 17284 15478 sw
tri 17366 15322 17522 15478 ne
rect 17522 15322 17678 15478
tri 17678 15322 17834 15478 sw
tri 17916 15322 18072 15478 ne
rect 18072 15322 18228 15478
tri 18228 15322 18384 15478 sw
tri 18466 15322 18622 15478 ne
rect 18622 15322 18778 15478
tri 18778 15322 18934 15478 sw
tri 19016 15322 19172 15478 ne
rect 19172 15322 19328 15478
tri 19328 15322 19484 15478 sw
tri 19566 15322 19722 15478 ne
rect 19722 15322 20300 15478
rect -2000 15185 234 15322
tri 234 15185 371 15322 sw
tri 472 15185 609 15322 ne
rect 609 15185 784 15322
tri 784 15185 921 15322 sw
tri 1022 15185 1159 15322 ne
rect 1159 15185 1334 15322
tri 1334 15185 1471 15322 sw
tri 1572 15185 1709 15322 ne
rect 1709 15185 1884 15322
tri 1884 15185 2021 15322 sw
tri 2122 15185 2259 15322 ne
rect 2259 15185 2434 15322
tri 2434 15185 2571 15322 sw
tri 2672 15185 2809 15322 ne
rect 2809 15185 2984 15322
tri 2984 15185 3121 15322 sw
tri 3222 15185 3359 15322 ne
rect 3359 15185 3534 15322
tri 3534 15185 3671 15322 sw
tri 3772 15185 3909 15322 ne
rect 3909 15185 4084 15322
tri 4084 15185 4221 15322 sw
tri 4322 15185 4459 15322 ne
rect 4459 15185 4634 15322
tri 4634 15185 4771 15322 sw
tri 4872 15185 5009 15322 ne
rect 5009 15185 5184 15322
tri 5184 15185 5321 15322 sw
tri 5422 15185 5559 15322 ne
rect 5559 15185 5734 15322
tri 5734 15185 5871 15322 sw
tri 5972 15185 6109 15322 ne
rect 6109 15185 6284 15322
tri 6284 15185 6421 15322 sw
tri 6522 15185 6659 15322 ne
rect 6659 15185 6834 15322
tri 6834 15185 6971 15322 sw
tri 7072 15185 7209 15322 ne
rect 7209 15185 7384 15322
tri 7384 15185 7521 15322 sw
tri 7622 15185 7759 15322 ne
rect 7759 15185 7934 15322
tri 7934 15185 8071 15322 sw
tri 8172 15185 8309 15322 ne
rect 8309 15185 8484 15322
tri 8484 15185 8621 15322 sw
tri 8722 15185 8859 15322 ne
rect 8859 15185 9034 15322
tri 9034 15185 9171 15322 sw
tri 9272 15185 9409 15322 ne
rect 9409 15185 9584 15322
tri 9584 15185 9721 15322 sw
tri 9822 15185 9959 15322 ne
rect 9959 15185 10134 15322
tri 10134 15185 10271 15322 sw
tri 10372 15185 10509 15322 ne
rect 10509 15185 10684 15322
tri 10684 15185 10821 15322 sw
tri 10922 15185 11059 15322 ne
rect 11059 15185 11234 15322
tri 11234 15185 11371 15322 sw
tri 11472 15185 11609 15322 ne
rect 11609 15185 11784 15322
tri 11784 15185 11921 15322 sw
tri 12022 15185 12159 15322 ne
rect 12159 15185 12334 15322
tri 12334 15185 12471 15322 sw
tri 12572 15185 12709 15322 ne
rect 12709 15185 12884 15322
tri 12884 15185 13021 15322 sw
tri 13122 15185 13259 15322 ne
rect 13259 15185 13434 15322
tri 13434 15185 13571 15322 sw
tri 13672 15185 13809 15322 ne
rect 13809 15185 13984 15322
tri 13984 15185 14121 15322 sw
tri 14222 15185 14359 15322 ne
rect 14359 15185 14534 15322
tri 14534 15185 14671 15322 sw
tri 14772 15185 14909 15322 ne
rect 14909 15185 15084 15322
tri 15084 15185 15221 15322 sw
tri 15322 15185 15459 15322 ne
rect 15459 15185 15634 15322
tri 15634 15185 15771 15322 sw
tri 15872 15185 16009 15322 ne
rect 16009 15185 16184 15322
tri 16184 15185 16321 15322 sw
tri 16422 15185 16559 15322 ne
rect 16559 15185 16734 15322
tri 16734 15185 16871 15322 sw
tri 16972 15185 17109 15322 ne
rect 17109 15185 17284 15322
tri 17284 15185 17421 15322 sw
tri 17522 15185 17659 15322 ne
rect 17659 15185 17834 15322
tri 17834 15185 17971 15322 sw
tri 18072 15185 18209 15322 ne
rect 18209 15185 18384 15322
tri 18384 15185 18521 15322 sw
tri 18622 15185 18759 15322 ne
rect 18759 15185 18934 15322
tri 18934 15185 19071 15322 sw
tri 19172 15185 19309 15322 ne
rect 19309 15185 19484 15322
tri 19484 15185 19621 15322 sw
rect -2000 15167 215 15185
rect -2000 14378 -1000 15167
tri 77 15065 179 15167 ne
rect 179 15065 215 15167
rect 335 15065 371 15185
tri 179 14928 316 15065 ne
rect 316 15010 371 15065
tri 371 15010 546 15185 sw
tri 609 15065 729 15185 ne
rect 729 15065 765 15185
rect 885 15065 921 15185
rect 316 14928 546 15010
tri 546 14928 628 15010 sw
tri 729 14928 866 15065 ne
rect 866 15010 921 15065
tri 921 15010 1096 15185 sw
tri 1159 15065 1279 15185 ne
rect 1279 15065 1315 15185
rect 1435 15065 1471 15185
rect 866 14928 1096 15010
tri 1096 14928 1178 15010 sw
tri 1279 14928 1416 15065 ne
rect 1416 15010 1471 15065
tri 1471 15010 1646 15185 sw
tri 1709 15065 1829 15185 ne
rect 1829 15065 1865 15185
rect 1985 15065 2021 15185
rect 1416 14928 1646 15010
tri 1646 14928 1728 15010 sw
tri 1829 14928 1966 15065 ne
rect 1966 15010 2021 15065
tri 2021 15010 2196 15185 sw
tri 2259 15065 2379 15185 ne
rect 2379 15065 2415 15185
rect 2535 15065 2571 15185
rect 1966 14928 2196 15010
tri 2196 14928 2278 15010 sw
tri 2379 14928 2516 15065 ne
rect 2516 15010 2571 15065
tri 2571 15010 2746 15185 sw
tri 2809 15065 2929 15185 ne
rect 2929 15065 2965 15185
rect 3085 15065 3121 15185
rect 2516 14928 2746 15010
tri 2746 14928 2828 15010 sw
tri 2929 14928 3066 15065 ne
rect 3066 15010 3121 15065
tri 3121 15010 3296 15185 sw
tri 3359 15065 3479 15185 ne
rect 3479 15065 3515 15185
rect 3635 15065 3671 15185
rect 3066 14928 3296 15010
tri 3296 14928 3378 15010 sw
tri 3479 14928 3616 15065 ne
rect 3616 15010 3671 15065
tri 3671 15010 3846 15185 sw
tri 3909 15065 4029 15185 ne
rect 4029 15065 4065 15185
rect 4185 15065 4221 15185
rect 3616 14928 3846 15010
tri 3846 14928 3928 15010 sw
tri 4029 14928 4166 15065 ne
rect 4166 15010 4221 15065
tri 4221 15010 4396 15185 sw
tri 4459 15065 4579 15185 ne
rect 4579 15065 4615 15185
rect 4735 15065 4771 15185
rect 4166 14928 4396 15010
tri 4396 14928 4478 15010 sw
tri 4579 14928 4716 15065 ne
rect 4716 15010 4771 15065
tri 4771 15010 4946 15185 sw
tri 5009 15065 5129 15185 ne
rect 5129 15065 5165 15185
rect 5285 15065 5321 15185
rect 4716 14928 4946 15010
tri 4946 14928 5028 15010 sw
tri 5129 14928 5266 15065 ne
rect 5266 15010 5321 15065
tri 5321 15010 5496 15185 sw
tri 5559 15065 5679 15185 ne
rect 5679 15065 5715 15185
rect 5835 15065 5871 15185
rect 5266 14928 5496 15010
tri 5496 14928 5578 15010 sw
tri 5679 14928 5816 15065 ne
rect 5816 15010 5871 15065
tri 5871 15010 6046 15185 sw
tri 6109 15065 6229 15185 ne
rect 6229 15065 6265 15185
rect 6385 15065 6421 15185
rect 5816 14928 6046 15010
tri 6046 14928 6128 15010 sw
tri 6229 14928 6366 15065 ne
rect 6366 15010 6421 15065
tri 6421 15010 6596 15185 sw
tri 6659 15065 6779 15185 ne
rect 6779 15065 6815 15185
rect 6935 15065 6971 15185
rect 6366 14928 6596 15010
tri 6596 14928 6678 15010 sw
tri 6779 14928 6916 15065 ne
rect 6916 15010 6971 15065
tri 6971 15010 7146 15185 sw
tri 7209 15065 7329 15185 ne
rect 7329 15065 7365 15185
rect 7485 15065 7521 15185
rect 6916 14928 7146 15010
tri 7146 14928 7228 15010 sw
tri 7329 14928 7466 15065 ne
rect 7466 15010 7521 15065
tri 7521 15010 7696 15185 sw
tri 7759 15065 7879 15185 ne
rect 7879 15065 7915 15185
rect 8035 15065 8071 15185
rect 7466 14928 7696 15010
tri 7696 14928 7778 15010 sw
tri 7879 14928 8016 15065 ne
rect 8016 15010 8071 15065
tri 8071 15010 8246 15185 sw
tri 8309 15065 8429 15185 ne
rect 8429 15065 8465 15185
rect 8585 15065 8621 15185
rect 8016 14928 8246 15010
tri 8246 14928 8328 15010 sw
tri 8429 14928 8566 15065 ne
rect 8566 15010 8621 15065
tri 8621 15010 8796 15185 sw
tri 8859 15065 8979 15185 ne
rect 8979 15065 9015 15185
rect 9135 15065 9171 15185
rect 8566 14928 8796 15010
tri 8796 14928 8878 15010 sw
tri 8979 14928 9116 15065 ne
rect 9116 15010 9171 15065
tri 9171 15010 9346 15185 sw
tri 9409 15065 9529 15185 ne
rect 9529 15065 9565 15185
rect 9685 15065 9721 15185
rect 9116 14928 9346 15010
tri 9346 14928 9428 15010 sw
tri 9529 14928 9666 15065 ne
rect 9666 15010 9721 15065
tri 9721 15010 9896 15185 sw
tri 9959 15065 10079 15185 ne
rect 10079 15065 10115 15185
rect 10235 15065 10271 15185
rect 9666 14928 9896 15010
tri 9896 14928 9978 15010 sw
tri 10079 14928 10216 15065 ne
rect 10216 15010 10271 15065
tri 10271 15010 10446 15185 sw
tri 10509 15065 10629 15185 ne
rect 10629 15065 10665 15185
rect 10785 15065 10821 15185
rect 10216 14928 10446 15010
tri 10446 14928 10528 15010 sw
tri 10629 14928 10766 15065 ne
rect 10766 15010 10821 15065
tri 10821 15010 10996 15185 sw
tri 11059 15065 11179 15185 ne
rect 11179 15065 11215 15185
rect 11335 15065 11371 15185
rect 10766 14928 10996 15010
tri 10996 14928 11078 15010 sw
tri 11179 14928 11316 15065 ne
rect 11316 15010 11371 15065
tri 11371 15010 11546 15185 sw
tri 11609 15065 11729 15185 ne
rect 11729 15065 11765 15185
rect 11885 15065 11921 15185
rect 11316 14928 11546 15010
tri 11546 14928 11628 15010 sw
tri 11729 14928 11866 15065 ne
rect 11866 15010 11921 15065
tri 11921 15010 12096 15185 sw
tri 12159 15065 12279 15185 ne
rect 12279 15065 12315 15185
rect 12435 15065 12471 15185
rect 11866 14928 12096 15010
tri 12096 14928 12178 15010 sw
tri 12279 14928 12416 15065 ne
rect 12416 15010 12471 15065
tri 12471 15010 12646 15185 sw
tri 12709 15065 12829 15185 ne
rect 12829 15065 12865 15185
rect 12985 15065 13021 15185
rect 12416 14928 12646 15010
tri 12646 14928 12728 15010 sw
tri 12829 14928 12966 15065 ne
rect 12966 15010 13021 15065
tri 13021 15010 13196 15185 sw
tri 13259 15065 13379 15185 ne
rect 13379 15065 13415 15185
rect 13535 15065 13571 15185
rect 12966 14928 13196 15010
tri 13196 14928 13278 15010 sw
tri 13379 14928 13516 15065 ne
rect 13516 15010 13571 15065
tri 13571 15010 13746 15185 sw
tri 13809 15065 13929 15185 ne
rect 13929 15065 13965 15185
rect 14085 15065 14121 15185
rect 13516 14928 13746 15010
tri 13746 14928 13828 15010 sw
tri 13929 14928 14066 15065 ne
rect 14066 15010 14121 15065
tri 14121 15010 14296 15185 sw
tri 14359 15065 14479 15185 ne
rect 14479 15065 14515 15185
rect 14635 15065 14671 15185
rect 14066 14928 14296 15010
tri 14296 14928 14378 15010 sw
tri 14479 14928 14616 15065 ne
rect 14616 15010 14671 15065
tri 14671 15010 14846 15185 sw
tri 14909 15065 15029 15185 ne
rect 15029 15065 15065 15185
rect 15185 15065 15221 15185
rect 14616 14928 14846 15010
tri 14846 14928 14928 15010 sw
tri 15029 14928 15166 15065 ne
rect 15166 15010 15221 15065
tri 15221 15010 15396 15185 sw
tri 15459 15065 15579 15185 ne
rect 15579 15065 15615 15185
rect 15735 15065 15771 15185
rect 15166 14928 15396 15010
tri 15396 14928 15478 15010 sw
tri 15579 14928 15716 15065 ne
rect 15716 15010 15771 15065
tri 15771 15010 15946 15185 sw
tri 16009 15065 16129 15185 ne
rect 16129 15065 16165 15185
rect 16285 15065 16321 15185
rect 15716 14928 15946 15010
tri 15946 14928 16028 15010 sw
tri 16129 14928 16266 15065 ne
rect 16266 15010 16321 15065
tri 16321 15010 16496 15185 sw
tri 16559 15065 16679 15185 ne
rect 16679 15065 16715 15185
rect 16835 15065 16871 15185
rect 16266 14928 16496 15010
tri 16496 14928 16578 15010 sw
tri 16679 14928 16816 15065 ne
rect 16816 15010 16871 15065
tri 16871 15010 17046 15185 sw
tri 17109 15065 17229 15185 ne
rect 17229 15065 17265 15185
rect 17385 15065 17421 15185
rect 16816 14928 17046 15010
tri 17046 14928 17128 15010 sw
tri 17229 14928 17366 15065 ne
rect 17366 15010 17421 15065
tri 17421 15010 17596 15185 sw
tri 17659 15065 17779 15185 ne
rect 17779 15065 17815 15185
rect 17935 15065 17971 15185
rect 17366 14928 17596 15010
tri 17596 14928 17678 15010 sw
tri 17779 14928 17916 15065 ne
rect 17916 15010 17971 15065
tri 17971 15010 18146 15185 sw
tri 18209 15065 18329 15185 ne
rect 18329 15065 18365 15185
rect 18485 15065 18521 15185
rect 17916 14928 18146 15010
tri 18146 14928 18228 15010 sw
tri 18329 14928 18466 15065 ne
rect 18466 15010 18521 15065
tri 18521 15010 18696 15185 sw
tri 18759 15065 18879 15185 ne
rect 18879 15065 18915 15185
rect 19035 15065 19071 15185
rect 18466 14928 18696 15010
tri 18696 14928 18778 15010 sw
tri 18879 14928 19016 15065 ne
rect 19016 15010 19071 15065
tri 19071 15010 19246 15185 sw
tri 19309 15065 19429 15185 ne
rect 19429 15065 19465 15185
rect 19585 15083 19621 15185
tri 19621 15083 19723 15185 sw
rect 20800 15083 21800 15872
rect 19585 15065 21800 15083
rect 19016 14928 19246 15010
tri 19246 14928 19328 15010 sw
tri 19429 14928 19566 15065 ne
rect 19566 14928 21800 15065
rect -500 14772 78 14928
tri 78 14772 234 14928 sw
tri 316 14772 472 14928 ne
rect 472 14772 628 14928
tri 628 14772 784 14928 sw
tri 866 14772 1022 14928 ne
rect 1022 14772 1178 14928
tri 1178 14772 1334 14928 sw
tri 1416 14772 1572 14928 ne
rect 1572 14772 1728 14928
tri 1728 14772 1884 14928 sw
tri 1966 14772 2122 14928 ne
rect 2122 14772 2278 14928
tri 2278 14772 2434 14928 sw
tri 2516 14772 2672 14928 ne
rect 2672 14772 2828 14928
tri 2828 14772 2984 14928 sw
tri 3066 14772 3222 14928 ne
rect 3222 14772 3378 14928
tri 3378 14772 3534 14928 sw
tri 3616 14772 3772 14928 ne
rect 3772 14772 3928 14928
tri 3928 14772 4084 14928 sw
tri 4166 14772 4322 14928 ne
rect 4322 14772 4478 14928
tri 4478 14772 4634 14928 sw
tri 4716 14772 4872 14928 ne
rect 4872 14772 5028 14928
tri 5028 14772 5184 14928 sw
tri 5266 14772 5422 14928 ne
rect 5422 14772 5578 14928
tri 5578 14772 5734 14928 sw
tri 5816 14772 5972 14928 ne
rect 5972 14772 6128 14928
tri 6128 14772 6284 14928 sw
tri 6366 14772 6522 14928 ne
rect 6522 14772 6678 14928
tri 6678 14772 6834 14928 sw
tri 6916 14772 7072 14928 ne
rect 7072 14772 7228 14928
tri 7228 14772 7384 14928 sw
tri 7466 14772 7622 14928 ne
rect 7622 14772 7778 14928
tri 7778 14772 7934 14928 sw
tri 8016 14772 8172 14928 ne
rect 8172 14772 8328 14928
tri 8328 14772 8484 14928 sw
tri 8566 14772 8722 14928 ne
rect 8722 14772 8878 14928
tri 8878 14772 9034 14928 sw
tri 9116 14772 9272 14928 ne
rect 9272 14772 9428 14928
tri 9428 14772 9584 14928 sw
tri 9666 14772 9822 14928 ne
rect 9822 14772 9978 14928
tri 9978 14772 10134 14928 sw
tri 10216 14772 10372 14928 ne
rect 10372 14772 10528 14928
tri 10528 14772 10684 14928 sw
tri 10766 14772 10922 14928 ne
rect 10922 14772 11078 14928
tri 11078 14772 11234 14928 sw
tri 11316 14772 11472 14928 ne
rect 11472 14772 11628 14928
tri 11628 14772 11784 14928 sw
tri 11866 14772 12022 14928 ne
rect 12022 14772 12178 14928
tri 12178 14772 12334 14928 sw
tri 12416 14772 12572 14928 ne
rect 12572 14772 12728 14928
tri 12728 14772 12884 14928 sw
tri 12966 14772 13122 14928 ne
rect 13122 14772 13278 14928
tri 13278 14772 13434 14928 sw
tri 13516 14772 13672 14928 ne
rect 13672 14772 13828 14928
tri 13828 14772 13984 14928 sw
tri 14066 14772 14222 14928 ne
rect 14222 14772 14378 14928
tri 14378 14772 14534 14928 sw
tri 14616 14772 14772 14928 ne
rect 14772 14772 14928 14928
tri 14928 14772 15084 14928 sw
tri 15166 14772 15322 14928 ne
rect 15322 14772 15478 14928
tri 15478 14772 15634 14928 sw
tri 15716 14772 15872 14928 ne
rect 15872 14772 16028 14928
tri 16028 14772 16184 14928 sw
tri 16266 14772 16422 14928 ne
rect 16422 14772 16578 14928
tri 16578 14772 16734 14928 sw
tri 16816 14772 16972 14928 ne
rect 16972 14772 17128 14928
tri 17128 14772 17284 14928 sw
tri 17366 14772 17522 14928 ne
rect 17522 14772 17678 14928
tri 17678 14772 17834 14928 sw
tri 17916 14772 18072 14928 ne
rect 18072 14772 18228 14928
tri 18228 14772 18384 14928 sw
tri 18466 14772 18622 14928 ne
rect 18622 14772 18778 14928
tri 18778 14772 18934 14928 sw
tri 19016 14772 19172 14928 ne
rect 19172 14772 19328 14928
tri 19328 14772 19484 14928 sw
tri 19566 14772 19722 14928 ne
rect 19722 14772 21800 14928
rect -500 14635 234 14772
tri 234 14635 371 14772 sw
tri 472 14635 609 14772 ne
rect 609 14635 784 14772
tri 784 14635 921 14772 sw
tri 1022 14635 1159 14772 ne
rect 1159 14635 1334 14772
tri 1334 14635 1471 14772 sw
tri 1572 14635 1709 14772 ne
rect 1709 14635 1884 14772
tri 1884 14635 2021 14772 sw
tri 2122 14635 2259 14772 ne
rect 2259 14635 2434 14772
tri 2434 14635 2571 14772 sw
tri 2672 14635 2809 14772 ne
rect 2809 14635 2984 14772
tri 2984 14635 3121 14772 sw
tri 3222 14635 3359 14772 ne
rect 3359 14635 3534 14772
tri 3534 14635 3671 14772 sw
tri 3772 14635 3909 14772 ne
rect 3909 14635 4084 14772
tri 4084 14635 4221 14772 sw
tri 4322 14635 4459 14772 ne
rect 4459 14635 4634 14772
tri 4634 14635 4771 14772 sw
tri 4872 14635 5009 14772 ne
rect 5009 14635 5184 14772
tri 5184 14635 5321 14772 sw
tri 5422 14635 5559 14772 ne
rect 5559 14635 5734 14772
tri 5734 14635 5871 14772 sw
tri 5972 14635 6109 14772 ne
rect 6109 14635 6284 14772
tri 6284 14635 6421 14772 sw
tri 6522 14635 6659 14772 ne
rect 6659 14635 6834 14772
tri 6834 14635 6971 14772 sw
tri 7072 14635 7209 14772 ne
rect 7209 14635 7384 14772
tri 7384 14635 7521 14772 sw
tri 7622 14635 7759 14772 ne
rect 7759 14635 7934 14772
tri 7934 14635 8071 14772 sw
tri 8172 14635 8309 14772 ne
rect 8309 14635 8484 14772
tri 8484 14635 8621 14772 sw
tri 8722 14635 8859 14772 ne
rect 8859 14635 9034 14772
tri 9034 14635 9171 14772 sw
tri 9272 14635 9409 14772 ne
rect 9409 14635 9584 14772
tri 9584 14635 9721 14772 sw
tri 9822 14635 9959 14772 ne
rect 9959 14635 10134 14772
tri 10134 14635 10271 14772 sw
tri 10372 14635 10509 14772 ne
rect 10509 14635 10684 14772
tri 10684 14635 10821 14772 sw
tri 10922 14635 11059 14772 ne
rect 11059 14635 11234 14772
tri 11234 14635 11371 14772 sw
tri 11472 14635 11609 14772 ne
rect 11609 14635 11784 14772
tri 11784 14635 11921 14772 sw
tri 12022 14635 12159 14772 ne
rect 12159 14635 12334 14772
tri 12334 14635 12471 14772 sw
tri 12572 14635 12709 14772 ne
rect 12709 14635 12884 14772
tri 12884 14635 13021 14772 sw
tri 13122 14635 13259 14772 ne
rect 13259 14635 13434 14772
tri 13434 14635 13571 14772 sw
tri 13672 14635 13809 14772 ne
rect 13809 14635 13984 14772
tri 13984 14635 14121 14772 sw
tri 14222 14635 14359 14772 ne
rect 14359 14635 14534 14772
tri 14534 14635 14671 14772 sw
tri 14772 14635 14909 14772 ne
rect 14909 14635 15084 14772
tri 15084 14635 15221 14772 sw
tri 15322 14635 15459 14772 ne
rect 15459 14635 15634 14772
tri 15634 14635 15771 14772 sw
tri 15872 14635 16009 14772 ne
rect 16009 14635 16184 14772
tri 16184 14635 16321 14772 sw
tri 16422 14635 16559 14772 ne
rect 16559 14635 16734 14772
tri 16734 14635 16871 14772 sw
tri 16972 14635 17109 14772 ne
rect 17109 14635 17284 14772
tri 17284 14635 17421 14772 sw
tri 17522 14635 17659 14772 ne
rect 17659 14635 17834 14772
tri 17834 14635 17971 14772 sw
tri 18072 14635 18209 14772 ne
rect 18209 14635 18384 14772
tri 18384 14635 18521 14772 sw
tri 18622 14635 18759 14772 ne
rect 18759 14635 18934 14772
tri 18934 14635 19071 14772 sw
tri 19172 14635 19309 14772 ne
rect 19309 14635 19484 14772
tri 19484 14635 19621 14772 sw
rect -500 14617 215 14635
tri 77 14515 179 14617 ne
rect 179 14515 215 14617
rect 335 14515 371 14635
tri 179 14378 316 14515 ne
rect 316 14460 371 14515
tri 371 14460 546 14635 sw
tri 609 14515 729 14635 ne
rect 729 14515 765 14635
rect 885 14515 921 14635
rect 316 14378 546 14460
tri 546 14378 628 14460 sw
tri 729 14378 866 14515 ne
rect 866 14460 921 14515
tri 921 14460 1096 14635 sw
tri 1159 14515 1279 14635 ne
rect 1279 14515 1315 14635
rect 1435 14515 1471 14635
rect 866 14378 1096 14460
tri 1096 14378 1178 14460 sw
tri 1279 14378 1416 14515 ne
rect 1416 14460 1471 14515
tri 1471 14460 1646 14635 sw
tri 1709 14515 1829 14635 ne
rect 1829 14515 1865 14635
rect 1985 14515 2021 14635
rect 1416 14378 1646 14460
tri 1646 14378 1728 14460 sw
tri 1829 14378 1966 14515 ne
rect 1966 14460 2021 14515
tri 2021 14460 2196 14635 sw
tri 2259 14515 2379 14635 ne
rect 2379 14515 2415 14635
rect 2535 14515 2571 14635
rect 1966 14378 2196 14460
tri 2196 14378 2278 14460 sw
tri 2379 14378 2516 14515 ne
rect 2516 14460 2571 14515
tri 2571 14460 2746 14635 sw
tri 2809 14515 2929 14635 ne
rect 2929 14515 2965 14635
rect 3085 14515 3121 14635
rect 2516 14378 2746 14460
tri 2746 14378 2828 14460 sw
tri 2929 14378 3066 14515 ne
rect 3066 14460 3121 14515
tri 3121 14460 3296 14635 sw
tri 3359 14515 3479 14635 ne
rect 3479 14515 3515 14635
rect 3635 14515 3671 14635
rect 3066 14378 3296 14460
tri 3296 14378 3378 14460 sw
tri 3479 14378 3616 14515 ne
rect 3616 14460 3671 14515
tri 3671 14460 3846 14635 sw
tri 3909 14515 4029 14635 ne
rect 4029 14515 4065 14635
rect 4185 14515 4221 14635
rect 3616 14378 3846 14460
tri 3846 14378 3928 14460 sw
tri 4029 14378 4166 14515 ne
rect 4166 14460 4221 14515
tri 4221 14460 4396 14635 sw
tri 4459 14515 4579 14635 ne
rect 4579 14515 4615 14635
rect 4735 14515 4771 14635
rect 4166 14378 4396 14460
tri 4396 14378 4478 14460 sw
tri 4579 14378 4716 14515 ne
rect 4716 14460 4771 14515
tri 4771 14460 4946 14635 sw
tri 5009 14515 5129 14635 ne
rect 5129 14515 5165 14635
rect 5285 14515 5321 14635
rect 4716 14378 4946 14460
tri 4946 14378 5028 14460 sw
tri 5129 14378 5266 14515 ne
rect 5266 14460 5321 14515
tri 5321 14460 5496 14635 sw
tri 5559 14515 5679 14635 ne
rect 5679 14515 5715 14635
rect 5835 14515 5871 14635
rect 5266 14378 5496 14460
tri 5496 14378 5578 14460 sw
tri 5679 14378 5816 14515 ne
rect 5816 14460 5871 14515
tri 5871 14460 6046 14635 sw
tri 6109 14515 6229 14635 ne
rect 6229 14515 6265 14635
rect 6385 14515 6421 14635
rect 5816 14378 6046 14460
tri 6046 14378 6128 14460 sw
tri 6229 14378 6366 14515 ne
rect 6366 14460 6421 14515
tri 6421 14460 6596 14635 sw
tri 6659 14515 6779 14635 ne
rect 6779 14515 6815 14635
rect 6935 14515 6971 14635
rect 6366 14378 6596 14460
tri 6596 14378 6678 14460 sw
tri 6779 14378 6916 14515 ne
rect 6916 14460 6971 14515
tri 6971 14460 7146 14635 sw
tri 7209 14515 7329 14635 ne
rect 7329 14515 7365 14635
rect 7485 14515 7521 14635
rect 6916 14378 7146 14460
tri 7146 14378 7228 14460 sw
tri 7329 14378 7466 14515 ne
rect 7466 14460 7521 14515
tri 7521 14460 7696 14635 sw
tri 7759 14515 7879 14635 ne
rect 7879 14515 7915 14635
rect 8035 14515 8071 14635
rect 7466 14378 7696 14460
tri 7696 14378 7778 14460 sw
tri 7879 14378 8016 14515 ne
rect 8016 14460 8071 14515
tri 8071 14460 8246 14635 sw
tri 8309 14515 8429 14635 ne
rect 8429 14515 8465 14635
rect 8585 14515 8621 14635
rect 8016 14378 8246 14460
tri 8246 14378 8328 14460 sw
tri 8429 14378 8566 14515 ne
rect 8566 14460 8621 14515
tri 8621 14460 8796 14635 sw
tri 8859 14515 8979 14635 ne
rect 8979 14515 9015 14635
rect 9135 14515 9171 14635
rect 8566 14378 8796 14460
tri 8796 14378 8878 14460 sw
tri 8979 14378 9116 14515 ne
rect 9116 14460 9171 14515
tri 9171 14460 9346 14635 sw
tri 9409 14515 9529 14635 ne
rect 9529 14515 9565 14635
rect 9685 14515 9721 14635
rect 9116 14378 9346 14460
tri 9346 14378 9428 14460 sw
tri 9529 14378 9666 14515 ne
rect 9666 14460 9721 14515
tri 9721 14460 9896 14635 sw
tri 9959 14515 10079 14635 ne
rect 10079 14515 10115 14635
rect 10235 14515 10271 14635
rect 9666 14378 9896 14460
tri 9896 14378 9978 14460 sw
tri 10079 14378 10216 14515 ne
rect 10216 14460 10271 14515
tri 10271 14460 10446 14635 sw
tri 10509 14515 10629 14635 ne
rect 10629 14515 10665 14635
rect 10785 14515 10821 14635
rect 10216 14378 10446 14460
tri 10446 14378 10528 14460 sw
tri 10629 14378 10766 14515 ne
rect 10766 14460 10821 14515
tri 10821 14460 10996 14635 sw
tri 11059 14515 11179 14635 ne
rect 11179 14515 11215 14635
rect 11335 14515 11371 14635
rect 10766 14378 10996 14460
tri 10996 14378 11078 14460 sw
tri 11179 14378 11316 14515 ne
rect 11316 14460 11371 14515
tri 11371 14460 11546 14635 sw
tri 11609 14515 11729 14635 ne
rect 11729 14515 11765 14635
rect 11885 14515 11921 14635
rect 11316 14378 11546 14460
tri 11546 14378 11628 14460 sw
tri 11729 14378 11866 14515 ne
rect 11866 14460 11921 14515
tri 11921 14460 12096 14635 sw
tri 12159 14515 12279 14635 ne
rect 12279 14515 12315 14635
rect 12435 14515 12471 14635
rect 11866 14378 12096 14460
tri 12096 14378 12178 14460 sw
tri 12279 14378 12416 14515 ne
rect 12416 14460 12471 14515
tri 12471 14460 12646 14635 sw
tri 12709 14515 12829 14635 ne
rect 12829 14515 12865 14635
rect 12985 14515 13021 14635
rect 12416 14378 12646 14460
tri 12646 14378 12728 14460 sw
tri 12829 14378 12966 14515 ne
rect 12966 14460 13021 14515
tri 13021 14460 13196 14635 sw
tri 13259 14515 13379 14635 ne
rect 13379 14515 13415 14635
rect 13535 14515 13571 14635
rect 12966 14378 13196 14460
tri 13196 14378 13278 14460 sw
tri 13379 14378 13516 14515 ne
rect 13516 14460 13571 14515
tri 13571 14460 13746 14635 sw
tri 13809 14515 13929 14635 ne
rect 13929 14515 13965 14635
rect 14085 14515 14121 14635
rect 13516 14378 13746 14460
tri 13746 14378 13828 14460 sw
tri 13929 14378 14066 14515 ne
rect 14066 14460 14121 14515
tri 14121 14460 14296 14635 sw
tri 14359 14515 14479 14635 ne
rect 14479 14515 14515 14635
rect 14635 14515 14671 14635
rect 14066 14378 14296 14460
tri 14296 14378 14378 14460 sw
tri 14479 14378 14616 14515 ne
rect 14616 14460 14671 14515
tri 14671 14460 14846 14635 sw
tri 14909 14515 15029 14635 ne
rect 15029 14515 15065 14635
rect 15185 14515 15221 14635
rect 14616 14378 14846 14460
tri 14846 14378 14928 14460 sw
tri 15029 14378 15166 14515 ne
rect 15166 14460 15221 14515
tri 15221 14460 15396 14635 sw
tri 15459 14515 15579 14635 ne
rect 15579 14515 15615 14635
rect 15735 14515 15771 14635
rect 15166 14378 15396 14460
tri 15396 14378 15478 14460 sw
tri 15579 14378 15716 14515 ne
rect 15716 14460 15771 14515
tri 15771 14460 15946 14635 sw
tri 16009 14515 16129 14635 ne
rect 16129 14515 16165 14635
rect 16285 14515 16321 14635
rect 15716 14378 15946 14460
tri 15946 14378 16028 14460 sw
tri 16129 14378 16266 14515 ne
rect 16266 14460 16321 14515
tri 16321 14460 16496 14635 sw
tri 16559 14515 16679 14635 ne
rect 16679 14515 16715 14635
rect 16835 14515 16871 14635
rect 16266 14378 16496 14460
tri 16496 14378 16578 14460 sw
tri 16679 14378 16816 14515 ne
rect 16816 14460 16871 14515
tri 16871 14460 17046 14635 sw
tri 17109 14515 17229 14635 ne
rect 17229 14515 17265 14635
rect 17385 14515 17421 14635
rect 16816 14378 17046 14460
tri 17046 14378 17128 14460 sw
tri 17229 14378 17366 14515 ne
rect 17366 14460 17421 14515
tri 17421 14460 17596 14635 sw
tri 17659 14515 17779 14635 ne
rect 17779 14515 17815 14635
rect 17935 14515 17971 14635
rect 17366 14378 17596 14460
tri 17596 14378 17678 14460 sw
tri 17779 14378 17916 14515 ne
rect 17916 14460 17971 14515
tri 17971 14460 18146 14635 sw
tri 18209 14515 18329 14635 ne
rect 18329 14515 18365 14635
rect 18485 14515 18521 14635
rect 17916 14378 18146 14460
tri 18146 14378 18228 14460 sw
tri 18329 14378 18466 14515 ne
rect 18466 14460 18521 14515
tri 18521 14460 18696 14635 sw
tri 18759 14515 18879 14635 ne
rect 18879 14515 18915 14635
rect 19035 14515 19071 14635
rect 18466 14378 18696 14460
tri 18696 14378 18778 14460 sw
tri 18879 14378 19016 14515 ne
rect 19016 14460 19071 14515
tri 19071 14460 19246 14635 sw
tri 19309 14515 19429 14635 ne
rect 19429 14515 19465 14635
rect 19585 14533 19621 14635
tri 19621 14533 19723 14635 sw
rect 19585 14515 20300 14533
rect 19016 14378 19246 14460
tri 19246 14378 19328 14460 sw
tri 19429 14378 19566 14515 ne
rect 19566 14378 20300 14515
rect -2000 14222 78 14378
tri 78 14222 234 14378 sw
tri 316 14222 472 14378 ne
rect 472 14222 628 14378
tri 628 14222 784 14378 sw
tri 866 14222 1022 14378 ne
rect 1022 14222 1178 14378
tri 1178 14222 1334 14378 sw
tri 1416 14222 1572 14378 ne
rect 1572 14222 1728 14378
tri 1728 14222 1884 14378 sw
tri 1966 14222 2122 14378 ne
rect 2122 14222 2278 14378
tri 2278 14222 2434 14378 sw
tri 2516 14222 2672 14378 ne
rect 2672 14222 2828 14378
tri 2828 14222 2984 14378 sw
tri 3066 14222 3222 14378 ne
rect 3222 14222 3378 14378
tri 3378 14222 3534 14378 sw
tri 3616 14222 3772 14378 ne
rect 3772 14222 3928 14378
tri 3928 14222 4084 14378 sw
tri 4166 14222 4322 14378 ne
rect 4322 14222 4478 14378
tri 4478 14222 4634 14378 sw
tri 4716 14222 4872 14378 ne
rect 4872 14222 5028 14378
tri 5028 14222 5184 14378 sw
tri 5266 14222 5422 14378 ne
rect 5422 14222 5578 14378
tri 5578 14222 5734 14378 sw
tri 5816 14222 5972 14378 ne
rect 5972 14222 6128 14378
tri 6128 14222 6284 14378 sw
tri 6366 14222 6522 14378 ne
rect 6522 14222 6678 14378
tri 6678 14222 6834 14378 sw
tri 6916 14222 7072 14378 ne
rect 7072 14222 7228 14378
tri 7228 14222 7384 14378 sw
tri 7466 14222 7622 14378 ne
rect 7622 14222 7778 14378
tri 7778 14222 7934 14378 sw
tri 8016 14222 8172 14378 ne
rect 8172 14222 8328 14378
tri 8328 14222 8484 14378 sw
tri 8566 14222 8722 14378 ne
rect 8722 14222 8878 14378
tri 8878 14222 9034 14378 sw
tri 9116 14222 9272 14378 ne
rect 9272 14222 9428 14378
tri 9428 14222 9584 14378 sw
tri 9666 14222 9822 14378 ne
rect 9822 14222 9978 14378
tri 9978 14222 10134 14378 sw
tri 10216 14222 10372 14378 ne
rect 10372 14222 10528 14378
tri 10528 14222 10684 14378 sw
tri 10766 14222 10922 14378 ne
rect 10922 14222 11078 14378
tri 11078 14222 11234 14378 sw
tri 11316 14222 11472 14378 ne
rect 11472 14222 11628 14378
tri 11628 14222 11784 14378 sw
tri 11866 14222 12022 14378 ne
rect 12022 14222 12178 14378
tri 12178 14222 12334 14378 sw
tri 12416 14222 12572 14378 ne
rect 12572 14222 12728 14378
tri 12728 14222 12884 14378 sw
tri 12966 14222 13122 14378 ne
rect 13122 14222 13278 14378
tri 13278 14222 13434 14378 sw
tri 13516 14222 13672 14378 ne
rect 13672 14222 13828 14378
tri 13828 14222 13984 14378 sw
tri 14066 14222 14222 14378 ne
rect 14222 14222 14378 14378
tri 14378 14222 14534 14378 sw
tri 14616 14222 14772 14378 ne
rect 14772 14222 14928 14378
tri 14928 14222 15084 14378 sw
tri 15166 14222 15322 14378 ne
rect 15322 14222 15478 14378
tri 15478 14222 15634 14378 sw
tri 15716 14222 15872 14378 ne
rect 15872 14222 16028 14378
tri 16028 14222 16184 14378 sw
tri 16266 14222 16422 14378 ne
rect 16422 14222 16578 14378
tri 16578 14222 16734 14378 sw
tri 16816 14222 16972 14378 ne
rect 16972 14222 17128 14378
tri 17128 14222 17284 14378 sw
tri 17366 14222 17522 14378 ne
rect 17522 14222 17678 14378
tri 17678 14222 17834 14378 sw
tri 17916 14222 18072 14378 ne
rect 18072 14222 18228 14378
tri 18228 14222 18384 14378 sw
tri 18466 14222 18622 14378 ne
rect 18622 14222 18778 14378
tri 18778 14222 18934 14378 sw
tri 19016 14222 19172 14378 ne
rect 19172 14222 19328 14378
tri 19328 14222 19484 14378 sw
tri 19566 14222 19722 14378 ne
rect 19722 14222 20300 14378
rect -2000 14085 234 14222
tri 234 14085 371 14222 sw
tri 472 14085 609 14222 ne
rect 609 14085 784 14222
tri 784 14085 921 14222 sw
tri 1022 14085 1159 14222 ne
rect 1159 14085 1334 14222
tri 1334 14085 1471 14222 sw
tri 1572 14085 1709 14222 ne
rect 1709 14085 1884 14222
tri 1884 14085 2021 14222 sw
tri 2122 14085 2259 14222 ne
rect 2259 14085 2434 14222
tri 2434 14085 2571 14222 sw
tri 2672 14085 2809 14222 ne
rect 2809 14085 2984 14222
tri 2984 14085 3121 14222 sw
tri 3222 14085 3359 14222 ne
rect 3359 14085 3534 14222
tri 3534 14085 3671 14222 sw
tri 3772 14085 3909 14222 ne
rect 3909 14085 4084 14222
tri 4084 14085 4221 14222 sw
tri 4322 14085 4459 14222 ne
rect 4459 14085 4634 14222
tri 4634 14085 4771 14222 sw
tri 4872 14085 5009 14222 ne
rect 5009 14085 5184 14222
tri 5184 14085 5321 14222 sw
tri 5422 14085 5559 14222 ne
rect 5559 14085 5734 14222
tri 5734 14085 5871 14222 sw
tri 5972 14085 6109 14222 ne
rect 6109 14085 6284 14222
tri 6284 14085 6421 14222 sw
tri 6522 14085 6659 14222 ne
rect 6659 14085 6834 14222
tri 6834 14085 6971 14222 sw
tri 7072 14085 7209 14222 ne
rect 7209 14085 7384 14222
tri 7384 14085 7521 14222 sw
tri 7622 14085 7759 14222 ne
rect 7759 14085 7934 14222
tri 7934 14085 8071 14222 sw
tri 8172 14085 8309 14222 ne
rect 8309 14085 8484 14222
tri 8484 14085 8621 14222 sw
tri 8722 14085 8859 14222 ne
rect 8859 14085 9034 14222
tri 9034 14085 9171 14222 sw
tri 9272 14085 9409 14222 ne
rect 9409 14085 9584 14222
tri 9584 14085 9721 14222 sw
tri 9822 14085 9959 14222 ne
rect 9959 14085 10134 14222
tri 10134 14085 10271 14222 sw
tri 10372 14085 10509 14222 ne
rect 10509 14085 10684 14222
tri 10684 14085 10821 14222 sw
tri 10922 14085 11059 14222 ne
rect 11059 14085 11234 14222
tri 11234 14085 11371 14222 sw
tri 11472 14085 11609 14222 ne
rect 11609 14085 11784 14222
tri 11784 14085 11921 14222 sw
tri 12022 14085 12159 14222 ne
rect 12159 14085 12334 14222
tri 12334 14085 12471 14222 sw
tri 12572 14085 12709 14222 ne
rect 12709 14085 12884 14222
tri 12884 14085 13021 14222 sw
tri 13122 14085 13259 14222 ne
rect 13259 14085 13434 14222
tri 13434 14085 13571 14222 sw
tri 13672 14085 13809 14222 ne
rect 13809 14085 13984 14222
tri 13984 14085 14121 14222 sw
tri 14222 14085 14359 14222 ne
rect 14359 14085 14534 14222
tri 14534 14085 14671 14222 sw
tri 14772 14085 14909 14222 ne
rect 14909 14085 15084 14222
tri 15084 14085 15221 14222 sw
tri 15322 14085 15459 14222 ne
rect 15459 14085 15634 14222
tri 15634 14085 15771 14222 sw
tri 15872 14085 16009 14222 ne
rect 16009 14085 16184 14222
tri 16184 14085 16321 14222 sw
tri 16422 14085 16559 14222 ne
rect 16559 14085 16734 14222
tri 16734 14085 16871 14222 sw
tri 16972 14085 17109 14222 ne
rect 17109 14085 17284 14222
tri 17284 14085 17421 14222 sw
tri 17522 14085 17659 14222 ne
rect 17659 14085 17834 14222
tri 17834 14085 17971 14222 sw
tri 18072 14085 18209 14222 ne
rect 18209 14085 18384 14222
tri 18384 14085 18521 14222 sw
tri 18622 14085 18759 14222 ne
rect 18759 14085 18934 14222
tri 18934 14085 19071 14222 sw
tri 19172 14085 19309 14222 ne
rect 19309 14085 19484 14222
tri 19484 14085 19621 14222 sw
rect -2000 14067 215 14085
rect -2000 13278 -1000 14067
tri 77 13965 179 14067 ne
rect 179 13965 215 14067
rect 335 13965 371 14085
tri 179 13828 316 13965 ne
rect 316 13910 371 13965
tri 371 13910 546 14085 sw
tri 609 13965 729 14085 ne
rect 729 13965 765 14085
rect 885 13965 921 14085
rect 316 13828 546 13910
tri 546 13828 628 13910 sw
tri 729 13828 866 13965 ne
rect 866 13910 921 13965
tri 921 13910 1096 14085 sw
tri 1159 13965 1279 14085 ne
rect 1279 13965 1315 14085
rect 1435 13965 1471 14085
rect 866 13828 1096 13910
tri 1096 13828 1178 13910 sw
tri 1279 13828 1416 13965 ne
rect 1416 13910 1471 13965
tri 1471 13910 1646 14085 sw
tri 1709 13965 1829 14085 ne
rect 1829 13965 1865 14085
rect 1985 13965 2021 14085
rect 1416 13828 1646 13910
tri 1646 13828 1728 13910 sw
tri 1829 13828 1966 13965 ne
rect 1966 13910 2021 13965
tri 2021 13910 2196 14085 sw
tri 2259 13965 2379 14085 ne
rect 2379 13965 2415 14085
rect 2535 13965 2571 14085
rect 1966 13828 2196 13910
tri 2196 13828 2278 13910 sw
tri 2379 13828 2516 13965 ne
rect 2516 13910 2571 13965
tri 2571 13910 2746 14085 sw
tri 2809 13965 2929 14085 ne
rect 2929 13965 2965 14085
rect 3085 13965 3121 14085
rect 2516 13828 2746 13910
tri 2746 13828 2828 13910 sw
tri 2929 13828 3066 13965 ne
rect 3066 13910 3121 13965
tri 3121 13910 3296 14085 sw
tri 3359 13965 3479 14085 ne
rect 3479 13965 3515 14085
rect 3635 13965 3671 14085
rect 3066 13828 3296 13910
tri 3296 13828 3378 13910 sw
tri 3479 13828 3616 13965 ne
rect 3616 13910 3671 13965
tri 3671 13910 3846 14085 sw
tri 3909 13965 4029 14085 ne
rect 4029 13965 4065 14085
rect 4185 13965 4221 14085
rect 3616 13828 3846 13910
tri 3846 13828 3928 13910 sw
tri 4029 13828 4166 13965 ne
rect 4166 13910 4221 13965
tri 4221 13910 4396 14085 sw
tri 4459 13965 4579 14085 ne
rect 4579 13965 4615 14085
rect 4735 13965 4771 14085
rect 4166 13828 4396 13910
tri 4396 13828 4478 13910 sw
tri 4579 13828 4716 13965 ne
rect 4716 13910 4771 13965
tri 4771 13910 4946 14085 sw
tri 5009 13965 5129 14085 ne
rect 5129 13965 5165 14085
rect 5285 13965 5321 14085
rect 4716 13828 4946 13910
tri 4946 13828 5028 13910 sw
tri 5129 13828 5266 13965 ne
rect 5266 13910 5321 13965
tri 5321 13910 5496 14085 sw
tri 5559 13965 5679 14085 ne
rect 5679 13965 5715 14085
rect 5835 13965 5871 14085
rect 5266 13828 5496 13910
tri 5496 13828 5578 13910 sw
tri 5679 13828 5816 13965 ne
rect 5816 13910 5871 13965
tri 5871 13910 6046 14085 sw
tri 6109 13965 6229 14085 ne
rect 6229 13965 6265 14085
rect 6385 13965 6421 14085
rect 5816 13828 6046 13910
tri 6046 13828 6128 13910 sw
tri 6229 13828 6366 13965 ne
rect 6366 13910 6421 13965
tri 6421 13910 6596 14085 sw
tri 6659 13965 6779 14085 ne
rect 6779 13965 6815 14085
rect 6935 13965 6971 14085
rect 6366 13828 6596 13910
tri 6596 13828 6678 13910 sw
tri 6779 13828 6916 13965 ne
rect 6916 13910 6971 13965
tri 6971 13910 7146 14085 sw
tri 7209 13965 7329 14085 ne
rect 7329 13965 7365 14085
rect 7485 13965 7521 14085
rect 6916 13828 7146 13910
tri 7146 13828 7228 13910 sw
tri 7329 13828 7466 13965 ne
rect 7466 13910 7521 13965
tri 7521 13910 7696 14085 sw
tri 7759 13965 7879 14085 ne
rect 7879 13965 7915 14085
rect 8035 13965 8071 14085
rect 7466 13828 7696 13910
tri 7696 13828 7778 13910 sw
tri 7879 13828 8016 13965 ne
rect 8016 13910 8071 13965
tri 8071 13910 8246 14085 sw
tri 8309 13965 8429 14085 ne
rect 8429 13965 8465 14085
rect 8585 13965 8621 14085
rect 8016 13828 8246 13910
tri 8246 13828 8328 13910 sw
tri 8429 13828 8566 13965 ne
rect 8566 13910 8621 13965
tri 8621 13910 8796 14085 sw
tri 8859 13965 8979 14085 ne
rect 8979 13965 9015 14085
rect 9135 13965 9171 14085
rect 8566 13828 8796 13910
tri 8796 13828 8878 13910 sw
tri 8979 13828 9116 13965 ne
rect 9116 13910 9171 13965
tri 9171 13910 9346 14085 sw
tri 9409 13965 9529 14085 ne
rect 9529 13965 9565 14085
rect 9685 13965 9721 14085
rect 9116 13828 9346 13910
tri 9346 13828 9428 13910 sw
tri 9529 13828 9666 13965 ne
rect 9666 13910 9721 13965
tri 9721 13910 9896 14085 sw
tri 9959 13965 10079 14085 ne
rect 10079 13965 10115 14085
rect 10235 13965 10271 14085
rect 9666 13828 9896 13910
tri 9896 13828 9978 13910 sw
tri 10079 13828 10216 13965 ne
rect 10216 13910 10271 13965
tri 10271 13910 10446 14085 sw
tri 10509 13965 10629 14085 ne
rect 10629 13965 10665 14085
rect 10785 13965 10821 14085
rect 10216 13828 10446 13910
tri 10446 13828 10528 13910 sw
tri 10629 13828 10766 13965 ne
rect 10766 13910 10821 13965
tri 10821 13910 10996 14085 sw
tri 11059 13965 11179 14085 ne
rect 11179 13965 11215 14085
rect 11335 13965 11371 14085
rect 10766 13828 10996 13910
tri 10996 13828 11078 13910 sw
tri 11179 13828 11316 13965 ne
rect 11316 13910 11371 13965
tri 11371 13910 11546 14085 sw
tri 11609 13965 11729 14085 ne
rect 11729 13965 11765 14085
rect 11885 13965 11921 14085
rect 11316 13828 11546 13910
tri 11546 13828 11628 13910 sw
tri 11729 13828 11866 13965 ne
rect 11866 13910 11921 13965
tri 11921 13910 12096 14085 sw
tri 12159 13965 12279 14085 ne
rect 12279 13965 12315 14085
rect 12435 13965 12471 14085
rect 11866 13828 12096 13910
tri 12096 13828 12178 13910 sw
tri 12279 13828 12416 13965 ne
rect 12416 13910 12471 13965
tri 12471 13910 12646 14085 sw
tri 12709 13965 12829 14085 ne
rect 12829 13965 12865 14085
rect 12985 13965 13021 14085
rect 12416 13828 12646 13910
tri 12646 13828 12728 13910 sw
tri 12829 13828 12966 13965 ne
rect 12966 13910 13021 13965
tri 13021 13910 13196 14085 sw
tri 13259 13965 13379 14085 ne
rect 13379 13965 13415 14085
rect 13535 13965 13571 14085
rect 12966 13828 13196 13910
tri 13196 13828 13278 13910 sw
tri 13379 13828 13516 13965 ne
rect 13516 13910 13571 13965
tri 13571 13910 13746 14085 sw
tri 13809 13965 13929 14085 ne
rect 13929 13965 13965 14085
rect 14085 13965 14121 14085
rect 13516 13828 13746 13910
tri 13746 13828 13828 13910 sw
tri 13929 13828 14066 13965 ne
rect 14066 13910 14121 13965
tri 14121 13910 14296 14085 sw
tri 14359 13965 14479 14085 ne
rect 14479 13965 14515 14085
rect 14635 13965 14671 14085
rect 14066 13828 14296 13910
tri 14296 13828 14378 13910 sw
tri 14479 13828 14616 13965 ne
rect 14616 13910 14671 13965
tri 14671 13910 14846 14085 sw
tri 14909 13965 15029 14085 ne
rect 15029 13965 15065 14085
rect 15185 13965 15221 14085
rect 14616 13828 14846 13910
tri 14846 13828 14928 13910 sw
tri 15029 13828 15166 13965 ne
rect 15166 13910 15221 13965
tri 15221 13910 15396 14085 sw
tri 15459 13965 15579 14085 ne
rect 15579 13965 15615 14085
rect 15735 13965 15771 14085
rect 15166 13828 15396 13910
tri 15396 13828 15478 13910 sw
tri 15579 13828 15716 13965 ne
rect 15716 13910 15771 13965
tri 15771 13910 15946 14085 sw
tri 16009 13965 16129 14085 ne
rect 16129 13965 16165 14085
rect 16285 13965 16321 14085
rect 15716 13828 15946 13910
tri 15946 13828 16028 13910 sw
tri 16129 13828 16266 13965 ne
rect 16266 13910 16321 13965
tri 16321 13910 16496 14085 sw
tri 16559 13965 16679 14085 ne
rect 16679 13965 16715 14085
rect 16835 13965 16871 14085
rect 16266 13828 16496 13910
tri 16496 13828 16578 13910 sw
tri 16679 13828 16816 13965 ne
rect 16816 13910 16871 13965
tri 16871 13910 17046 14085 sw
tri 17109 13965 17229 14085 ne
rect 17229 13965 17265 14085
rect 17385 13965 17421 14085
rect 16816 13828 17046 13910
tri 17046 13828 17128 13910 sw
tri 17229 13828 17366 13965 ne
rect 17366 13910 17421 13965
tri 17421 13910 17596 14085 sw
tri 17659 13965 17779 14085 ne
rect 17779 13965 17815 14085
rect 17935 13965 17971 14085
rect 17366 13828 17596 13910
tri 17596 13828 17678 13910 sw
tri 17779 13828 17916 13965 ne
rect 17916 13910 17971 13965
tri 17971 13910 18146 14085 sw
tri 18209 13965 18329 14085 ne
rect 18329 13965 18365 14085
rect 18485 13965 18521 14085
rect 17916 13828 18146 13910
tri 18146 13828 18228 13910 sw
tri 18329 13828 18466 13965 ne
rect 18466 13910 18521 13965
tri 18521 13910 18696 14085 sw
tri 18759 13965 18879 14085 ne
rect 18879 13965 18915 14085
rect 19035 13965 19071 14085
rect 18466 13828 18696 13910
tri 18696 13828 18778 13910 sw
tri 18879 13828 19016 13965 ne
rect 19016 13910 19071 13965
tri 19071 13910 19246 14085 sw
tri 19309 13965 19429 14085 ne
rect 19429 13965 19465 14085
rect 19585 13983 19621 14085
tri 19621 13983 19723 14085 sw
rect 20800 13983 21800 14772
rect 19585 13965 21800 13983
rect 19016 13828 19246 13910
tri 19246 13828 19328 13910 sw
tri 19429 13828 19566 13965 ne
rect 19566 13828 21800 13965
rect -500 13672 78 13828
tri 78 13672 234 13828 sw
tri 316 13672 472 13828 ne
rect 472 13672 628 13828
tri 628 13672 784 13828 sw
tri 866 13672 1022 13828 ne
rect 1022 13672 1178 13828
tri 1178 13672 1334 13828 sw
tri 1416 13672 1572 13828 ne
rect 1572 13672 1728 13828
tri 1728 13672 1884 13828 sw
tri 1966 13672 2122 13828 ne
rect 2122 13672 2278 13828
tri 2278 13672 2434 13828 sw
tri 2516 13672 2672 13828 ne
rect 2672 13672 2828 13828
tri 2828 13672 2984 13828 sw
tri 3066 13672 3222 13828 ne
rect 3222 13672 3378 13828
tri 3378 13672 3534 13828 sw
tri 3616 13672 3772 13828 ne
rect 3772 13672 3928 13828
tri 3928 13672 4084 13828 sw
tri 4166 13672 4322 13828 ne
rect 4322 13672 4478 13828
tri 4478 13672 4634 13828 sw
tri 4716 13672 4872 13828 ne
rect 4872 13672 5028 13828
tri 5028 13672 5184 13828 sw
tri 5266 13672 5422 13828 ne
rect 5422 13672 5578 13828
tri 5578 13672 5734 13828 sw
tri 5816 13672 5972 13828 ne
rect 5972 13672 6128 13828
tri 6128 13672 6284 13828 sw
tri 6366 13672 6522 13828 ne
rect 6522 13672 6678 13828
tri 6678 13672 6834 13828 sw
tri 6916 13672 7072 13828 ne
rect 7072 13672 7228 13828
tri 7228 13672 7384 13828 sw
tri 7466 13672 7622 13828 ne
rect 7622 13672 7778 13828
tri 7778 13672 7934 13828 sw
tri 8016 13672 8172 13828 ne
rect 8172 13672 8328 13828
tri 8328 13672 8484 13828 sw
tri 8566 13672 8722 13828 ne
rect 8722 13672 8878 13828
tri 8878 13672 9034 13828 sw
tri 9116 13672 9272 13828 ne
rect 9272 13672 9428 13828
tri 9428 13672 9584 13828 sw
tri 9666 13672 9822 13828 ne
rect 9822 13672 9978 13828
tri 9978 13672 10134 13828 sw
tri 10216 13672 10372 13828 ne
rect 10372 13672 10528 13828
tri 10528 13672 10684 13828 sw
tri 10766 13672 10922 13828 ne
rect 10922 13672 11078 13828
tri 11078 13672 11234 13828 sw
tri 11316 13672 11472 13828 ne
rect 11472 13672 11628 13828
tri 11628 13672 11784 13828 sw
tri 11866 13672 12022 13828 ne
rect 12022 13672 12178 13828
tri 12178 13672 12334 13828 sw
tri 12416 13672 12572 13828 ne
rect 12572 13672 12728 13828
tri 12728 13672 12884 13828 sw
tri 12966 13672 13122 13828 ne
rect 13122 13672 13278 13828
tri 13278 13672 13434 13828 sw
tri 13516 13672 13672 13828 ne
rect 13672 13672 13828 13828
tri 13828 13672 13984 13828 sw
tri 14066 13672 14222 13828 ne
rect 14222 13672 14378 13828
tri 14378 13672 14534 13828 sw
tri 14616 13672 14772 13828 ne
rect 14772 13672 14928 13828
tri 14928 13672 15084 13828 sw
tri 15166 13672 15322 13828 ne
rect 15322 13672 15478 13828
tri 15478 13672 15634 13828 sw
tri 15716 13672 15872 13828 ne
rect 15872 13672 16028 13828
tri 16028 13672 16184 13828 sw
tri 16266 13672 16422 13828 ne
rect 16422 13672 16578 13828
tri 16578 13672 16734 13828 sw
tri 16816 13672 16972 13828 ne
rect 16972 13672 17128 13828
tri 17128 13672 17284 13828 sw
tri 17366 13672 17522 13828 ne
rect 17522 13672 17678 13828
tri 17678 13672 17834 13828 sw
tri 17916 13672 18072 13828 ne
rect 18072 13672 18228 13828
tri 18228 13672 18384 13828 sw
tri 18466 13672 18622 13828 ne
rect 18622 13672 18778 13828
tri 18778 13672 18934 13828 sw
tri 19016 13672 19172 13828 ne
rect 19172 13672 19328 13828
tri 19328 13672 19484 13828 sw
tri 19566 13672 19722 13828 ne
rect 19722 13672 21800 13828
rect -500 13535 234 13672
tri 234 13535 371 13672 sw
tri 472 13535 609 13672 ne
rect 609 13535 784 13672
tri 784 13535 921 13672 sw
tri 1022 13535 1159 13672 ne
rect 1159 13535 1334 13672
tri 1334 13535 1471 13672 sw
tri 1572 13535 1709 13672 ne
rect 1709 13535 1884 13672
tri 1884 13535 2021 13672 sw
tri 2122 13535 2259 13672 ne
rect 2259 13535 2434 13672
tri 2434 13535 2571 13672 sw
tri 2672 13535 2809 13672 ne
rect 2809 13535 2984 13672
tri 2984 13535 3121 13672 sw
tri 3222 13535 3359 13672 ne
rect 3359 13535 3534 13672
tri 3534 13535 3671 13672 sw
tri 3772 13535 3909 13672 ne
rect 3909 13535 4084 13672
tri 4084 13535 4221 13672 sw
tri 4322 13535 4459 13672 ne
rect 4459 13535 4634 13672
tri 4634 13535 4771 13672 sw
tri 4872 13535 5009 13672 ne
rect 5009 13535 5184 13672
tri 5184 13535 5321 13672 sw
tri 5422 13535 5559 13672 ne
rect 5559 13535 5734 13672
tri 5734 13535 5871 13672 sw
tri 5972 13535 6109 13672 ne
rect 6109 13535 6284 13672
tri 6284 13535 6421 13672 sw
tri 6522 13535 6659 13672 ne
rect 6659 13535 6834 13672
tri 6834 13535 6971 13672 sw
tri 7072 13535 7209 13672 ne
rect 7209 13535 7384 13672
tri 7384 13535 7521 13672 sw
tri 7622 13535 7759 13672 ne
rect 7759 13535 7934 13672
tri 7934 13535 8071 13672 sw
tri 8172 13535 8309 13672 ne
rect 8309 13535 8484 13672
tri 8484 13535 8621 13672 sw
tri 8722 13535 8859 13672 ne
rect 8859 13535 9034 13672
tri 9034 13535 9171 13672 sw
tri 9272 13535 9409 13672 ne
rect 9409 13535 9584 13672
tri 9584 13535 9721 13672 sw
tri 9822 13535 9959 13672 ne
rect 9959 13535 10134 13672
tri 10134 13535 10271 13672 sw
tri 10372 13535 10509 13672 ne
rect 10509 13535 10684 13672
tri 10684 13535 10821 13672 sw
tri 10922 13535 11059 13672 ne
rect 11059 13535 11234 13672
tri 11234 13535 11371 13672 sw
tri 11472 13535 11609 13672 ne
rect 11609 13535 11784 13672
tri 11784 13535 11921 13672 sw
tri 12022 13535 12159 13672 ne
rect 12159 13535 12334 13672
tri 12334 13535 12471 13672 sw
tri 12572 13535 12709 13672 ne
rect 12709 13535 12884 13672
tri 12884 13535 13021 13672 sw
tri 13122 13535 13259 13672 ne
rect 13259 13535 13434 13672
tri 13434 13535 13571 13672 sw
tri 13672 13535 13809 13672 ne
rect 13809 13535 13984 13672
tri 13984 13535 14121 13672 sw
tri 14222 13535 14359 13672 ne
rect 14359 13535 14534 13672
tri 14534 13535 14671 13672 sw
tri 14772 13535 14909 13672 ne
rect 14909 13535 15084 13672
tri 15084 13535 15221 13672 sw
tri 15322 13535 15459 13672 ne
rect 15459 13535 15634 13672
tri 15634 13535 15771 13672 sw
tri 15872 13535 16009 13672 ne
rect 16009 13535 16184 13672
tri 16184 13535 16321 13672 sw
tri 16422 13535 16559 13672 ne
rect 16559 13535 16734 13672
tri 16734 13535 16871 13672 sw
tri 16972 13535 17109 13672 ne
rect 17109 13535 17284 13672
tri 17284 13535 17421 13672 sw
tri 17522 13535 17659 13672 ne
rect 17659 13535 17834 13672
tri 17834 13535 17971 13672 sw
tri 18072 13535 18209 13672 ne
rect 18209 13535 18384 13672
tri 18384 13535 18521 13672 sw
tri 18622 13535 18759 13672 ne
rect 18759 13535 18934 13672
tri 18934 13535 19071 13672 sw
tri 19172 13535 19309 13672 ne
rect 19309 13535 19484 13672
tri 19484 13535 19621 13672 sw
rect -500 13517 215 13535
tri 77 13415 179 13517 ne
rect 179 13415 215 13517
rect 335 13415 371 13535
tri 179 13278 316 13415 ne
rect 316 13360 371 13415
tri 371 13360 546 13535 sw
tri 609 13415 729 13535 ne
rect 729 13415 765 13535
rect 885 13415 921 13535
rect 316 13278 546 13360
tri 546 13278 628 13360 sw
tri 729 13278 866 13415 ne
rect 866 13360 921 13415
tri 921 13360 1096 13535 sw
tri 1159 13415 1279 13535 ne
rect 1279 13415 1315 13535
rect 1435 13415 1471 13535
rect 866 13278 1096 13360
tri 1096 13278 1178 13360 sw
tri 1279 13278 1416 13415 ne
rect 1416 13360 1471 13415
tri 1471 13360 1646 13535 sw
tri 1709 13415 1829 13535 ne
rect 1829 13415 1865 13535
rect 1985 13415 2021 13535
rect 1416 13278 1646 13360
tri 1646 13278 1728 13360 sw
tri 1829 13278 1966 13415 ne
rect 1966 13360 2021 13415
tri 2021 13360 2196 13535 sw
tri 2259 13415 2379 13535 ne
rect 2379 13415 2415 13535
rect 2535 13415 2571 13535
rect 1966 13278 2196 13360
tri 2196 13278 2278 13360 sw
tri 2379 13278 2516 13415 ne
rect 2516 13360 2571 13415
tri 2571 13360 2746 13535 sw
tri 2809 13415 2929 13535 ne
rect 2929 13415 2965 13535
rect 3085 13415 3121 13535
rect 2516 13278 2746 13360
tri 2746 13278 2828 13360 sw
tri 2929 13278 3066 13415 ne
rect 3066 13360 3121 13415
tri 3121 13360 3296 13535 sw
tri 3359 13415 3479 13535 ne
rect 3479 13415 3515 13535
rect 3635 13415 3671 13535
rect 3066 13278 3296 13360
tri 3296 13278 3378 13360 sw
tri 3479 13278 3616 13415 ne
rect 3616 13360 3671 13415
tri 3671 13360 3846 13535 sw
tri 3909 13415 4029 13535 ne
rect 4029 13415 4065 13535
rect 4185 13415 4221 13535
rect 3616 13278 3846 13360
tri 3846 13278 3928 13360 sw
tri 4029 13278 4166 13415 ne
rect 4166 13360 4221 13415
tri 4221 13360 4396 13535 sw
tri 4459 13415 4579 13535 ne
rect 4579 13415 4615 13535
rect 4735 13415 4771 13535
rect 4166 13278 4396 13360
tri 4396 13278 4478 13360 sw
tri 4579 13278 4716 13415 ne
rect 4716 13360 4771 13415
tri 4771 13360 4946 13535 sw
tri 5009 13415 5129 13535 ne
rect 5129 13415 5165 13535
rect 5285 13415 5321 13535
rect 4716 13278 4946 13360
tri 4946 13278 5028 13360 sw
tri 5129 13278 5266 13415 ne
rect 5266 13360 5321 13415
tri 5321 13360 5496 13535 sw
tri 5559 13415 5679 13535 ne
rect 5679 13415 5715 13535
rect 5835 13415 5871 13535
rect 5266 13278 5496 13360
tri 5496 13278 5578 13360 sw
tri 5679 13278 5816 13415 ne
rect 5816 13360 5871 13415
tri 5871 13360 6046 13535 sw
tri 6109 13415 6229 13535 ne
rect 6229 13415 6265 13535
rect 6385 13415 6421 13535
rect 5816 13278 6046 13360
tri 6046 13278 6128 13360 sw
tri 6229 13278 6366 13415 ne
rect 6366 13360 6421 13415
tri 6421 13360 6596 13535 sw
tri 6659 13415 6779 13535 ne
rect 6779 13415 6815 13535
rect 6935 13415 6971 13535
rect 6366 13278 6596 13360
tri 6596 13278 6678 13360 sw
tri 6779 13278 6916 13415 ne
rect 6916 13360 6971 13415
tri 6971 13360 7146 13535 sw
tri 7209 13415 7329 13535 ne
rect 7329 13415 7365 13535
rect 7485 13415 7521 13535
rect 6916 13278 7146 13360
tri 7146 13278 7228 13360 sw
tri 7329 13278 7466 13415 ne
rect 7466 13360 7521 13415
tri 7521 13360 7696 13535 sw
tri 7759 13415 7879 13535 ne
rect 7879 13415 7915 13535
rect 8035 13415 8071 13535
rect 7466 13278 7696 13360
tri 7696 13278 7778 13360 sw
tri 7879 13278 8016 13415 ne
rect 8016 13360 8071 13415
tri 8071 13360 8246 13535 sw
tri 8309 13415 8429 13535 ne
rect 8429 13415 8465 13535
rect 8585 13415 8621 13535
rect 8016 13278 8246 13360
tri 8246 13278 8328 13360 sw
tri 8429 13278 8566 13415 ne
rect 8566 13360 8621 13415
tri 8621 13360 8796 13535 sw
tri 8859 13415 8979 13535 ne
rect 8979 13415 9015 13535
rect 9135 13415 9171 13535
rect 8566 13278 8796 13360
tri 8796 13278 8878 13360 sw
tri 8979 13278 9116 13415 ne
rect 9116 13360 9171 13415
tri 9171 13360 9346 13535 sw
tri 9409 13415 9529 13535 ne
rect 9529 13415 9565 13535
rect 9685 13415 9721 13535
rect 9116 13278 9346 13360
tri 9346 13278 9428 13360 sw
tri 9529 13278 9666 13415 ne
rect 9666 13360 9721 13415
tri 9721 13360 9896 13535 sw
tri 9959 13415 10079 13535 ne
rect 10079 13415 10115 13535
rect 10235 13415 10271 13535
rect 9666 13278 9896 13360
tri 9896 13278 9978 13360 sw
tri 10079 13278 10216 13415 ne
rect 10216 13360 10271 13415
tri 10271 13360 10446 13535 sw
tri 10509 13415 10629 13535 ne
rect 10629 13415 10665 13535
rect 10785 13415 10821 13535
rect 10216 13278 10446 13360
tri 10446 13278 10528 13360 sw
tri 10629 13278 10766 13415 ne
rect 10766 13360 10821 13415
tri 10821 13360 10996 13535 sw
tri 11059 13415 11179 13535 ne
rect 11179 13415 11215 13535
rect 11335 13415 11371 13535
rect 10766 13278 10996 13360
tri 10996 13278 11078 13360 sw
tri 11179 13278 11316 13415 ne
rect 11316 13360 11371 13415
tri 11371 13360 11546 13535 sw
tri 11609 13415 11729 13535 ne
rect 11729 13415 11765 13535
rect 11885 13415 11921 13535
rect 11316 13278 11546 13360
tri 11546 13278 11628 13360 sw
tri 11729 13278 11866 13415 ne
rect 11866 13360 11921 13415
tri 11921 13360 12096 13535 sw
tri 12159 13415 12279 13535 ne
rect 12279 13415 12315 13535
rect 12435 13415 12471 13535
rect 11866 13278 12096 13360
tri 12096 13278 12178 13360 sw
tri 12279 13278 12416 13415 ne
rect 12416 13360 12471 13415
tri 12471 13360 12646 13535 sw
tri 12709 13415 12829 13535 ne
rect 12829 13415 12865 13535
rect 12985 13415 13021 13535
rect 12416 13278 12646 13360
tri 12646 13278 12728 13360 sw
tri 12829 13278 12966 13415 ne
rect 12966 13360 13021 13415
tri 13021 13360 13196 13535 sw
tri 13259 13415 13379 13535 ne
rect 13379 13415 13415 13535
rect 13535 13415 13571 13535
rect 12966 13278 13196 13360
tri 13196 13278 13278 13360 sw
tri 13379 13278 13516 13415 ne
rect 13516 13360 13571 13415
tri 13571 13360 13746 13535 sw
tri 13809 13415 13929 13535 ne
rect 13929 13415 13965 13535
rect 14085 13415 14121 13535
rect 13516 13278 13746 13360
tri 13746 13278 13828 13360 sw
tri 13929 13278 14066 13415 ne
rect 14066 13360 14121 13415
tri 14121 13360 14296 13535 sw
tri 14359 13415 14479 13535 ne
rect 14479 13415 14515 13535
rect 14635 13415 14671 13535
rect 14066 13278 14296 13360
tri 14296 13278 14378 13360 sw
tri 14479 13278 14616 13415 ne
rect 14616 13360 14671 13415
tri 14671 13360 14846 13535 sw
tri 14909 13415 15029 13535 ne
rect 15029 13415 15065 13535
rect 15185 13415 15221 13535
rect 14616 13278 14846 13360
tri 14846 13278 14928 13360 sw
tri 15029 13278 15166 13415 ne
rect 15166 13360 15221 13415
tri 15221 13360 15396 13535 sw
tri 15459 13415 15579 13535 ne
rect 15579 13415 15615 13535
rect 15735 13415 15771 13535
rect 15166 13278 15396 13360
tri 15396 13278 15478 13360 sw
tri 15579 13278 15716 13415 ne
rect 15716 13360 15771 13415
tri 15771 13360 15946 13535 sw
tri 16009 13415 16129 13535 ne
rect 16129 13415 16165 13535
rect 16285 13415 16321 13535
rect 15716 13278 15946 13360
tri 15946 13278 16028 13360 sw
tri 16129 13278 16266 13415 ne
rect 16266 13360 16321 13415
tri 16321 13360 16496 13535 sw
tri 16559 13415 16679 13535 ne
rect 16679 13415 16715 13535
rect 16835 13415 16871 13535
rect 16266 13278 16496 13360
tri 16496 13278 16578 13360 sw
tri 16679 13278 16816 13415 ne
rect 16816 13360 16871 13415
tri 16871 13360 17046 13535 sw
tri 17109 13415 17229 13535 ne
rect 17229 13415 17265 13535
rect 17385 13415 17421 13535
rect 16816 13278 17046 13360
tri 17046 13278 17128 13360 sw
tri 17229 13278 17366 13415 ne
rect 17366 13360 17421 13415
tri 17421 13360 17596 13535 sw
tri 17659 13415 17779 13535 ne
rect 17779 13415 17815 13535
rect 17935 13415 17971 13535
rect 17366 13278 17596 13360
tri 17596 13278 17678 13360 sw
tri 17779 13278 17916 13415 ne
rect 17916 13360 17971 13415
tri 17971 13360 18146 13535 sw
tri 18209 13415 18329 13535 ne
rect 18329 13415 18365 13535
rect 18485 13415 18521 13535
rect 17916 13278 18146 13360
tri 18146 13278 18228 13360 sw
tri 18329 13278 18466 13415 ne
rect 18466 13360 18521 13415
tri 18521 13360 18696 13535 sw
tri 18759 13415 18879 13535 ne
rect 18879 13415 18915 13535
rect 19035 13415 19071 13535
rect 18466 13278 18696 13360
tri 18696 13278 18778 13360 sw
tri 18879 13278 19016 13415 ne
rect 19016 13360 19071 13415
tri 19071 13360 19246 13535 sw
tri 19309 13415 19429 13535 ne
rect 19429 13415 19465 13535
rect 19585 13433 19621 13535
tri 19621 13433 19723 13535 sw
rect 19585 13415 20300 13433
rect 19016 13278 19246 13360
tri 19246 13278 19328 13360 sw
tri 19429 13278 19566 13415 ne
rect 19566 13278 20300 13415
rect -2000 13122 78 13278
tri 78 13122 234 13278 sw
tri 316 13122 472 13278 ne
rect 472 13122 628 13278
tri 628 13122 784 13278 sw
tri 866 13122 1022 13278 ne
rect 1022 13122 1178 13278
tri 1178 13122 1334 13278 sw
tri 1416 13122 1572 13278 ne
rect 1572 13122 1728 13278
tri 1728 13122 1884 13278 sw
tri 1966 13122 2122 13278 ne
rect 2122 13122 2278 13278
tri 2278 13122 2434 13278 sw
tri 2516 13122 2672 13278 ne
rect 2672 13122 2828 13278
tri 2828 13122 2984 13278 sw
tri 3066 13122 3222 13278 ne
rect 3222 13122 3378 13278
tri 3378 13122 3534 13278 sw
tri 3616 13122 3772 13278 ne
rect 3772 13122 3928 13278
tri 3928 13122 4084 13278 sw
tri 4166 13122 4322 13278 ne
rect 4322 13122 4478 13278
tri 4478 13122 4634 13278 sw
tri 4716 13122 4872 13278 ne
rect 4872 13122 5028 13278
tri 5028 13122 5184 13278 sw
tri 5266 13122 5422 13278 ne
rect 5422 13122 5578 13278
tri 5578 13122 5734 13278 sw
tri 5816 13122 5972 13278 ne
rect 5972 13122 6128 13278
tri 6128 13122 6284 13278 sw
tri 6366 13122 6522 13278 ne
rect 6522 13122 6678 13278
tri 6678 13122 6834 13278 sw
tri 6916 13122 7072 13278 ne
rect 7072 13122 7228 13278
tri 7228 13122 7384 13278 sw
tri 7466 13122 7622 13278 ne
rect 7622 13122 7778 13278
tri 7778 13122 7934 13278 sw
tri 8016 13122 8172 13278 ne
rect 8172 13122 8328 13278
tri 8328 13122 8484 13278 sw
tri 8566 13122 8722 13278 ne
rect 8722 13122 8878 13278
tri 8878 13122 9034 13278 sw
tri 9116 13122 9272 13278 ne
rect 9272 13122 9428 13278
tri 9428 13122 9584 13278 sw
tri 9666 13122 9822 13278 ne
rect 9822 13122 9978 13278
tri 9978 13122 10134 13278 sw
tri 10216 13122 10372 13278 ne
rect 10372 13122 10528 13278
tri 10528 13122 10684 13278 sw
tri 10766 13122 10922 13278 ne
rect 10922 13122 11078 13278
tri 11078 13122 11234 13278 sw
tri 11316 13122 11472 13278 ne
rect 11472 13122 11628 13278
tri 11628 13122 11784 13278 sw
tri 11866 13122 12022 13278 ne
rect 12022 13122 12178 13278
tri 12178 13122 12334 13278 sw
tri 12416 13122 12572 13278 ne
rect 12572 13122 12728 13278
tri 12728 13122 12884 13278 sw
tri 12966 13122 13122 13278 ne
rect 13122 13122 13278 13278
tri 13278 13122 13434 13278 sw
tri 13516 13122 13672 13278 ne
rect 13672 13122 13828 13278
tri 13828 13122 13984 13278 sw
tri 14066 13122 14222 13278 ne
rect 14222 13122 14378 13278
tri 14378 13122 14534 13278 sw
tri 14616 13122 14772 13278 ne
rect 14772 13122 14928 13278
tri 14928 13122 15084 13278 sw
tri 15166 13122 15322 13278 ne
rect 15322 13122 15478 13278
tri 15478 13122 15634 13278 sw
tri 15716 13122 15872 13278 ne
rect 15872 13122 16028 13278
tri 16028 13122 16184 13278 sw
tri 16266 13122 16422 13278 ne
rect 16422 13122 16578 13278
tri 16578 13122 16734 13278 sw
tri 16816 13122 16972 13278 ne
rect 16972 13122 17128 13278
tri 17128 13122 17284 13278 sw
tri 17366 13122 17522 13278 ne
rect 17522 13122 17678 13278
tri 17678 13122 17834 13278 sw
tri 17916 13122 18072 13278 ne
rect 18072 13122 18228 13278
tri 18228 13122 18384 13278 sw
tri 18466 13122 18622 13278 ne
rect 18622 13122 18778 13278
tri 18778 13122 18934 13278 sw
tri 19016 13122 19172 13278 ne
rect 19172 13122 19328 13278
tri 19328 13122 19484 13278 sw
tri 19566 13122 19722 13278 ne
rect 19722 13122 20300 13278
rect -2000 12985 234 13122
tri 234 12985 371 13122 sw
tri 472 12985 609 13122 ne
rect 609 12985 784 13122
tri 784 12985 921 13122 sw
tri 1022 12985 1159 13122 ne
rect 1159 12985 1334 13122
tri 1334 12985 1471 13122 sw
tri 1572 12985 1709 13122 ne
rect 1709 12985 1884 13122
tri 1884 12985 2021 13122 sw
tri 2122 12985 2259 13122 ne
rect 2259 12985 2434 13122
tri 2434 12985 2571 13122 sw
tri 2672 12985 2809 13122 ne
rect 2809 12985 2984 13122
tri 2984 12985 3121 13122 sw
tri 3222 12985 3359 13122 ne
rect 3359 12985 3534 13122
tri 3534 12985 3671 13122 sw
tri 3772 12985 3909 13122 ne
rect 3909 12985 4084 13122
tri 4084 12985 4221 13122 sw
tri 4322 12985 4459 13122 ne
rect 4459 12985 4634 13122
tri 4634 12985 4771 13122 sw
tri 4872 12985 5009 13122 ne
rect 5009 12985 5184 13122
tri 5184 12985 5321 13122 sw
tri 5422 12985 5559 13122 ne
rect 5559 12985 5734 13122
tri 5734 12985 5871 13122 sw
tri 5972 12985 6109 13122 ne
rect 6109 12985 6284 13122
tri 6284 12985 6421 13122 sw
tri 6522 12985 6659 13122 ne
rect 6659 12985 6834 13122
tri 6834 12985 6971 13122 sw
tri 7072 12985 7209 13122 ne
rect 7209 12985 7384 13122
tri 7384 12985 7521 13122 sw
tri 7622 12985 7759 13122 ne
rect 7759 12985 7934 13122
tri 7934 12985 8071 13122 sw
tri 8172 12985 8309 13122 ne
rect 8309 12985 8484 13122
tri 8484 12985 8621 13122 sw
tri 8722 12985 8859 13122 ne
rect 8859 12985 9034 13122
tri 9034 12985 9171 13122 sw
tri 9272 12985 9409 13122 ne
rect 9409 12985 9584 13122
tri 9584 12985 9721 13122 sw
tri 9822 12985 9959 13122 ne
rect 9959 12985 10134 13122
tri 10134 12985 10271 13122 sw
tri 10372 12985 10509 13122 ne
rect 10509 12985 10684 13122
tri 10684 12985 10821 13122 sw
tri 10922 12985 11059 13122 ne
rect 11059 12985 11234 13122
tri 11234 12985 11371 13122 sw
tri 11472 12985 11609 13122 ne
rect 11609 12985 11784 13122
tri 11784 12985 11921 13122 sw
tri 12022 12985 12159 13122 ne
rect 12159 12985 12334 13122
tri 12334 12985 12471 13122 sw
tri 12572 12985 12709 13122 ne
rect 12709 12985 12884 13122
tri 12884 12985 13021 13122 sw
tri 13122 12985 13259 13122 ne
rect 13259 12985 13434 13122
tri 13434 12985 13571 13122 sw
tri 13672 12985 13809 13122 ne
rect 13809 12985 13984 13122
tri 13984 12985 14121 13122 sw
tri 14222 12985 14359 13122 ne
rect 14359 12985 14534 13122
tri 14534 12985 14671 13122 sw
tri 14772 12985 14909 13122 ne
rect 14909 12985 15084 13122
tri 15084 12985 15221 13122 sw
tri 15322 12985 15459 13122 ne
rect 15459 12985 15634 13122
tri 15634 12985 15771 13122 sw
tri 15872 12985 16009 13122 ne
rect 16009 12985 16184 13122
tri 16184 12985 16321 13122 sw
tri 16422 12985 16559 13122 ne
rect 16559 12985 16734 13122
tri 16734 12985 16871 13122 sw
tri 16972 12985 17109 13122 ne
rect 17109 12985 17284 13122
tri 17284 12985 17421 13122 sw
tri 17522 12985 17659 13122 ne
rect 17659 12985 17834 13122
tri 17834 12985 17971 13122 sw
tri 18072 12985 18209 13122 ne
rect 18209 12985 18384 13122
tri 18384 12985 18521 13122 sw
tri 18622 12985 18759 13122 ne
rect 18759 12985 18934 13122
tri 18934 12985 19071 13122 sw
tri 19172 12985 19309 13122 ne
rect 19309 12985 19484 13122
tri 19484 12985 19621 13122 sw
rect -2000 12967 215 12985
rect -2000 12178 -1000 12967
tri 77 12865 179 12967 ne
rect 179 12865 215 12967
rect 335 12865 371 12985
tri 179 12728 316 12865 ne
rect 316 12810 371 12865
tri 371 12810 546 12985 sw
tri 609 12865 729 12985 ne
rect 729 12865 765 12985
rect 885 12865 921 12985
rect 316 12728 546 12810
tri 546 12728 628 12810 sw
tri 729 12728 866 12865 ne
rect 866 12810 921 12865
tri 921 12810 1096 12985 sw
tri 1159 12865 1279 12985 ne
rect 1279 12865 1315 12985
rect 1435 12865 1471 12985
rect 866 12728 1096 12810
tri 1096 12728 1178 12810 sw
tri 1279 12728 1416 12865 ne
rect 1416 12810 1471 12865
tri 1471 12810 1646 12985 sw
tri 1709 12865 1829 12985 ne
rect 1829 12865 1865 12985
rect 1985 12865 2021 12985
rect 1416 12728 1646 12810
tri 1646 12728 1728 12810 sw
tri 1829 12728 1966 12865 ne
rect 1966 12810 2021 12865
tri 2021 12810 2196 12985 sw
tri 2259 12865 2379 12985 ne
rect 2379 12865 2415 12985
rect 2535 12865 2571 12985
rect 1966 12728 2196 12810
tri 2196 12728 2278 12810 sw
tri 2379 12728 2516 12865 ne
rect 2516 12810 2571 12865
tri 2571 12810 2746 12985 sw
tri 2809 12865 2929 12985 ne
rect 2929 12865 2965 12985
rect 3085 12865 3121 12985
rect 2516 12728 2746 12810
tri 2746 12728 2828 12810 sw
tri 2929 12728 3066 12865 ne
rect 3066 12810 3121 12865
tri 3121 12810 3296 12985 sw
tri 3359 12865 3479 12985 ne
rect 3479 12865 3515 12985
rect 3635 12865 3671 12985
rect 3066 12728 3296 12810
tri 3296 12728 3378 12810 sw
tri 3479 12728 3616 12865 ne
rect 3616 12810 3671 12865
tri 3671 12810 3846 12985 sw
tri 3909 12865 4029 12985 ne
rect 4029 12865 4065 12985
rect 4185 12865 4221 12985
rect 3616 12728 3846 12810
tri 3846 12728 3928 12810 sw
tri 4029 12728 4166 12865 ne
rect 4166 12810 4221 12865
tri 4221 12810 4396 12985 sw
tri 4459 12865 4579 12985 ne
rect 4579 12865 4615 12985
rect 4735 12865 4771 12985
rect 4166 12728 4396 12810
tri 4396 12728 4478 12810 sw
tri 4579 12728 4716 12865 ne
rect 4716 12810 4771 12865
tri 4771 12810 4946 12985 sw
tri 5009 12865 5129 12985 ne
rect 5129 12865 5165 12985
rect 5285 12865 5321 12985
rect 4716 12728 4946 12810
tri 4946 12728 5028 12810 sw
tri 5129 12728 5266 12865 ne
rect 5266 12810 5321 12865
tri 5321 12810 5496 12985 sw
tri 5559 12865 5679 12985 ne
rect 5679 12865 5715 12985
rect 5835 12865 5871 12985
rect 5266 12728 5496 12810
tri 5496 12728 5578 12810 sw
tri 5679 12728 5816 12865 ne
rect 5816 12810 5871 12865
tri 5871 12810 6046 12985 sw
tri 6109 12865 6229 12985 ne
rect 6229 12865 6265 12985
rect 6385 12865 6421 12985
rect 5816 12728 6046 12810
tri 6046 12728 6128 12810 sw
tri 6229 12728 6366 12865 ne
rect 6366 12810 6421 12865
tri 6421 12810 6596 12985 sw
tri 6659 12865 6779 12985 ne
rect 6779 12865 6815 12985
rect 6935 12865 6971 12985
rect 6366 12728 6596 12810
tri 6596 12728 6678 12810 sw
tri 6779 12728 6916 12865 ne
rect 6916 12810 6971 12865
tri 6971 12810 7146 12985 sw
tri 7209 12865 7329 12985 ne
rect 7329 12865 7365 12985
rect 7485 12865 7521 12985
rect 6916 12728 7146 12810
tri 7146 12728 7228 12810 sw
tri 7329 12728 7466 12865 ne
rect 7466 12810 7521 12865
tri 7521 12810 7696 12985 sw
tri 7759 12865 7879 12985 ne
rect 7879 12865 7915 12985
rect 8035 12865 8071 12985
rect 7466 12728 7696 12810
tri 7696 12728 7778 12810 sw
tri 7879 12728 8016 12865 ne
rect 8016 12810 8071 12865
tri 8071 12810 8246 12985 sw
tri 8309 12865 8429 12985 ne
rect 8429 12865 8465 12985
rect 8585 12865 8621 12985
rect 8016 12728 8246 12810
tri 8246 12728 8328 12810 sw
tri 8429 12728 8566 12865 ne
rect 8566 12810 8621 12865
tri 8621 12810 8796 12985 sw
tri 8859 12865 8979 12985 ne
rect 8979 12865 9015 12985
rect 9135 12865 9171 12985
rect 8566 12728 8796 12810
tri 8796 12728 8878 12810 sw
tri 8979 12728 9116 12865 ne
rect 9116 12810 9171 12865
tri 9171 12810 9346 12985 sw
tri 9409 12865 9529 12985 ne
rect 9529 12865 9565 12985
rect 9685 12865 9721 12985
rect 9116 12728 9346 12810
tri 9346 12728 9428 12810 sw
tri 9529 12728 9666 12865 ne
rect 9666 12810 9721 12865
tri 9721 12810 9896 12985 sw
tri 9959 12865 10079 12985 ne
rect 10079 12865 10115 12985
rect 10235 12865 10271 12985
rect 9666 12728 9896 12810
tri 9896 12728 9978 12810 sw
tri 10079 12728 10216 12865 ne
rect 10216 12810 10271 12865
tri 10271 12810 10446 12985 sw
tri 10509 12865 10629 12985 ne
rect 10629 12865 10665 12985
rect 10785 12865 10821 12985
rect 10216 12728 10446 12810
tri 10446 12728 10528 12810 sw
tri 10629 12728 10766 12865 ne
rect 10766 12810 10821 12865
tri 10821 12810 10996 12985 sw
tri 11059 12865 11179 12985 ne
rect 11179 12865 11215 12985
rect 11335 12865 11371 12985
rect 10766 12728 10996 12810
tri 10996 12728 11078 12810 sw
tri 11179 12728 11316 12865 ne
rect 11316 12810 11371 12865
tri 11371 12810 11546 12985 sw
tri 11609 12865 11729 12985 ne
rect 11729 12865 11765 12985
rect 11885 12865 11921 12985
rect 11316 12728 11546 12810
tri 11546 12728 11628 12810 sw
tri 11729 12728 11866 12865 ne
rect 11866 12810 11921 12865
tri 11921 12810 12096 12985 sw
tri 12159 12865 12279 12985 ne
rect 12279 12865 12315 12985
rect 12435 12865 12471 12985
rect 11866 12728 12096 12810
tri 12096 12728 12178 12810 sw
tri 12279 12728 12416 12865 ne
rect 12416 12810 12471 12865
tri 12471 12810 12646 12985 sw
tri 12709 12865 12829 12985 ne
rect 12829 12865 12865 12985
rect 12985 12865 13021 12985
rect 12416 12728 12646 12810
tri 12646 12728 12728 12810 sw
tri 12829 12728 12966 12865 ne
rect 12966 12810 13021 12865
tri 13021 12810 13196 12985 sw
tri 13259 12865 13379 12985 ne
rect 13379 12865 13415 12985
rect 13535 12865 13571 12985
rect 12966 12728 13196 12810
tri 13196 12728 13278 12810 sw
tri 13379 12728 13516 12865 ne
rect 13516 12810 13571 12865
tri 13571 12810 13746 12985 sw
tri 13809 12865 13929 12985 ne
rect 13929 12865 13965 12985
rect 14085 12865 14121 12985
rect 13516 12728 13746 12810
tri 13746 12728 13828 12810 sw
tri 13929 12728 14066 12865 ne
rect 14066 12810 14121 12865
tri 14121 12810 14296 12985 sw
tri 14359 12865 14479 12985 ne
rect 14479 12865 14515 12985
rect 14635 12865 14671 12985
rect 14066 12728 14296 12810
tri 14296 12728 14378 12810 sw
tri 14479 12728 14616 12865 ne
rect 14616 12810 14671 12865
tri 14671 12810 14846 12985 sw
tri 14909 12865 15029 12985 ne
rect 15029 12865 15065 12985
rect 15185 12865 15221 12985
rect 14616 12728 14846 12810
tri 14846 12728 14928 12810 sw
tri 15029 12728 15166 12865 ne
rect 15166 12810 15221 12865
tri 15221 12810 15396 12985 sw
tri 15459 12865 15579 12985 ne
rect 15579 12865 15615 12985
rect 15735 12865 15771 12985
rect 15166 12728 15396 12810
tri 15396 12728 15478 12810 sw
tri 15579 12728 15716 12865 ne
rect 15716 12810 15771 12865
tri 15771 12810 15946 12985 sw
tri 16009 12865 16129 12985 ne
rect 16129 12865 16165 12985
rect 16285 12865 16321 12985
rect 15716 12728 15946 12810
tri 15946 12728 16028 12810 sw
tri 16129 12728 16266 12865 ne
rect 16266 12810 16321 12865
tri 16321 12810 16496 12985 sw
tri 16559 12865 16679 12985 ne
rect 16679 12865 16715 12985
rect 16835 12865 16871 12985
rect 16266 12728 16496 12810
tri 16496 12728 16578 12810 sw
tri 16679 12728 16816 12865 ne
rect 16816 12810 16871 12865
tri 16871 12810 17046 12985 sw
tri 17109 12865 17229 12985 ne
rect 17229 12865 17265 12985
rect 17385 12865 17421 12985
rect 16816 12728 17046 12810
tri 17046 12728 17128 12810 sw
tri 17229 12728 17366 12865 ne
rect 17366 12810 17421 12865
tri 17421 12810 17596 12985 sw
tri 17659 12865 17779 12985 ne
rect 17779 12865 17815 12985
rect 17935 12865 17971 12985
rect 17366 12728 17596 12810
tri 17596 12728 17678 12810 sw
tri 17779 12728 17916 12865 ne
rect 17916 12810 17971 12865
tri 17971 12810 18146 12985 sw
tri 18209 12865 18329 12985 ne
rect 18329 12865 18365 12985
rect 18485 12865 18521 12985
rect 17916 12728 18146 12810
tri 18146 12728 18228 12810 sw
tri 18329 12728 18466 12865 ne
rect 18466 12810 18521 12865
tri 18521 12810 18696 12985 sw
tri 18759 12865 18879 12985 ne
rect 18879 12865 18915 12985
rect 19035 12865 19071 12985
rect 18466 12728 18696 12810
tri 18696 12728 18778 12810 sw
tri 18879 12728 19016 12865 ne
rect 19016 12810 19071 12865
tri 19071 12810 19246 12985 sw
tri 19309 12865 19429 12985 ne
rect 19429 12865 19465 12985
rect 19585 12883 19621 12985
tri 19621 12883 19723 12985 sw
rect 20800 12883 21800 13672
rect 19585 12865 21800 12883
rect 19016 12728 19246 12810
tri 19246 12728 19328 12810 sw
tri 19429 12728 19566 12865 ne
rect 19566 12728 21800 12865
rect -500 12572 78 12728
tri 78 12572 234 12728 sw
tri 316 12572 472 12728 ne
rect 472 12572 628 12728
tri 628 12572 784 12728 sw
tri 866 12572 1022 12728 ne
rect 1022 12572 1178 12728
tri 1178 12572 1334 12728 sw
tri 1416 12572 1572 12728 ne
rect 1572 12572 1728 12728
tri 1728 12572 1884 12728 sw
tri 1966 12572 2122 12728 ne
rect 2122 12572 2278 12728
tri 2278 12572 2434 12728 sw
tri 2516 12572 2672 12728 ne
rect 2672 12572 2828 12728
tri 2828 12572 2984 12728 sw
tri 3066 12572 3222 12728 ne
rect 3222 12572 3378 12728
tri 3378 12572 3534 12728 sw
tri 3616 12572 3772 12728 ne
rect 3772 12572 3928 12728
tri 3928 12572 4084 12728 sw
tri 4166 12572 4322 12728 ne
rect 4322 12572 4478 12728
tri 4478 12572 4634 12728 sw
tri 4716 12572 4872 12728 ne
rect 4872 12572 5028 12728
tri 5028 12572 5184 12728 sw
tri 5266 12572 5422 12728 ne
rect 5422 12572 5578 12728
tri 5578 12572 5734 12728 sw
tri 5816 12572 5972 12728 ne
rect 5972 12572 6128 12728
tri 6128 12572 6284 12728 sw
tri 6366 12572 6522 12728 ne
rect 6522 12572 6678 12728
tri 6678 12572 6834 12728 sw
tri 6916 12572 7072 12728 ne
rect 7072 12572 7228 12728
tri 7228 12572 7384 12728 sw
tri 7466 12572 7622 12728 ne
rect 7622 12572 7778 12728
tri 7778 12572 7934 12728 sw
tri 8016 12572 8172 12728 ne
rect 8172 12572 8328 12728
tri 8328 12572 8484 12728 sw
tri 8566 12572 8722 12728 ne
rect 8722 12572 8878 12728
tri 8878 12572 9034 12728 sw
tri 9116 12572 9272 12728 ne
rect 9272 12572 9428 12728
tri 9428 12572 9584 12728 sw
tri 9666 12572 9822 12728 ne
rect 9822 12572 9978 12728
tri 9978 12572 10134 12728 sw
tri 10216 12572 10372 12728 ne
rect 10372 12572 10528 12728
tri 10528 12572 10684 12728 sw
tri 10766 12572 10922 12728 ne
rect 10922 12572 11078 12728
tri 11078 12572 11234 12728 sw
tri 11316 12572 11472 12728 ne
rect 11472 12572 11628 12728
tri 11628 12572 11784 12728 sw
tri 11866 12572 12022 12728 ne
rect 12022 12572 12178 12728
tri 12178 12572 12334 12728 sw
tri 12416 12572 12572 12728 ne
rect 12572 12572 12728 12728
tri 12728 12572 12884 12728 sw
tri 12966 12572 13122 12728 ne
rect 13122 12572 13278 12728
tri 13278 12572 13434 12728 sw
tri 13516 12572 13672 12728 ne
rect 13672 12572 13828 12728
tri 13828 12572 13984 12728 sw
tri 14066 12572 14222 12728 ne
rect 14222 12572 14378 12728
tri 14378 12572 14534 12728 sw
tri 14616 12572 14772 12728 ne
rect 14772 12572 14928 12728
tri 14928 12572 15084 12728 sw
tri 15166 12572 15322 12728 ne
rect 15322 12572 15478 12728
tri 15478 12572 15634 12728 sw
tri 15716 12572 15872 12728 ne
rect 15872 12572 16028 12728
tri 16028 12572 16184 12728 sw
tri 16266 12572 16422 12728 ne
rect 16422 12572 16578 12728
tri 16578 12572 16734 12728 sw
tri 16816 12572 16972 12728 ne
rect 16972 12572 17128 12728
tri 17128 12572 17284 12728 sw
tri 17366 12572 17522 12728 ne
rect 17522 12572 17678 12728
tri 17678 12572 17834 12728 sw
tri 17916 12572 18072 12728 ne
rect 18072 12572 18228 12728
tri 18228 12572 18384 12728 sw
tri 18466 12572 18622 12728 ne
rect 18622 12572 18778 12728
tri 18778 12572 18934 12728 sw
tri 19016 12572 19172 12728 ne
rect 19172 12572 19328 12728
tri 19328 12572 19484 12728 sw
tri 19566 12572 19722 12728 ne
rect 19722 12572 21800 12728
rect -500 12435 234 12572
tri 234 12435 371 12572 sw
tri 472 12435 609 12572 ne
rect 609 12435 784 12572
tri 784 12435 921 12572 sw
tri 1022 12435 1159 12572 ne
rect 1159 12435 1334 12572
tri 1334 12435 1471 12572 sw
tri 1572 12435 1709 12572 ne
rect 1709 12435 1884 12572
tri 1884 12435 2021 12572 sw
tri 2122 12435 2259 12572 ne
rect 2259 12435 2434 12572
tri 2434 12435 2571 12572 sw
tri 2672 12435 2809 12572 ne
rect 2809 12435 2984 12572
tri 2984 12435 3121 12572 sw
tri 3222 12435 3359 12572 ne
rect 3359 12435 3534 12572
tri 3534 12435 3671 12572 sw
tri 3772 12435 3909 12572 ne
rect 3909 12435 4084 12572
tri 4084 12435 4221 12572 sw
tri 4322 12435 4459 12572 ne
rect 4459 12435 4634 12572
tri 4634 12435 4771 12572 sw
tri 4872 12435 5009 12572 ne
rect 5009 12435 5184 12572
tri 5184 12435 5321 12572 sw
tri 5422 12435 5559 12572 ne
rect 5559 12435 5734 12572
tri 5734 12435 5871 12572 sw
tri 5972 12435 6109 12572 ne
rect 6109 12435 6284 12572
tri 6284 12435 6421 12572 sw
tri 6522 12435 6659 12572 ne
rect 6659 12435 6834 12572
tri 6834 12435 6971 12572 sw
tri 7072 12435 7209 12572 ne
rect 7209 12435 7384 12572
tri 7384 12435 7521 12572 sw
tri 7622 12435 7759 12572 ne
rect 7759 12435 7934 12572
tri 7934 12435 8071 12572 sw
tri 8172 12435 8309 12572 ne
rect 8309 12435 8484 12572
tri 8484 12435 8621 12572 sw
tri 8722 12435 8859 12572 ne
rect 8859 12435 9034 12572
tri 9034 12435 9171 12572 sw
tri 9272 12435 9409 12572 ne
rect 9409 12435 9584 12572
tri 9584 12435 9721 12572 sw
tri 9822 12435 9959 12572 ne
rect 9959 12435 10134 12572
tri 10134 12435 10271 12572 sw
tri 10372 12435 10509 12572 ne
rect 10509 12435 10684 12572
tri 10684 12435 10821 12572 sw
tri 10922 12435 11059 12572 ne
rect 11059 12435 11234 12572
tri 11234 12435 11371 12572 sw
tri 11472 12435 11609 12572 ne
rect 11609 12435 11784 12572
tri 11784 12435 11921 12572 sw
tri 12022 12435 12159 12572 ne
rect 12159 12435 12334 12572
tri 12334 12435 12471 12572 sw
tri 12572 12435 12709 12572 ne
rect 12709 12435 12884 12572
tri 12884 12435 13021 12572 sw
tri 13122 12435 13259 12572 ne
rect 13259 12435 13434 12572
tri 13434 12435 13571 12572 sw
tri 13672 12435 13809 12572 ne
rect 13809 12435 13984 12572
tri 13984 12435 14121 12572 sw
tri 14222 12435 14359 12572 ne
rect 14359 12435 14534 12572
tri 14534 12435 14671 12572 sw
tri 14772 12435 14909 12572 ne
rect 14909 12435 15084 12572
tri 15084 12435 15221 12572 sw
tri 15322 12435 15459 12572 ne
rect 15459 12435 15634 12572
tri 15634 12435 15771 12572 sw
tri 15872 12435 16009 12572 ne
rect 16009 12435 16184 12572
tri 16184 12435 16321 12572 sw
tri 16422 12435 16559 12572 ne
rect 16559 12435 16734 12572
tri 16734 12435 16871 12572 sw
tri 16972 12435 17109 12572 ne
rect 17109 12435 17284 12572
tri 17284 12435 17421 12572 sw
tri 17522 12435 17659 12572 ne
rect 17659 12435 17834 12572
tri 17834 12435 17971 12572 sw
tri 18072 12435 18209 12572 ne
rect 18209 12435 18384 12572
tri 18384 12435 18521 12572 sw
tri 18622 12435 18759 12572 ne
rect 18759 12435 18934 12572
tri 18934 12435 19071 12572 sw
tri 19172 12435 19309 12572 ne
rect 19309 12435 19484 12572
tri 19484 12435 19621 12572 sw
rect -500 12417 215 12435
tri 77 12315 179 12417 ne
rect 179 12315 215 12417
rect 335 12315 371 12435
tri 179 12178 316 12315 ne
rect 316 12260 371 12315
tri 371 12260 546 12435 sw
tri 609 12315 729 12435 ne
rect 729 12315 765 12435
rect 885 12315 921 12435
rect 316 12178 546 12260
tri 546 12178 628 12260 sw
tri 729 12178 866 12315 ne
rect 866 12260 921 12315
tri 921 12260 1096 12435 sw
tri 1159 12315 1279 12435 ne
rect 1279 12315 1315 12435
rect 1435 12315 1471 12435
rect 866 12178 1096 12260
tri 1096 12178 1178 12260 sw
tri 1279 12178 1416 12315 ne
rect 1416 12260 1471 12315
tri 1471 12260 1646 12435 sw
tri 1709 12315 1829 12435 ne
rect 1829 12315 1865 12435
rect 1985 12315 2021 12435
rect 1416 12178 1646 12260
tri 1646 12178 1728 12260 sw
tri 1829 12178 1966 12315 ne
rect 1966 12260 2021 12315
tri 2021 12260 2196 12435 sw
tri 2259 12315 2379 12435 ne
rect 2379 12315 2415 12435
rect 2535 12315 2571 12435
rect 1966 12178 2196 12260
tri 2196 12178 2278 12260 sw
tri 2379 12178 2516 12315 ne
rect 2516 12260 2571 12315
tri 2571 12260 2746 12435 sw
tri 2809 12315 2929 12435 ne
rect 2929 12315 2965 12435
rect 3085 12315 3121 12435
rect 2516 12178 2746 12260
tri 2746 12178 2828 12260 sw
tri 2929 12178 3066 12315 ne
rect 3066 12260 3121 12315
tri 3121 12260 3296 12435 sw
tri 3359 12315 3479 12435 ne
rect 3479 12315 3515 12435
rect 3635 12315 3671 12435
rect 3066 12178 3296 12260
tri 3296 12178 3378 12260 sw
tri 3479 12178 3616 12315 ne
rect 3616 12260 3671 12315
tri 3671 12260 3846 12435 sw
tri 3909 12315 4029 12435 ne
rect 4029 12315 4065 12435
rect 4185 12315 4221 12435
rect 3616 12178 3846 12260
tri 3846 12178 3928 12260 sw
tri 4029 12178 4166 12315 ne
rect 4166 12260 4221 12315
tri 4221 12260 4396 12435 sw
tri 4459 12315 4579 12435 ne
rect 4579 12315 4615 12435
rect 4735 12315 4771 12435
rect 4166 12178 4396 12260
tri 4396 12178 4478 12260 sw
tri 4579 12178 4716 12315 ne
rect 4716 12260 4771 12315
tri 4771 12260 4946 12435 sw
tri 5009 12315 5129 12435 ne
rect 5129 12315 5165 12435
rect 5285 12315 5321 12435
rect 4716 12178 4946 12260
tri 4946 12178 5028 12260 sw
tri 5129 12178 5266 12315 ne
rect 5266 12260 5321 12315
tri 5321 12260 5496 12435 sw
tri 5559 12315 5679 12435 ne
rect 5679 12315 5715 12435
rect 5835 12315 5871 12435
rect 5266 12178 5496 12260
tri 5496 12178 5578 12260 sw
tri 5679 12178 5816 12315 ne
rect 5816 12260 5871 12315
tri 5871 12260 6046 12435 sw
tri 6109 12315 6229 12435 ne
rect 6229 12315 6265 12435
rect 6385 12315 6421 12435
rect 5816 12178 6046 12260
tri 6046 12178 6128 12260 sw
tri 6229 12178 6366 12315 ne
rect 6366 12260 6421 12315
tri 6421 12260 6596 12435 sw
tri 6659 12315 6779 12435 ne
rect 6779 12315 6815 12435
rect 6935 12315 6971 12435
rect 6366 12178 6596 12260
tri 6596 12178 6678 12260 sw
tri 6779 12178 6916 12315 ne
rect 6916 12260 6971 12315
tri 6971 12260 7146 12435 sw
tri 7209 12315 7329 12435 ne
rect 7329 12315 7365 12435
rect 7485 12315 7521 12435
rect 6916 12178 7146 12260
tri 7146 12178 7228 12260 sw
tri 7329 12178 7466 12315 ne
rect 7466 12260 7521 12315
tri 7521 12260 7696 12435 sw
tri 7759 12315 7879 12435 ne
rect 7879 12315 7915 12435
rect 8035 12315 8071 12435
rect 7466 12178 7696 12260
tri 7696 12178 7778 12260 sw
tri 7879 12178 8016 12315 ne
rect 8016 12260 8071 12315
tri 8071 12260 8246 12435 sw
tri 8309 12315 8429 12435 ne
rect 8429 12315 8465 12435
rect 8585 12315 8621 12435
rect 8016 12178 8246 12260
tri 8246 12178 8328 12260 sw
tri 8429 12178 8566 12315 ne
rect 8566 12260 8621 12315
tri 8621 12260 8796 12435 sw
tri 8859 12315 8979 12435 ne
rect 8979 12315 9015 12435
rect 9135 12315 9171 12435
rect 8566 12178 8796 12260
tri 8796 12178 8878 12260 sw
tri 8979 12178 9116 12315 ne
rect 9116 12260 9171 12315
tri 9171 12260 9346 12435 sw
tri 9409 12315 9529 12435 ne
rect 9529 12315 9565 12435
rect 9685 12315 9721 12435
rect 9116 12178 9346 12260
tri 9346 12178 9428 12260 sw
tri 9529 12178 9666 12315 ne
rect 9666 12260 9721 12315
tri 9721 12260 9896 12435 sw
tri 9959 12315 10079 12435 ne
rect 10079 12315 10115 12435
rect 10235 12315 10271 12435
rect 9666 12178 9896 12260
tri 9896 12178 9978 12260 sw
tri 10079 12178 10216 12315 ne
rect 10216 12260 10271 12315
tri 10271 12260 10446 12435 sw
tri 10509 12315 10629 12435 ne
rect 10629 12315 10665 12435
rect 10785 12315 10821 12435
rect 10216 12178 10446 12260
tri 10446 12178 10528 12260 sw
tri 10629 12178 10766 12315 ne
rect 10766 12260 10821 12315
tri 10821 12260 10996 12435 sw
tri 11059 12315 11179 12435 ne
rect 11179 12315 11215 12435
rect 11335 12315 11371 12435
rect 10766 12178 10996 12260
tri 10996 12178 11078 12260 sw
tri 11179 12178 11316 12315 ne
rect 11316 12260 11371 12315
tri 11371 12260 11546 12435 sw
tri 11609 12315 11729 12435 ne
rect 11729 12315 11765 12435
rect 11885 12315 11921 12435
rect 11316 12178 11546 12260
tri 11546 12178 11628 12260 sw
tri 11729 12178 11866 12315 ne
rect 11866 12260 11921 12315
tri 11921 12260 12096 12435 sw
tri 12159 12315 12279 12435 ne
rect 12279 12315 12315 12435
rect 12435 12315 12471 12435
rect 11866 12178 12096 12260
tri 12096 12178 12178 12260 sw
tri 12279 12178 12416 12315 ne
rect 12416 12260 12471 12315
tri 12471 12260 12646 12435 sw
tri 12709 12315 12829 12435 ne
rect 12829 12315 12865 12435
rect 12985 12315 13021 12435
rect 12416 12178 12646 12260
tri 12646 12178 12728 12260 sw
tri 12829 12178 12966 12315 ne
rect 12966 12260 13021 12315
tri 13021 12260 13196 12435 sw
tri 13259 12315 13379 12435 ne
rect 13379 12315 13415 12435
rect 13535 12315 13571 12435
rect 12966 12178 13196 12260
tri 13196 12178 13278 12260 sw
tri 13379 12178 13516 12315 ne
rect 13516 12260 13571 12315
tri 13571 12260 13746 12435 sw
tri 13809 12315 13929 12435 ne
rect 13929 12315 13965 12435
rect 14085 12315 14121 12435
rect 13516 12178 13746 12260
tri 13746 12178 13828 12260 sw
tri 13929 12178 14066 12315 ne
rect 14066 12260 14121 12315
tri 14121 12260 14296 12435 sw
tri 14359 12315 14479 12435 ne
rect 14479 12315 14515 12435
rect 14635 12315 14671 12435
rect 14066 12178 14296 12260
tri 14296 12178 14378 12260 sw
tri 14479 12178 14616 12315 ne
rect 14616 12260 14671 12315
tri 14671 12260 14846 12435 sw
tri 14909 12315 15029 12435 ne
rect 15029 12315 15065 12435
rect 15185 12315 15221 12435
rect 14616 12178 14846 12260
tri 14846 12178 14928 12260 sw
tri 15029 12178 15166 12315 ne
rect 15166 12260 15221 12315
tri 15221 12260 15396 12435 sw
tri 15459 12315 15579 12435 ne
rect 15579 12315 15615 12435
rect 15735 12315 15771 12435
rect 15166 12178 15396 12260
tri 15396 12178 15478 12260 sw
tri 15579 12178 15716 12315 ne
rect 15716 12260 15771 12315
tri 15771 12260 15946 12435 sw
tri 16009 12315 16129 12435 ne
rect 16129 12315 16165 12435
rect 16285 12315 16321 12435
rect 15716 12178 15946 12260
tri 15946 12178 16028 12260 sw
tri 16129 12178 16266 12315 ne
rect 16266 12260 16321 12315
tri 16321 12260 16496 12435 sw
tri 16559 12315 16679 12435 ne
rect 16679 12315 16715 12435
rect 16835 12315 16871 12435
rect 16266 12178 16496 12260
tri 16496 12178 16578 12260 sw
tri 16679 12178 16816 12315 ne
rect 16816 12260 16871 12315
tri 16871 12260 17046 12435 sw
tri 17109 12315 17229 12435 ne
rect 17229 12315 17265 12435
rect 17385 12315 17421 12435
rect 16816 12178 17046 12260
tri 17046 12178 17128 12260 sw
tri 17229 12178 17366 12315 ne
rect 17366 12260 17421 12315
tri 17421 12260 17596 12435 sw
tri 17659 12315 17779 12435 ne
rect 17779 12315 17815 12435
rect 17935 12315 17971 12435
rect 17366 12178 17596 12260
tri 17596 12178 17678 12260 sw
tri 17779 12178 17916 12315 ne
rect 17916 12260 17971 12315
tri 17971 12260 18146 12435 sw
tri 18209 12315 18329 12435 ne
rect 18329 12315 18365 12435
rect 18485 12315 18521 12435
rect 17916 12178 18146 12260
tri 18146 12178 18228 12260 sw
tri 18329 12178 18466 12315 ne
rect 18466 12260 18521 12315
tri 18521 12260 18696 12435 sw
tri 18759 12315 18879 12435 ne
rect 18879 12315 18915 12435
rect 19035 12315 19071 12435
rect 18466 12178 18696 12260
tri 18696 12178 18778 12260 sw
tri 18879 12178 19016 12315 ne
rect 19016 12260 19071 12315
tri 19071 12260 19246 12435 sw
tri 19309 12315 19429 12435 ne
rect 19429 12315 19465 12435
rect 19585 12333 19621 12435
tri 19621 12333 19723 12435 sw
rect 19585 12315 20300 12333
rect 19016 12178 19246 12260
tri 19246 12178 19328 12260 sw
tri 19429 12178 19566 12315 ne
rect 19566 12178 20300 12315
rect -2000 12022 78 12178
tri 78 12022 234 12178 sw
tri 316 12022 472 12178 ne
rect 472 12022 628 12178
tri 628 12022 784 12178 sw
tri 866 12022 1022 12178 ne
rect 1022 12022 1178 12178
tri 1178 12022 1334 12178 sw
tri 1416 12022 1572 12178 ne
rect 1572 12022 1728 12178
tri 1728 12022 1884 12178 sw
tri 1966 12022 2122 12178 ne
rect 2122 12022 2278 12178
tri 2278 12022 2434 12178 sw
tri 2516 12022 2672 12178 ne
rect 2672 12022 2828 12178
tri 2828 12022 2984 12178 sw
tri 3066 12022 3222 12178 ne
rect 3222 12022 3378 12178
tri 3378 12022 3534 12178 sw
tri 3616 12022 3772 12178 ne
rect 3772 12022 3928 12178
tri 3928 12022 4084 12178 sw
tri 4166 12022 4322 12178 ne
rect 4322 12022 4478 12178
tri 4478 12022 4634 12178 sw
tri 4716 12022 4872 12178 ne
rect 4872 12022 5028 12178
tri 5028 12022 5184 12178 sw
tri 5266 12022 5422 12178 ne
rect 5422 12022 5578 12178
tri 5578 12022 5734 12178 sw
tri 5816 12022 5972 12178 ne
rect 5972 12022 6128 12178
tri 6128 12022 6284 12178 sw
tri 6366 12022 6522 12178 ne
rect 6522 12022 6678 12178
tri 6678 12022 6834 12178 sw
tri 6916 12022 7072 12178 ne
rect 7072 12022 7228 12178
tri 7228 12022 7384 12178 sw
tri 7466 12022 7622 12178 ne
rect 7622 12022 7778 12178
tri 7778 12022 7934 12178 sw
tri 8016 12022 8172 12178 ne
rect 8172 12022 8328 12178
tri 8328 12022 8484 12178 sw
tri 8566 12022 8722 12178 ne
rect 8722 12022 8878 12178
tri 8878 12022 9034 12178 sw
tri 9116 12022 9272 12178 ne
rect 9272 12022 9428 12178
tri 9428 12022 9584 12178 sw
tri 9666 12022 9822 12178 ne
rect 9822 12022 9978 12178
tri 9978 12022 10134 12178 sw
tri 10216 12022 10372 12178 ne
rect 10372 12022 10528 12178
tri 10528 12022 10684 12178 sw
tri 10766 12022 10922 12178 ne
rect 10922 12022 11078 12178
tri 11078 12022 11234 12178 sw
tri 11316 12022 11472 12178 ne
rect 11472 12022 11628 12178
tri 11628 12022 11784 12178 sw
tri 11866 12022 12022 12178 ne
rect 12022 12022 12178 12178
tri 12178 12022 12334 12178 sw
tri 12416 12022 12572 12178 ne
rect 12572 12022 12728 12178
tri 12728 12022 12884 12178 sw
tri 12966 12022 13122 12178 ne
rect 13122 12022 13278 12178
tri 13278 12022 13434 12178 sw
tri 13516 12022 13672 12178 ne
rect 13672 12022 13828 12178
tri 13828 12022 13984 12178 sw
tri 14066 12022 14222 12178 ne
rect 14222 12022 14378 12178
tri 14378 12022 14534 12178 sw
tri 14616 12022 14772 12178 ne
rect 14772 12022 14928 12178
tri 14928 12022 15084 12178 sw
tri 15166 12022 15322 12178 ne
rect 15322 12022 15478 12178
tri 15478 12022 15634 12178 sw
tri 15716 12022 15872 12178 ne
rect 15872 12022 16028 12178
tri 16028 12022 16184 12178 sw
tri 16266 12022 16422 12178 ne
rect 16422 12022 16578 12178
tri 16578 12022 16734 12178 sw
tri 16816 12022 16972 12178 ne
rect 16972 12022 17128 12178
tri 17128 12022 17284 12178 sw
tri 17366 12022 17522 12178 ne
rect 17522 12022 17678 12178
tri 17678 12022 17834 12178 sw
tri 17916 12022 18072 12178 ne
rect 18072 12022 18228 12178
tri 18228 12022 18384 12178 sw
tri 18466 12022 18622 12178 ne
rect 18622 12022 18778 12178
tri 18778 12022 18934 12178 sw
tri 19016 12022 19172 12178 ne
rect 19172 12022 19328 12178
tri 19328 12022 19484 12178 sw
tri 19566 12022 19722 12178 ne
rect 19722 12022 20300 12178
rect -2000 11885 234 12022
tri 234 11885 371 12022 sw
tri 472 11885 609 12022 ne
rect 609 11885 784 12022
tri 784 11885 921 12022 sw
tri 1022 11885 1159 12022 ne
rect 1159 11885 1334 12022
tri 1334 11885 1471 12022 sw
tri 1572 11885 1709 12022 ne
rect 1709 11885 1884 12022
tri 1884 11885 2021 12022 sw
tri 2122 11885 2259 12022 ne
rect 2259 11885 2434 12022
tri 2434 11885 2571 12022 sw
tri 2672 11885 2809 12022 ne
rect 2809 11885 2984 12022
tri 2984 11885 3121 12022 sw
tri 3222 11885 3359 12022 ne
rect 3359 11885 3534 12022
tri 3534 11885 3671 12022 sw
tri 3772 11885 3909 12022 ne
rect 3909 11885 4084 12022
tri 4084 11885 4221 12022 sw
tri 4322 11885 4459 12022 ne
rect 4459 11885 4634 12022
tri 4634 11885 4771 12022 sw
tri 4872 11885 5009 12022 ne
rect 5009 11885 5184 12022
tri 5184 11885 5321 12022 sw
tri 5422 11885 5559 12022 ne
rect 5559 11885 5734 12022
tri 5734 11885 5871 12022 sw
tri 5972 11885 6109 12022 ne
rect 6109 11885 6284 12022
tri 6284 11885 6421 12022 sw
tri 6522 11885 6659 12022 ne
rect 6659 11885 6834 12022
tri 6834 11885 6971 12022 sw
tri 7072 11885 7209 12022 ne
rect 7209 11885 7384 12022
tri 7384 11885 7521 12022 sw
tri 7622 11885 7759 12022 ne
rect 7759 11885 7934 12022
tri 7934 11885 8071 12022 sw
tri 8172 11885 8309 12022 ne
rect 8309 11885 8484 12022
tri 8484 11885 8621 12022 sw
tri 8722 11885 8859 12022 ne
rect 8859 11885 9034 12022
tri 9034 11885 9171 12022 sw
tri 9272 11885 9409 12022 ne
rect 9409 11885 9584 12022
tri 9584 11885 9721 12022 sw
tri 9822 11885 9959 12022 ne
rect 9959 11885 10134 12022
tri 10134 11885 10271 12022 sw
tri 10372 11885 10509 12022 ne
rect 10509 11885 10684 12022
tri 10684 11885 10821 12022 sw
tri 10922 11885 11059 12022 ne
rect 11059 11885 11234 12022
tri 11234 11885 11371 12022 sw
tri 11472 11885 11609 12022 ne
rect 11609 11885 11784 12022
tri 11784 11885 11921 12022 sw
tri 12022 11885 12159 12022 ne
rect 12159 11885 12334 12022
tri 12334 11885 12471 12022 sw
tri 12572 11885 12709 12022 ne
rect 12709 11885 12884 12022
tri 12884 11885 13021 12022 sw
tri 13122 11885 13259 12022 ne
rect 13259 11885 13434 12022
tri 13434 11885 13571 12022 sw
tri 13672 11885 13809 12022 ne
rect 13809 11885 13984 12022
tri 13984 11885 14121 12022 sw
tri 14222 11885 14359 12022 ne
rect 14359 11885 14534 12022
tri 14534 11885 14671 12022 sw
tri 14772 11885 14909 12022 ne
rect 14909 11885 15084 12022
tri 15084 11885 15221 12022 sw
tri 15322 11885 15459 12022 ne
rect 15459 11885 15634 12022
tri 15634 11885 15771 12022 sw
tri 15872 11885 16009 12022 ne
rect 16009 11885 16184 12022
tri 16184 11885 16321 12022 sw
tri 16422 11885 16559 12022 ne
rect 16559 11885 16734 12022
tri 16734 11885 16871 12022 sw
tri 16972 11885 17109 12022 ne
rect 17109 11885 17284 12022
tri 17284 11885 17421 12022 sw
tri 17522 11885 17659 12022 ne
rect 17659 11885 17834 12022
tri 17834 11885 17971 12022 sw
tri 18072 11885 18209 12022 ne
rect 18209 11885 18384 12022
tri 18384 11885 18521 12022 sw
tri 18622 11885 18759 12022 ne
rect 18759 11885 18934 12022
tri 18934 11885 19071 12022 sw
tri 19172 11885 19309 12022 ne
rect 19309 11885 19484 12022
tri 19484 11885 19621 12022 sw
rect -2000 11867 215 11885
rect -2000 11078 -1000 11867
tri 77 11765 179 11867 ne
rect 179 11765 215 11867
rect 335 11765 371 11885
tri 179 11628 316 11765 ne
rect 316 11710 371 11765
tri 371 11710 546 11885 sw
tri 609 11765 729 11885 ne
rect 729 11765 765 11885
rect 885 11765 921 11885
rect 316 11628 546 11710
tri 546 11628 628 11710 sw
tri 729 11628 866 11765 ne
rect 866 11710 921 11765
tri 921 11710 1096 11885 sw
tri 1159 11765 1279 11885 ne
rect 1279 11765 1315 11885
rect 1435 11765 1471 11885
rect 866 11628 1096 11710
tri 1096 11628 1178 11710 sw
tri 1279 11628 1416 11765 ne
rect 1416 11710 1471 11765
tri 1471 11710 1646 11885 sw
tri 1709 11765 1829 11885 ne
rect 1829 11765 1865 11885
rect 1985 11765 2021 11885
rect 1416 11628 1646 11710
tri 1646 11628 1728 11710 sw
tri 1829 11628 1966 11765 ne
rect 1966 11710 2021 11765
tri 2021 11710 2196 11885 sw
tri 2259 11765 2379 11885 ne
rect 2379 11765 2415 11885
rect 2535 11765 2571 11885
rect 1966 11628 2196 11710
tri 2196 11628 2278 11710 sw
tri 2379 11628 2516 11765 ne
rect 2516 11710 2571 11765
tri 2571 11710 2746 11885 sw
tri 2809 11765 2929 11885 ne
rect 2929 11765 2965 11885
rect 3085 11765 3121 11885
rect 2516 11628 2746 11710
tri 2746 11628 2828 11710 sw
tri 2929 11628 3066 11765 ne
rect 3066 11710 3121 11765
tri 3121 11710 3296 11885 sw
tri 3359 11765 3479 11885 ne
rect 3479 11765 3515 11885
rect 3635 11765 3671 11885
rect 3066 11628 3296 11710
tri 3296 11628 3378 11710 sw
tri 3479 11628 3616 11765 ne
rect 3616 11710 3671 11765
tri 3671 11710 3846 11885 sw
tri 3909 11765 4029 11885 ne
rect 4029 11765 4065 11885
rect 4185 11765 4221 11885
rect 3616 11628 3846 11710
tri 3846 11628 3928 11710 sw
tri 4029 11628 4166 11765 ne
rect 4166 11710 4221 11765
tri 4221 11710 4396 11885 sw
tri 4459 11765 4579 11885 ne
rect 4579 11765 4615 11885
rect 4735 11765 4771 11885
rect 4166 11628 4396 11710
tri 4396 11628 4478 11710 sw
tri 4579 11628 4716 11765 ne
rect 4716 11710 4771 11765
tri 4771 11710 4946 11885 sw
tri 5009 11765 5129 11885 ne
rect 5129 11765 5165 11885
rect 5285 11765 5321 11885
rect 4716 11628 4946 11710
tri 4946 11628 5028 11710 sw
tri 5129 11628 5266 11765 ne
rect 5266 11710 5321 11765
tri 5321 11710 5496 11885 sw
tri 5559 11765 5679 11885 ne
rect 5679 11765 5715 11885
rect 5835 11765 5871 11885
rect 5266 11628 5496 11710
tri 5496 11628 5578 11710 sw
tri 5679 11628 5816 11765 ne
rect 5816 11710 5871 11765
tri 5871 11710 6046 11885 sw
tri 6109 11765 6229 11885 ne
rect 6229 11765 6265 11885
rect 6385 11765 6421 11885
rect 5816 11628 6046 11710
tri 6046 11628 6128 11710 sw
tri 6229 11628 6366 11765 ne
rect 6366 11710 6421 11765
tri 6421 11710 6596 11885 sw
tri 6659 11765 6779 11885 ne
rect 6779 11765 6815 11885
rect 6935 11765 6971 11885
rect 6366 11628 6596 11710
tri 6596 11628 6678 11710 sw
tri 6779 11628 6916 11765 ne
rect 6916 11710 6971 11765
tri 6971 11710 7146 11885 sw
tri 7209 11765 7329 11885 ne
rect 7329 11765 7365 11885
rect 7485 11765 7521 11885
rect 6916 11628 7146 11710
tri 7146 11628 7228 11710 sw
tri 7329 11628 7466 11765 ne
rect 7466 11710 7521 11765
tri 7521 11710 7696 11885 sw
tri 7759 11765 7879 11885 ne
rect 7879 11765 7915 11885
rect 8035 11765 8071 11885
rect 7466 11628 7696 11710
tri 7696 11628 7778 11710 sw
tri 7879 11628 8016 11765 ne
rect 8016 11710 8071 11765
tri 8071 11710 8246 11885 sw
tri 8309 11765 8429 11885 ne
rect 8429 11765 8465 11885
rect 8585 11765 8621 11885
rect 8016 11628 8246 11710
tri 8246 11628 8328 11710 sw
tri 8429 11628 8566 11765 ne
rect 8566 11710 8621 11765
tri 8621 11710 8796 11885 sw
tri 8859 11765 8979 11885 ne
rect 8979 11765 9015 11885
rect 9135 11765 9171 11885
rect 8566 11628 8796 11710
tri 8796 11628 8878 11710 sw
tri 8979 11628 9116 11765 ne
rect 9116 11710 9171 11765
tri 9171 11710 9346 11885 sw
tri 9409 11765 9529 11885 ne
rect 9529 11765 9565 11885
rect 9685 11765 9721 11885
rect 9116 11628 9346 11710
tri 9346 11628 9428 11710 sw
tri 9529 11628 9666 11765 ne
rect 9666 11710 9721 11765
tri 9721 11710 9896 11885 sw
tri 9959 11765 10079 11885 ne
rect 10079 11765 10115 11885
rect 10235 11765 10271 11885
rect 9666 11628 9896 11710
tri 9896 11628 9978 11710 sw
tri 10079 11628 10216 11765 ne
rect 10216 11710 10271 11765
tri 10271 11710 10446 11885 sw
tri 10509 11765 10629 11885 ne
rect 10629 11765 10665 11885
rect 10785 11765 10821 11885
rect 10216 11628 10446 11710
tri 10446 11628 10528 11710 sw
tri 10629 11628 10766 11765 ne
rect 10766 11710 10821 11765
tri 10821 11710 10996 11885 sw
tri 11059 11765 11179 11885 ne
rect 11179 11765 11215 11885
rect 11335 11765 11371 11885
rect 10766 11628 10996 11710
tri 10996 11628 11078 11710 sw
tri 11179 11628 11316 11765 ne
rect 11316 11710 11371 11765
tri 11371 11710 11546 11885 sw
tri 11609 11765 11729 11885 ne
rect 11729 11765 11765 11885
rect 11885 11765 11921 11885
rect 11316 11628 11546 11710
tri 11546 11628 11628 11710 sw
tri 11729 11628 11866 11765 ne
rect 11866 11710 11921 11765
tri 11921 11710 12096 11885 sw
tri 12159 11765 12279 11885 ne
rect 12279 11765 12315 11885
rect 12435 11765 12471 11885
rect 11866 11628 12096 11710
tri 12096 11628 12178 11710 sw
tri 12279 11628 12416 11765 ne
rect 12416 11710 12471 11765
tri 12471 11710 12646 11885 sw
tri 12709 11765 12829 11885 ne
rect 12829 11765 12865 11885
rect 12985 11765 13021 11885
rect 12416 11628 12646 11710
tri 12646 11628 12728 11710 sw
tri 12829 11628 12966 11765 ne
rect 12966 11710 13021 11765
tri 13021 11710 13196 11885 sw
tri 13259 11765 13379 11885 ne
rect 13379 11765 13415 11885
rect 13535 11765 13571 11885
rect 12966 11628 13196 11710
tri 13196 11628 13278 11710 sw
tri 13379 11628 13516 11765 ne
rect 13516 11710 13571 11765
tri 13571 11710 13746 11885 sw
tri 13809 11765 13929 11885 ne
rect 13929 11765 13965 11885
rect 14085 11765 14121 11885
rect 13516 11628 13746 11710
tri 13746 11628 13828 11710 sw
tri 13929 11628 14066 11765 ne
rect 14066 11710 14121 11765
tri 14121 11710 14296 11885 sw
tri 14359 11765 14479 11885 ne
rect 14479 11765 14515 11885
rect 14635 11765 14671 11885
rect 14066 11628 14296 11710
tri 14296 11628 14378 11710 sw
tri 14479 11628 14616 11765 ne
rect 14616 11710 14671 11765
tri 14671 11710 14846 11885 sw
tri 14909 11765 15029 11885 ne
rect 15029 11765 15065 11885
rect 15185 11765 15221 11885
rect 14616 11628 14846 11710
tri 14846 11628 14928 11710 sw
tri 15029 11628 15166 11765 ne
rect 15166 11710 15221 11765
tri 15221 11710 15396 11885 sw
tri 15459 11765 15579 11885 ne
rect 15579 11765 15615 11885
rect 15735 11765 15771 11885
rect 15166 11628 15396 11710
tri 15396 11628 15478 11710 sw
tri 15579 11628 15716 11765 ne
rect 15716 11710 15771 11765
tri 15771 11710 15946 11885 sw
tri 16009 11765 16129 11885 ne
rect 16129 11765 16165 11885
rect 16285 11765 16321 11885
rect 15716 11628 15946 11710
tri 15946 11628 16028 11710 sw
tri 16129 11628 16266 11765 ne
rect 16266 11710 16321 11765
tri 16321 11710 16496 11885 sw
tri 16559 11765 16679 11885 ne
rect 16679 11765 16715 11885
rect 16835 11765 16871 11885
rect 16266 11628 16496 11710
tri 16496 11628 16578 11710 sw
tri 16679 11628 16816 11765 ne
rect 16816 11710 16871 11765
tri 16871 11710 17046 11885 sw
tri 17109 11765 17229 11885 ne
rect 17229 11765 17265 11885
rect 17385 11765 17421 11885
rect 16816 11628 17046 11710
tri 17046 11628 17128 11710 sw
tri 17229 11628 17366 11765 ne
rect 17366 11710 17421 11765
tri 17421 11710 17596 11885 sw
tri 17659 11765 17779 11885 ne
rect 17779 11765 17815 11885
rect 17935 11765 17971 11885
rect 17366 11628 17596 11710
tri 17596 11628 17678 11710 sw
tri 17779 11628 17916 11765 ne
rect 17916 11710 17971 11765
tri 17971 11710 18146 11885 sw
tri 18209 11765 18329 11885 ne
rect 18329 11765 18365 11885
rect 18485 11765 18521 11885
rect 17916 11628 18146 11710
tri 18146 11628 18228 11710 sw
tri 18329 11628 18466 11765 ne
rect 18466 11710 18521 11765
tri 18521 11710 18696 11885 sw
tri 18759 11765 18879 11885 ne
rect 18879 11765 18915 11885
rect 19035 11765 19071 11885
rect 18466 11628 18696 11710
tri 18696 11628 18778 11710 sw
tri 18879 11628 19016 11765 ne
rect 19016 11710 19071 11765
tri 19071 11710 19246 11885 sw
tri 19309 11765 19429 11885 ne
rect 19429 11765 19465 11885
rect 19585 11783 19621 11885
tri 19621 11783 19723 11885 sw
rect 20800 11783 21800 12572
rect 19585 11765 21800 11783
rect 19016 11628 19246 11710
tri 19246 11628 19328 11710 sw
tri 19429 11628 19566 11765 ne
rect 19566 11628 21800 11765
rect -500 11472 78 11628
tri 78 11472 234 11628 sw
tri 316 11472 472 11628 ne
rect 472 11472 628 11628
tri 628 11472 784 11628 sw
tri 866 11472 1022 11628 ne
rect 1022 11472 1178 11628
tri 1178 11472 1334 11628 sw
tri 1416 11472 1572 11628 ne
rect 1572 11472 1728 11628
tri 1728 11472 1884 11628 sw
tri 1966 11472 2122 11628 ne
rect 2122 11472 2278 11628
tri 2278 11472 2434 11628 sw
tri 2516 11472 2672 11628 ne
rect 2672 11472 2828 11628
tri 2828 11472 2984 11628 sw
tri 3066 11472 3222 11628 ne
rect 3222 11472 3378 11628
tri 3378 11472 3534 11628 sw
tri 3616 11472 3772 11628 ne
rect 3772 11472 3928 11628
tri 3928 11472 4084 11628 sw
tri 4166 11472 4322 11628 ne
rect 4322 11472 4478 11628
tri 4478 11472 4634 11628 sw
tri 4716 11472 4872 11628 ne
rect 4872 11472 5028 11628
tri 5028 11472 5184 11628 sw
tri 5266 11472 5422 11628 ne
rect 5422 11472 5578 11628
tri 5578 11472 5734 11628 sw
tri 5816 11472 5972 11628 ne
rect 5972 11472 6128 11628
tri 6128 11472 6284 11628 sw
tri 6366 11472 6522 11628 ne
rect 6522 11472 6678 11628
tri 6678 11472 6834 11628 sw
tri 6916 11472 7072 11628 ne
rect 7072 11472 7228 11628
tri 7228 11472 7384 11628 sw
tri 7466 11472 7622 11628 ne
rect 7622 11472 7778 11628
tri 7778 11472 7934 11628 sw
tri 8016 11472 8172 11628 ne
rect 8172 11472 8328 11628
tri 8328 11472 8484 11628 sw
tri 8566 11472 8722 11628 ne
rect 8722 11472 8878 11628
tri 8878 11472 9034 11628 sw
tri 9116 11472 9272 11628 ne
rect 9272 11472 9428 11628
tri 9428 11472 9584 11628 sw
tri 9666 11472 9822 11628 ne
rect 9822 11472 9978 11628
tri 9978 11472 10134 11628 sw
tri 10216 11472 10372 11628 ne
rect 10372 11472 10528 11628
tri 10528 11472 10684 11628 sw
tri 10766 11472 10922 11628 ne
rect 10922 11472 11078 11628
tri 11078 11472 11234 11628 sw
tri 11316 11472 11472 11628 ne
rect 11472 11472 11628 11628
tri 11628 11472 11784 11628 sw
tri 11866 11472 12022 11628 ne
rect 12022 11472 12178 11628
tri 12178 11472 12334 11628 sw
tri 12416 11472 12572 11628 ne
rect 12572 11472 12728 11628
tri 12728 11472 12884 11628 sw
tri 12966 11472 13122 11628 ne
rect 13122 11472 13278 11628
tri 13278 11472 13434 11628 sw
tri 13516 11472 13672 11628 ne
rect 13672 11472 13828 11628
tri 13828 11472 13984 11628 sw
tri 14066 11472 14222 11628 ne
rect 14222 11472 14378 11628
tri 14378 11472 14534 11628 sw
tri 14616 11472 14772 11628 ne
rect 14772 11472 14928 11628
tri 14928 11472 15084 11628 sw
tri 15166 11472 15322 11628 ne
rect 15322 11472 15478 11628
tri 15478 11472 15634 11628 sw
tri 15716 11472 15872 11628 ne
rect 15872 11472 16028 11628
tri 16028 11472 16184 11628 sw
tri 16266 11472 16422 11628 ne
rect 16422 11472 16578 11628
tri 16578 11472 16734 11628 sw
tri 16816 11472 16972 11628 ne
rect 16972 11472 17128 11628
tri 17128 11472 17284 11628 sw
tri 17366 11472 17522 11628 ne
rect 17522 11472 17678 11628
tri 17678 11472 17834 11628 sw
tri 17916 11472 18072 11628 ne
rect 18072 11472 18228 11628
tri 18228 11472 18384 11628 sw
tri 18466 11472 18622 11628 ne
rect 18622 11472 18778 11628
tri 18778 11472 18934 11628 sw
tri 19016 11472 19172 11628 ne
rect 19172 11472 19328 11628
tri 19328 11472 19484 11628 sw
tri 19566 11472 19722 11628 ne
rect 19722 11472 21800 11628
rect -500 11335 234 11472
tri 234 11335 371 11472 sw
tri 472 11335 609 11472 ne
rect 609 11335 784 11472
tri 784 11335 921 11472 sw
tri 1022 11335 1159 11472 ne
rect 1159 11335 1334 11472
tri 1334 11335 1471 11472 sw
tri 1572 11335 1709 11472 ne
rect 1709 11335 1884 11472
tri 1884 11335 2021 11472 sw
tri 2122 11335 2259 11472 ne
rect 2259 11335 2434 11472
tri 2434 11335 2571 11472 sw
tri 2672 11335 2809 11472 ne
rect 2809 11335 2984 11472
tri 2984 11335 3121 11472 sw
tri 3222 11335 3359 11472 ne
rect 3359 11335 3534 11472
tri 3534 11335 3671 11472 sw
tri 3772 11335 3909 11472 ne
rect 3909 11335 4084 11472
tri 4084 11335 4221 11472 sw
tri 4322 11335 4459 11472 ne
rect 4459 11335 4634 11472
tri 4634 11335 4771 11472 sw
tri 4872 11335 5009 11472 ne
rect 5009 11335 5184 11472
tri 5184 11335 5321 11472 sw
tri 5422 11335 5559 11472 ne
rect 5559 11335 5734 11472
tri 5734 11335 5871 11472 sw
tri 5972 11335 6109 11472 ne
rect 6109 11335 6284 11472
tri 6284 11335 6421 11472 sw
tri 6522 11335 6659 11472 ne
rect 6659 11335 6834 11472
tri 6834 11335 6971 11472 sw
tri 7072 11335 7209 11472 ne
rect 7209 11335 7384 11472
tri 7384 11335 7521 11472 sw
tri 7622 11335 7759 11472 ne
rect 7759 11335 7934 11472
tri 7934 11335 8071 11472 sw
tri 8172 11335 8309 11472 ne
rect 8309 11335 8484 11472
tri 8484 11335 8621 11472 sw
tri 8722 11335 8859 11472 ne
rect 8859 11335 9034 11472
tri 9034 11335 9171 11472 sw
tri 9272 11335 9409 11472 ne
rect 9409 11335 9584 11472
tri 9584 11335 9721 11472 sw
tri 9822 11335 9959 11472 ne
rect 9959 11335 10134 11472
tri 10134 11335 10271 11472 sw
tri 10372 11335 10509 11472 ne
rect 10509 11335 10684 11472
tri 10684 11335 10821 11472 sw
tri 10922 11335 11059 11472 ne
rect 11059 11335 11234 11472
tri 11234 11335 11371 11472 sw
tri 11472 11335 11609 11472 ne
rect 11609 11335 11784 11472
tri 11784 11335 11921 11472 sw
tri 12022 11335 12159 11472 ne
rect 12159 11335 12334 11472
tri 12334 11335 12471 11472 sw
tri 12572 11335 12709 11472 ne
rect 12709 11335 12884 11472
tri 12884 11335 13021 11472 sw
tri 13122 11335 13259 11472 ne
rect 13259 11335 13434 11472
tri 13434 11335 13571 11472 sw
tri 13672 11335 13809 11472 ne
rect 13809 11335 13984 11472
tri 13984 11335 14121 11472 sw
tri 14222 11335 14359 11472 ne
rect 14359 11335 14534 11472
tri 14534 11335 14671 11472 sw
tri 14772 11335 14909 11472 ne
rect 14909 11335 15084 11472
tri 15084 11335 15221 11472 sw
tri 15322 11335 15459 11472 ne
rect 15459 11335 15634 11472
tri 15634 11335 15771 11472 sw
tri 15872 11335 16009 11472 ne
rect 16009 11335 16184 11472
tri 16184 11335 16321 11472 sw
tri 16422 11335 16559 11472 ne
rect 16559 11335 16734 11472
tri 16734 11335 16871 11472 sw
tri 16972 11335 17109 11472 ne
rect 17109 11335 17284 11472
tri 17284 11335 17421 11472 sw
tri 17522 11335 17659 11472 ne
rect 17659 11335 17834 11472
tri 17834 11335 17971 11472 sw
tri 18072 11335 18209 11472 ne
rect 18209 11335 18384 11472
tri 18384 11335 18521 11472 sw
tri 18622 11335 18759 11472 ne
rect 18759 11335 18934 11472
tri 18934 11335 19071 11472 sw
tri 19172 11335 19309 11472 ne
rect 19309 11335 19484 11472
tri 19484 11335 19621 11472 sw
rect -500 11317 215 11335
tri 77 11215 179 11317 ne
rect 179 11215 215 11317
rect 335 11215 371 11335
tri 179 11078 316 11215 ne
rect 316 11160 371 11215
tri 371 11160 546 11335 sw
tri 609 11215 729 11335 ne
rect 729 11215 765 11335
rect 885 11215 921 11335
rect 316 11078 546 11160
tri 546 11078 628 11160 sw
tri 729 11078 866 11215 ne
rect 866 11160 921 11215
tri 921 11160 1096 11335 sw
tri 1159 11215 1279 11335 ne
rect 1279 11215 1315 11335
rect 1435 11215 1471 11335
rect 866 11078 1096 11160
tri 1096 11078 1178 11160 sw
tri 1279 11078 1416 11215 ne
rect 1416 11160 1471 11215
tri 1471 11160 1646 11335 sw
tri 1709 11215 1829 11335 ne
rect 1829 11215 1865 11335
rect 1985 11215 2021 11335
rect 1416 11078 1646 11160
tri 1646 11078 1728 11160 sw
tri 1829 11078 1966 11215 ne
rect 1966 11160 2021 11215
tri 2021 11160 2196 11335 sw
tri 2259 11215 2379 11335 ne
rect 2379 11215 2415 11335
rect 2535 11215 2571 11335
rect 1966 11078 2196 11160
tri 2196 11078 2278 11160 sw
tri 2379 11078 2516 11215 ne
rect 2516 11160 2571 11215
tri 2571 11160 2746 11335 sw
tri 2809 11215 2929 11335 ne
rect 2929 11215 2965 11335
rect 3085 11215 3121 11335
rect 2516 11078 2746 11160
tri 2746 11078 2828 11160 sw
tri 2929 11078 3066 11215 ne
rect 3066 11160 3121 11215
tri 3121 11160 3296 11335 sw
tri 3359 11215 3479 11335 ne
rect 3479 11215 3515 11335
rect 3635 11215 3671 11335
rect 3066 11078 3296 11160
tri 3296 11078 3378 11160 sw
tri 3479 11078 3616 11215 ne
rect 3616 11160 3671 11215
tri 3671 11160 3846 11335 sw
tri 3909 11215 4029 11335 ne
rect 4029 11215 4065 11335
rect 4185 11215 4221 11335
rect 3616 11078 3846 11160
tri 3846 11078 3928 11160 sw
tri 4029 11078 4166 11215 ne
rect 4166 11160 4221 11215
tri 4221 11160 4396 11335 sw
tri 4459 11215 4579 11335 ne
rect 4579 11215 4615 11335
rect 4735 11215 4771 11335
rect 4166 11078 4396 11160
tri 4396 11078 4478 11160 sw
tri 4579 11078 4716 11215 ne
rect 4716 11160 4771 11215
tri 4771 11160 4946 11335 sw
tri 5009 11215 5129 11335 ne
rect 5129 11215 5165 11335
rect 5285 11215 5321 11335
rect 4716 11078 4946 11160
tri 4946 11078 5028 11160 sw
tri 5129 11078 5266 11215 ne
rect 5266 11160 5321 11215
tri 5321 11160 5496 11335 sw
tri 5559 11215 5679 11335 ne
rect 5679 11215 5715 11335
rect 5835 11215 5871 11335
rect 5266 11078 5496 11160
tri 5496 11078 5578 11160 sw
tri 5679 11078 5816 11215 ne
rect 5816 11160 5871 11215
tri 5871 11160 6046 11335 sw
tri 6109 11215 6229 11335 ne
rect 6229 11215 6265 11335
rect 6385 11215 6421 11335
rect 5816 11078 6046 11160
tri 6046 11078 6128 11160 sw
tri 6229 11078 6366 11215 ne
rect 6366 11160 6421 11215
tri 6421 11160 6596 11335 sw
tri 6659 11215 6779 11335 ne
rect 6779 11215 6815 11335
rect 6935 11215 6971 11335
rect 6366 11078 6596 11160
tri 6596 11078 6678 11160 sw
tri 6779 11078 6916 11215 ne
rect 6916 11160 6971 11215
tri 6971 11160 7146 11335 sw
tri 7209 11215 7329 11335 ne
rect 7329 11215 7365 11335
rect 7485 11215 7521 11335
rect 6916 11078 7146 11160
tri 7146 11078 7228 11160 sw
tri 7329 11078 7466 11215 ne
rect 7466 11160 7521 11215
tri 7521 11160 7696 11335 sw
tri 7759 11215 7879 11335 ne
rect 7879 11215 7915 11335
rect 8035 11215 8071 11335
rect 7466 11078 7696 11160
tri 7696 11078 7778 11160 sw
tri 7879 11078 8016 11215 ne
rect 8016 11160 8071 11215
tri 8071 11160 8246 11335 sw
tri 8309 11215 8429 11335 ne
rect 8429 11215 8465 11335
rect 8585 11215 8621 11335
rect 8016 11078 8246 11160
tri 8246 11078 8328 11160 sw
tri 8429 11078 8566 11215 ne
rect 8566 11160 8621 11215
tri 8621 11160 8796 11335 sw
tri 8859 11215 8979 11335 ne
rect 8979 11215 9015 11335
rect 9135 11215 9171 11335
rect 8566 11078 8796 11160
tri 8796 11078 8878 11160 sw
tri 8979 11078 9116 11215 ne
rect 9116 11160 9171 11215
tri 9171 11160 9346 11335 sw
tri 9409 11215 9529 11335 ne
rect 9529 11215 9565 11335
rect 9685 11215 9721 11335
rect 9116 11078 9346 11160
tri 9346 11078 9428 11160 sw
tri 9529 11078 9666 11215 ne
rect 9666 11160 9721 11215
tri 9721 11160 9896 11335 sw
tri 9959 11215 10079 11335 ne
rect 10079 11215 10115 11335
rect 10235 11215 10271 11335
rect 9666 11078 9896 11160
tri 9896 11078 9978 11160 sw
tri 10079 11078 10216 11215 ne
rect 10216 11160 10271 11215
tri 10271 11160 10446 11335 sw
tri 10509 11215 10629 11335 ne
rect 10629 11215 10665 11335
rect 10785 11215 10821 11335
rect 10216 11078 10446 11160
tri 10446 11078 10528 11160 sw
tri 10629 11078 10766 11215 ne
rect 10766 11160 10821 11215
tri 10821 11160 10996 11335 sw
tri 11059 11215 11179 11335 ne
rect 11179 11215 11215 11335
rect 11335 11215 11371 11335
rect 10766 11078 10996 11160
tri 10996 11078 11078 11160 sw
tri 11179 11078 11316 11215 ne
rect 11316 11160 11371 11215
tri 11371 11160 11546 11335 sw
tri 11609 11215 11729 11335 ne
rect 11729 11215 11765 11335
rect 11885 11215 11921 11335
rect 11316 11078 11546 11160
tri 11546 11078 11628 11160 sw
tri 11729 11078 11866 11215 ne
rect 11866 11160 11921 11215
tri 11921 11160 12096 11335 sw
tri 12159 11215 12279 11335 ne
rect 12279 11215 12315 11335
rect 12435 11215 12471 11335
rect 11866 11078 12096 11160
tri 12096 11078 12178 11160 sw
tri 12279 11078 12416 11215 ne
rect 12416 11160 12471 11215
tri 12471 11160 12646 11335 sw
tri 12709 11215 12829 11335 ne
rect 12829 11215 12865 11335
rect 12985 11215 13021 11335
rect 12416 11078 12646 11160
tri 12646 11078 12728 11160 sw
tri 12829 11078 12966 11215 ne
rect 12966 11160 13021 11215
tri 13021 11160 13196 11335 sw
tri 13259 11215 13379 11335 ne
rect 13379 11215 13415 11335
rect 13535 11215 13571 11335
rect 12966 11078 13196 11160
tri 13196 11078 13278 11160 sw
tri 13379 11078 13516 11215 ne
rect 13516 11160 13571 11215
tri 13571 11160 13746 11335 sw
tri 13809 11215 13929 11335 ne
rect 13929 11215 13965 11335
rect 14085 11215 14121 11335
rect 13516 11078 13746 11160
tri 13746 11078 13828 11160 sw
tri 13929 11078 14066 11215 ne
rect 14066 11160 14121 11215
tri 14121 11160 14296 11335 sw
tri 14359 11215 14479 11335 ne
rect 14479 11215 14515 11335
rect 14635 11215 14671 11335
rect 14066 11078 14296 11160
tri 14296 11078 14378 11160 sw
tri 14479 11078 14616 11215 ne
rect 14616 11160 14671 11215
tri 14671 11160 14846 11335 sw
tri 14909 11215 15029 11335 ne
rect 15029 11215 15065 11335
rect 15185 11215 15221 11335
rect 14616 11078 14846 11160
tri 14846 11078 14928 11160 sw
tri 15029 11078 15166 11215 ne
rect 15166 11160 15221 11215
tri 15221 11160 15396 11335 sw
tri 15459 11215 15579 11335 ne
rect 15579 11215 15615 11335
rect 15735 11215 15771 11335
rect 15166 11078 15396 11160
tri 15396 11078 15478 11160 sw
tri 15579 11078 15716 11215 ne
rect 15716 11160 15771 11215
tri 15771 11160 15946 11335 sw
tri 16009 11215 16129 11335 ne
rect 16129 11215 16165 11335
rect 16285 11215 16321 11335
rect 15716 11078 15946 11160
tri 15946 11078 16028 11160 sw
tri 16129 11078 16266 11215 ne
rect 16266 11160 16321 11215
tri 16321 11160 16496 11335 sw
tri 16559 11215 16679 11335 ne
rect 16679 11215 16715 11335
rect 16835 11215 16871 11335
rect 16266 11078 16496 11160
tri 16496 11078 16578 11160 sw
tri 16679 11078 16816 11215 ne
rect 16816 11160 16871 11215
tri 16871 11160 17046 11335 sw
tri 17109 11215 17229 11335 ne
rect 17229 11215 17265 11335
rect 17385 11215 17421 11335
rect 16816 11078 17046 11160
tri 17046 11078 17128 11160 sw
tri 17229 11078 17366 11215 ne
rect 17366 11160 17421 11215
tri 17421 11160 17596 11335 sw
tri 17659 11215 17779 11335 ne
rect 17779 11215 17815 11335
rect 17935 11215 17971 11335
rect 17366 11078 17596 11160
tri 17596 11078 17678 11160 sw
tri 17779 11078 17916 11215 ne
rect 17916 11160 17971 11215
tri 17971 11160 18146 11335 sw
tri 18209 11215 18329 11335 ne
rect 18329 11215 18365 11335
rect 18485 11215 18521 11335
rect 17916 11078 18146 11160
tri 18146 11078 18228 11160 sw
tri 18329 11078 18466 11215 ne
rect 18466 11160 18521 11215
tri 18521 11160 18696 11335 sw
tri 18759 11215 18879 11335 ne
rect 18879 11215 18915 11335
rect 19035 11215 19071 11335
rect 18466 11078 18696 11160
tri 18696 11078 18778 11160 sw
tri 18879 11078 19016 11215 ne
rect 19016 11160 19071 11215
tri 19071 11160 19246 11335 sw
tri 19309 11215 19429 11335 ne
rect 19429 11215 19465 11335
rect 19585 11233 19621 11335
tri 19621 11233 19723 11335 sw
rect 19585 11215 20300 11233
rect 19016 11078 19246 11160
tri 19246 11078 19328 11160 sw
tri 19429 11078 19566 11215 ne
rect 19566 11078 20300 11215
rect -2000 10922 78 11078
tri 78 10922 234 11078 sw
tri 316 10922 472 11078 ne
rect 472 10922 628 11078
tri 628 10922 784 11078 sw
tri 866 10922 1022 11078 ne
rect 1022 10922 1178 11078
tri 1178 10922 1334 11078 sw
tri 1416 10922 1572 11078 ne
rect 1572 10922 1728 11078
tri 1728 10922 1884 11078 sw
tri 1966 10922 2122 11078 ne
rect 2122 10922 2278 11078
tri 2278 10922 2434 11078 sw
tri 2516 10922 2672 11078 ne
rect 2672 10922 2828 11078
tri 2828 10922 2984 11078 sw
tri 3066 10922 3222 11078 ne
rect 3222 10922 3378 11078
tri 3378 10922 3534 11078 sw
tri 3616 10922 3772 11078 ne
rect 3772 10922 3928 11078
tri 3928 10922 4084 11078 sw
tri 4166 10922 4322 11078 ne
rect 4322 10922 4478 11078
tri 4478 10922 4634 11078 sw
tri 4716 10922 4872 11078 ne
rect 4872 10922 5028 11078
tri 5028 10922 5184 11078 sw
tri 5266 10922 5422 11078 ne
rect 5422 10922 5578 11078
tri 5578 10922 5734 11078 sw
tri 5816 10922 5972 11078 ne
rect 5972 10922 6128 11078
tri 6128 10922 6284 11078 sw
tri 6366 10922 6522 11078 ne
rect 6522 10922 6678 11078
tri 6678 10922 6834 11078 sw
tri 6916 10922 7072 11078 ne
rect 7072 10922 7228 11078
tri 7228 10922 7384 11078 sw
tri 7466 10922 7622 11078 ne
rect 7622 10922 7778 11078
tri 7778 10922 7934 11078 sw
tri 8016 10922 8172 11078 ne
rect 8172 10922 8328 11078
tri 8328 10922 8484 11078 sw
tri 8566 10922 8722 11078 ne
rect 8722 10922 8878 11078
tri 8878 10922 9034 11078 sw
tri 9116 10922 9272 11078 ne
rect 9272 10922 9428 11078
tri 9428 10922 9584 11078 sw
tri 9666 10922 9822 11078 ne
rect 9822 10922 9978 11078
tri 9978 10922 10134 11078 sw
tri 10216 10922 10372 11078 ne
rect 10372 10922 10528 11078
tri 10528 10922 10684 11078 sw
tri 10766 10922 10922 11078 ne
rect 10922 10922 11078 11078
tri 11078 10922 11234 11078 sw
tri 11316 10922 11472 11078 ne
rect 11472 10922 11628 11078
tri 11628 10922 11784 11078 sw
tri 11866 10922 12022 11078 ne
rect 12022 10922 12178 11078
tri 12178 10922 12334 11078 sw
tri 12416 10922 12572 11078 ne
rect 12572 10922 12728 11078
tri 12728 10922 12884 11078 sw
tri 12966 10922 13122 11078 ne
rect 13122 10922 13278 11078
tri 13278 10922 13434 11078 sw
tri 13516 10922 13672 11078 ne
rect 13672 10922 13828 11078
tri 13828 10922 13984 11078 sw
tri 14066 10922 14222 11078 ne
rect 14222 10922 14378 11078
tri 14378 10922 14534 11078 sw
tri 14616 10922 14772 11078 ne
rect 14772 10922 14928 11078
tri 14928 10922 15084 11078 sw
tri 15166 10922 15322 11078 ne
rect 15322 10922 15478 11078
tri 15478 10922 15634 11078 sw
tri 15716 10922 15872 11078 ne
rect 15872 10922 16028 11078
tri 16028 10922 16184 11078 sw
tri 16266 10922 16422 11078 ne
rect 16422 10922 16578 11078
tri 16578 10922 16734 11078 sw
tri 16816 10922 16972 11078 ne
rect 16972 10922 17128 11078
tri 17128 10922 17284 11078 sw
tri 17366 10922 17522 11078 ne
rect 17522 10922 17678 11078
tri 17678 10922 17834 11078 sw
tri 17916 10922 18072 11078 ne
rect 18072 10922 18228 11078
tri 18228 10922 18384 11078 sw
tri 18466 10922 18622 11078 ne
rect 18622 10922 18778 11078
tri 18778 10922 18934 11078 sw
tri 19016 10922 19172 11078 ne
rect 19172 10922 19328 11078
tri 19328 10922 19484 11078 sw
tri 19566 10922 19722 11078 ne
rect 19722 10922 20300 11078
rect -2000 10785 234 10922
tri 234 10785 371 10922 sw
tri 472 10785 609 10922 ne
rect 609 10785 784 10922
tri 784 10785 921 10922 sw
tri 1022 10785 1159 10922 ne
rect 1159 10785 1334 10922
tri 1334 10785 1471 10922 sw
tri 1572 10785 1709 10922 ne
rect 1709 10785 1884 10922
tri 1884 10785 2021 10922 sw
tri 2122 10785 2259 10922 ne
rect 2259 10785 2434 10922
tri 2434 10785 2571 10922 sw
tri 2672 10785 2809 10922 ne
rect 2809 10785 2984 10922
tri 2984 10785 3121 10922 sw
tri 3222 10785 3359 10922 ne
rect 3359 10785 3534 10922
tri 3534 10785 3671 10922 sw
tri 3772 10785 3909 10922 ne
rect 3909 10785 4084 10922
tri 4084 10785 4221 10922 sw
tri 4322 10785 4459 10922 ne
rect 4459 10785 4634 10922
tri 4634 10785 4771 10922 sw
tri 4872 10785 5009 10922 ne
rect 5009 10785 5184 10922
tri 5184 10785 5321 10922 sw
tri 5422 10785 5559 10922 ne
rect 5559 10785 5734 10922
tri 5734 10785 5871 10922 sw
tri 5972 10785 6109 10922 ne
rect 6109 10785 6284 10922
tri 6284 10785 6421 10922 sw
tri 6522 10785 6659 10922 ne
rect 6659 10785 6834 10922
tri 6834 10785 6971 10922 sw
tri 7072 10785 7209 10922 ne
rect 7209 10785 7384 10922
tri 7384 10785 7521 10922 sw
tri 7622 10785 7759 10922 ne
rect 7759 10785 7934 10922
tri 7934 10785 8071 10922 sw
tri 8172 10785 8309 10922 ne
rect 8309 10785 8484 10922
tri 8484 10785 8621 10922 sw
tri 8722 10785 8859 10922 ne
rect 8859 10785 9034 10922
tri 9034 10785 9171 10922 sw
tri 9272 10785 9409 10922 ne
rect 9409 10785 9584 10922
tri 9584 10785 9721 10922 sw
tri 9822 10785 9959 10922 ne
rect 9959 10785 10134 10922
tri 10134 10785 10271 10922 sw
tri 10372 10785 10509 10922 ne
rect 10509 10785 10684 10922
tri 10684 10785 10821 10922 sw
tri 10922 10785 11059 10922 ne
rect 11059 10785 11234 10922
tri 11234 10785 11371 10922 sw
tri 11472 10785 11609 10922 ne
rect 11609 10785 11784 10922
tri 11784 10785 11921 10922 sw
tri 12022 10785 12159 10922 ne
rect 12159 10785 12334 10922
tri 12334 10785 12471 10922 sw
tri 12572 10785 12709 10922 ne
rect 12709 10785 12884 10922
tri 12884 10785 13021 10922 sw
tri 13122 10785 13259 10922 ne
rect 13259 10785 13434 10922
tri 13434 10785 13571 10922 sw
tri 13672 10785 13809 10922 ne
rect 13809 10785 13984 10922
tri 13984 10785 14121 10922 sw
tri 14222 10785 14359 10922 ne
rect 14359 10785 14534 10922
tri 14534 10785 14671 10922 sw
tri 14772 10785 14909 10922 ne
rect 14909 10785 15084 10922
tri 15084 10785 15221 10922 sw
tri 15322 10785 15459 10922 ne
rect 15459 10785 15634 10922
tri 15634 10785 15771 10922 sw
tri 15872 10785 16009 10922 ne
rect 16009 10785 16184 10922
tri 16184 10785 16321 10922 sw
tri 16422 10785 16559 10922 ne
rect 16559 10785 16734 10922
tri 16734 10785 16871 10922 sw
tri 16972 10785 17109 10922 ne
rect 17109 10785 17284 10922
tri 17284 10785 17421 10922 sw
tri 17522 10785 17659 10922 ne
rect 17659 10785 17834 10922
tri 17834 10785 17971 10922 sw
tri 18072 10785 18209 10922 ne
rect 18209 10785 18384 10922
tri 18384 10785 18521 10922 sw
tri 18622 10785 18759 10922 ne
rect 18759 10785 18934 10922
tri 18934 10785 19071 10922 sw
tri 19172 10785 19309 10922 ne
rect 19309 10785 19484 10922
tri 19484 10785 19621 10922 sw
rect -2000 10767 215 10785
rect -2000 9978 -1000 10767
tri 77 10665 179 10767 ne
rect 179 10665 215 10767
rect 335 10665 371 10785
tri 179 10528 316 10665 ne
rect 316 10610 371 10665
tri 371 10610 546 10785 sw
tri 609 10665 729 10785 ne
rect 729 10665 765 10785
rect 885 10665 921 10785
rect 316 10528 546 10610
tri 546 10528 628 10610 sw
tri 729 10528 866 10665 ne
rect 866 10610 921 10665
tri 921 10610 1096 10785 sw
tri 1159 10665 1279 10785 ne
rect 1279 10665 1315 10785
rect 1435 10665 1471 10785
rect 866 10528 1096 10610
tri 1096 10528 1178 10610 sw
tri 1279 10528 1416 10665 ne
rect 1416 10610 1471 10665
tri 1471 10610 1646 10785 sw
tri 1709 10665 1829 10785 ne
rect 1829 10665 1865 10785
rect 1985 10665 2021 10785
rect 1416 10528 1646 10610
tri 1646 10528 1728 10610 sw
tri 1829 10528 1966 10665 ne
rect 1966 10610 2021 10665
tri 2021 10610 2196 10785 sw
tri 2259 10665 2379 10785 ne
rect 2379 10665 2415 10785
rect 2535 10665 2571 10785
rect 1966 10528 2196 10610
tri 2196 10528 2278 10610 sw
tri 2379 10528 2516 10665 ne
rect 2516 10610 2571 10665
tri 2571 10610 2746 10785 sw
tri 2809 10665 2929 10785 ne
rect 2929 10665 2965 10785
rect 3085 10665 3121 10785
rect 2516 10528 2746 10610
tri 2746 10528 2828 10610 sw
tri 2929 10528 3066 10665 ne
rect 3066 10610 3121 10665
tri 3121 10610 3296 10785 sw
tri 3359 10665 3479 10785 ne
rect 3479 10665 3515 10785
rect 3635 10665 3671 10785
rect 3066 10528 3296 10610
tri 3296 10528 3378 10610 sw
tri 3479 10528 3616 10665 ne
rect 3616 10610 3671 10665
tri 3671 10610 3846 10785 sw
tri 3909 10665 4029 10785 ne
rect 4029 10665 4065 10785
rect 4185 10665 4221 10785
rect 3616 10528 3846 10610
tri 3846 10528 3928 10610 sw
tri 4029 10528 4166 10665 ne
rect 4166 10610 4221 10665
tri 4221 10610 4396 10785 sw
tri 4459 10665 4579 10785 ne
rect 4579 10665 4615 10785
rect 4735 10665 4771 10785
rect 4166 10528 4396 10610
tri 4396 10528 4478 10610 sw
tri 4579 10528 4716 10665 ne
rect 4716 10610 4771 10665
tri 4771 10610 4946 10785 sw
tri 5009 10665 5129 10785 ne
rect 5129 10665 5165 10785
rect 5285 10665 5321 10785
rect 4716 10528 4946 10610
tri 4946 10528 5028 10610 sw
tri 5129 10528 5266 10665 ne
rect 5266 10610 5321 10665
tri 5321 10610 5496 10785 sw
tri 5559 10665 5679 10785 ne
rect 5679 10665 5715 10785
rect 5835 10665 5871 10785
rect 5266 10528 5496 10610
tri 5496 10528 5578 10610 sw
tri 5679 10528 5816 10665 ne
rect 5816 10610 5871 10665
tri 5871 10610 6046 10785 sw
tri 6109 10665 6229 10785 ne
rect 6229 10665 6265 10785
rect 6385 10665 6421 10785
rect 5816 10528 6046 10610
tri 6046 10528 6128 10610 sw
tri 6229 10528 6366 10665 ne
rect 6366 10610 6421 10665
tri 6421 10610 6596 10785 sw
tri 6659 10665 6779 10785 ne
rect 6779 10665 6815 10785
rect 6935 10665 6971 10785
rect 6366 10528 6596 10610
tri 6596 10528 6678 10610 sw
tri 6779 10528 6916 10665 ne
rect 6916 10610 6971 10665
tri 6971 10610 7146 10785 sw
tri 7209 10665 7329 10785 ne
rect 7329 10665 7365 10785
rect 7485 10665 7521 10785
rect 6916 10528 7146 10610
tri 7146 10528 7228 10610 sw
tri 7329 10528 7466 10665 ne
rect 7466 10610 7521 10665
tri 7521 10610 7696 10785 sw
tri 7759 10665 7879 10785 ne
rect 7879 10665 7915 10785
rect 8035 10665 8071 10785
rect 7466 10528 7696 10610
tri 7696 10528 7778 10610 sw
tri 7879 10528 8016 10665 ne
rect 8016 10610 8071 10665
tri 8071 10610 8246 10785 sw
tri 8309 10665 8429 10785 ne
rect 8429 10665 8465 10785
rect 8585 10665 8621 10785
rect 8016 10528 8246 10610
tri 8246 10528 8328 10610 sw
tri 8429 10528 8566 10665 ne
rect 8566 10610 8621 10665
tri 8621 10610 8796 10785 sw
tri 8859 10665 8979 10785 ne
rect 8979 10665 9015 10785
rect 9135 10665 9171 10785
rect 8566 10528 8796 10610
tri 8796 10528 8878 10610 sw
tri 8979 10528 9116 10665 ne
rect 9116 10610 9171 10665
tri 9171 10610 9346 10785 sw
tri 9409 10665 9529 10785 ne
rect 9529 10665 9565 10785
rect 9685 10665 9721 10785
rect 9116 10528 9346 10610
tri 9346 10528 9428 10610 sw
tri 9529 10528 9666 10665 ne
rect 9666 10610 9721 10665
tri 9721 10610 9896 10785 sw
tri 9959 10665 10079 10785 ne
rect 10079 10665 10115 10785
rect 10235 10665 10271 10785
rect 9666 10528 9896 10610
tri 9896 10528 9978 10610 sw
tri 10079 10528 10216 10665 ne
rect 10216 10610 10271 10665
tri 10271 10610 10446 10785 sw
tri 10509 10665 10629 10785 ne
rect 10629 10665 10665 10785
rect 10785 10665 10821 10785
rect 10216 10528 10446 10610
tri 10446 10528 10528 10610 sw
tri 10629 10528 10766 10665 ne
rect 10766 10610 10821 10665
tri 10821 10610 10996 10785 sw
tri 11059 10665 11179 10785 ne
rect 11179 10665 11215 10785
rect 11335 10665 11371 10785
rect 10766 10528 10996 10610
tri 10996 10528 11078 10610 sw
tri 11179 10528 11316 10665 ne
rect 11316 10610 11371 10665
tri 11371 10610 11546 10785 sw
tri 11609 10665 11729 10785 ne
rect 11729 10665 11765 10785
rect 11885 10665 11921 10785
rect 11316 10528 11546 10610
tri 11546 10528 11628 10610 sw
tri 11729 10528 11866 10665 ne
rect 11866 10610 11921 10665
tri 11921 10610 12096 10785 sw
tri 12159 10665 12279 10785 ne
rect 12279 10665 12315 10785
rect 12435 10665 12471 10785
rect 11866 10528 12096 10610
tri 12096 10528 12178 10610 sw
tri 12279 10528 12416 10665 ne
rect 12416 10610 12471 10665
tri 12471 10610 12646 10785 sw
tri 12709 10665 12829 10785 ne
rect 12829 10665 12865 10785
rect 12985 10665 13021 10785
rect 12416 10528 12646 10610
tri 12646 10528 12728 10610 sw
tri 12829 10528 12966 10665 ne
rect 12966 10610 13021 10665
tri 13021 10610 13196 10785 sw
tri 13259 10665 13379 10785 ne
rect 13379 10665 13415 10785
rect 13535 10665 13571 10785
rect 12966 10528 13196 10610
tri 13196 10528 13278 10610 sw
tri 13379 10528 13516 10665 ne
rect 13516 10610 13571 10665
tri 13571 10610 13746 10785 sw
tri 13809 10665 13929 10785 ne
rect 13929 10665 13965 10785
rect 14085 10665 14121 10785
rect 13516 10528 13746 10610
tri 13746 10528 13828 10610 sw
tri 13929 10528 14066 10665 ne
rect 14066 10610 14121 10665
tri 14121 10610 14296 10785 sw
tri 14359 10665 14479 10785 ne
rect 14479 10665 14515 10785
rect 14635 10665 14671 10785
rect 14066 10528 14296 10610
tri 14296 10528 14378 10610 sw
tri 14479 10528 14616 10665 ne
rect 14616 10610 14671 10665
tri 14671 10610 14846 10785 sw
tri 14909 10665 15029 10785 ne
rect 15029 10665 15065 10785
rect 15185 10665 15221 10785
rect 14616 10528 14846 10610
tri 14846 10528 14928 10610 sw
tri 15029 10528 15166 10665 ne
rect 15166 10610 15221 10665
tri 15221 10610 15396 10785 sw
tri 15459 10665 15579 10785 ne
rect 15579 10665 15615 10785
rect 15735 10665 15771 10785
rect 15166 10528 15396 10610
tri 15396 10528 15478 10610 sw
tri 15579 10528 15716 10665 ne
rect 15716 10610 15771 10665
tri 15771 10610 15946 10785 sw
tri 16009 10665 16129 10785 ne
rect 16129 10665 16165 10785
rect 16285 10665 16321 10785
rect 15716 10528 15946 10610
tri 15946 10528 16028 10610 sw
tri 16129 10528 16266 10665 ne
rect 16266 10610 16321 10665
tri 16321 10610 16496 10785 sw
tri 16559 10665 16679 10785 ne
rect 16679 10665 16715 10785
rect 16835 10665 16871 10785
rect 16266 10528 16496 10610
tri 16496 10528 16578 10610 sw
tri 16679 10528 16816 10665 ne
rect 16816 10610 16871 10665
tri 16871 10610 17046 10785 sw
tri 17109 10665 17229 10785 ne
rect 17229 10665 17265 10785
rect 17385 10665 17421 10785
rect 16816 10528 17046 10610
tri 17046 10528 17128 10610 sw
tri 17229 10528 17366 10665 ne
rect 17366 10610 17421 10665
tri 17421 10610 17596 10785 sw
tri 17659 10665 17779 10785 ne
rect 17779 10665 17815 10785
rect 17935 10665 17971 10785
rect 17366 10528 17596 10610
tri 17596 10528 17678 10610 sw
tri 17779 10528 17916 10665 ne
rect 17916 10610 17971 10665
tri 17971 10610 18146 10785 sw
tri 18209 10665 18329 10785 ne
rect 18329 10665 18365 10785
rect 18485 10665 18521 10785
rect 17916 10528 18146 10610
tri 18146 10528 18228 10610 sw
tri 18329 10528 18466 10665 ne
rect 18466 10610 18521 10665
tri 18521 10610 18696 10785 sw
tri 18759 10665 18879 10785 ne
rect 18879 10665 18915 10785
rect 19035 10665 19071 10785
rect 18466 10528 18696 10610
tri 18696 10528 18778 10610 sw
tri 18879 10528 19016 10665 ne
rect 19016 10610 19071 10665
tri 19071 10610 19246 10785 sw
tri 19309 10665 19429 10785 ne
rect 19429 10665 19465 10785
rect 19585 10683 19621 10785
tri 19621 10683 19723 10785 sw
rect 20800 10683 21800 11472
rect 19585 10665 21800 10683
rect 19016 10528 19246 10610
tri 19246 10528 19328 10610 sw
tri 19429 10528 19566 10665 ne
rect 19566 10528 21800 10665
rect -500 10372 78 10528
tri 78 10372 234 10528 sw
tri 316 10372 472 10528 ne
rect 472 10372 628 10528
tri 628 10372 784 10528 sw
tri 866 10372 1022 10528 ne
rect 1022 10372 1178 10528
tri 1178 10372 1334 10528 sw
tri 1416 10372 1572 10528 ne
rect 1572 10372 1728 10528
tri 1728 10372 1884 10528 sw
tri 1966 10372 2122 10528 ne
rect 2122 10372 2278 10528
tri 2278 10372 2434 10528 sw
tri 2516 10372 2672 10528 ne
rect 2672 10372 2828 10528
tri 2828 10372 2984 10528 sw
tri 3066 10372 3222 10528 ne
rect 3222 10372 3378 10528
tri 3378 10372 3534 10528 sw
tri 3616 10372 3772 10528 ne
rect 3772 10372 3928 10528
tri 3928 10372 4084 10528 sw
tri 4166 10372 4322 10528 ne
rect 4322 10372 4478 10528
tri 4478 10372 4634 10528 sw
tri 4716 10372 4872 10528 ne
rect 4872 10372 5028 10528
tri 5028 10372 5184 10528 sw
tri 5266 10372 5422 10528 ne
rect 5422 10372 5578 10528
tri 5578 10372 5734 10528 sw
tri 5816 10372 5972 10528 ne
rect 5972 10372 6128 10528
tri 6128 10372 6284 10528 sw
tri 6366 10372 6522 10528 ne
rect 6522 10372 6678 10528
tri 6678 10372 6834 10528 sw
tri 6916 10372 7072 10528 ne
rect 7072 10372 7228 10528
tri 7228 10372 7384 10528 sw
tri 7466 10372 7622 10528 ne
rect 7622 10372 7778 10528
tri 7778 10372 7934 10528 sw
tri 8016 10372 8172 10528 ne
rect 8172 10372 8328 10528
tri 8328 10372 8484 10528 sw
tri 8566 10372 8722 10528 ne
rect 8722 10372 8878 10528
tri 8878 10372 9034 10528 sw
tri 9116 10372 9272 10528 ne
rect 9272 10372 9428 10528
tri 9428 10372 9584 10528 sw
tri 9666 10372 9822 10528 ne
rect 9822 10372 9978 10528
tri 9978 10372 10134 10528 sw
tri 10216 10372 10372 10528 ne
rect 10372 10372 10528 10528
tri 10528 10372 10684 10528 sw
tri 10766 10372 10922 10528 ne
rect 10922 10372 11078 10528
tri 11078 10372 11234 10528 sw
tri 11316 10372 11472 10528 ne
rect 11472 10372 11628 10528
tri 11628 10372 11784 10528 sw
tri 11866 10372 12022 10528 ne
rect 12022 10372 12178 10528
tri 12178 10372 12334 10528 sw
tri 12416 10372 12572 10528 ne
rect 12572 10372 12728 10528
tri 12728 10372 12884 10528 sw
tri 12966 10372 13122 10528 ne
rect 13122 10372 13278 10528
tri 13278 10372 13434 10528 sw
tri 13516 10372 13672 10528 ne
rect 13672 10372 13828 10528
tri 13828 10372 13984 10528 sw
tri 14066 10372 14222 10528 ne
rect 14222 10372 14378 10528
tri 14378 10372 14534 10528 sw
tri 14616 10372 14772 10528 ne
rect 14772 10372 14928 10528
tri 14928 10372 15084 10528 sw
tri 15166 10372 15322 10528 ne
rect 15322 10372 15478 10528
tri 15478 10372 15634 10528 sw
tri 15716 10372 15872 10528 ne
rect 15872 10372 16028 10528
tri 16028 10372 16184 10528 sw
tri 16266 10372 16422 10528 ne
rect 16422 10372 16578 10528
tri 16578 10372 16734 10528 sw
tri 16816 10372 16972 10528 ne
rect 16972 10372 17128 10528
tri 17128 10372 17284 10528 sw
tri 17366 10372 17522 10528 ne
rect 17522 10372 17678 10528
tri 17678 10372 17834 10528 sw
tri 17916 10372 18072 10528 ne
rect 18072 10372 18228 10528
tri 18228 10372 18384 10528 sw
tri 18466 10372 18622 10528 ne
rect 18622 10372 18778 10528
tri 18778 10372 18934 10528 sw
tri 19016 10372 19172 10528 ne
rect 19172 10372 19328 10528
tri 19328 10372 19484 10528 sw
tri 19566 10372 19722 10528 ne
rect 19722 10372 21800 10528
rect -500 10235 234 10372
tri 234 10235 371 10372 sw
tri 472 10235 609 10372 ne
rect 609 10235 784 10372
tri 784 10235 921 10372 sw
tri 1022 10235 1159 10372 ne
rect 1159 10235 1334 10372
tri 1334 10235 1471 10372 sw
tri 1572 10235 1709 10372 ne
rect 1709 10235 1884 10372
tri 1884 10235 2021 10372 sw
tri 2122 10235 2259 10372 ne
rect 2259 10235 2434 10372
tri 2434 10235 2571 10372 sw
tri 2672 10235 2809 10372 ne
rect 2809 10235 2984 10372
tri 2984 10235 3121 10372 sw
tri 3222 10235 3359 10372 ne
rect 3359 10235 3534 10372
tri 3534 10235 3671 10372 sw
tri 3772 10235 3909 10372 ne
rect 3909 10235 4084 10372
tri 4084 10235 4221 10372 sw
tri 4322 10235 4459 10372 ne
rect 4459 10235 4634 10372
tri 4634 10235 4771 10372 sw
tri 4872 10235 5009 10372 ne
rect 5009 10235 5184 10372
tri 5184 10235 5321 10372 sw
tri 5422 10235 5559 10372 ne
rect 5559 10235 5734 10372
tri 5734 10235 5871 10372 sw
tri 5972 10235 6109 10372 ne
rect 6109 10235 6284 10372
tri 6284 10235 6421 10372 sw
tri 6522 10235 6659 10372 ne
rect 6659 10235 6834 10372
tri 6834 10235 6971 10372 sw
tri 7072 10235 7209 10372 ne
rect 7209 10235 7384 10372
tri 7384 10235 7521 10372 sw
tri 7622 10235 7759 10372 ne
rect 7759 10235 7934 10372
tri 7934 10235 8071 10372 sw
tri 8172 10235 8309 10372 ne
rect 8309 10235 8484 10372
tri 8484 10235 8621 10372 sw
tri 8722 10235 8859 10372 ne
rect 8859 10235 9034 10372
tri 9034 10235 9171 10372 sw
tri 9272 10235 9409 10372 ne
rect 9409 10235 9584 10372
tri 9584 10235 9721 10372 sw
tri 9822 10235 9959 10372 ne
rect 9959 10235 10134 10372
tri 10134 10235 10271 10372 sw
tri 10372 10235 10509 10372 ne
rect 10509 10235 10684 10372
tri 10684 10235 10821 10372 sw
tri 10922 10235 11059 10372 ne
rect 11059 10235 11234 10372
tri 11234 10235 11371 10372 sw
tri 11472 10235 11609 10372 ne
rect 11609 10235 11784 10372
tri 11784 10235 11921 10372 sw
tri 12022 10235 12159 10372 ne
rect 12159 10235 12334 10372
tri 12334 10235 12471 10372 sw
tri 12572 10235 12709 10372 ne
rect 12709 10235 12884 10372
tri 12884 10235 13021 10372 sw
tri 13122 10235 13259 10372 ne
rect 13259 10235 13434 10372
tri 13434 10235 13571 10372 sw
tri 13672 10235 13809 10372 ne
rect 13809 10235 13984 10372
tri 13984 10235 14121 10372 sw
tri 14222 10235 14359 10372 ne
rect 14359 10235 14534 10372
tri 14534 10235 14671 10372 sw
tri 14772 10235 14909 10372 ne
rect 14909 10235 15084 10372
tri 15084 10235 15221 10372 sw
tri 15322 10235 15459 10372 ne
rect 15459 10235 15634 10372
tri 15634 10235 15771 10372 sw
tri 15872 10235 16009 10372 ne
rect 16009 10235 16184 10372
tri 16184 10235 16321 10372 sw
tri 16422 10235 16559 10372 ne
rect 16559 10235 16734 10372
tri 16734 10235 16871 10372 sw
tri 16972 10235 17109 10372 ne
rect 17109 10235 17284 10372
tri 17284 10235 17421 10372 sw
tri 17522 10235 17659 10372 ne
rect 17659 10235 17834 10372
tri 17834 10235 17971 10372 sw
tri 18072 10235 18209 10372 ne
rect 18209 10235 18384 10372
tri 18384 10235 18521 10372 sw
tri 18622 10235 18759 10372 ne
rect 18759 10235 18934 10372
tri 18934 10235 19071 10372 sw
tri 19172 10235 19309 10372 ne
rect 19309 10235 19484 10372
tri 19484 10235 19621 10372 sw
rect -500 10217 215 10235
tri 77 10115 179 10217 ne
rect 179 10115 215 10217
rect 335 10115 371 10235
tri 179 9978 316 10115 ne
rect 316 10060 371 10115
tri 371 10060 546 10235 sw
tri 609 10115 729 10235 ne
rect 729 10115 765 10235
rect 885 10115 921 10235
rect 316 9978 546 10060
tri 546 9978 628 10060 sw
tri 729 9978 866 10115 ne
rect 866 10060 921 10115
tri 921 10060 1096 10235 sw
tri 1159 10115 1279 10235 ne
rect 1279 10115 1315 10235
rect 1435 10115 1471 10235
rect 866 9978 1096 10060
tri 1096 9978 1178 10060 sw
tri 1279 9978 1416 10115 ne
rect 1416 10060 1471 10115
tri 1471 10060 1646 10235 sw
tri 1709 10115 1829 10235 ne
rect 1829 10115 1865 10235
rect 1985 10115 2021 10235
rect 1416 9978 1646 10060
tri 1646 9978 1728 10060 sw
tri 1829 9978 1966 10115 ne
rect 1966 10060 2021 10115
tri 2021 10060 2196 10235 sw
tri 2259 10115 2379 10235 ne
rect 2379 10115 2415 10235
rect 2535 10115 2571 10235
rect 1966 9978 2196 10060
tri 2196 9978 2278 10060 sw
tri 2379 9978 2516 10115 ne
rect 2516 10060 2571 10115
tri 2571 10060 2746 10235 sw
tri 2809 10115 2929 10235 ne
rect 2929 10115 2965 10235
rect 3085 10115 3121 10235
rect 2516 9978 2746 10060
tri 2746 9978 2828 10060 sw
tri 2929 9978 3066 10115 ne
rect 3066 10060 3121 10115
tri 3121 10060 3296 10235 sw
tri 3359 10115 3479 10235 ne
rect 3479 10115 3515 10235
rect 3635 10115 3671 10235
rect 3066 9978 3296 10060
tri 3296 9978 3378 10060 sw
tri 3479 9978 3616 10115 ne
rect 3616 10060 3671 10115
tri 3671 10060 3846 10235 sw
tri 3909 10115 4029 10235 ne
rect 4029 10115 4065 10235
rect 4185 10115 4221 10235
rect 3616 9978 3846 10060
tri 3846 9978 3928 10060 sw
tri 4029 9978 4166 10115 ne
rect 4166 10060 4221 10115
tri 4221 10060 4396 10235 sw
tri 4459 10115 4579 10235 ne
rect 4579 10115 4615 10235
rect 4735 10115 4771 10235
rect 4166 9978 4396 10060
tri 4396 9978 4478 10060 sw
tri 4579 9978 4716 10115 ne
rect 4716 10060 4771 10115
tri 4771 10060 4946 10235 sw
tri 5009 10115 5129 10235 ne
rect 5129 10115 5165 10235
rect 5285 10115 5321 10235
rect 4716 9978 4946 10060
tri 4946 9978 5028 10060 sw
tri 5129 9978 5266 10115 ne
rect 5266 10060 5321 10115
tri 5321 10060 5496 10235 sw
tri 5559 10115 5679 10235 ne
rect 5679 10115 5715 10235
rect 5835 10115 5871 10235
rect 5266 9978 5496 10060
tri 5496 9978 5578 10060 sw
tri 5679 9978 5816 10115 ne
rect 5816 10060 5871 10115
tri 5871 10060 6046 10235 sw
tri 6109 10115 6229 10235 ne
rect 6229 10115 6265 10235
rect 6385 10115 6421 10235
rect 5816 9978 6046 10060
tri 6046 9978 6128 10060 sw
tri 6229 9978 6366 10115 ne
rect 6366 10060 6421 10115
tri 6421 10060 6596 10235 sw
tri 6659 10115 6779 10235 ne
rect 6779 10115 6815 10235
rect 6935 10115 6971 10235
rect 6366 9978 6596 10060
tri 6596 9978 6678 10060 sw
tri 6779 9978 6916 10115 ne
rect 6916 10060 6971 10115
tri 6971 10060 7146 10235 sw
tri 7209 10115 7329 10235 ne
rect 7329 10115 7365 10235
rect 7485 10115 7521 10235
rect 6916 9978 7146 10060
tri 7146 9978 7228 10060 sw
tri 7329 9978 7466 10115 ne
rect 7466 10060 7521 10115
tri 7521 10060 7696 10235 sw
tri 7759 10115 7879 10235 ne
rect 7879 10115 7915 10235
rect 8035 10115 8071 10235
rect 7466 9978 7696 10060
tri 7696 9978 7778 10060 sw
tri 7879 9978 8016 10115 ne
rect 8016 10060 8071 10115
tri 8071 10060 8246 10235 sw
tri 8309 10115 8429 10235 ne
rect 8429 10115 8465 10235
rect 8585 10115 8621 10235
rect 8016 9978 8246 10060
tri 8246 9978 8328 10060 sw
tri 8429 9978 8566 10115 ne
rect 8566 10060 8621 10115
tri 8621 10060 8796 10235 sw
tri 8859 10115 8979 10235 ne
rect 8979 10115 9015 10235
rect 9135 10115 9171 10235
rect 8566 9978 8796 10060
tri 8796 9978 8878 10060 sw
tri 8979 9978 9116 10115 ne
rect 9116 10060 9171 10115
tri 9171 10060 9346 10235 sw
tri 9409 10115 9529 10235 ne
rect 9529 10115 9565 10235
rect 9685 10115 9721 10235
rect 9116 9978 9346 10060
tri 9346 9978 9428 10060 sw
tri 9529 9978 9666 10115 ne
rect 9666 10060 9721 10115
tri 9721 10060 9896 10235 sw
tri 9959 10115 10079 10235 ne
rect 10079 10115 10115 10235
rect 10235 10115 10271 10235
rect 9666 9978 9896 10060
tri 9896 9978 9978 10060 sw
tri 10079 9978 10216 10115 ne
rect 10216 10060 10271 10115
tri 10271 10060 10446 10235 sw
tri 10509 10115 10629 10235 ne
rect 10629 10115 10665 10235
rect 10785 10115 10821 10235
rect 10216 9978 10446 10060
tri 10446 9978 10528 10060 sw
tri 10629 9978 10766 10115 ne
rect 10766 10060 10821 10115
tri 10821 10060 10996 10235 sw
tri 11059 10115 11179 10235 ne
rect 11179 10115 11215 10235
rect 11335 10115 11371 10235
rect 10766 9978 10996 10060
tri 10996 9978 11078 10060 sw
tri 11179 9978 11316 10115 ne
rect 11316 10060 11371 10115
tri 11371 10060 11546 10235 sw
tri 11609 10115 11729 10235 ne
rect 11729 10115 11765 10235
rect 11885 10115 11921 10235
rect 11316 9978 11546 10060
tri 11546 9978 11628 10060 sw
tri 11729 9978 11866 10115 ne
rect 11866 10060 11921 10115
tri 11921 10060 12096 10235 sw
tri 12159 10115 12279 10235 ne
rect 12279 10115 12315 10235
rect 12435 10115 12471 10235
rect 11866 9978 12096 10060
tri 12096 9978 12178 10060 sw
tri 12279 9978 12416 10115 ne
rect 12416 10060 12471 10115
tri 12471 10060 12646 10235 sw
tri 12709 10115 12829 10235 ne
rect 12829 10115 12865 10235
rect 12985 10115 13021 10235
rect 12416 9978 12646 10060
tri 12646 9978 12728 10060 sw
tri 12829 9978 12966 10115 ne
rect 12966 10060 13021 10115
tri 13021 10060 13196 10235 sw
tri 13259 10115 13379 10235 ne
rect 13379 10115 13415 10235
rect 13535 10115 13571 10235
rect 12966 9978 13196 10060
tri 13196 9978 13278 10060 sw
tri 13379 9978 13516 10115 ne
rect 13516 10060 13571 10115
tri 13571 10060 13746 10235 sw
tri 13809 10115 13929 10235 ne
rect 13929 10115 13965 10235
rect 14085 10115 14121 10235
rect 13516 9978 13746 10060
tri 13746 9978 13828 10060 sw
tri 13929 9978 14066 10115 ne
rect 14066 10060 14121 10115
tri 14121 10060 14296 10235 sw
tri 14359 10115 14479 10235 ne
rect 14479 10115 14515 10235
rect 14635 10115 14671 10235
rect 14066 9978 14296 10060
tri 14296 9978 14378 10060 sw
tri 14479 9978 14616 10115 ne
rect 14616 10060 14671 10115
tri 14671 10060 14846 10235 sw
tri 14909 10115 15029 10235 ne
rect 15029 10115 15065 10235
rect 15185 10115 15221 10235
rect 14616 9978 14846 10060
tri 14846 9978 14928 10060 sw
tri 15029 9978 15166 10115 ne
rect 15166 10060 15221 10115
tri 15221 10060 15396 10235 sw
tri 15459 10115 15579 10235 ne
rect 15579 10115 15615 10235
rect 15735 10115 15771 10235
rect 15166 9978 15396 10060
tri 15396 9978 15478 10060 sw
tri 15579 9978 15716 10115 ne
rect 15716 10060 15771 10115
tri 15771 10060 15946 10235 sw
tri 16009 10115 16129 10235 ne
rect 16129 10115 16165 10235
rect 16285 10115 16321 10235
rect 15716 9978 15946 10060
tri 15946 9978 16028 10060 sw
tri 16129 9978 16266 10115 ne
rect 16266 10060 16321 10115
tri 16321 10060 16496 10235 sw
tri 16559 10115 16679 10235 ne
rect 16679 10115 16715 10235
rect 16835 10115 16871 10235
rect 16266 9978 16496 10060
tri 16496 9978 16578 10060 sw
tri 16679 9978 16816 10115 ne
rect 16816 10060 16871 10115
tri 16871 10060 17046 10235 sw
tri 17109 10115 17229 10235 ne
rect 17229 10115 17265 10235
rect 17385 10115 17421 10235
rect 16816 9978 17046 10060
tri 17046 9978 17128 10060 sw
tri 17229 9978 17366 10115 ne
rect 17366 10060 17421 10115
tri 17421 10060 17596 10235 sw
tri 17659 10115 17779 10235 ne
rect 17779 10115 17815 10235
rect 17935 10115 17971 10235
rect 17366 9978 17596 10060
tri 17596 9978 17678 10060 sw
tri 17779 9978 17916 10115 ne
rect 17916 10060 17971 10115
tri 17971 10060 18146 10235 sw
tri 18209 10115 18329 10235 ne
rect 18329 10115 18365 10235
rect 18485 10115 18521 10235
rect 17916 9978 18146 10060
tri 18146 9978 18228 10060 sw
tri 18329 9978 18466 10115 ne
rect 18466 10060 18521 10115
tri 18521 10060 18696 10235 sw
tri 18759 10115 18879 10235 ne
rect 18879 10115 18915 10235
rect 19035 10115 19071 10235
rect 18466 9978 18696 10060
tri 18696 9978 18778 10060 sw
tri 18879 9978 19016 10115 ne
rect 19016 10060 19071 10115
tri 19071 10060 19246 10235 sw
tri 19309 10115 19429 10235 ne
rect 19429 10115 19465 10235
rect 19585 10133 19621 10235
tri 19621 10133 19723 10235 sw
rect 19585 10115 20300 10133
rect 19016 9978 19246 10060
tri 19246 9978 19328 10060 sw
tri 19429 9978 19566 10115 ne
rect 19566 9978 20300 10115
rect -2000 9822 78 9978
tri 78 9822 234 9978 sw
tri 316 9822 472 9978 ne
rect 472 9822 628 9978
tri 628 9822 784 9978 sw
tri 866 9822 1022 9978 ne
rect 1022 9822 1178 9978
tri 1178 9822 1334 9978 sw
tri 1416 9822 1572 9978 ne
rect 1572 9822 1728 9978
tri 1728 9822 1884 9978 sw
tri 1966 9822 2122 9978 ne
rect 2122 9822 2278 9978
tri 2278 9822 2434 9978 sw
tri 2516 9822 2672 9978 ne
rect 2672 9822 2828 9978
tri 2828 9822 2984 9978 sw
tri 3066 9822 3222 9978 ne
rect 3222 9822 3378 9978
tri 3378 9822 3534 9978 sw
tri 3616 9822 3772 9978 ne
rect 3772 9822 3928 9978
tri 3928 9822 4084 9978 sw
tri 4166 9822 4322 9978 ne
rect 4322 9822 4478 9978
tri 4478 9822 4634 9978 sw
tri 4716 9822 4872 9978 ne
rect 4872 9822 5028 9978
tri 5028 9822 5184 9978 sw
tri 5266 9822 5422 9978 ne
rect 5422 9822 5578 9978
tri 5578 9822 5734 9978 sw
tri 5816 9822 5972 9978 ne
rect 5972 9822 6128 9978
tri 6128 9822 6284 9978 sw
tri 6366 9822 6522 9978 ne
rect 6522 9822 6678 9978
tri 6678 9822 6834 9978 sw
tri 6916 9822 7072 9978 ne
rect 7072 9822 7228 9978
tri 7228 9822 7384 9978 sw
tri 7466 9822 7622 9978 ne
rect 7622 9822 7778 9978
tri 7778 9822 7934 9978 sw
tri 8016 9822 8172 9978 ne
rect 8172 9822 8328 9978
tri 8328 9822 8484 9978 sw
tri 8566 9822 8722 9978 ne
rect 8722 9822 8878 9978
tri 8878 9822 9034 9978 sw
tri 9116 9822 9272 9978 ne
rect 9272 9822 9428 9978
tri 9428 9822 9584 9978 sw
tri 9666 9822 9822 9978 ne
rect 9822 9822 9978 9978
tri 9978 9822 10134 9978 sw
tri 10216 9822 10372 9978 ne
rect 10372 9822 10528 9978
tri 10528 9822 10684 9978 sw
tri 10766 9822 10922 9978 ne
rect 10922 9822 11078 9978
tri 11078 9822 11234 9978 sw
tri 11316 9822 11472 9978 ne
rect 11472 9822 11628 9978
tri 11628 9822 11784 9978 sw
tri 11866 9822 12022 9978 ne
rect 12022 9822 12178 9978
tri 12178 9822 12334 9978 sw
tri 12416 9822 12572 9978 ne
rect 12572 9822 12728 9978
tri 12728 9822 12884 9978 sw
tri 12966 9822 13122 9978 ne
rect 13122 9822 13278 9978
tri 13278 9822 13434 9978 sw
tri 13516 9822 13672 9978 ne
rect 13672 9822 13828 9978
tri 13828 9822 13984 9978 sw
tri 14066 9822 14222 9978 ne
rect 14222 9822 14378 9978
tri 14378 9822 14534 9978 sw
tri 14616 9822 14772 9978 ne
rect 14772 9822 14928 9978
tri 14928 9822 15084 9978 sw
tri 15166 9822 15322 9978 ne
rect 15322 9822 15478 9978
tri 15478 9822 15634 9978 sw
tri 15716 9822 15872 9978 ne
rect 15872 9822 16028 9978
tri 16028 9822 16184 9978 sw
tri 16266 9822 16422 9978 ne
rect 16422 9822 16578 9978
tri 16578 9822 16734 9978 sw
tri 16816 9822 16972 9978 ne
rect 16972 9822 17128 9978
tri 17128 9822 17284 9978 sw
tri 17366 9822 17522 9978 ne
rect 17522 9822 17678 9978
tri 17678 9822 17834 9978 sw
tri 17916 9822 18072 9978 ne
rect 18072 9822 18228 9978
tri 18228 9822 18384 9978 sw
tri 18466 9822 18622 9978 ne
rect 18622 9822 18778 9978
tri 18778 9822 18934 9978 sw
tri 19016 9822 19172 9978 ne
rect 19172 9822 19328 9978
tri 19328 9822 19484 9978 sw
tri 19566 9822 19722 9978 ne
rect 19722 9822 20300 9978
rect -2000 9685 234 9822
tri 234 9685 371 9822 sw
tri 472 9685 609 9822 ne
rect 609 9685 784 9822
tri 784 9685 921 9822 sw
tri 1022 9685 1159 9822 ne
rect 1159 9685 1334 9822
tri 1334 9685 1471 9822 sw
tri 1572 9685 1709 9822 ne
rect 1709 9685 1884 9822
tri 1884 9685 2021 9822 sw
tri 2122 9685 2259 9822 ne
rect 2259 9685 2434 9822
tri 2434 9685 2571 9822 sw
tri 2672 9685 2809 9822 ne
rect 2809 9685 2984 9822
tri 2984 9685 3121 9822 sw
tri 3222 9685 3359 9822 ne
rect 3359 9685 3534 9822
tri 3534 9685 3671 9822 sw
tri 3772 9685 3909 9822 ne
rect 3909 9685 4084 9822
tri 4084 9685 4221 9822 sw
tri 4322 9685 4459 9822 ne
rect 4459 9685 4634 9822
tri 4634 9685 4771 9822 sw
tri 4872 9685 5009 9822 ne
rect 5009 9685 5184 9822
tri 5184 9685 5321 9822 sw
tri 5422 9685 5559 9822 ne
rect 5559 9685 5734 9822
tri 5734 9685 5871 9822 sw
tri 5972 9685 6109 9822 ne
rect 6109 9685 6284 9822
tri 6284 9685 6421 9822 sw
tri 6522 9685 6659 9822 ne
rect 6659 9685 6834 9822
tri 6834 9685 6971 9822 sw
tri 7072 9685 7209 9822 ne
rect 7209 9685 7384 9822
tri 7384 9685 7521 9822 sw
tri 7622 9685 7759 9822 ne
rect 7759 9685 7934 9822
tri 7934 9685 8071 9822 sw
tri 8172 9685 8309 9822 ne
rect 8309 9685 8484 9822
tri 8484 9685 8621 9822 sw
tri 8722 9685 8859 9822 ne
rect 8859 9685 9034 9822
tri 9034 9685 9171 9822 sw
tri 9272 9685 9409 9822 ne
rect 9409 9685 9584 9822
tri 9584 9685 9721 9822 sw
tri 9822 9685 9959 9822 ne
rect 9959 9685 10134 9822
tri 10134 9685 10271 9822 sw
tri 10372 9685 10509 9822 ne
rect 10509 9685 10684 9822
tri 10684 9685 10821 9822 sw
tri 10922 9685 11059 9822 ne
rect 11059 9685 11234 9822
tri 11234 9685 11371 9822 sw
tri 11472 9685 11609 9822 ne
rect 11609 9685 11784 9822
tri 11784 9685 11921 9822 sw
tri 12022 9685 12159 9822 ne
rect 12159 9685 12334 9822
tri 12334 9685 12471 9822 sw
tri 12572 9685 12709 9822 ne
rect 12709 9685 12884 9822
tri 12884 9685 13021 9822 sw
tri 13122 9685 13259 9822 ne
rect 13259 9685 13434 9822
tri 13434 9685 13571 9822 sw
tri 13672 9685 13809 9822 ne
rect 13809 9685 13984 9822
tri 13984 9685 14121 9822 sw
tri 14222 9685 14359 9822 ne
rect 14359 9685 14534 9822
tri 14534 9685 14671 9822 sw
tri 14772 9685 14909 9822 ne
rect 14909 9685 15084 9822
tri 15084 9685 15221 9822 sw
tri 15322 9685 15459 9822 ne
rect 15459 9685 15634 9822
tri 15634 9685 15771 9822 sw
tri 15872 9685 16009 9822 ne
rect 16009 9685 16184 9822
tri 16184 9685 16321 9822 sw
tri 16422 9685 16559 9822 ne
rect 16559 9685 16734 9822
tri 16734 9685 16871 9822 sw
tri 16972 9685 17109 9822 ne
rect 17109 9685 17284 9822
tri 17284 9685 17421 9822 sw
tri 17522 9685 17659 9822 ne
rect 17659 9685 17834 9822
tri 17834 9685 17971 9822 sw
tri 18072 9685 18209 9822 ne
rect 18209 9685 18384 9822
tri 18384 9685 18521 9822 sw
tri 18622 9685 18759 9822 ne
rect 18759 9685 18934 9822
tri 18934 9685 19071 9822 sw
tri 19172 9685 19309 9822 ne
rect 19309 9685 19484 9822
tri 19484 9685 19621 9822 sw
rect -2000 9667 215 9685
rect -2000 8878 -1000 9667
tri 77 9565 179 9667 ne
rect 179 9565 215 9667
rect 335 9565 371 9685
tri 179 9428 316 9565 ne
rect 316 9510 371 9565
tri 371 9510 546 9685 sw
tri 609 9565 729 9685 ne
rect 729 9565 765 9685
rect 885 9565 921 9685
rect 316 9428 546 9510
tri 546 9428 628 9510 sw
tri 729 9428 866 9565 ne
rect 866 9510 921 9565
tri 921 9510 1096 9685 sw
tri 1159 9565 1279 9685 ne
rect 1279 9565 1315 9685
rect 1435 9565 1471 9685
rect 866 9428 1096 9510
tri 1096 9428 1178 9510 sw
tri 1279 9428 1416 9565 ne
rect 1416 9510 1471 9565
tri 1471 9510 1646 9685 sw
tri 1709 9565 1829 9685 ne
rect 1829 9565 1865 9685
rect 1985 9565 2021 9685
rect 1416 9428 1646 9510
tri 1646 9428 1728 9510 sw
tri 1829 9428 1966 9565 ne
rect 1966 9510 2021 9565
tri 2021 9510 2196 9685 sw
tri 2259 9565 2379 9685 ne
rect 2379 9565 2415 9685
rect 2535 9565 2571 9685
rect 1966 9428 2196 9510
tri 2196 9428 2278 9510 sw
tri 2379 9428 2516 9565 ne
rect 2516 9510 2571 9565
tri 2571 9510 2746 9685 sw
tri 2809 9565 2929 9685 ne
rect 2929 9565 2965 9685
rect 3085 9565 3121 9685
rect 2516 9428 2746 9510
tri 2746 9428 2828 9510 sw
tri 2929 9428 3066 9565 ne
rect 3066 9510 3121 9565
tri 3121 9510 3296 9685 sw
tri 3359 9565 3479 9685 ne
rect 3479 9565 3515 9685
rect 3635 9565 3671 9685
rect 3066 9428 3296 9510
tri 3296 9428 3378 9510 sw
tri 3479 9428 3616 9565 ne
rect 3616 9510 3671 9565
tri 3671 9510 3846 9685 sw
tri 3909 9565 4029 9685 ne
rect 4029 9565 4065 9685
rect 4185 9565 4221 9685
rect 3616 9428 3846 9510
tri 3846 9428 3928 9510 sw
tri 4029 9428 4166 9565 ne
rect 4166 9510 4221 9565
tri 4221 9510 4396 9685 sw
tri 4459 9565 4579 9685 ne
rect 4579 9565 4615 9685
rect 4735 9565 4771 9685
rect 4166 9428 4396 9510
tri 4396 9428 4478 9510 sw
tri 4579 9428 4716 9565 ne
rect 4716 9510 4771 9565
tri 4771 9510 4946 9685 sw
tri 5009 9565 5129 9685 ne
rect 5129 9565 5165 9685
rect 5285 9565 5321 9685
rect 4716 9428 4946 9510
tri 4946 9428 5028 9510 sw
tri 5129 9428 5266 9565 ne
rect 5266 9510 5321 9565
tri 5321 9510 5496 9685 sw
tri 5559 9565 5679 9685 ne
rect 5679 9565 5715 9685
rect 5835 9565 5871 9685
rect 5266 9428 5496 9510
tri 5496 9428 5578 9510 sw
tri 5679 9428 5816 9565 ne
rect 5816 9510 5871 9565
tri 5871 9510 6046 9685 sw
tri 6109 9565 6229 9685 ne
rect 6229 9565 6265 9685
rect 6385 9565 6421 9685
rect 5816 9428 6046 9510
tri 6046 9428 6128 9510 sw
tri 6229 9428 6366 9565 ne
rect 6366 9510 6421 9565
tri 6421 9510 6596 9685 sw
tri 6659 9565 6779 9685 ne
rect 6779 9565 6815 9685
rect 6935 9565 6971 9685
rect 6366 9428 6596 9510
tri 6596 9428 6678 9510 sw
tri 6779 9428 6916 9565 ne
rect 6916 9510 6971 9565
tri 6971 9510 7146 9685 sw
tri 7209 9565 7329 9685 ne
rect 7329 9565 7365 9685
rect 7485 9565 7521 9685
rect 6916 9428 7146 9510
tri 7146 9428 7228 9510 sw
tri 7329 9428 7466 9565 ne
rect 7466 9510 7521 9565
tri 7521 9510 7696 9685 sw
tri 7759 9565 7879 9685 ne
rect 7879 9565 7915 9685
rect 8035 9565 8071 9685
rect 7466 9428 7696 9510
tri 7696 9428 7778 9510 sw
tri 7879 9428 8016 9565 ne
rect 8016 9510 8071 9565
tri 8071 9510 8246 9685 sw
tri 8309 9565 8429 9685 ne
rect 8429 9565 8465 9685
rect 8585 9565 8621 9685
rect 8016 9428 8246 9510
tri 8246 9428 8328 9510 sw
tri 8429 9428 8566 9565 ne
rect 8566 9510 8621 9565
tri 8621 9510 8796 9685 sw
tri 8859 9565 8979 9685 ne
rect 8979 9565 9015 9685
rect 9135 9565 9171 9685
rect 8566 9428 8796 9510
tri 8796 9428 8878 9510 sw
tri 8979 9428 9116 9565 ne
rect 9116 9510 9171 9565
tri 9171 9510 9346 9685 sw
tri 9409 9565 9529 9685 ne
rect 9529 9565 9565 9685
rect 9685 9565 9721 9685
rect 9116 9428 9346 9510
tri 9346 9428 9428 9510 sw
tri 9529 9428 9666 9565 ne
rect 9666 9510 9721 9565
tri 9721 9510 9896 9685 sw
tri 9959 9565 10079 9685 ne
rect 10079 9565 10115 9685
rect 10235 9565 10271 9685
rect 9666 9428 9896 9510
tri 9896 9428 9978 9510 sw
tri 10079 9428 10216 9565 ne
rect 10216 9510 10271 9565
tri 10271 9510 10446 9685 sw
tri 10509 9565 10629 9685 ne
rect 10629 9565 10665 9685
rect 10785 9565 10821 9685
rect 10216 9428 10446 9510
tri 10446 9428 10528 9510 sw
tri 10629 9428 10766 9565 ne
rect 10766 9510 10821 9565
tri 10821 9510 10996 9685 sw
tri 11059 9565 11179 9685 ne
rect 11179 9565 11215 9685
rect 11335 9565 11371 9685
rect 10766 9428 10996 9510
tri 10996 9428 11078 9510 sw
tri 11179 9428 11316 9565 ne
rect 11316 9510 11371 9565
tri 11371 9510 11546 9685 sw
tri 11609 9565 11729 9685 ne
rect 11729 9565 11765 9685
rect 11885 9565 11921 9685
rect 11316 9428 11546 9510
tri 11546 9428 11628 9510 sw
tri 11729 9428 11866 9565 ne
rect 11866 9510 11921 9565
tri 11921 9510 12096 9685 sw
tri 12159 9565 12279 9685 ne
rect 12279 9565 12315 9685
rect 12435 9565 12471 9685
rect 11866 9428 12096 9510
tri 12096 9428 12178 9510 sw
tri 12279 9428 12416 9565 ne
rect 12416 9510 12471 9565
tri 12471 9510 12646 9685 sw
tri 12709 9565 12829 9685 ne
rect 12829 9565 12865 9685
rect 12985 9565 13021 9685
rect 12416 9428 12646 9510
tri 12646 9428 12728 9510 sw
tri 12829 9428 12966 9565 ne
rect 12966 9510 13021 9565
tri 13021 9510 13196 9685 sw
tri 13259 9565 13379 9685 ne
rect 13379 9565 13415 9685
rect 13535 9565 13571 9685
rect 12966 9428 13196 9510
tri 13196 9428 13278 9510 sw
tri 13379 9428 13516 9565 ne
rect 13516 9510 13571 9565
tri 13571 9510 13746 9685 sw
tri 13809 9565 13929 9685 ne
rect 13929 9565 13965 9685
rect 14085 9565 14121 9685
rect 13516 9428 13746 9510
tri 13746 9428 13828 9510 sw
tri 13929 9428 14066 9565 ne
rect 14066 9510 14121 9565
tri 14121 9510 14296 9685 sw
tri 14359 9565 14479 9685 ne
rect 14479 9565 14515 9685
rect 14635 9565 14671 9685
rect 14066 9428 14296 9510
tri 14296 9428 14378 9510 sw
tri 14479 9428 14616 9565 ne
rect 14616 9510 14671 9565
tri 14671 9510 14846 9685 sw
tri 14909 9565 15029 9685 ne
rect 15029 9565 15065 9685
rect 15185 9565 15221 9685
rect 14616 9428 14846 9510
tri 14846 9428 14928 9510 sw
tri 15029 9428 15166 9565 ne
rect 15166 9510 15221 9565
tri 15221 9510 15396 9685 sw
tri 15459 9565 15579 9685 ne
rect 15579 9565 15615 9685
rect 15735 9565 15771 9685
rect 15166 9428 15396 9510
tri 15396 9428 15478 9510 sw
tri 15579 9428 15716 9565 ne
rect 15716 9510 15771 9565
tri 15771 9510 15946 9685 sw
tri 16009 9565 16129 9685 ne
rect 16129 9565 16165 9685
rect 16285 9565 16321 9685
rect 15716 9428 15946 9510
tri 15946 9428 16028 9510 sw
tri 16129 9428 16266 9565 ne
rect 16266 9510 16321 9565
tri 16321 9510 16496 9685 sw
tri 16559 9565 16679 9685 ne
rect 16679 9565 16715 9685
rect 16835 9565 16871 9685
rect 16266 9428 16496 9510
tri 16496 9428 16578 9510 sw
tri 16679 9428 16816 9565 ne
rect 16816 9510 16871 9565
tri 16871 9510 17046 9685 sw
tri 17109 9565 17229 9685 ne
rect 17229 9565 17265 9685
rect 17385 9565 17421 9685
rect 16816 9428 17046 9510
tri 17046 9428 17128 9510 sw
tri 17229 9428 17366 9565 ne
rect 17366 9510 17421 9565
tri 17421 9510 17596 9685 sw
tri 17659 9565 17779 9685 ne
rect 17779 9565 17815 9685
rect 17935 9565 17971 9685
rect 17366 9428 17596 9510
tri 17596 9428 17678 9510 sw
tri 17779 9428 17916 9565 ne
rect 17916 9510 17971 9565
tri 17971 9510 18146 9685 sw
tri 18209 9565 18329 9685 ne
rect 18329 9565 18365 9685
rect 18485 9565 18521 9685
rect 17916 9428 18146 9510
tri 18146 9428 18228 9510 sw
tri 18329 9428 18466 9565 ne
rect 18466 9510 18521 9565
tri 18521 9510 18696 9685 sw
tri 18759 9565 18879 9685 ne
rect 18879 9565 18915 9685
rect 19035 9565 19071 9685
rect 18466 9428 18696 9510
tri 18696 9428 18778 9510 sw
tri 18879 9428 19016 9565 ne
rect 19016 9510 19071 9565
tri 19071 9510 19246 9685 sw
tri 19309 9565 19429 9685 ne
rect 19429 9565 19465 9685
rect 19585 9583 19621 9685
tri 19621 9583 19723 9685 sw
rect 20800 9583 21800 10372
rect 19585 9565 21800 9583
rect 19016 9428 19246 9510
tri 19246 9428 19328 9510 sw
tri 19429 9428 19566 9565 ne
rect 19566 9428 21800 9565
rect -500 9272 78 9428
tri 78 9272 234 9428 sw
tri 316 9272 472 9428 ne
rect 472 9272 628 9428
tri 628 9272 784 9428 sw
tri 866 9272 1022 9428 ne
rect 1022 9272 1178 9428
tri 1178 9272 1334 9428 sw
tri 1416 9272 1572 9428 ne
rect 1572 9272 1728 9428
tri 1728 9272 1884 9428 sw
tri 1966 9272 2122 9428 ne
rect 2122 9272 2278 9428
tri 2278 9272 2434 9428 sw
tri 2516 9272 2672 9428 ne
rect 2672 9272 2828 9428
tri 2828 9272 2984 9428 sw
tri 3066 9272 3222 9428 ne
rect 3222 9272 3378 9428
tri 3378 9272 3534 9428 sw
tri 3616 9272 3772 9428 ne
rect 3772 9272 3928 9428
tri 3928 9272 4084 9428 sw
tri 4166 9272 4322 9428 ne
rect 4322 9272 4478 9428
tri 4478 9272 4634 9428 sw
tri 4716 9272 4872 9428 ne
rect 4872 9272 5028 9428
tri 5028 9272 5184 9428 sw
tri 5266 9272 5422 9428 ne
rect 5422 9272 5578 9428
tri 5578 9272 5734 9428 sw
tri 5816 9272 5972 9428 ne
rect 5972 9272 6128 9428
tri 6128 9272 6284 9428 sw
tri 6366 9272 6522 9428 ne
rect 6522 9272 6678 9428
tri 6678 9272 6834 9428 sw
tri 6916 9272 7072 9428 ne
rect 7072 9272 7228 9428
tri 7228 9272 7384 9428 sw
tri 7466 9272 7622 9428 ne
rect 7622 9272 7778 9428
tri 7778 9272 7934 9428 sw
tri 8016 9272 8172 9428 ne
rect 8172 9272 8328 9428
tri 8328 9272 8484 9428 sw
tri 8566 9272 8722 9428 ne
rect 8722 9272 8878 9428
tri 8878 9272 9034 9428 sw
tri 9116 9272 9272 9428 ne
rect 9272 9272 9428 9428
tri 9428 9272 9584 9428 sw
tri 9666 9272 9822 9428 ne
rect 9822 9272 9978 9428
tri 9978 9272 10134 9428 sw
tri 10216 9272 10372 9428 ne
rect 10372 9272 10528 9428
tri 10528 9272 10684 9428 sw
tri 10766 9272 10922 9428 ne
rect 10922 9272 11078 9428
tri 11078 9272 11234 9428 sw
tri 11316 9272 11472 9428 ne
rect 11472 9272 11628 9428
tri 11628 9272 11784 9428 sw
tri 11866 9272 12022 9428 ne
rect 12022 9272 12178 9428
tri 12178 9272 12334 9428 sw
tri 12416 9272 12572 9428 ne
rect 12572 9272 12728 9428
tri 12728 9272 12884 9428 sw
tri 12966 9272 13122 9428 ne
rect 13122 9272 13278 9428
tri 13278 9272 13434 9428 sw
tri 13516 9272 13672 9428 ne
rect 13672 9272 13828 9428
tri 13828 9272 13984 9428 sw
tri 14066 9272 14222 9428 ne
rect 14222 9272 14378 9428
tri 14378 9272 14534 9428 sw
tri 14616 9272 14772 9428 ne
rect 14772 9272 14928 9428
tri 14928 9272 15084 9428 sw
tri 15166 9272 15322 9428 ne
rect 15322 9272 15478 9428
tri 15478 9272 15634 9428 sw
tri 15716 9272 15872 9428 ne
rect 15872 9272 16028 9428
tri 16028 9272 16184 9428 sw
tri 16266 9272 16422 9428 ne
rect 16422 9272 16578 9428
tri 16578 9272 16734 9428 sw
tri 16816 9272 16972 9428 ne
rect 16972 9272 17128 9428
tri 17128 9272 17284 9428 sw
tri 17366 9272 17522 9428 ne
rect 17522 9272 17678 9428
tri 17678 9272 17834 9428 sw
tri 17916 9272 18072 9428 ne
rect 18072 9272 18228 9428
tri 18228 9272 18384 9428 sw
tri 18466 9272 18622 9428 ne
rect 18622 9272 18778 9428
tri 18778 9272 18934 9428 sw
tri 19016 9272 19172 9428 ne
rect 19172 9272 19328 9428
tri 19328 9272 19484 9428 sw
tri 19566 9272 19722 9428 ne
rect 19722 9272 21800 9428
rect -500 9135 234 9272
tri 234 9135 371 9272 sw
tri 472 9135 609 9272 ne
rect 609 9135 784 9272
tri 784 9135 921 9272 sw
tri 1022 9135 1159 9272 ne
rect 1159 9135 1334 9272
tri 1334 9135 1471 9272 sw
tri 1572 9135 1709 9272 ne
rect 1709 9135 1884 9272
tri 1884 9135 2021 9272 sw
tri 2122 9135 2259 9272 ne
rect 2259 9135 2434 9272
tri 2434 9135 2571 9272 sw
tri 2672 9135 2809 9272 ne
rect 2809 9135 2984 9272
tri 2984 9135 3121 9272 sw
tri 3222 9135 3359 9272 ne
rect 3359 9135 3534 9272
tri 3534 9135 3671 9272 sw
tri 3772 9135 3909 9272 ne
rect 3909 9135 4084 9272
tri 4084 9135 4221 9272 sw
tri 4322 9135 4459 9272 ne
rect 4459 9135 4634 9272
tri 4634 9135 4771 9272 sw
tri 4872 9135 5009 9272 ne
rect 5009 9135 5184 9272
tri 5184 9135 5321 9272 sw
tri 5422 9135 5559 9272 ne
rect 5559 9135 5734 9272
tri 5734 9135 5871 9272 sw
tri 5972 9135 6109 9272 ne
rect 6109 9135 6284 9272
tri 6284 9135 6421 9272 sw
tri 6522 9135 6659 9272 ne
rect 6659 9135 6834 9272
tri 6834 9135 6971 9272 sw
tri 7072 9135 7209 9272 ne
rect 7209 9135 7384 9272
tri 7384 9135 7521 9272 sw
tri 7622 9135 7759 9272 ne
rect 7759 9135 7934 9272
tri 7934 9135 8071 9272 sw
tri 8172 9135 8309 9272 ne
rect 8309 9135 8484 9272
tri 8484 9135 8621 9272 sw
tri 8722 9135 8859 9272 ne
rect 8859 9135 9034 9272
tri 9034 9135 9171 9272 sw
tri 9272 9135 9409 9272 ne
rect 9409 9135 9584 9272
tri 9584 9135 9721 9272 sw
tri 9822 9135 9959 9272 ne
rect 9959 9135 10134 9272
tri 10134 9135 10271 9272 sw
tri 10372 9135 10509 9272 ne
rect 10509 9135 10684 9272
tri 10684 9135 10821 9272 sw
tri 10922 9135 11059 9272 ne
rect 11059 9135 11234 9272
tri 11234 9135 11371 9272 sw
tri 11472 9135 11609 9272 ne
rect 11609 9135 11784 9272
tri 11784 9135 11921 9272 sw
tri 12022 9135 12159 9272 ne
rect 12159 9135 12334 9272
tri 12334 9135 12471 9272 sw
tri 12572 9135 12709 9272 ne
rect 12709 9135 12884 9272
tri 12884 9135 13021 9272 sw
tri 13122 9135 13259 9272 ne
rect 13259 9135 13434 9272
tri 13434 9135 13571 9272 sw
tri 13672 9135 13809 9272 ne
rect 13809 9135 13984 9272
tri 13984 9135 14121 9272 sw
tri 14222 9135 14359 9272 ne
rect 14359 9135 14534 9272
tri 14534 9135 14671 9272 sw
tri 14772 9135 14909 9272 ne
rect 14909 9135 15084 9272
tri 15084 9135 15221 9272 sw
tri 15322 9135 15459 9272 ne
rect 15459 9135 15634 9272
tri 15634 9135 15771 9272 sw
tri 15872 9135 16009 9272 ne
rect 16009 9135 16184 9272
tri 16184 9135 16321 9272 sw
tri 16422 9135 16559 9272 ne
rect 16559 9135 16734 9272
tri 16734 9135 16871 9272 sw
tri 16972 9135 17109 9272 ne
rect 17109 9135 17284 9272
tri 17284 9135 17421 9272 sw
tri 17522 9135 17659 9272 ne
rect 17659 9135 17834 9272
tri 17834 9135 17971 9272 sw
tri 18072 9135 18209 9272 ne
rect 18209 9135 18384 9272
tri 18384 9135 18521 9272 sw
tri 18622 9135 18759 9272 ne
rect 18759 9135 18934 9272
tri 18934 9135 19071 9272 sw
tri 19172 9135 19309 9272 ne
rect 19309 9135 19484 9272
tri 19484 9135 19621 9272 sw
rect -500 9117 215 9135
tri 77 9015 179 9117 ne
rect 179 9015 215 9117
rect 335 9015 371 9135
tri 179 8878 316 9015 ne
rect 316 8960 371 9015
tri 371 8960 546 9135 sw
tri 609 9015 729 9135 ne
rect 729 9015 765 9135
rect 885 9015 921 9135
rect 316 8878 546 8960
tri 546 8878 628 8960 sw
tri 729 8878 866 9015 ne
rect 866 8960 921 9015
tri 921 8960 1096 9135 sw
tri 1159 9015 1279 9135 ne
rect 1279 9015 1315 9135
rect 1435 9015 1471 9135
rect 866 8878 1096 8960
tri 1096 8878 1178 8960 sw
tri 1279 8878 1416 9015 ne
rect 1416 8960 1471 9015
tri 1471 8960 1646 9135 sw
tri 1709 9015 1829 9135 ne
rect 1829 9015 1865 9135
rect 1985 9015 2021 9135
rect 1416 8878 1646 8960
tri 1646 8878 1728 8960 sw
tri 1829 8878 1966 9015 ne
rect 1966 8960 2021 9015
tri 2021 8960 2196 9135 sw
tri 2259 9015 2379 9135 ne
rect 2379 9015 2415 9135
rect 2535 9015 2571 9135
rect 1966 8878 2196 8960
tri 2196 8878 2278 8960 sw
tri 2379 8878 2516 9015 ne
rect 2516 8960 2571 9015
tri 2571 8960 2746 9135 sw
tri 2809 9015 2929 9135 ne
rect 2929 9015 2965 9135
rect 3085 9015 3121 9135
rect 2516 8878 2746 8960
tri 2746 8878 2828 8960 sw
tri 2929 8878 3066 9015 ne
rect 3066 8960 3121 9015
tri 3121 8960 3296 9135 sw
tri 3359 9015 3479 9135 ne
rect 3479 9015 3515 9135
rect 3635 9015 3671 9135
rect 3066 8878 3296 8960
tri 3296 8878 3378 8960 sw
tri 3479 8878 3616 9015 ne
rect 3616 8960 3671 9015
tri 3671 8960 3846 9135 sw
tri 3909 9015 4029 9135 ne
rect 4029 9015 4065 9135
rect 4185 9015 4221 9135
rect 3616 8878 3846 8960
tri 3846 8878 3928 8960 sw
tri 4029 8878 4166 9015 ne
rect 4166 8960 4221 9015
tri 4221 8960 4396 9135 sw
tri 4459 9015 4579 9135 ne
rect 4579 9015 4615 9135
rect 4735 9015 4771 9135
rect 4166 8878 4396 8960
tri 4396 8878 4478 8960 sw
tri 4579 8878 4716 9015 ne
rect 4716 8960 4771 9015
tri 4771 8960 4946 9135 sw
tri 5009 9015 5129 9135 ne
rect 5129 9015 5165 9135
rect 5285 9015 5321 9135
rect 4716 8878 4946 8960
tri 4946 8878 5028 8960 sw
tri 5129 8878 5266 9015 ne
rect 5266 8960 5321 9015
tri 5321 8960 5496 9135 sw
tri 5559 9015 5679 9135 ne
rect 5679 9015 5715 9135
rect 5835 9015 5871 9135
rect 5266 8878 5496 8960
tri 5496 8878 5578 8960 sw
tri 5679 8878 5816 9015 ne
rect 5816 8960 5871 9015
tri 5871 8960 6046 9135 sw
tri 6109 9015 6229 9135 ne
rect 6229 9015 6265 9135
rect 6385 9015 6421 9135
rect 5816 8878 6046 8960
tri 6046 8878 6128 8960 sw
tri 6229 8878 6366 9015 ne
rect 6366 8960 6421 9015
tri 6421 8960 6596 9135 sw
tri 6659 9015 6779 9135 ne
rect 6779 9015 6815 9135
rect 6935 9015 6971 9135
rect 6366 8878 6596 8960
tri 6596 8878 6678 8960 sw
tri 6779 8878 6916 9015 ne
rect 6916 8960 6971 9015
tri 6971 8960 7146 9135 sw
tri 7209 9015 7329 9135 ne
rect 7329 9015 7365 9135
rect 7485 9015 7521 9135
rect 6916 8878 7146 8960
tri 7146 8878 7228 8960 sw
tri 7329 8878 7466 9015 ne
rect 7466 8960 7521 9015
tri 7521 8960 7696 9135 sw
tri 7759 9015 7879 9135 ne
rect 7879 9015 7915 9135
rect 8035 9015 8071 9135
rect 7466 8878 7696 8960
tri 7696 8878 7778 8960 sw
tri 7879 8878 8016 9015 ne
rect 8016 8960 8071 9015
tri 8071 8960 8246 9135 sw
tri 8309 9015 8429 9135 ne
rect 8429 9015 8465 9135
rect 8585 9015 8621 9135
rect 8016 8878 8246 8960
tri 8246 8878 8328 8960 sw
tri 8429 8878 8566 9015 ne
rect 8566 8960 8621 9015
tri 8621 8960 8796 9135 sw
tri 8859 9015 8979 9135 ne
rect 8979 9015 9015 9135
rect 9135 9015 9171 9135
rect 8566 8878 8796 8960
tri 8796 8878 8878 8960 sw
tri 8979 8878 9116 9015 ne
rect 9116 8960 9171 9015
tri 9171 8960 9346 9135 sw
tri 9409 9015 9529 9135 ne
rect 9529 9015 9565 9135
rect 9685 9015 9721 9135
rect 9116 8878 9346 8960
tri 9346 8878 9428 8960 sw
tri 9529 8878 9666 9015 ne
rect 9666 8960 9721 9015
tri 9721 8960 9896 9135 sw
tri 9959 9015 10079 9135 ne
rect 10079 9015 10115 9135
rect 10235 9015 10271 9135
rect 9666 8878 9896 8960
tri 9896 8878 9978 8960 sw
tri 10079 8878 10216 9015 ne
rect 10216 8960 10271 9015
tri 10271 8960 10446 9135 sw
tri 10509 9015 10629 9135 ne
rect 10629 9015 10665 9135
rect 10785 9015 10821 9135
rect 10216 8878 10446 8960
tri 10446 8878 10528 8960 sw
tri 10629 8878 10766 9015 ne
rect 10766 8960 10821 9015
tri 10821 8960 10996 9135 sw
tri 11059 9015 11179 9135 ne
rect 11179 9015 11215 9135
rect 11335 9015 11371 9135
rect 10766 8878 10996 8960
tri 10996 8878 11078 8960 sw
tri 11179 8878 11316 9015 ne
rect 11316 8960 11371 9015
tri 11371 8960 11546 9135 sw
tri 11609 9015 11729 9135 ne
rect 11729 9015 11765 9135
rect 11885 9015 11921 9135
rect 11316 8878 11546 8960
tri 11546 8878 11628 8960 sw
tri 11729 8878 11866 9015 ne
rect 11866 8960 11921 9015
tri 11921 8960 12096 9135 sw
tri 12159 9015 12279 9135 ne
rect 12279 9015 12315 9135
rect 12435 9015 12471 9135
rect 11866 8878 12096 8960
tri 12096 8878 12178 8960 sw
tri 12279 8878 12416 9015 ne
rect 12416 8960 12471 9015
tri 12471 8960 12646 9135 sw
tri 12709 9015 12829 9135 ne
rect 12829 9015 12865 9135
rect 12985 9015 13021 9135
rect 12416 8878 12646 8960
tri 12646 8878 12728 8960 sw
tri 12829 8878 12966 9015 ne
rect 12966 8960 13021 9015
tri 13021 8960 13196 9135 sw
tri 13259 9015 13379 9135 ne
rect 13379 9015 13415 9135
rect 13535 9015 13571 9135
rect 12966 8878 13196 8960
tri 13196 8878 13278 8960 sw
tri 13379 8878 13516 9015 ne
rect 13516 8960 13571 9015
tri 13571 8960 13746 9135 sw
tri 13809 9015 13929 9135 ne
rect 13929 9015 13965 9135
rect 14085 9015 14121 9135
rect 13516 8878 13746 8960
tri 13746 8878 13828 8960 sw
tri 13929 8878 14066 9015 ne
rect 14066 8960 14121 9015
tri 14121 8960 14296 9135 sw
tri 14359 9015 14479 9135 ne
rect 14479 9015 14515 9135
rect 14635 9015 14671 9135
rect 14066 8878 14296 8960
tri 14296 8878 14378 8960 sw
tri 14479 8878 14616 9015 ne
rect 14616 8960 14671 9015
tri 14671 8960 14846 9135 sw
tri 14909 9015 15029 9135 ne
rect 15029 9015 15065 9135
rect 15185 9015 15221 9135
rect 14616 8878 14846 8960
tri 14846 8878 14928 8960 sw
tri 15029 8878 15166 9015 ne
rect 15166 8960 15221 9015
tri 15221 8960 15396 9135 sw
tri 15459 9015 15579 9135 ne
rect 15579 9015 15615 9135
rect 15735 9015 15771 9135
rect 15166 8878 15396 8960
tri 15396 8878 15478 8960 sw
tri 15579 8878 15716 9015 ne
rect 15716 8960 15771 9015
tri 15771 8960 15946 9135 sw
tri 16009 9015 16129 9135 ne
rect 16129 9015 16165 9135
rect 16285 9015 16321 9135
rect 15716 8878 15946 8960
tri 15946 8878 16028 8960 sw
tri 16129 8878 16266 9015 ne
rect 16266 8960 16321 9015
tri 16321 8960 16496 9135 sw
tri 16559 9015 16679 9135 ne
rect 16679 9015 16715 9135
rect 16835 9015 16871 9135
rect 16266 8878 16496 8960
tri 16496 8878 16578 8960 sw
tri 16679 8878 16816 9015 ne
rect 16816 8960 16871 9015
tri 16871 8960 17046 9135 sw
tri 17109 9015 17229 9135 ne
rect 17229 9015 17265 9135
rect 17385 9015 17421 9135
rect 16816 8878 17046 8960
tri 17046 8878 17128 8960 sw
tri 17229 8878 17366 9015 ne
rect 17366 8960 17421 9015
tri 17421 8960 17596 9135 sw
tri 17659 9015 17779 9135 ne
rect 17779 9015 17815 9135
rect 17935 9015 17971 9135
rect 17366 8878 17596 8960
tri 17596 8878 17678 8960 sw
tri 17779 8878 17916 9015 ne
rect 17916 8960 17971 9015
tri 17971 8960 18146 9135 sw
tri 18209 9015 18329 9135 ne
rect 18329 9015 18365 9135
rect 18485 9015 18521 9135
rect 17916 8878 18146 8960
tri 18146 8878 18228 8960 sw
tri 18329 8878 18466 9015 ne
rect 18466 8960 18521 9015
tri 18521 8960 18696 9135 sw
tri 18759 9015 18879 9135 ne
rect 18879 9015 18915 9135
rect 19035 9015 19071 9135
rect 18466 8878 18696 8960
tri 18696 8878 18778 8960 sw
tri 18879 8878 19016 9015 ne
rect 19016 8960 19071 9015
tri 19071 8960 19246 9135 sw
tri 19309 9015 19429 9135 ne
rect 19429 9015 19465 9135
rect 19585 9033 19621 9135
tri 19621 9033 19723 9135 sw
rect 19585 9015 20300 9033
rect 19016 8878 19246 8960
tri 19246 8878 19328 8960 sw
tri 19429 8878 19566 9015 ne
rect 19566 8878 20300 9015
rect -2000 8722 78 8878
tri 78 8722 234 8878 sw
tri 316 8722 472 8878 ne
rect 472 8722 628 8878
tri 628 8722 784 8878 sw
tri 866 8722 1022 8878 ne
rect 1022 8722 1178 8878
tri 1178 8722 1334 8878 sw
tri 1416 8722 1572 8878 ne
rect 1572 8722 1728 8878
tri 1728 8722 1884 8878 sw
tri 1966 8722 2122 8878 ne
rect 2122 8722 2278 8878
tri 2278 8722 2434 8878 sw
tri 2516 8722 2672 8878 ne
rect 2672 8722 2828 8878
tri 2828 8722 2984 8878 sw
tri 3066 8722 3222 8878 ne
rect 3222 8722 3378 8878
tri 3378 8722 3534 8878 sw
tri 3616 8722 3772 8878 ne
rect 3772 8722 3928 8878
tri 3928 8722 4084 8878 sw
tri 4166 8722 4322 8878 ne
rect 4322 8722 4478 8878
tri 4478 8722 4634 8878 sw
tri 4716 8722 4872 8878 ne
rect 4872 8722 5028 8878
tri 5028 8722 5184 8878 sw
tri 5266 8722 5422 8878 ne
rect 5422 8722 5578 8878
tri 5578 8722 5734 8878 sw
tri 5816 8722 5972 8878 ne
rect 5972 8722 6128 8878
tri 6128 8722 6284 8878 sw
tri 6366 8722 6522 8878 ne
rect 6522 8722 6678 8878
tri 6678 8722 6834 8878 sw
tri 6916 8722 7072 8878 ne
rect 7072 8722 7228 8878
tri 7228 8722 7384 8878 sw
tri 7466 8722 7622 8878 ne
rect 7622 8722 7778 8878
tri 7778 8722 7934 8878 sw
tri 8016 8722 8172 8878 ne
rect 8172 8722 8328 8878
tri 8328 8722 8484 8878 sw
tri 8566 8722 8722 8878 ne
rect 8722 8722 8878 8878
tri 8878 8722 9034 8878 sw
tri 9116 8722 9272 8878 ne
rect 9272 8722 9428 8878
tri 9428 8722 9584 8878 sw
tri 9666 8722 9822 8878 ne
rect 9822 8722 9978 8878
tri 9978 8722 10134 8878 sw
tri 10216 8722 10372 8878 ne
rect 10372 8722 10528 8878
tri 10528 8722 10684 8878 sw
tri 10766 8722 10922 8878 ne
rect 10922 8722 11078 8878
tri 11078 8722 11234 8878 sw
tri 11316 8722 11472 8878 ne
rect 11472 8722 11628 8878
tri 11628 8722 11784 8878 sw
tri 11866 8722 12022 8878 ne
rect 12022 8722 12178 8878
tri 12178 8722 12334 8878 sw
tri 12416 8722 12572 8878 ne
rect 12572 8722 12728 8878
tri 12728 8722 12884 8878 sw
tri 12966 8722 13122 8878 ne
rect 13122 8722 13278 8878
tri 13278 8722 13434 8878 sw
tri 13516 8722 13672 8878 ne
rect 13672 8722 13828 8878
tri 13828 8722 13984 8878 sw
tri 14066 8722 14222 8878 ne
rect 14222 8722 14378 8878
tri 14378 8722 14534 8878 sw
tri 14616 8722 14772 8878 ne
rect 14772 8722 14928 8878
tri 14928 8722 15084 8878 sw
tri 15166 8722 15322 8878 ne
rect 15322 8722 15478 8878
tri 15478 8722 15634 8878 sw
tri 15716 8722 15872 8878 ne
rect 15872 8722 16028 8878
tri 16028 8722 16184 8878 sw
tri 16266 8722 16422 8878 ne
rect 16422 8722 16578 8878
tri 16578 8722 16734 8878 sw
tri 16816 8722 16972 8878 ne
rect 16972 8722 17128 8878
tri 17128 8722 17284 8878 sw
tri 17366 8722 17522 8878 ne
rect 17522 8722 17678 8878
tri 17678 8722 17834 8878 sw
tri 17916 8722 18072 8878 ne
rect 18072 8722 18228 8878
tri 18228 8722 18384 8878 sw
tri 18466 8722 18622 8878 ne
rect 18622 8722 18778 8878
tri 18778 8722 18934 8878 sw
tri 19016 8722 19172 8878 ne
rect 19172 8722 19328 8878
tri 19328 8722 19484 8878 sw
tri 19566 8722 19722 8878 ne
rect 19722 8722 20300 8878
rect -2000 8585 234 8722
tri 234 8585 371 8722 sw
tri 472 8585 609 8722 ne
rect 609 8585 784 8722
tri 784 8585 921 8722 sw
tri 1022 8585 1159 8722 ne
rect 1159 8585 1334 8722
tri 1334 8585 1471 8722 sw
tri 1572 8585 1709 8722 ne
rect 1709 8585 1884 8722
tri 1884 8585 2021 8722 sw
tri 2122 8585 2259 8722 ne
rect 2259 8585 2434 8722
tri 2434 8585 2571 8722 sw
tri 2672 8585 2809 8722 ne
rect 2809 8585 2984 8722
tri 2984 8585 3121 8722 sw
tri 3222 8585 3359 8722 ne
rect 3359 8585 3534 8722
tri 3534 8585 3671 8722 sw
tri 3772 8585 3909 8722 ne
rect 3909 8585 4084 8722
tri 4084 8585 4221 8722 sw
tri 4322 8585 4459 8722 ne
rect 4459 8585 4634 8722
tri 4634 8585 4771 8722 sw
tri 4872 8585 5009 8722 ne
rect 5009 8585 5184 8722
tri 5184 8585 5321 8722 sw
tri 5422 8585 5559 8722 ne
rect 5559 8585 5734 8722
tri 5734 8585 5871 8722 sw
tri 5972 8585 6109 8722 ne
rect 6109 8585 6284 8722
tri 6284 8585 6421 8722 sw
tri 6522 8585 6659 8722 ne
rect 6659 8585 6834 8722
tri 6834 8585 6971 8722 sw
tri 7072 8585 7209 8722 ne
rect 7209 8585 7384 8722
tri 7384 8585 7521 8722 sw
tri 7622 8585 7759 8722 ne
rect 7759 8585 7934 8722
tri 7934 8585 8071 8722 sw
tri 8172 8585 8309 8722 ne
rect 8309 8585 8484 8722
tri 8484 8585 8621 8722 sw
tri 8722 8585 8859 8722 ne
rect 8859 8585 9034 8722
tri 9034 8585 9171 8722 sw
tri 9272 8585 9409 8722 ne
rect 9409 8585 9584 8722
tri 9584 8585 9721 8722 sw
tri 9822 8585 9959 8722 ne
rect 9959 8585 10134 8722
tri 10134 8585 10271 8722 sw
tri 10372 8585 10509 8722 ne
rect 10509 8585 10684 8722
tri 10684 8585 10821 8722 sw
tri 10922 8585 11059 8722 ne
rect 11059 8585 11234 8722
tri 11234 8585 11371 8722 sw
tri 11472 8585 11609 8722 ne
rect 11609 8585 11784 8722
tri 11784 8585 11921 8722 sw
tri 12022 8585 12159 8722 ne
rect 12159 8585 12334 8722
tri 12334 8585 12471 8722 sw
tri 12572 8585 12709 8722 ne
rect 12709 8585 12884 8722
tri 12884 8585 13021 8722 sw
tri 13122 8585 13259 8722 ne
rect 13259 8585 13434 8722
tri 13434 8585 13571 8722 sw
tri 13672 8585 13809 8722 ne
rect 13809 8585 13984 8722
tri 13984 8585 14121 8722 sw
tri 14222 8585 14359 8722 ne
rect 14359 8585 14534 8722
tri 14534 8585 14671 8722 sw
tri 14772 8585 14909 8722 ne
rect 14909 8585 15084 8722
tri 15084 8585 15221 8722 sw
tri 15322 8585 15459 8722 ne
rect 15459 8585 15634 8722
tri 15634 8585 15771 8722 sw
tri 15872 8585 16009 8722 ne
rect 16009 8585 16184 8722
tri 16184 8585 16321 8722 sw
tri 16422 8585 16559 8722 ne
rect 16559 8585 16734 8722
tri 16734 8585 16871 8722 sw
tri 16972 8585 17109 8722 ne
rect 17109 8585 17284 8722
tri 17284 8585 17421 8722 sw
tri 17522 8585 17659 8722 ne
rect 17659 8585 17834 8722
tri 17834 8585 17971 8722 sw
tri 18072 8585 18209 8722 ne
rect 18209 8585 18384 8722
tri 18384 8585 18521 8722 sw
tri 18622 8585 18759 8722 ne
rect 18759 8585 18934 8722
tri 18934 8585 19071 8722 sw
tri 19172 8585 19309 8722 ne
rect 19309 8585 19484 8722
tri 19484 8585 19621 8722 sw
rect -2000 8567 215 8585
rect -2000 7778 -1000 8567
tri 77 8465 179 8567 ne
rect 179 8465 215 8567
rect 335 8465 371 8585
tri 179 8328 316 8465 ne
rect 316 8410 371 8465
tri 371 8410 546 8585 sw
tri 609 8465 729 8585 ne
rect 729 8465 765 8585
rect 885 8465 921 8585
rect 316 8328 546 8410
tri 546 8328 628 8410 sw
tri 729 8328 866 8465 ne
rect 866 8410 921 8465
tri 921 8410 1096 8585 sw
tri 1159 8465 1279 8585 ne
rect 1279 8465 1315 8585
rect 1435 8465 1471 8585
rect 866 8328 1096 8410
tri 1096 8328 1178 8410 sw
tri 1279 8328 1416 8465 ne
rect 1416 8410 1471 8465
tri 1471 8410 1646 8585 sw
tri 1709 8465 1829 8585 ne
rect 1829 8465 1865 8585
rect 1985 8465 2021 8585
rect 1416 8328 1646 8410
tri 1646 8328 1728 8410 sw
tri 1829 8328 1966 8465 ne
rect 1966 8410 2021 8465
tri 2021 8410 2196 8585 sw
tri 2259 8465 2379 8585 ne
rect 2379 8465 2415 8585
rect 2535 8465 2571 8585
rect 1966 8328 2196 8410
tri 2196 8328 2278 8410 sw
tri 2379 8328 2516 8465 ne
rect 2516 8410 2571 8465
tri 2571 8410 2746 8585 sw
tri 2809 8465 2929 8585 ne
rect 2929 8465 2965 8585
rect 3085 8465 3121 8585
rect 2516 8328 2746 8410
tri 2746 8328 2828 8410 sw
tri 2929 8328 3066 8465 ne
rect 3066 8410 3121 8465
tri 3121 8410 3296 8585 sw
tri 3359 8465 3479 8585 ne
rect 3479 8465 3515 8585
rect 3635 8465 3671 8585
rect 3066 8328 3296 8410
tri 3296 8328 3378 8410 sw
tri 3479 8328 3616 8465 ne
rect 3616 8410 3671 8465
tri 3671 8410 3846 8585 sw
tri 3909 8465 4029 8585 ne
rect 4029 8465 4065 8585
rect 4185 8465 4221 8585
rect 3616 8328 3846 8410
tri 3846 8328 3928 8410 sw
tri 4029 8328 4166 8465 ne
rect 4166 8410 4221 8465
tri 4221 8410 4396 8585 sw
tri 4459 8465 4579 8585 ne
rect 4579 8465 4615 8585
rect 4735 8465 4771 8585
rect 4166 8328 4396 8410
tri 4396 8328 4478 8410 sw
tri 4579 8328 4716 8465 ne
rect 4716 8410 4771 8465
tri 4771 8410 4946 8585 sw
tri 5009 8465 5129 8585 ne
rect 5129 8465 5165 8585
rect 5285 8465 5321 8585
rect 4716 8328 4946 8410
tri 4946 8328 5028 8410 sw
tri 5129 8328 5266 8465 ne
rect 5266 8410 5321 8465
tri 5321 8410 5496 8585 sw
tri 5559 8465 5679 8585 ne
rect 5679 8465 5715 8585
rect 5835 8465 5871 8585
rect 5266 8328 5496 8410
tri 5496 8328 5578 8410 sw
tri 5679 8328 5816 8465 ne
rect 5816 8410 5871 8465
tri 5871 8410 6046 8585 sw
tri 6109 8465 6229 8585 ne
rect 6229 8465 6265 8585
rect 6385 8465 6421 8585
rect 5816 8328 6046 8410
tri 6046 8328 6128 8410 sw
tri 6229 8328 6366 8465 ne
rect 6366 8410 6421 8465
tri 6421 8410 6596 8585 sw
tri 6659 8465 6779 8585 ne
rect 6779 8465 6815 8585
rect 6935 8465 6971 8585
rect 6366 8328 6596 8410
tri 6596 8328 6678 8410 sw
tri 6779 8328 6916 8465 ne
rect 6916 8410 6971 8465
tri 6971 8410 7146 8585 sw
tri 7209 8465 7329 8585 ne
rect 7329 8465 7365 8585
rect 7485 8465 7521 8585
rect 6916 8328 7146 8410
tri 7146 8328 7228 8410 sw
tri 7329 8328 7466 8465 ne
rect 7466 8410 7521 8465
tri 7521 8410 7696 8585 sw
tri 7759 8465 7879 8585 ne
rect 7879 8465 7915 8585
rect 8035 8465 8071 8585
rect 7466 8328 7696 8410
tri 7696 8328 7778 8410 sw
tri 7879 8328 8016 8465 ne
rect 8016 8410 8071 8465
tri 8071 8410 8246 8585 sw
tri 8309 8465 8429 8585 ne
rect 8429 8465 8465 8585
rect 8585 8465 8621 8585
rect 8016 8328 8246 8410
tri 8246 8328 8328 8410 sw
tri 8429 8328 8566 8465 ne
rect 8566 8410 8621 8465
tri 8621 8410 8796 8585 sw
tri 8859 8465 8979 8585 ne
rect 8979 8465 9015 8585
rect 9135 8465 9171 8585
rect 8566 8328 8796 8410
tri 8796 8328 8878 8410 sw
tri 8979 8328 9116 8465 ne
rect 9116 8410 9171 8465
tri 9171 8410 9346 8585 sw
tri 9409 8465 9529 8585 ne
rect 9529 8465 9565 8585
rect 9685 8465 9721 8585
rect 9116 8328 9346 8410
tri 9346 8328 9428 8410 sw
tri 9529 8328 9666 8465 ne
rect 9666 8410 9721 8465
tri 9721 8410 9896 8585 sw
tri 9959 8465 10079 8585 ne
rect 10079 8465 10115 8585
rect 10235 8465 10271 8585
rect 9666 8328 9896 8410
tri 9896 8328 9978 8410 sw
tri 10079 8328 10216 8465 ne
rect 10216 8410 10271 8465
tri 10271 8410 10446 8585 sw
tri 10509 8465 10629 8585 ne
rect 10629 8465 10665 8585
rect 10785 8465 10821 8585
rect 10216 8328 10446 8410
tri 10446 8328 10528 8410 sw
tri 10629 8328 10766 8465 ne
rect 10766 8410 10821 8465
tri 10821 8410 10996 8585 sw
tri 11059 8465 11179 8585 ne
rect 11179 8465 11215 8585
rect 11335 8465 11371 8585
rect 10766 8328 10996 8410
tri 10996 8328 11078 8410 sw
tri 11179 8328 11316 8465 ne
rect 11316 8410 11371 8465
tri 11371 8410 11546 8585 sw
tri 11609 8465 11729 8585 ne
rect 11729 8465 11765 8585
rect 11885 8465 11921 8585
rect 11316 8328 11546 8410
tri 11546 8328 11628 8410 sw
tri 11729 8328 11866 8465 ne
rect 11866 8410 11921 8465
tri 11921 8410 12096 8585 sw
tri 12159 8465 12279 8585 ne
rect 12279 8465 12315 8585
rect 12435 8465 12471 8585
rect 11866 8328 12096 8410
tri 12096 8328 12178 8410 sw
tri 12279 8328 12416 8465 ne
rect 12416 8410 12471 8465
tri 12471 8410 12646 8585 sw
tri 12709 8465 12829 8585 ne
rect 12829 8465 12865 8585
rect 12985 8465 13021 8585
rect 12416 8328 12646 8410
tri 12646 8328 12728 8410 sw
tri 12829 8328 12966 8465 ne
rect 12966 8410 13021 8465
tri 13021 8410 13196 8585 sw
tri 13259 8465 13379 8585 ne
rect 13379 8465 13415 8585
rect 13535 8465 13571 8585
rect 12966 8328 13196 8410
tri 13196 8328 13278 8410 sw
tri 13379 8328 13516 8465 ne
rect 13516 8410 13571 8465
tri 13571 8410 13746 8585 sw
tri 13809 8465 13929 8585 ne
rect 13929 8465 13965 8585
rect 14085 8465 14121 8585
rect 13516 8328 13746 8410
tri 13746 8328 13828 8410 sw
tri 13929 8328 14066 8465 ne
rect 14066 8410 14121 8465
tri 14121 8410 14296 8585 sw
tri 14359 8465 14479 8585 ne
rect 14479 8465 14515 8585
rect 14635 8465 14671 8585
rect 14066 8328 14296 8410
tri 14296 8328 14378 8410 sw
tri 14479 8328 14616 8465 ne
rect 14616 8410 14671 8465
tri 14671 8410 14846 8585 sw
tri 14909 8465 15029 8585 ne
rect 15029 8465 15065 8585
rect 15185 8465 15221 8585
rect 14616 8328 14846 8410
tri 14846 8328 14928 8410 sw
tri 15029 8328 15166 8465 ne
rect 15166 8410 15221 8465
tri 15221 8410 15396 8585 sw
tri 15459 8465 15579 8585 ne
rect 15579 8465 15615 8585
rect 15735 8465 15771 8585
rect 15166 8328 15396 8410
tri 15396 8328 15478 8410 sw
tri 15579 8328 15716 8465 ne
rect 15716 8410 15771 8465
tri 15771 8410 15946 8585 sw
tri 16009 8465 16129 8585 ne
rect 16129 8465 16165 8585
rect 16285 8465 16321 8585
rect 15716 8328 15946 8410
tri 15946 8328 16028 8410 sw
tri 16129 8328 16266 8465 ne
rect 16266 8410 16321 8465
tri 16321 8410 16496 8585 sw
tri 16559 8465 16679 8585 ne
rect 16679 8465 16715 8585
rect 16835 8465 16871 8585
rect 16266 8328 16496 8410
tri 16496 8328 16578 8410 sw
tri 16679 8328 16816 8465 ne
rect 16816 8410 16871 8465
tri 16871 8410 17046 8585 sw
tri 17109 8465 17229 8585 ne
rect 17229 8465 17265 8585
rect 17385 8465 17421 8585
rect 16816 8328 17046 8410
tri 17046 8328 17128 8410 sw
tri 17229 8328 17366 8465 ne
rect 17366 8410 17421 8465
tri 17421 8410 17596 8585 sw
tri 17659 8465 17779 8585 ne
rect 17779 8465 17815 8585
rect 17935 8465 17971 8585
rect 17366 8328 17596 8410
tri 17596 8328 17678 8410 sw
tri 17779 8328 17916 8465 ne
rect 17916 8410 17971 8465
tri 17971 8410 18146 8585 sw
tri 18209 8465 18329 8585 ne
rect 18329 8465 18365 8585
rect 18485 8465 18521 8585
rect 17916 8328 18146 8410
tri 18146 8328 18228 8410 sw
tri 18329 8328 18466 8465 ne
rect 18466 8410 18521 8465
tri 18521 8410 18696 8585 sw
tri 18759 8465 18879 8585 ne
rect 18879 8465 18915 8585
rect 19035 8465 19071 8585
rect 18466 8328 18696 8410
tri 18696 8328 18778 8410 sw
tri 18879 8328 19016 8465 ne
rect 19016 8410 19071 8465
tri 19071 8410 19246 8585 sw
tri 19309 8465 19429 8585 ne
rect 19429 8465 19465 8585
rect 19585 8483 19621 8585
tri 19621 8483 19723 8585 sw
rect 20800 8483 21800 9272
rect 19585 8465 21800 8483
rect 19016 8328 19246 8410
tri 19246 8328 19328 8410 sw
tri 19429 8328 19566 8465 ne
rect 19566 8328 21800 8465
rect -500 8172 78 8328
tri 78 8172 234 8328 sw
tri 316 8172 472 8328 ne
rect 472 8172 628 8328
tri 628 8172 784 8328 sw
tri 866 8172 1022 8328 ne
rect 1022 8172 1178 8328
tri 1178 8172 1334 8328 sw
tri 1416 8172 1572 8328 ne
rect 1572 8172 1728 8328
tri 1728 8172 1884 8328 sw
tri 1966 8172 2122 8328 ne
rect 2122 8172 2278 8328
tri 2278 8172 2434 8328 sw
tri 2516 8172 2672 8328 ne
rect 2672 8172 2828 8328
tri 2828 8172 2984 8328 sw
tri 3066 8172 3222 8328 ne
rect 3222 8172 3378 8328
tri 3378 8172 3534 8328 sw
tri 3616 8172 3772 8328 ne
rect 3772 8172 3928 8328
tri 3928 8172 4084 8328 sw
tri 4166 8172 4322 8328 ne
rect 4322 8172 4478 8328
tri 4478 8172 4634 8328 sw
tri 4716 8172 4872 8328 ne
rect 4872 8172 5028 8328
tri 5028 8172 5184 8328 sw
tri 5266 8172 5422 8328 ne
rect 5422 8172 5578 8328
tri 5578 8172 5734 8328 sw
tri 5816 8172 5972 8328 ne
rect 5972 8172 6128 8328
tri 6128 8172 6284 8328 sw
tri 6366 8172 6522 8328 ne
rect 6522 8172 6678 8328
tri 6678 8172 6834 8328 sw
tri 6916 8172 7072 8328 ne
rect 7072 8172 7228 8328
tri 7228 8172 7384 8328 sw
tri 7466 8172 7622 8328 ne
rect 7622 8172 7778 8328
tri 7778 8172 7934 8328 sw
tri 8016 8172 8172 8328 ne
rect 8172 8172 8328 8328
tri 8328 8172 8484 8328 sw
tri 8566 8172 8722 8328 ne
rect 8722 8172 8878 8328
tri 8878 8172 9034 8328 sw
tri 9116 8172 9272 8328 ne
rect 9272 8172 9428 8328
tri 9428 8172 9584 8328 sw
tri 9666 8172 9822 8328 ne
rect 9822 8172 9978 8328
tri 9978 8172 10134 8328 sw
tri 10216 8172 10372 8328 ne
rect 10372 8172 10528 8328
tri 10528 8172 10684 8328 sw
tri 10766 8172 10922 8328 ne
rect 10922 8172 11078 8328
tri 11078 8172 11234 8328 sw
tri 11316 8172 11472 8328 ne
rect 11472 8172 11628 8328
tri 11628 8172 11784 8328 sw
tri 11866 8172 12022 8328 ne
rect 12022 8172 12178 8328
tri 12178 8172 12334 8328 sw
tri 12416 8172 12572 8328 ne
rect 12572 8172 12728 8328
tri 12728 8172 12884 8328 sw
tri 12966 8172 13122 8328 ne
rect 13122 8172 13278 8328
tri 13278 8172 13434 8328 sw
tri 13516 8172 13672 8328 ne
rect 13672 8172 13828 8328
tri 13828 8172 13984 8328 sw
tri 14066 8172 14222 8328 ne
rect 14222 8172 14378 8328
tri 14378 8172 14534 8328 sw
tri 14616 8172 14772 8328 ne
rect 14772 8172 14928 8328
tri 14928 8172 15084 8328 sw
tri 15166 8172 15322 8328 ne
rect 15322 8172 15478 8328
tri 15478 8172 15634 8328 sw
tri 15716 8172 15872 8328 ne
rect 15872 8172 16028 8328
tri 16028 8172 16184 8328 sw
tri 16266 8172 16422 8328 ne
rect 16422 8172 16578 8328
tri 16578 8172 16734 8328 sw
tri 16816 8172 16972 8328 ne
rect 16972 8172 17128 8328
tri 17128 8172 17284 8328 sw
tri 17366 8172 17522 8328 ne
rect 17522 8172 17678 8328
tri 17678 8172 17834 8328 sw
tri 17916 8172 18072 8328 ne
rect 18072 8172 18228 8328
tri 18228 8172 18384 8328 sw
tri 18466 8172 18622 8328 ne
rect 18622 8172 18778 8328
tri 18778 8172 18934 8328 sw
tri 19016 8172 19172 8328 ne
rect 19172 8172 19328 8328
tri 19328 8172 19484 8328 sw
tri 19566 8172 19722 8328 ne
rect 19722 8172 21800 8328
rect -500 8035 234 8172
tri 234 8035 371 8172 sw
tri 472 8035 609 8172 ne
rect 609 8035 784 8172
tri 784 8035 921 8172 sw
tri 1022 8035 1159 8172 ne
rect 1159 8035 1334 8172
tri 1334 8035 1471 8172 sw
tri 1572 8035 1709 8172 ne
rect 1709 8035 1884 8172
tri 1884 8035 2021 8172 sw
tri 2122 8035 2259 8172 ne
rect 2259 8035 2434 8172
tri 2434 8035 2571 8172 sw
tri 2672 8035 2809 8172 ne
rect 2809 8035 2984 8172
tri 2984 8035 3121 8172 sw
tri 3222 8035 3359 8172 ne
rect 3359 8035 3534 8172
tri 3534 8035 3671 8172 sw
tri 3772 8035 3909 8172 ne
rect 3909 8035 4084 8172
tri 4084 8035 4221 8172 sw
tri 4322 8035 4459 8172 ne
rect 4459 8035 4634 8172
tri 4634 8035 4771 8172 sw
tri 4872 8035 5009 8172 ne
rect 5009 8035 5184 8172
tri 5184 8035 5321 8172 sw
tri 5422 8035 5559 8172 ne
rect 5559 8035 5734 8172
tri 5734 8035 5871 8172 sw
tri 5972 8035 6109 8172 ne
rect 6109 8035 6284 8172
tri 6284 8035 6421 8172 sw
tri 6522 8035 6659 8172 ne
rect 6659 8035 6834 8172
tri 6834 8035 6971 8172 sw
tri 7072 8035 7209 8172 ne
rect 7209 8035 7384 8172
tri 7384 8035 7521 8172 sw
tri 7622 8035 7759 8172 ne
rect 7759 8035 7934 8172
tri 7934 8035 8071 8172 sw
tri 8172 8035 8309 8172 ne
rect 8309 8035 8484 8172
tri 8484 8035 8621 8172 sw
tri 8722 8035 8859 8172 ne
rect 8859 8035 9034 8172
tri 9034 8035 9171 8172 sw
tri 9272 8035 9409 8172 ne
rect 9409 8035 9584 8172
tri 9584 8035 9721 8172 sw
tri 9822 8035 9959 8172 ne
rect 9959 8035 10134 8172
tri 10134 8035 10271 8172 sw
tri 10372 8035 10509 8172 ne
rect 10509 8035 10684 8172
tri 10684 8035 10821 8172 sw
tri 10922 8035 11059 8172 ne
rect 11059 8035 11234 8172
tri 11234 8035 11371 8172 sw
tri 11472 8035 11609 8172 ne
rect 11609 8035 11784 8172
tri 11784 8035 11921 8172 sw
tri 12022 8035 12159 8172 ne
rect 12159 8035 12334 8172
tri 12334 8035 12471 8172 sw
tri 12572 8035 12709 8172 ne
rect 12709 8035 12884 8172
tri 12884 8035 13021 8172 sw
tri 13122 8035 13259 8172 ne
rect 13259 8035 13434 8172
tri 13434 8035 13571 8172 sw
tri 13672 8035 13809 8172 ne
rect 13809 8035 13984 8172
tri 13984 8035 14121 8172 sw
tri 14222 8035 14359 8172 ne
rect 14359 8035 14534 8172
tri 14534 8035 14671 8172 sw
tri 14772 8035 14909 8172 ne
rect 14909 8035 15084 8172
tri 15084 8035 15221 8172 sw
tri 15322 8035 15459 8172 ne
rect 15459 8035 15634 8172
tri 15634 8035 15771 8172 sw
tri 15872 8035 16009 8172 ne
rect 16009 8035 16184 8172
tri 16184 8035 16321 8172 sw
tri 16422 8035 16559 8172 ne
rect 16559 8035 16734 8172
tri 16734 8035 16871 8172 sw
tri 16972 8035 17109 8172 ne
rect 17109 8035 17284 8172
tri 17284 8035 17421 8172 sw
tri 17522 8035 17659 8172 ne
rect 17659 8035 17834 8172
tri 17834 8035 17971 8172 sw
tri 18072 8035 18209 8172 ne
rect 18209 8035 18384 8172
tri 18384 8035 18521 8172 sw
tri 18622 8035 18759 8172 ne
rect 18759 8035 18934 8172
tri 18934 8035 19071 8172 sw
tri 19172 8035 19309 8172 ne
rect 19309 8035 19484 8172
tri 19484 8035 19621 8172 sw
rect -500 8017 215 8035
tri 77 7915 179 8017 ne
rect 179 7915 215 8017
rect 335 7915 371 8035
tri 179 7778 316 7915 ne
rect 316 7860 371 7915
tri 371 7860 546 8035 sw
tri 609 7915 729 8035 ne
rect 729 7915 765 8035
rect 885 7915 921 8035
rect 316 7778 546 7860
tri 546 7778 628 7860 sw
tri 729 7778 866 7915 ne
rect 866 7860 921 7915
tri 921 7860 1096 8035 sw
tri 1159 7915 1279 8035 ne
rect 1279 7915 1315 8035
rect 1435 7915 1471 8035
rect 866 7778 1096 7860
tri 1096 7778 1178 7860 sw
tri 1279 7778 1416 7915 ne
rect 1416 7860 1471 7915
tri 1471 7860 1646 8035 sw
tri 1709 7915 1829 8035 ne
rect 1829 7915 1865 8035
rect 1985 7915 2021 8035
rect 1416 7778 1646 7860
tri 1646 7778 1728 7860 sw
tri 1829 7778 1966 7915 ne
rect 1966 7860 2021 7915
tri 2021 7860 2196 8035 sw
tri 2259 7915 2379 8035 ne
rect 2379 7915 2415 8035
rect 2535 7915 2571 8035
rect 1966 7778 2196 7860
tri 2196 7778 2278 7860 sw
tri 2379 7778 2516 7915 ne
rect 2516 7860 2571 7915
tri 2571 7860 2746 8035 sw
tri 2809 7915 2929 8035 ne
rect 2929 7915 2965 8035
rect 3085 7915 3121 8035
rect 2516 7778 2746 7860
tri 2746 7778 2828 7860 sw
tri 2929 7778 3066 7915 ne
rect 3066 7860 3121 7915
tri 3121 7860 3296 8035 sw
tri 3359 7915 3479 8035 ne
rect 3479 7915 3515 8035
rect 3635 7915 3671 8035
rect 3066 7778 3296 7860
tri 3296 7778 3378 7860 sw
tri 3479 7778 3616 7915 ne
rect 3616 7860 3671 7915
tri 3671 7860 3846 8035 sw
tri 3909 7915 4029 8035 ne
rect 4029 7915 4065 8035
rect 4185 7915 4221 8035
rect 3616 7778 3846 7860
tri 3846 7778 3928 7860 sw
tri 4029 7778 4166 7915 ne
rect 4166 7860 4221 7915
tri 4221 7860 4396 8035 sw
tri 4459 7915 4579 8035 ne
rect 4579 7915 4615 8035
rect 4735 7915 4771 8035
rect 4166 7778 4396 7860
tri 4396 7778 4478 7860 sw
tri 4579 7778 4716 7915 ne
rect 4716 7860 4771 7915
tri 4771 7860 4946 8035 sw
tri 5009 7915 5129 8035 ne
rect 5129 7915 5165 8035
rect 5285 7915 5321 8035
rect 4716 7778 4946 7860
tri 4946 7778 5028 7860 sw
tri 5129 7778 5266 7915 ne
rect 5266 7860 5321 7915
tri 5321 7860 5496 8035 sw
tri 5559 7915 5679 8035 ne
rect 5679 7915 5715 8035
rect 5835 7915 5871 8035
rect 5266 7778 5496 7860
tri 5496 7778 5578 7860 sw
tri 5679 7778 5816 7915 ne
rect 5816 7860 5871 7915
tri 5871 7860 6046 8035 sw
tri 6109 7915 6229 8035 ne
rect 6229 7915 6265 8035
rect 6385 7915 6421 8035
rect 5816 7778 6046 7860
tri 6046 7778 6128 7860 sw
tri 6229 7778 6366 7915 ne
rect 6366 7860 6421 7915
tri 6421 7860 6596 8035 sw
tri 6659 7915 6779 8035 ne
rect 6779 7915 6815 8035
rect 6935 7915 6971 8035
rect 6366 7778 6596 7860
tri 6596 7778 6678 7860 sw
tri 6779 7778 6916 7915 ne
rect 6916 7860 6971 7915
tri 6971 7860 7146 8035 sw
tri 7209 7915 7329 8035 ne
rect 7329 7915 7365 8035
rect 7485 7915 7521 8035
rect 6916 7778 7146 7860
tri 7146 7778 7228 7860 sw
tri 7329 7778 7466 7915 ne
rect 7466 7860 7521 7915
tri 7521 7860 7696 8035 sw
tri 7759 7915 7879 8035 ne
rect 7879 7915 7915 8035
rect 8035 7915 8071 8035
rect 7466 7778 7696 7860
tri 7696 7778 7778 7860 sw
tri 7879 7778 8016 7915 ne
rect 8016 7860 8071 7915
tri 8071 7860 8246 8035 sw
tri 8309 7915 8429 8035 ne
rect 8429 7915 8465 8035
rect 8585 7915 8621 8035
rect 8016 7778 8246 7860
tri 8246 7778 8328 7860 sw
tri 8429 7778 8566 7915 ne
rect 8566 7860 8621 7915
tri 8621 7860 8796 8035 sw
tri 8859 7915 8979 8035 ne
rect 8979 7915 9015 8035
rect 9135 7915 9171 8035
rect 8566 7778 8796 7860
tri 8796 7778 8878 7860 sw
tri 8979 7778 9116 7915 ne
rect 9116 7860 9171 7915
tri 9171 7860 9346 8035 sw
tri 9409 7915 9529 8035 ne
rect 9529 7915 9565 8035
rect 9685 7915 9721 8035
rect 9116 7778 9346 7860
tri 9346 7778 9428 7860 sw
tri 9529 7778 9666 7915 ne
rect 9666 7860 9721 7915
tri 9721 7860 9896 8035 sw
tri 9959 7915 10079 8035 ne
rect 10079 7915 10115 8035
rect 10235 7915 10271 8035
rect 9666 7778 9896 7860
tri 9896 7778 9978 7860 sw
tri 10079 7778 10216 7915 ne
rect 10216 7860 10271 7915
tri 10271 7860 10446 8035 sw
tri 10509 7915 10629 8035 ne
rect 10629 7915 10665 8035
rect 10785 7915 10821 8035
rect 10216 7778 10446 7860
tri 10446 7778 10528 7860 sw
tri 10629 7778 10766 7915 ne
rect 10766 7860 10821 7915
tri 10821 7860 10996 8035 sw
tri 11059 7915 11179 8035 ne
rect 11179 7915 11215 8035
rect 11335 7915 11371 8035
rect 10766 7778 10996 7860
tri 10996 7778 11078 7860 sw
tri 11179 7778 11316 7915 ne
rect 11316 7860 11371 7915
tri 11371 7860 11546 8035 sw
tri 11609 7915 11729 8035 ne
rect 11729 7915 11765 8035
rect 11885 7915 11921 8035
rect 11316 7778 11546 7860
tri 11546 7778 11628 7860 sw
tri 11729 7778 11866 7915 ne
rect 11866 7860 11921 7915
tri 11921 7860 12096 8035 sw
tri 12159 7915 12279 8035 ne
rect 12279 7915 12315 8035
rect 12435 7915 12471 8035
rect 11866 7778 12096 7860
tri 12096 7778 12178 7860 sw
tri 12279 7778 12416 7915 ne
rect 12416 7860 12471 7915
tri 12471 7860 12646 8035 sw
tri 12709 7915 12829 8035 ne
rect 12829 7915 12865 8035
rect 12985 7915 13021 8035
rect 12416 7778 12646 7860
tri 12646 7778 12728 7860 sw
tri 12829 7778 12966 7915 ne
rect 12966 7860 13021 7915
tri 13021 7860 13196 8035 sw
tri 13259 7915 13379 8035 ne
rect 13379 7915 13415 8035
rect 13535 7915 13571 8035
rect 12966 7778 13196 7860
tri 13196 7778 13278 7860 sw
tri 13379 7778 13516 7915 ne
rect 13516 7860 13571 7915
tri 13571 7860 13746 8035 sw
tri 13809 7915 13929 8035 ne
rect 13929 7915 13965 8035
rect 14085 7915 14121 8035
rect 13516 7778 13746 7860
tri 13746 7778 13828 7860 sw
tri 13929 7778 14066 7915 ne
rect 14066 7860 14121 7915
tri 14121 7860 14296 8035 sw
tri 14359 7915 14479 8035 ne
rect 14479 7915 14515 8035
rect 14635 7915 14671 8035
rect 14066 7778 14296 7860
tri 14296 7778 14378 7860 sw
tri 14479 7778 14616 7915 ne
rect 14616 7860 14671 7915
tri 14671 7860 14846 8035 sw
tri 14909 7915 15029 8035 ne
rect 15029 7915 15065 8035
rect 15185 7915 15221 8035
rect 14616 7778 14846 7860
tri 14846 7778 14928 7860 sw
tri 15029 7778 15166 7915 ne
rect 15166 7860 15221 7915
tri 15221 7860 15396 8035 sw
tri 15459 7915 15579 8035 ne
rect 15579 7915 15615 8035
rect 15735 7915 15771 8035
rect 15166 7778 15396 7860
tri 15396 7778 15478 7860 sw
tri 15579 7778 15716 7915 ne
rect 15716 7860 15771 7915
tri 15771 7860 15946 8035 sw
tri 16009 7915 16129 8035 ne
rect 16129 7915 16165 8035
rect 16285 7915 16321 8035
rect 15716 7778 15946 7860
tri 15946 7778 16028 7860 sw
tri 16129 7778 16266 7915 ne
rect 16266 7860 16321 7915
tri 16321 7860 16496 8035 sw
tri 16559 7915 16679 8035 ne
rect 16679 7915 16715 8035
rect 16835 7915 16871 8035
rect 16266 7778 16496 7860
tri 16496 7778 16578 7860 sw
tri 16679 7778 16816 7915 ne
rect 16816 7860 16871 7915
tri 16871 7860 17046 8035 sw
tri 17109 7915 17229 8035 ne
rect 17229 7915 17265 8035
rect 17385 7915 17421 8035
rect 16816 7778 17046 7860
tri 17046 7778 17128 7860 sw
tri 17229 7778 17366 7915 ne
rect 17366 7860 17421 7915
tri 17421 7860 17596 8035 sw
tri 17659 7915 17779 8035 ne
rect 17779 7915 17815 8035
rect 17935 7915 17971 8035
rect 17366 7778 17596 7860
tri 17596 7778 17678 7860 sw
tri 17779 7778 17916 7915 ne
rect 17916 7860 17971 7915
tri 17971 7860 18146 8035 sw
tri 18209 7915 18329 8035 ne
rect 18329 7915 18365 8035
rect 18485 7915 18521 8035
rect 17916 7778 18146 7860
tri 18146 7778 18228 7860 sw
tri 18329 7778 18466 7915 ne
rect 18466 7860 18521 7915
tri 18521 7860 18696 8035 sw
tri 18759 7915 18879 8035 ne
rect 18879 7915 18915 8035
rect 19035 7915 19071 8035
rect 18466 7778 18696 7860
tri 18696 7778 18778 7860 sw
tri 18879 7778 19016 7915 ne
rect 19016 7860 19071 7915
tri 19071 7860 19246 8035 sw
tri 19309 7915 19429 8035 ne
rect 19429 7915 19465 8035
rect 19585 7933 19621 8035
tri 19621 7933 19723 8035 sw
rect 19585 7915 20300 7933
rect 19016 7778 19246 7860
tri 19246 7778 19328 7860 sw
tri 19429 7778 19566 7915 ne
rect 19566 7778 20300 7915
rect -2000 7622 78 7778
tri 78 7622 234 7778 sw
tri 316 7622 472 7778 ne
rect 472 7622 628 7778
tri 628 7622 784 7778 sw
tri 866 7622 1022 7778 ne
rect 1022 7622 1178 7778
tri 1178 7622 1334 7778 sw
tri 1416 7622 1572 7778 ne
rect 1572 7622 1728 7778
tri 1728 7622 1884 7778 sw
tri 1966 7622 2122 7778 ne
rect 2122 7622 2278 7778
tri 2278 7622 2434 7778 sw
tri 2516 7622 2672 7778 ne
rect 2672 7622 2828 7778
tri 2828 7622 2984 7778 sw
tri 3066 7622 3222 7778 ne
rect 3222 7622 3378 7778
tri 3378 7622 3534 7778 sw
tri 3616 7622 3772 7778 ne
rect 3772 7622 3928 7778
tri 3928 7622 4084 7778 sw
tri 4166 7622 4322 7778 ne
rect 4322 7622 4478 7778
tri 4478 7622 4634 7778 sw
tri 4716 7622 4872 7778 ne
rect 4872 7622 5028 7778
tri 5028 7622 5184 7778 sw
tri 5266 7622 5422 7778 ne
rect 5422 7622 5578 7778
tri 5578 7622 5734 7778 sw
tri 5816 7622 5972 7778 ne
rect 5972 7622 6128 7778
tri 6128 7622 6284 7778 sw
tri 6366 7622 6522 7778 ne
rect 6522 7622 6678 7778
tri 6678 7622 6834 7778 sw
tri 6916 7622 7072 7778 ne
rect 7072 7622 7228 7778
tri 7228 7622 7384 7778 sw
tri 7466 7622 7622 7778 ne
rect 7622 7622 7778 7778
tri 7778 7622 7934 7778 sw
tri 8016 7622 8172 7778 ne
rect 8172 7622 8328 7778
tri 8328 7622 8484 7778 sw
tri 8566 7622 8722 7778 ne
rect 8722 7622 8878 7778
tri 8878 7622 9034 7778 sw
tri 9116 7622 9272 7778 ne
rect 9272 7622 9428 7778
tri 9428 7622 9584 7778 sw
tri 9666 7622 9822 7778 ne
rect 9822 7622 9978 7778
tri 9978 7622 10134 7778 sw
tri 10216 7622 10372 7778 ne
rect 10372 7622 10528 7778
tri 10528 7622 10684 7778 sw
tri 10766 7622 10922 7778 ne
rect 10922 7622 11078 7778
tri 11078 7622 11234 7778 sw
tri 11316 7622 11472 7778 ne
rect 11472 7622 11628 7778
tri 11628 7622 11784 7778 sw
tri 11866 7622 12022 7778 ne
rect 12022 7622 12178 7778
tri 12178 7622 12334 7778 sw
tri 12416 7622 12572 7778 ne
rect 12572 7622 12728 7778
tri 12728 7622 12884 7778 sw
tri 12966 7622 13122 7778 ne
rect 13122 7622 13278 7778
tri 13278 7622 13434 7778 sw
tri 13516 7622 13672 7778 ne
rect 13672 7622 13828 7778
tri 13828 7622 13984 7778 sw
tri 14066 7622 14222 7778 ne
rect 14222 7622 14378 7778
tri 14378 7622 14534 7778 sw
tri 14616 7622 14772 7778 ne
rect 14772 7622 14928 7778
tri 14928 7622 15084 7778 sw
tri 15166 7622 15322 7778 ne
rect 15322 7622 15478 7778
tri 15478 7622 15634 7778 sw
tri 15716 7622 15872 7778 ne
rect 15872 7622 16028 7778
tri 16028 7622 16184 7778 sw
tri 16266 7622 16422 7778 ne
rect 16422 7622 16578 7778
tri 16578 7622 16734 7778 sw
tri 16816 7622 16972 7778 ne
rect 16972 7622 17128 7778
tri 17128 7622 17284 7778 sw
tri 17366 7622 17522 7778 ne
rect 17522 7622 17678 7778
tri 17678 7622 17834 7778 sw
tri 17916 7622 18072 7778 ne
rect 18072 7622 18228 7778
tri 18228 7622 18384 7778 sw
tri 18466 7622 18622 7778 ne
rect 18622 7622 18778 7778
tri 18778 7622 18934 7778 sw
tri 19016 7622 19172 7778 ne
rect 19172 7622 19328 7778
tri 19328 7622 19484 7778 sw
tri 19566 7622 19722 7778 ne
rect 19722 7622 20300 7778
rect -2000 7485 234 7622
tri 234 7485 371 7622 sw
tri 472 7485 609 7622 ne
rect 609 7485 784 7622
tri 784 7485 921 7622 sw
tri 1022 7485 1159 7622 ne
rect 1159 7485 1334 7622
tri 1334 7485 1471 7622 sw
tri 1572 7485 1709 7622 ne
rect 1709 7485 1884 7622
tri 1884 7485 2021 7622 sw
tri 2122 7485 2259 7622 ne
rect 2259 7485 2434 7622
tri 2434 7485 2571 7622 sw
tri 2672 7485 2809 7622 ne
rect 2809 7485 2984 7622
tri 2984 7485 3121 7622 sw
tri 3222 7485 3359 7622 ne
rect 3359 7485 3534 7622
tri 3534 7485 3671 7622 sw
tri 3772 7485 3909 7622 ne
rect 3909 7485 4084 7622
tri 4084 7485 4221 7622 sw
tri 4322 7485 4459 7622 ne
rect 4459 7485 4634 7622
tri 4634 7485 4771 7622 sw
tri 4872 7485 5009 7622 ne
rect 5009 7485 5184 7622
tri 5184 7485 5321 7622 sw
tri 5422 7485 5559 7622 ne
rect 5559 7485 5734 7622
tri 5734 7485 5871 7622 sw
tri 5972 7485 6109 7622 ne
rect 6109 7485 6284 7622
tri 6284 7485 6421 7622 sw
tri 6522 7485 6659 7622 ne
rect 6659 7485 6834 7622
tri 6834 7485 6971 7622 sw
tri 7072 7485 7209 7622 ne
rect 7209 7485 7384 7622
tri 7384 7485 7521 7622 sw
tri 7622 7485 7759 7622 ne
rect 7759 7485 7934 7622
tri 7934 7485 8071 7622 sw
tri 8172 7485 8309 7622 ne
rect 8309 7485 8484 7622
tri 8484 7485 8621 7622 sw
tri 8722 7485 8859 7622 ne
rect 8859 7485 9034 7622
tri 9034 7485 9171 7622 sw
tri 9272 7485 9409 7622 ne
rect 9409 7485 9584 7622
tri 9584 7485 9721 7622 sw
tri 9822 7485 9959 7622 ne
rect 9959 7485 10134 7622
tri 10134 7485 10271 7622 sw
tri 10372 7485 10509 7622 ne
rect 10509 7485 10684 7622
tri 10684 7485 10821 7622 sw
tri 10922 7485 11059 7622 ne
rect 11059 7485 11234 7622
tri 11234 7485 11371 7622 sw
tri 11472 7485 11609 7622 ne
rect 11609 7485 11784 7622
tri 11784 7485 11921 7622 sw
tri 12022 7485 12159 7622 ne
rect 12159 7485 12334 7622
tri 12334 7485 12471 7622 sw
tri 12572 7485 12709 7622 ne
rect 12709 7485 12884 7622
tri 12884 7485 13021 7622 sw
tri 13122 7485 13259 7622 ne
rect 13259 7485 13434 7622
tri 13434 7485 13571 7622 sw
tri 13672 7485 13809 7622 ne
rect 13809 7485 13984 7622
tri 13984 7485 14121 7622 sw
tri 14222 7485 14359 7622 ne
rect 14359 7485 14534 7622
tri 14534 7485 14671 7622 sw
tri 14772 7485 14909 7622 ne
rect 14909 7485 15084 7622
tri 15084 7485 15221 7622 sw
tri 15322 7485 15459 7622 ne
rect 15459 7485 15634 7622
tri 15634 7485 15771 7622 sw
tri 15872 7485 16009 7622 ne
rect 16009 7485 16184 7622
tri 16184 7485 16321 7622 sw
tri 16422 7485 16559 7622 ne
rect 16559 7485 16734 7622
tri 16734 7485 16871 7622 sw
tri 16972 7485 17109 7622 ne
rect 17109 7485 17284 7622
tri 17284 7485 17421 7622 sw
tri 17522 7485 17659 7622 ne
rect 17659 7485 17834 7622
tri 17834 7485 17971 7622 sw
tri 18072 7485 18209 7622 ne
rect 18209 7485 18384 7622
tri 18384 7485 18521 7622 sw
tri 18622 7485 18759 7622 ne
rect 18759 7485 18934 7622
tri 18934 7485 19071 7622 sw
tri 19172 7485 19309 7622 ne
rect 19309 7485 19484 7622
tri 19484 7485 19621 7622 sw
rect -2000 7467 215 7485
rect -2000 6678 -1000 7467
tri 77 7365 179 7467 ne
rect 179 7365 215 7467
rect 335 7365 371 7485
tri 179 7228 316 7365 ne
rect 316 7310 371 7365
tri 371 7310 546 7485 sw
tri 609 7365 729 7485 ne
rect 729 7365 765 7485
rect 885 7365 921 7485
rect 316 7228 546 7310
tri 546 7228 628 7310 sw
tri 729 7228 866 7365 ne
rect 866 7310 921 7365
tri 921 7310 1096 7485 sw
tri 1159 7365 1279 7485 ne
rect 1279 7365 1315 7485
rect 1435 7365 1471 7485
rect 866 7228 1096 7310
tri 1096 7228 1178 7310 sw
tri 1279 7228 1416 7365 ne
rect 1416 7310 1471 7365
tri 1471 7310 1646 7485 sw
tri 1709 7365 1829 7485 ne
rect 1829 7365 1865 7485
rect 1985 7365 2021 7485
rect 1416 7228 1646 7310
tri 1646 7228 1728 7310 sw
tri 1829 7228 1966 7365 ne
rect 1966 7310 2021 7365
tri 2021 7310 2196 7485 sw
tri 2259 7365 2379 7485 ne
rect 2379 7365 2415 7485
rect 2535 7365 2571 7485
rect 1966 7228 2196 7310
tri 2196 7228 2278 7310 sw
tri 2379 7228 2516 7365 ne
rect 2516 7310 2571 7365
tri 2571 7310 2746 7485 sw
tri 2809 7365 2929 7485 ne
rect 2929 7365 2965 7485
rect 3085 7365 3121 7485
rect 2516 7228 2746 7310
tri 2746 7228 2828 7310 sw
tri 2929 7228 3066 7365 ne
rect 3066 7310 3121 7365
tri 3121 7310 3296 7485 sw
tri 3359 7365 3479 7485 ne
rect 3479 7365 3515 7485
rect 3635 7365 3671 7485
rect 3066 7228 3296 7310
tri 3296 7228 3378 7310 sw
tri 3479 7228 3616 7365 ne
rect 3616 7310 3671 7365
tri 3671 7310 3846 7485 sw
tri 3909 7365 4029 7485 ne
rect 4029 7365 4065 7485
rect 4185 7365 4221 7485
rect 3616 7228 3846 7310
tri 3846 7228 3928 7310 sw
tri 4029 7228 4166 7365 ne
rect 4166 7310 4221 7365
tri 4221 7310 4396 7485 sw
tri 4459 7365 4579 7485 ne
rect 4579 7365 4615 7485
rect 4735 7365 4771 7485
rect 4166 7228 4396 7310
tri 4396 7228 4478 7310 sw
tri 4579 7228 4716 7365 ne
rect 4716 7310 4771 7365
tri 4771 7310 4946 7485 sw
tri 5009 7365 5129 7485 ne
rect 5129 7365 5165 7485
rect 5285 7365 5321 7485
rect 4716 7228 4946 7310
tri 4946 7228 5028 7310 sw
tri 5129 7228 5266 7365 ne
rect 5266 7310 5321 7365
tri 5321 7310 5496 7485 sw
tri 5559 7365 5679 7485 ne
rect 5679 7365 5715 7485
rect 5835 7365 5871 7485
rect 5266 7228 5496 7310
tri 5496 7228 5578 7310 sw
tri 5679 7228 5816 7365 ne
rect 5816 7310 5871 7365
tri 5871 7310 6046 7485 sw
tri 6109 7365 6229 7485 ne
rect 6229 7365 6265 7485
rect 6385 7365 6421 7485
rect 5816 7228 6046 7310
tri 6046 7228 6128 7310 sw
tri 6229 7228 6366 7365 ne
rect 6366 7310 6421 7365
tri 6421 7310 6596 7485 sw
tri 6659 7365 6779 7485 ne
rect 6779 7365 6815 7485
rect 6935 7365 6971 7485
rect 6366 7228 6596 7310
tri 6596 7228 6678 7310 sw
tri 6779 7228 6916 7365 ne
rect 6916 7310 6971 7365
tri 6971 7310 7146 7485 sw
tri 7209 7365 7329 7485 ne
rect 7329 7365 7365 7485
rect 7485 7365 7521 7485
rect 6916 7228 7146 7310
tri 7146 7228 7228 7310 sw
tri 7329 7228 7466 7365 ne
rect 7466 7310 7521 7365
tri 7521 7310 7696 7485 sw
tri 7759 7365 7879 7485 ne
rect 7879 7365 7915 7485
rect 8035 7365 8071 7485
rect 7466 7228 7696 7310
tri 7696 7228 7778 7310 sw
tri 7879 7228 8016 7365 ne
rect 8016 7310 8071 7365
tri 8071 7310 8246 7485 sw
tri 8309 7365 8429 7485 ne
rect 8429 7365 8465 7485
rect 8585 7365 8621 7485
rect 8016 7228 8246 7310
tri 8246 7228 8328 7310 sw
tri 8429 7228 8566 7365 ne
rect 8566 7310 8621 7365
tri 8621 7310 8796 7485 sw
tri 8859 7365 8979 7485 ne
rect 8979 7365 9015 7485
rect 9135 7365 9171 7485
rect 8566 7228 8796 7310
tri 8796 7228 8878 7310 sw
tri 8979 7228 9116 7365 ne
rect 9116 7310 9171 7365
tri 9171 7310 9346 7485 sw
tri 9409 7365 9529 7485 ne
rect 9529 7365 9565 7485
rect 9685 7365 9721 7485
rect 9116 7228 9346 7310
tri 9346 7228 9428 7310 sw
tri 9529 7228 9666 7365 ne
rect 9666 7310 9721 7365
tri 9721 7310 9896 7485 sw
tri 9959 7365 10079 7485 ne
rect 10079 7365 10115 7485
rect 10235 7365 10271 7485
rect 9666 7228 9896 7310
tri 9896 7228 9978 7310 sw
tri 10079 7228 10216 7365 ne
rect 10216 7310 10271 7365
tri 10271 7310 10446 7485 sw
tri 10509 7365 10629 7485 ne
rect 10629 7365 10665 7485
rect 10785 7365 10821 7485
rect 10216 7228 10446 7310
tri 10446 7228 10528 7310 sw
tri 10629 7228 10766 7365 ne
rect 10766 7310 10821 7365
tri 10821 7310 10996 7485 sw
tri 11059 7365 11179 7485 ne
rect 11179 7365 11215 7485
rect 11335 7365 11371 7485
rect 10766 7228 10996 7310
tri 10996 7228 11078 7310 sw
tri 11179 7228 11316 7365 ne
rect 11316 7310 11371 7365
tri 11371 7310 11546 7485 sw
tri 11609 7365 11729 7485 ne
rect 11729 7365 11765 7485
rect 11885 7365 11921 7485
rect 11316 7228 11546 7310
tri 11546 7228 11628 7310 sw
tri 11729 7228 11866 7365 ne
rect 11866 7310 11921 7365
tri 11921 7310 12096 7485 sw
tri 12159 7365 12279 7485 ne
rect 12279 7365 12315 7485
rect 12435 7365 12471 7485
rect 11866 7228 12096 7310
tri 12096 7228 12178 7310 sw
tri 12279 7228 12416 7365 ne
rect 12416 7310 12471 7365
tri 12471 7310 12646 7485 sw
tri 12709 7365 12829 7485 ne
rect 12829 7365 12865 7485
rect 12985 7365 13021 7485
rect 12416 7228 12646 7310
tri 12646 7228 12728 7310 sw
tri 12829 7228 12966 7365 ne
rect 12966 7310 13021 7365
tri 13021 7310 13196 7485 sw
tri 13259 7365 13379 7485 ne
rect 13379 7365 13415 7485
rect 13535 7365 13571 7485
rect 12966 7228 13196 7310
tri 13196 7228 13278 7310 sw
tri 13379 7228 13516 7365 ne
rect 13516 7310 13571 7365
tri 13571 7310 13746 7485 sw
tri 13809 7365 13929 7485 ne
rect 13929 7365 13965 7485
rect 14085 7365 14121 7485
rect 13516 7228 13746 7310
tri 13746 7228 13828 7310 sw
tri 13929 7228 14066 7365 ne
rect 14066 7310 14121 7365
tri 14121 7310 14296 7485 sw
tri 14359 7365 14479 7485 ne
rect 14479 7365 14515 7485
rect 14635 7365 14671 7485
rect 14066 7228 14296 7310
tri 14296 7228 14378 7310 sw
tri 14479 7228 14616 7365 ne
rect 14616 7310 14671 7365
tri 14671 7310 14846 7485 sw
tri 14909 7365 15029 7485 ne
rect 15029 7365 15065 7485
rect 15185 7365 15221 7485
rect 14616 7228 14846 7310
tri 14846 7228 14928 7310 sw
tri 15029 7228 15166 7365 ne
rect 15166 7310 15221 7365
tri 15221 7310 15396 7485 sw
tri 15459 7365 15579 7485 ne
rect 15579 7365 15615 7485
rect 15735 7365 15771 7485
rect 15166 7228 15396 7310
tri 15396 7228 15478 7310 sw
tri 15579 7228 15716 7365 ne
rect 15716 7310 15771 7365
tri 15771 7310 15946 7485 sw
tri 16009 7365 16129 7485 ne
rect 16129 7365 16165 7485
rect 16285 7365 16321 7485
rect 15716 7228 15946 7310
tri 15946 7228 16028 7310 sw
tri 16129 7228 16266 7365 ne
rect 16266 7310 16321 7365
tri 16321 7310 16496 7485 sw
tri 16559 7365 16679 7485 ne
rect 16679 7365 16715 7485
rect 16835 7365 16871 7485
rect 16266 7228 16496 7310
tri 16496 7228 16578 7310 sw
tri 16679 7228 16816 7365 ne
rect 16816 7310 16871 7365
tri 16871 7310 17046 7485 sw
tri 17109 7365 17229 7485 ne
rect 17229 7365 17265 7485
rect 17385 7365 17421 7485
rect 16816 7228 17046 7310
tri 17046 7228 17128 7310 sw
tri 17229 7228 17366 7365 ne
rect 17366 7310 17421 7365
tri 17421 7310 17596 7485 sw
tri 17659 7365 17779 7485 ne
rect 17779 7365 17815 7485
rect 17935 7365 17971 7485
rect 17366 7228 17596 7310
tri 17596 7228 17678 7310 sw
tri 17779 7228 17916 7365 ne
rect 17916 7310 17971 7365
tri 17971 7310 18146 7485 sw
tri 18209 7365 18329 7485 ne
rect 18329 7365 18365 7485
rect 18485 7365 18521 7485
rect 17916 7228 18146 7310
tri 18146 7228 18228 7310 sw
tri 18329 7228 18466 7365 ne
rect 18466 7310 18521 7365
tri 18521 7310 18696 7485 sw
tri 18759 7365 18879 7485 ne
rect 18879 7365 18915 7485
rect 19035 7365 19071 7485
rect 18466 7228 18696 7310
tri 18696 7228 18778 7310 sw
tri 18879 7228 19016 7365 ne
rect 19016 7310 19071 7365
tri 19071 7310 19246 7485 sw
tri 19309 7365 19429 7485 ne
rect 19429 7365 19465 7485
rect 19585 7383 19621 7485
tri 19621 7383 19723 7485 sw
rect 20800 7383 21800 8172
rect 19585 7365 21800 7383
rect 19016 7228 19246 7310
tri 19246 7228 19328 7310 sw
tri 19429 7228 19566 7365 ne
rect 19566 7228 21800 7365
rect -500 7072 78 7228
tri 78 7072 234 7228 sw
tri 316 7072 472 7228 ne
rect 472 7072 628 7228
tri 628 7072 784 7228 sw
tri 866 7072 1022 7228 ne
rect 1022 7072 1178 7228
tri 1178 7072 1334 7228 sw
tri 1416 7072 1572 7228 ne
rect 1572 7072 1728 7228
tri 1728 7072 1884 7228 sw
tri 1966 7072 2122 7228 ne
rect 2122 7072 2278 7228
tri 2278 7072 2434 7228 sw
tri 2516 7072 2672 7228 ne
rect 2672 7072 2828 7228
tri 2828 7072 2984 7228 sw
tri 3066 7072 3222 7228 ne
rect 3222 7072 3378 7228
tri 3378 7072 3534 7228 sw
tri 3616 7072 3772 7228 ne
rect 3772 7072 3928 7228
tri 3928 7072 4084 7228 sw
tri 4166 7072 4322 7228 ne
rect 4322 7072 4478 7228
tri 4478 7072 4634 7228 sw
tri 4716 7072 4872 7228 ne
rect 4872 7072 5028 7228
tri 5028 7072 5184 7228 sw
tri 5266 7072 5422 7228 ne
rect 5422 7072 5578 7228
tri 5578 7072 5734 7228 sw
tri 5816 7072 5972 7228 ne
rect 5972 7072 6128 7228
tri 6128 7072 6284 7228 sw
tri 6366 7072 6522 7228 ne
rect 6522 7072 6678 7228
tri 6678 7072 6834 7228 sw
tri 6916 7072 7072 7228 ne
rect 7072 7072 7228 7228
tri 7228 7072 7384 7228 sw
tri 7466 7072 7622 7228 ne
rect 7622 7072 7778 7228
tri 7778 7072 7934 7228 sw
tri 8016 7072 8172 7228 ne
rect 8172 7072 8328 7228
tri 8328 7072 8484 7228 sw
tri 8566 7072 8722 7228 ne
rect 8722 7072 8878 7228
tri 8878 7072 9034 7228 sw
tri 9116 7072 9272 7228 ne
rect 9272 7072 9428 7228
tri 9428 7072 9584 7228 sw
tri 9666 7072 9822 7228 ne
rect 9822 7072 9978 7228
tri 9978 7072 10134 7228 sw
tri 10216 7072 10372 7228 ne
rect 10372 7072 10528 7228
tri 10528 7072 10684 7228 sw
tri 10766 7072 10922 7228 ne
rect 10922 7072 11078 7228
tri 11078 7072 11234 7228 sw
tri 11316 7072 11472 7228 ne
rect 11472 7072 11628 7228
tri 11628 7072 11784 7228 sw
tri 11866 7072 12022 7228 ne
rect 12022 7072 12178 7228
tri 12178 7072 12334 7228 sw
tri 12416 7072 12572 7228 ne
rect 12572 7072 12728 7228
tri 12728 7072 12884 7228 sw
tri 12966 7072 13122 7228 ne
rect 13122 7072 13278 7228
tri 13278 7072 13434 7228 sw
tri 13516 7072 13672 7228 ne
rect 13672 7072 13828 7228
tri 13828 7072 13984 7228 sw
tri 14066 7072 14222 7228 ne
rect 14222 7072 14378 7228
tri 14378 7072 14534 7228 sw
tri 14616 7072 14772 7228 ne
rect 14772 7072 14928 7228
tri 14928 7072 15084 7228 sw
tri 15166 7072 15322 7228 ne
rect 15322 7072 15478 7228
tri 15478 7072 15634 7228 sw
tri 15716 7072 15872 7228 ne
rect 15872 7072 16028 7228
tri 16028 7072 16184 7228 sw
tri 16266 7072 16422 7228 ne
rect 16422 7072 16578 7228
tri 16578 7072 16734 7228 sw
tri 16816 7072 16972 7228 ne
rect 16972 7072 17128 7228
tri 17128 7072 17284 7228 sw
tri 17366 7072 17522 7228 ne
rect 17522 7072 17678 7228
tri 17678 7072 17834 7228 sw
tri 17916 7072 18072 7228 ne
rect 18072 7072 18228 7228
tri 18228 7072 18384 7228 sw
tri 18466 7072 18622 7228 ne
rect 18622 7072 18778 7228
tri 18778 7072 18934 7228 sw
tri 19016 7072 19172 7228 ne
rect 19172 7072 19328 7228
tri 19328 7072 19484 7228 sw
tri 19566 7072 19722 7228 ne
rect 19722 7072 21800 7228
rect -500 6935 234 7072
tri 234 6935 371 7072 sw
tri 472 6935 609 7072 ne
rect 609 6935 784 7072
tri 784 6935 921 7072 sw
tri 1022 6935 1159 7072 ne
rect 1159 6935 1334 7072
tri 1334 6935 1471 7072 sw
tri 1572 6935 1709 7072 ne
rect 1709 6935 1884 7072
tri 1884 6935 2021 7072 sw
tri 2122 6935 2259 7072 ne
rect 2259 6935 2434 7072
tri 2434 6935 2571 7072 sw
tri 2672 6935 2809 7072 ne
rect 2809 6935 2984 7072
tri 2984 6935 3121 7072 sw
tri 3222 6935 3359 7072 ne
rect 3359 6935 3534 7072
tri 3534 6935 3671 7072 sw
tri 3772 6935 3909 7072 ne
rect 3909 6935 4084 7072
tri 4084 6935 4221 7072 sw
tri 4322 6935 4459 7072 ne
rect 4459 6935 4634 7072
tri 4634 6935 4771 7072 sw
tri 4872 6935 5009 7072 ne
rect 5009 6935 5184 7072
tri 5184 6935 5321 7072 sw
tri 5422 6935 5559 7072 ne
rect 5559 6935 5734 7072
tri 5734 6935 5871 7072 sw
tri 5972 6935 6109 7072 ne
rect 6109 6935 6284 7072
tri 6284 6935 6421 7072 sw
tri 6522 6935 6659 7072 ne
rect 6659 6935 6834 7072
tri 6834 6935 6971 7072 sw
tri 7072 6935 7209 7072 ne
rect 7209 6935 7384 7072
tri 7384 6935 7521 7072 sw
tri 7622 6935 7759 7072 ne
rect 7759 6935 7934 7072
tri 7934 6935 8071 7072 sw
tri 8172 6935 8309 7072 ne
rect 8309 6935 8484 7072
tri 8484 6935 8621 7072 sw
tri 8722 6935 8859 7072 ne
rect 8859 6935 9034 7072
tri 9034 6935 9171 7072 sw
tri 9272 6935 9409 7072 ne
rect 9409 6935 9584 7072
tri 9584 6935 9721 7072 sw
tri 9822 6935 9959 7072 ne
rect 9959 6935 10134 7072
tri 10134 6935 10271 7072 sw
tri 10372 6935 10509 7072 ne
rect 10509 6935 10684 7072
tri 10684 6935 10821 7072 sw
tri 10922 6935 11059 7072 ne
rect 11059 6935 11234 7072
tri 11234 6935 11371 7072 sw
tri 11472 6935 11609 7072 ne
rect 11609 6935 11784 7072
tri 11784 6935 11921 7072 sw
tri 12022 6935 12159 7072 ne
rect 12159 6935 12334 7072
tri 12334 6935 12471 7072 sw
tri 12572 6935 12709 7072 ne
rect 12709 6935 12884 7072
tri 12884 6935 13021 7072 sw
tri 13122 6935 13259 7072 ne
rect 13259 6935 13434 7072
tri 13434 6935 13571 7072 sw
tri 13672 6935 13809 7072 ne
rect 13809 6935 13984 7072
tri 13984 6935 14121 7072 sw
tri 14222 6935 14359 7072 ne
rect 14359 6935 14534 7072
tri 14534 6935 14671 7072 sw
tri 14772 6935 14909 7072 ne
rect 14909 6935 15084 7072
tri 15084 6935 15221 7072 sw
tri 15322 6935 15459 7072 ne
rect 15459 6935 15634 7072
tri 15634 6935 15771 7072 sw
tri 15872 6935 16009 7072 ne
rect 16009 6935 16184 7072
tri 16184 6935 16321 7072 sw
tri 16422 6935 16559 7072 ne
rect 16559 6935 16734 7072
tri 16734 6935 16871 7072 sw
tri 16972 6935 17109 7072 ne
rect 17109 6935 17284 7072
tri 17284 6935 17421 7072 sw
tri 17522 6935 17659 7072 ne
rect 17659 6935 17834 7072
tri 17834 6935 17971 7072 sw
tri 18072 6935 18209 7072 ne
rect 18209 6935 18384 7072
tri 18384 6935 18521 7072 sw
tri 18622 6935 18759 7072 ne
rect 18759 6935 18934 7072
tri 18934 6935 19071 7072 sw
tri 19172 6935 19309 7072 ne
rect 19309 6935 19484 7072
tri 19484 6935 19621 7072 sw
rect -500 6917 215 6935
tri 77 6815 179 6917 ne
rect 179 6815 215 6917
rect 335 6815 371 6935
tri 179 6678 316 6815 ne
rect 316 6760 371 6815
tri 371 6760 546 6935 sw
tri 609 6815 729 6935 ne
rect 729 6815 765 6935
rect 885 6815 921 6935
rect 316 6678 546 6760
tri 546 6678 628 6760 sw
tri 729 6678 866 6815 ne
rect 866 6760 921 6815
tri 921 6760 1096 6935 sw
tri 1159 6815 1279 6935 ne
rect 1279 6815 1315 6935
rect 1435 6815 1471 6935
rect 866 6678 1096 6760
tri 1096 6678 1178 6760 sw
tri 1279 6678 1416 6815 ne
rect 1416 6760 1471 6815
tri 1471 6760 1646 6935 sw
tri 1709 6815 1829 6935 ne
rect 1829 6815 1865 6935
rect 1985 6815 2021 6935
rect 1416 6678 1646 6760
tri 1646 6678 1728 6760 sw
tri 1829 6678 1966 6815 ne
rect 1966 6760 2021 6815
tri 2021 6760 2196 6935 sw
tri 2259 6815 2379 6935 ne
rect 2379 6815 2415 6935
rect 2535 6815 2571 6935
rect 1966 6678 2196 6760
tri 2196 6678 2278 6760 sw
tri 2379 6678 2516 6815 ne
rect 2516 6760 2571 6815
tri 2571 6760 2746 6935 sw
tri 2809 6815 2929 6935 ne
rect 2929 6815 2965 6935
rect 3085 6815 3121 6935
rect 2516 6678 2746 6760
tri 2746 6678 2828 6760 sw
tri 2929 6678 3066 6815 ne
rect 3066 6760 3121 6815
tri 3121 6760 3296 6935 sw
tri 3359 6815 3479 6935 ne
rect 3479 6815 3515 6935
rect 3635 6815 3671 6935
rect 3066 6678 3296 6760
tri 3296 6678 3378 6760 sw
tri 3479 6678 3616 6815 ne
rect 3616 6760 3671 6815
tri 3671 6760 3846 6935 sw
tri 3909 6815 4029 6935 ne
rect 4029 6815 4065 6935
rect 4185 6815 4221 6935
rect 3616 6678 3846 6760
tri 3846 6678 3928 6760 sw
tri 4029 6678 4166 6815 ne
rect 4166 6760 4221 6815
tri 4221 6760 4396 6935 sw
tri 4459 6815 4579 6935 ne
rect 4579 6815 4615 6935
rect 4735 6815 4771 6935
rect 4166 6678 4396 6760
tri 4396 6678 4478 6760 sw
tri 4579 6678 4716 6815 ne
rect 4716 6760 4771 6815
tri 4771 6760 4946 6935 sw
tri 5009 6815 5129 6935 ne
rect 5129 6815 5165 6935
rect 5285 6815 5321 6935
rect 4716 6678 4946 6760
tri 4946 6678 5028 6760 sw
tri 5129 6678 5266 6815 ne
rect 5266 6760 5321 6815
tri 5321 6760 5496 6935 sw
tri 5559 6815 5679 6935 ne
rect 5679 6815 5715 6935
rect 5835 6815 5871 6935
rect 5266 6678 5496 6760
tri 5496 6678 5578 6760 sw
tri 5679 6678 5816 6815 ne
rect 5816 6760 5871 6815
tri 5871 6760 6046 6935 sw
tri 6109 6815 6229 6935 ne
rect 6229 6815 6265 6935
rect 6385 6815 6421 6935
rect 5816 6678 6046 6760
tri 6046 6678 6128 6760 sw
tri 6229 6678 6366 6815 ne
rect 6366 6760 6421 6815
tri 6421 6760 6596 6935 sw
tri 6659 6815 6779 6935 ne
rect 6779 6815 6815 6935
rect 6935 6815 6971 6935
rect 6366 6678 6596 6760
tri 6596 6678 6678 6760 sw
tri 6779 6678 6916 6815 ne
rect 6916 6760 6971 6815
tri 6971 6760 7146 6935 sw
tri 7209 6815 7329 6935 ne
rect 7329 6815 7365 6935
rect 7485 6815 7521 6935
rect 6916 6678 7146 6760
tri 7146 6678 7228 6760 sw
tri 7329 6678 7466 6815 ne
rect 7466 6760 7521 6815
tri 7521 6760 7696 6935 sw
tri 7759 6815 7879 6935 ne
rect 7879 6815 7915 6935
rect 8035 6815 8071 6935
rect 7466 6678 7696 6760
tri 7696 6678 7778 6760 sw
tri 7879 6678 8016 6815 ne
rect 8016 6760 8071 6815
tri 8071 6760 8246 6935 sw
tri 8309 6815 8429 6935 ne
rect 8429 6815 8465 6935
rect 8585 6815 8621 6935
rect 8016 6678 8246 6760
tri 8246 6678 8328 6760 sw
tri 8429 6678 8566 6815 ne
rect 8566 6760 8621 6815
tri 8621 6760 8796 6935 sw
tri 8859 6815 8979 6935 ne
rect 8979 6815 9015 6935
rect 9135 6815 9171 6935
rect 8566 6678 8796 6760
tri 8796 6678 8878 6760 sw
tri 8979 6678 9116 6815 ne
rect 9116 6760 9171 6815
tri 9171 6760 9346 6935 sw
tri 9409 6815 9529 6935 ne
rect 9529 6815 9565 6935
rect 9685 6815 9721 6935
rect 9116 6678 9346 6760
tri 9346 6678 9428 6760 sw
tri 9529 6678 9666 6815 ne
rect 9666 6760 9721 6815
tri 9721 6760 9896 6935 sw
tri 9959 6815 10079 6935 ne
rect 10079 6815 10115 6935
rect 10235 6815 10271 6935
rect 9666 6678 9896 6760
tri 9896 6678 9978 6760 sw
tri 10079 6678 10216 6815 ne
rect 10216 6760 10271 6815
tri 10271 6760 10446 6935 sw
tri 10509 6815 10629 6935 ne
rect 10629 6815 10665 6935
rect 10785 6815 10821 6935
rect 10216 6678 10446 6760
tri 10446 6678 10528 6760 sw
tri 10629 6678 10766 6815 ne
rect 10766 6760 10821 6815
tri 10821 6760 10996 6935 sw
tri 11059 6815 11179 6935 ne
rect 11179 6815 11215 6935
rect 11335 6815 11371 6935
rect 10766 6678 10996 6760
tri 10996 6678 11078 6760 sw
tri 11179 6678 11316 6815 ne
rect 11316 6760 11371 6815
tri 11371 6760 11546 6935 sw
tri 11609 6815 11729 6935 ne
rect 11729 6815 11765 6935
rect 11885 6815 11921 6935
rect 11316 6678 11546 6760
tri 11546 6678 11628 6760 sw
tri 11729 6678 11866 6815 ne
rect 11866 6760 11921 6815
tri 11921 6760 12096 6935 sw
tri 12159 6815 12279 6935 ne
rect 12279 6815 12315 6935
rect 12435 6815 12471 6935
rect 11866 6678 12096 6760
tri 12096 6678 12178 6760 sw
tri 12279 6678 12416 6815 ne
rect 12416 6760 12471 6815
tri 12471 6760 12646 6935 sw
tri 12709 6815 12829 6935 ne
rect 12829 6815 12865 6935
rect 12985 6815 13021 6935
rect 12416 6678 12646 6760
tri 12646 6678 12728 6760 sw
tri 12829 6678 12966 6815 ne
rect 12966 6760 13021 6815
tri 13021 6760 13196 6935 sw
tri 13259 6815 13379 6935 ne
rect 13379 6815 13415 6935
rect 13535 6815 13571 6935
rect 12966 6678 13196 6760
tri 13196 6678 13278 6760 sw
tri 13379 6678 13516 6815 ne
rect 13516 6760 13571 6815
tri 13571 6760 13746 6935 sw
tri 13809 6815 13929 6935 ne
rect 13929 6815 13965 6935
rect 14085 6815 14121 6935
rect 13516 6678 13746 6760
tri 13746 6678 13828 6760 sw
tri 13929 6678 14066 6815 ne
rect 14066 6760 14121 6815
tri 14121 6760 14296 6935 sw
tri 14359 6815 14479 6935 ne
rect 14479 6815 14515 6935
rect 14635 6815 14671 6935
rect 14066 6678 14296 6760
tri 14296 6678 14378 6760 sw
tri 14479 6678 14616 6815 ne
rect 14616 6760 14671 6815
tri 14671 6760 14846 6935 sw
tri 14909 6815 15029 6935 ne
rect 15029 6815 15065 6935
rect 15185 6815 15221 6935
rect 14616 6678 14846 6760
tri 14846 6678 14928 6760 sw
tri 15029 6678 15166 6815 ne
rect 15166 6760 15221 6815
tri 15221 6760 15396 6935 sw
tri 15459 6815 15579 6935 ne
rect 15579 6815 15615 6935
rect 15735 6815 15771 6935
rect 15166 6678 15396 6760
tri 15396 6678 15478 6760 sw
tri 15579 6678 15716 6815 ne
rect 15716 6760 15771 6815
tri 15771 6760 15946 6935 sw
tri 16009 6815 16129 6935 ne
rect 16129 6815 16165 6935
rect 16285 6815 16321 6935
rect 15716 6678 15946 6760
tri 15946 6678 16028 6760 sw
tri 16129 6678 16266 6815 ne
rect 16266 6760 16321 6815
tri 16321 6760 16496 6935 sw
tri 16559 6815 16679 6935 ne
rect 16679 6815 16715 6935
rect 16835 6815 16871 6935
rect 16266 6678 16496 6760
tri 16496 6678 16578 6760 sw
tri 16679 6678 16816 6815 ne
rect 16816 6760 16871 6815
tri 16871 6760 17046 6935 sw
tri 17109 6815 17229 6935 ne
rect 17229 6815 17265 6935
rect 17385 6815 17421 6935
rect 16816 6678 17046 6760
tri 17046 6678 17128 6760 sw
tri 17229 6678 17366 6815 ne
rect 17366 6760 17421 6815
tri 17421 6760 17596 6935 sw
tri 17659 6815 17779 6935 ne
rect 17779 6815 17815 6935
rect 17935 6815 17971 6935
rect 17366 6678 17596 6760
tri 17596 6678 17678 6760 sw
tri 17779 6678 17916 6815 ne
rect 17916 6760 17971 6815
tri 17971 6760 18146 6935 sw
tri 18209 6815 18329 6935 ne
rect 18329 6815 18365 6935
rect 18485 6815 18521 6935
rect 17916 6678 18146 6760
tri 18146 6678 18228 6760 sw
tri 18329 6678 18466 6815 ne
rect 18466 6760 18521 6815
tri 18521 6760 18696 6935 sw
tri 18759 6815 18879 6935 ne
rect 18879 6815 18915 6935
rect 19035 6815 19071 6935
rect 18466 6678 18696 6760
tri 18696 6678 18778 6760 sw
tri 18879 6678 19016 6815 ne
rect 19016 6760 19071 6815
tri 19071 6760 19246 6935 sw
tri 19309 6815 19429 6935 ne
rect 19429 6815 19465 6935
rect 19585 6833 19621 6935
tri 19621 6833 19723 6935 sw
rect 19585 6815 20300 6833
rect 19016 6678 19246 6760
tri 19246 6678 19328 6760 sw
tri 19429 6678 19566 6815 ne
rect 19566 6678 20300 6815
rect -2000 6522 78 6678
tri 78 6522 234 6678 sw
tri 316 6522 472 6678 ne
rect 472 6522 628 6678
tri 628 6522 784 6678 sw
tri 866 6522 1022 6678 ne
rect 1022 6522 1178 6678
tri 1178 6522 1334 6678 sw
tri 1416 6522 1572 6678 ne
rect 1572 6522 1728 6678
tri 1728 6522 1884 6678 sw
tri 1966 6522 2122 6678 ne
rect 2122 6522 2278 6678
tri 2278 6522 2434 6678 sw
tri 2516 6522 2672 6678 ne
rect 2672 6522 2828 6678
tri 2828 6522 2984 6678 sw
tri 3066 6522 3222 6678 ne
rect 3222 6522 3378 6678
tri 3378 6522 3534 6678 sw
tri 3616 6522 3772 6678 ne
rect 3772 6522 3928 6678
tri 3928 6522 4084 6678 sw
tri 4166 6522 4322 6678 ne
rect 4322 6522 4478 6678
tri 4478 6522 4634 6678 sw
tri 4716 6522 4872 6678 ne
rect 4872 6522 5028 6678
tri 5028 6522 5184 6678 sw
tri 5266 6522 5422 6678 ne
rect 5422 6522 5578 6678
tri 5578 6522 5734 6678 sw
tri 5816 6522 5972 6678 ne
rect 5972 6522 6128 6678
tri 6128 6522 6284 6678 sw
tri 6366 6522 6522 6678 ne
rect 6522 6522 6678 6678
tri 6678 6522 6834 6678 sw
tri 6916 6522 7072 6678 ne
rect 7072 6522 7228 6678
tri 7228 6522 7384 6678 sw
tri 7466 6522 7622 6678 ne
rect 7622 6522 7778 6678
tri 7778 6522 7934 6678 sw
tri 8016 6522 8172 6678 ne
rect 8172 6522 8328 6678
tri 8328 6522 8484 6678 sw
tri 8566 6522 8722 6678 ne
rect 8722 6522 8878 6678
tri 8878 6522 9034 6678 sw
tri 9116 6522 9272 6678 ne
rect 9272 6522 9428 6678
tri 9428 6522 9584 6678 sw
tri 9666 6522 9822 6678 ne
rect 9822 6522 9978 6678
tri 9978 6522 10134 6678 sw
tri 10216 6522 10372 6678 ne
rect 10372 6522 10528 6678
tri 10528 6522 10684 6678 sw
tri 10766 6522 10922 6678 ne
rect 10922 6522 11078 6678
tri 11078 6522 11234 6678 sw
tri 11316 6522 11472 6678 ne
rect 11472 6522 11628 6678
tri 11628 6522 11784 6678 sw
tri 11866 6522 12022 6678 ne
rect 12022 6522 12178 6678
tri 12178 6522 12334 6678 sw
tri 12416 6522 12572 6678 ne
rect 12572 6522 12728 6678
tri 12728 6522 12884 6678 sw
tri 12966 6522 13122 6678 ne
rect 13122 6522 13278 6678
tri 13278 6522 13434 6678 sw
tri 13516 6522 13672 6678 ne
rect 13672 6522 13828 6678
tri 13828 6522 13984 6678 sw
tri 14066 6522 14222 6678 ne
rect 14222 6522 14378 6678
tri 14378 6522 14534 6678 sw
tri 14616 6522 14772 6678 ne
rect 14772 6522 14928 6678
tri 14928 6522 15084 6678 sw
tri 15166 6522 15322 6678 ne
rect 15322 6522 15478 6678
tri 15478 6522 15634 6678 sw
tri 15716 6522 15872 6678 ne
rect 15872 6522 16028 6678
tri 16028 6522 16184 6678 sw
tri 16266 6522 16422 6678 ne
rect 16422 6522 16578 6678
tri 16578 6522 16734 6678 sw
tri 16816 6522 16972 6678 ne
rect 16972 6522 17128 6678
tri 17128 6522 17284 6678 sw
tri 17366 6522 17522 6678 ne
rect 17522 6522 17678 6678
tri 17678 6522 17834 6678 sw
tri 17916 6522 18072 6678 ne
rect 18072 6522 18228 6678
tri 18228 6522 18384 6678 sw
tri 18466 6522 18622 6678 ne
rect 18622 6522 18778 6678
tri 18778 6522 18934 6678 sw
tri 19016 6522 19172 6678 ne
rect 19172 6522 19328 6678
tri 19328 6522 19484 6678 sw
tri 19566 6522 19722 6678 ne
rect 19722 6522 20300 6678
rect -2000 6385 234 6522
tri 234 6385 371 6522 sw
tri 472 6385 609 6522 ne
rect 609 6385 784 6522
tri 784 6385 921 6522 sw
tri 1022 6385 1159 6522 ne
rect 1159 6385 1334 6522
tri 1334 6385 1471 6522 sw
tri 1572 6385 1709 6522 ne
rect 1709 6385 1884 6522
tri 1884 6385 2021 6522 sw
tri 2122 6385 2259 6522 ne
rect 2259 6385 2434 6522
tri 2434 6385 2571 6522 sw
tri 2672 6385 2809 6522 ne
rect 2809 6385 2984 6522
tri 2984 6385 3121 6522 sw
tri 3222 6385 3359 6522 ne
rect 3359 6385 3534 6522
tri 3534 6385 3671 6522 sw
tri 3772 6385 3909 6522 ne
rect 3909 6385 4084 6522
tri 4084 6385 4221 6522 sw
tri 4322 6385 4459 6522 ne
rect 4459 6385 4634 6522
tri 4634 6385 4771 6522 sw
tri 4872 6385 5009 6522 ne
rect 5009 6385 5184 6522
tri 5184 6385 5321 6522 sw
tri 5422 6385 5559 6522 ne
rect 5559 6385 5734 6522
tri 5734 6385 5871 6522 sw
tri 5972 6385 6109 6522 ne
rect 6109 6385 6284 6522
tri 6284 6385 6421 6522 sw
tri 6522 6385 6659 6522 ne
rect 6659 6385 6834 6522
tri 6834 6385 6971 6522 sw
tri 7072 6385 7209 6522 ne
rect 7209 6385 7384 6522
tri 7384 6385 7521 6522 sw
tri 7622 6385 7759 6522 ne
rect 7759 6385 7934 6522
tri 7934 6385 8071 6522 sw
tri 8172 6385 8309 6522 ne
rect 8309 6385 8484 6522
tri 8484 6385 8621 6522 sw
tri 8722 6385 8859 6522 ne
rect 8859 6385 9034 6522
tri 9034 6385 9171 6522 sw
tri 9272 6385 9409 6522 ne
rect 9409 6385 9584 6522
tri 9584 6385 9721 6522 sw
tri 9822 6385 9959 6522 ne
rect 9959 6385 10134 6522
tri 10134 6385 10271 6522 sw
tri 10372 6385 10509 6522 ne
rect 10509 6385 10684 6522
tri 10684 6385 10821 6522 sw
tri 10922 6385 11059 6522 ne
rect 11059 6385 11234 6522
tri 11234 6385 11371 6522 sw
tri 11472 6385 11609 6522 ne
rect 11609 6385 11784 6522
tri 11784 6385 11921 6522 sw
tri 12022 6385 12159 6522 ne
rect 12159 6385 12334 6522
tri 12334 6385 12471 6522 sw
tri 12572 6385 12709 6522 ne
rect 12709 6385 12884 6522
tri 12884 6385 13021 6522 sw
tri 13122 6385 13259 6522 ne
rect 13259 6385 13434 6522
tri 13434 6385 13571 6522 sw
tri 13672 6385 13809 6522 ne
rect 13809 6385 13984 6522
tri 13984 6385 14121 6522 sw
tri 14222 6385 14359 6522 ne
rect 14359 6385 14534 6522
tri 14534 6385 14671 6522 sw
tri 14772 6385 14909 6522 ne
rect 14909 6385 15084 6522
tri 15084 6385 15221 6522 sw
tri 15322 6385 15459 6522 ne
rect 15459 6385 15634 6522
tri 15634 6385 15771 6522 sw
tri 15872 6385 16009 6522 ne
rect 16009 6385 16184 6522
tri 16184 6385 16321 6522 sw
tri 16422 6385 16559 6522 ne
rect 16559 6385 16734 6522
tri 16734 6385 16871 6522 sw
tri 16972 6385 17109 6522 ne
rect 17109 6385 17284 6522
tri 17284 6385 17421 6522 sw
tri 17522 6385 17659 6522 ne
rect 17659 6385 17834 6522
tri 17834 6385 17971 6522 sw
tri 18072 6385 18209 6522 ne
rect 18209 6385 18384 6522
tri 18384 6385 18521 6522 sw
tri 18622 6385 18759 6522 ne
rect 18759 6385 18934 6522
tri 18934 6385 19071 6522 sw
tri 19172 6385 19309 6522 ne
rect 19309 6385 19484 6522
tri 19484 6385 19621 6522 sw
rect -2000 6367 215 6385
rect -2000 5578 -1000 6367
tri 77 6265 179 6367 ne
rect 179 6265 215 6367
rect 335 6265 371 6385
tri 179 6128 316 6265 ne
rect 316 6210 371 6265
tri 371 6210 546 6385 sw
tri 609 6265 729 6385 ne
rect 729 6265 765 6385
rect 885 6265 921 6385
rect 316 6128 546 6210
tri 546 6128 628 6210 sw
tri 729 6128 866 6265 ne
rect 866 6210 921 6265
tri 921 6210 1096 6385 sw
tri 1159 6265 1279 6385 ne
rect 1279 6265 1315 6385
rect 1435 6265 1471 6385
rect 866 6128 1096 6210
tri 1096 6128 1178 6210 sw
tri 1279 6128 1416 6265 ne
rect 1416 6210 1471 6265
tri 1471 6210 1646 6385 sw
tri 1709 6265 1829 6385 ne
rect 1829 6265 1865 6385
rect 1985 6265 2021 6385
rect 1416 6128 1646 6210
tri 1646 6128 1728 6210 sw
tri 1829 6128 1966 6265 ne
rect 1966 6210 2021 6265
tri 2021 6210 2196 6385 sw
tri 2259 6265 2379 6385 ne
rect 2379 6265 2415 6385
rect 2535 6265 2571 6385
rect 1966 6128 2196 6210
tri 2196 6128 2278 6210 sw
tri 2379 6128 2516 6265 ne
rect 2516 6210 2571 6265
tri 2571 6210 2746 6385 sw
tri 2809 6265 2929 6385 ne
rect 2929 6265 2965 6385
rect 3085 6265 3121 6385
rect 2516 6128 2746 6210
tri 2746 6128 2828 6210 sw
tri 2929 6128 3066 6265 ne
rect 3066 6210 3121 6265
tri 3121 6210 3296 6385 sw
tri 3359 6265 3479 6385 ne
rect 3479 6265 3515 6385
rect 3635 6265 3671 6385
rect 3066 6128 3296 6210
tri 3296 6128 3378 6210 sw
tri 3479 6128 3616 6265 ne
rect 3616 6210 3671 6265
tri 3671 6210 3846 6385 sw
tri 3909 6265 4029 6385 ne
rect 4029 6265 4065 6385
rect 4185 6265 4221 6385
rect 3616 6128 3846 6210
tri 3846 6128 3928 6210 sw
tri 4029 6128 4166 6265 ne
rect 4166 6210 4221 6265
tri 4221 6210 4396 6385 sw
tri 4459 6265 4579 6385 ne
rect 4579 6265 4615 6385
rect 4735 6265 4771 6385
rect 4166 6128 4396 6210
tri 4396 6128 4478 6210 sw
tri 4579 6128 4716 6265 ne
rect 4716 6210 4771 6265
tri 4771 6210 4946 6385 sw
tri 5009 6265 5129 6385 ne
rect 5129 6265 5165 6385
rect 5285 6265 5321 6385
rect 4716 6128 4946 6210
tri 4946 6128 5028 6210 sw
tri 5129 6128 5266 6265 ne
rect 5266 6210 5321 6265
tri 5321 6210 5496 6385 sw
tri 5559 6265 5679 6385 ne
rect 5679 6265 5715 6385
rect 5835 6265 5871 6385
rect 5266 6128 5496 6210
tri 5496 6128 5578 6210 sw
tri 5679 6128 5816 6265 ne
rect 5816 6210 5871 6265
tri 5871 6210 6046 6385 sw
tri 6109 6265 6229 6385 ne
rect 6229 6265 6265 6385
rect 6385 6265 6421 6385
rect 5816 6128 6046 6210
tri 6046 6128 6128 6210 sw
tri 6229 6128 6366 6265 ne
rect 6366 6210 6421 6265
tri 6421 6210 6596 6385 sw
tri 6659 6265 6779 6385 ne
rect 6779 6265 6815 6385
rect 6935 6265 6971 6385
rect 6366 6128 6596 6210
tri 6596 6128 6678 6210 sw
tri 6779 6128 6916 6265 ne
rect 6916 6210 6971 6265
tri 6971 6210 7146 6385 sw
tri 7209 6265 7329 6385 ne
rect 7329 6265 7365 6385
rect 7485 6265 7521 6385
rect 6916 6128 7146 6210
tri 7146 6128 7228 6210 sw
tri 7329 6128 7466 6265 ne
rect 7466 6210 7521 6265
tri 7521 6210 7696 6385 sw
tri 7759 6265 7879 6385 ne
rect 7879 6265 7915 6385
rect 8035 6265 8071 6385
rect 7466 6128 7696 6210
tri 7696 6128 7778 6210 sw
tri 7879 6128 8016 6265 ne
rect 8016 6210 8071 6265
tri 8071 6210 8246 6385 sw
tri 8309 6265 8429 6385 ne
rect 8429 6265 8465 6385
rect 8585 6265 8621 6385
rect 8016 6128 8246 6210
tri 8246 6128 8328 6210 sw
tri 8429 6128 8566 6265 ne
rect 8566 6210 8621 6265
tri 8621 6210 8796 6385 sw
tri 8859 6265 8979 6385 ne
rect 8979 6265 9015 6385
rect 9135 6265 9171 6385
rect 8566 6128 8796 6210
tri 8796 6128 8878 6210 sw
tri 8979 6128 9116 6265 ne
rect 9116 6210 9171 6265
tri 9171 6210 9346 6385 sw
tri 9409 6265 9529 6385 ne
rect 9529 6265 9565 6385
rect 9685 6265 9721 6385
rect 9116 6128 9346 6210
tri 9346 6128 9428 6210 sw
tri 9529 6128 9666 6265 ne
rect 9666 6210 9721 6265
tri 9721 6210 9896 6385 sw
tri 9959 6265 10079 6385 ne
rect 10079 6265 10115 6385
rect 10235 6265 10271 6385
rect 9666 6128 9896 6210
tri 9896 6128 9978 6210 sw
tri 10079 6128 10216 6265 ne
rect 10216 6210 10271 6265
tri 10271 6210 10446 6385 sw
tri 10509 6265 10629 6385 ne
rect 10629 6265 10665 6385
rect 10785 6265 10821 6385
rect 10216 6128 10446 6210
tri 10446 6128 10528 6210 sw
tri 10629 6128 10766 6265 ne
rect 10766 6210 10821 6265
tri 10821 6210 10996 6385 sw
tri 11059 6265 11179 6385 ne
rect 11179 6265 11215 6385
rect 11335 6265 11371 6385
rect 10766 6128 10996 6210
tri 10996 6128 11078 6210 sw
tri 11179 6128 11316 6265 ne
rect 11316 6210 11371 6265
tri 11371 6210 11546 6385 sw
tri 11609 6265 11729 6385 ne
rect 11729 6265 11765 6385
rect 11885 6265 11921 6385
rect 11316 6128 11546 6210
tri 11546 6128 11628 6210 sw
tri 11729 6128 11866 6265 ne
rect 11866 6210 11921 6265
tri 11921 6210 12096 6385 sw
tri 12159 6265 12279 6385 ne
rect 12279 6265 12315 6385
rect 12435 6265 12471 6385
rect 11866 6128 12096 6210
tri 12096 6128 12178 6210 sw
tri 12279 6128 12416 6265 ne
rect 12416 6210 12471 6265
tri 12471 6210 12646 6385 sw
tri 12709 6265 12829 6385 ne
rect 12829 6265 12865 6385
rect 12985 6265 13021 6385
rect 12416 6128 12646 6210
tri 12646 6128 12728 6210 sw
tri 12829 6128 12966 6265 ne
rect 12966 6210 13021 6265
tri 13021 6210 13196 6385 sw
tri 13259 6265 13379 6385 ne
rect 13379 6265 13415 6385
rect 13535 6265 13571 6385
rect 12966 6128 13196 6210
tri 13196 6128 13278 6210 sw
tri 13379 6128 13516 6265 ne
rect 13516 6210 13571 6265
tri 13571 6210 13746 6385 sw
tri 13809 6265 13929 6385 ne
rect 13929 6265 13965 6385
rect 14085 6265 14121 6385
rect 13516 6128 13746 6210
tri 13746 6128 13828 6210 sw
tri 13929 6128 14066 6265 ne
rect 14066 6210 14121 6265
tri 14121 6210 14296 6385 sw
tri 14359 6265 14479 6385 ne
rect 14479 6265 14515 6385
rect 14635 6265 14671 6385
rect 14066 6128 14296 6210
tri 14296 6128 14378 6210 sw
tri 14479 6128 14616 6265 ne
rect 14616 6210 14671 6265
tri 14671 6210 14846 6385 sw
tri 14909 6265 15029 6385 ne
rect 15029 6265 15065 6385
rect 15185 6265 15221 6385
rect 14616 6128 14846 6210
tri 14846 6128 14928 6210 sw
tri 15029 6128 15166 6265 ne
rect 15166 6210 15221 6265
tri 15221 6210 15396 6385 sw
tri 15459 6265 15579 6385 ne
rect 15579 6265 15615 6385
rect 15735 6265 15771 6385
rect 15166 6128 15396 6210
tri 15396 6128 15478 6210 sw
tri 15579 6128 15716 6265 ne
rect 15716 6210 15771 6265
tri 15771 6210 15946 6385 sw
tri 16009 6265 16129 6385 ne
rect 16129 6265 16165 6385
rect 16285 6265 16321 6385
rect 15716 6128 15946 6210
tri 15946 6128 16028 6210 sw
tri 16129 6128 16266 6265 ne
rect 16266 6210 16321 6265
tri 16321 6210 16496 6385 sw
tri 16559 6265 16679 6385 ne
rect 16679 6265 16715 6385
rect 16835 6265 16871 6385
rect 16266 6128 16496 6210
tri 16496 6128 16578 6210 sw
tri 16679 6128 16816 6265 ne
rect 16816 6210 16871 6265
tri 16871 6210 17046 6385 sw
tri 17109 6265 17229 6385 ne
rect 17229 6265 17265 6385
rect 17385 6265 17421 6385
rect 16816 6128 17046 6210
tri 17046 6128 17128 6210 sw
tri 17229 6128 17366 6265 ne
rect 17366 6210 17421 6265
tri 17421 6210 17596 6385 sw
tri 17659 6265 17779 6385 ne
rect 17779 6265 17815 6385
rect 17935 6265 17971 6385
rect 17366 6128 17596 6210
tri 17596 6128 17678 6210 sw
tri 17779 6128 17916 6265 ne
rect 17916 6210 17971 6265
tri 17971 6210 18146 6385 sw
tri 18209 6265 18329 6385 ne
rect 18329 6265 18365 6385
rect 18485 6265 18521 6385
rect 17916 6128 18146 6210
tri 18146 6128 18228 6210 sw
tri 18329 6128 18466 6265 ne
rect 18466 6210 18521 6265
tri 18521 6210 18696 6385 sw
tri 18759 6265 18879 6385 ne
rect 18879 6265 18915 6385
rect 19035 6265 19071 6385
rect 18466 6128 18696 6210
tri 18696 6128 18778 6210 sw
tri 18879 6128 19016 6265 ne
rect 19016 6210 19071 6265
tri 19071 6210 19246 6385 sw
tri 19309 6265 19429 6385 ne
rect 19429 6265 19465 6385
rect 19585 6283 19621 6385
tri 19621 6283 19723 6385 sw
rect 20800 6283 21800 7072
rect 19585 6265 21800 6283
rect 19016 6128 19246 6210
tri 19246 6128 19328 6210 sw
tri 19429 6128 19566 6265 ne
rect 19566 6128 21800 6265
rect -500 5972 78 6128
tri 78 5972 234 6128 sw
tri 316 5972 472 6128 ne
rect 472 5972 628 6128
tri 628 5972 784 6128 sw
tri 866 5972 1022 6128 ne
rect 1022 5972 1178 6128
tri 1178 5972 1334 6128 sw
tri 1416 5972 1572 6128 ne
rect 1572 5972 1728 6128
tri 1728 5972 1884 6128 sw
tri 1966 5972 2122 6128 ne
rect 2122 5972 2278 6128
tri 2278 5972 2434 6128 sw
tri 2516 5972 2672 6128 ne
rect 2672 5972 2828 6128
tri 2828 5972 2984 6128 sw
tri 3066 5972 3222 6128 ne
rect 3222 5972 3378 6128
tri 3378 5972 3534 6128 sw
tri 3616 5972 3772 6128 ne
rect 3772 5972 3928 6128
tri 3928 5972 4084 6128 sw
tri 4166 5972 4322 6128 ne
rect 4322 5972 4478 6128
tri 4478 5972 4634 6128 sw
tri 4716 5972 4872 6128 ne
rect 4872 5972 5028 6128
tri 5028 5972 5184 6128 sw
tri 5266 5972 5422 6128 ne
rect 5422 5972 5578 6128
tri 5578 5972 5734 6128 sw
tri 5816 5972 5972 6128 ne
rect 5972 5972 6128 6128
tri 6128 5972 6284 6128 sw
tri 6366 5972 6522 6128 ne
rect 6522 5972 6678 6128
tri 6678 5972 6834 6128 sw
tri 6916 5972 7072 6128 ne
rect 7072 5972 7228 6128
tri 7228 5972 7384 6128 sw
tri 7466 5972 7622 6128 ne
rect 7622 5972 7778 6128
tri 7778 5972 7934 6128 sw
tri 8016 5972 8172 6128 ne
rect 8172 5972 8328 6128
tri 8328 5972 8484 6128 sw
tri 8566 5972 8722 6128 ne
rect 8722 5972 8878 6128
tri 8878 5972 9034 6128 sw
tri 9116 5972 9272 6128 ne
rect 9272 5972 9428 6128
tri 9428 5972 9584 6128 sw
tri 9666 5972 9822 6128 ne
rect 9822 5972 9978 6128
tri 9978 5972 10134 6128 sw
tri 10216 5972 10372 6128 ne
rect 10372 5972 10528 6128
tri 10528 5972 10684 6128 sw
tri 10766 5972 10922 6128 ne
rect 10922 5972 11078 6128
tri 11078 5972 11234 6128 sw
tri 11316 5972 11472 6128 ne
rect 11472 5972 11628 6128
tri 11628 5972 11784 6128 sw
tri 11866 5972 12022 6128 ne
rect 12022 5972 12178 6128
tri 12178 5972 12334 6128 sw
tri 12416 5972 12572 6128 ne
rect 12572 5972 12728 6128
tri 12728 5972 12884 6128 sw
tri 12966 5972 13122 6128 ne
rect 13122 5972 13278 6128
tri 13278 5972 13434 6128 sw
tri 13516 5972 13672 6128 ne
rect 13672 5972 13828 6128
tri 13828 5972 13984 6128 sw
tri 14066 5972 14222 6128 ne
rect 14222 5972 14378 6128
tri 14378 5972 14534 6128 sw
tri 14616 5972 14772 6128 ne
rect 14772 5972 14928 6128
tri 14928 5972 15084 6128 sw
tri 15166 5972 15322 6128 ne
rect 15322 5972 15478 6128
tri 15478 5972 15634 6128 sw
tri 15716 5972 15872 6128 ne
rect 15872 5972 16028 6128
tri 16028 5972 16184 6128 sw
tri 16266 5972 16422 6128 ne
rect 16422 5972 16578 6128
tri 16578 5972 16734 6128 sw
tri 16816 5972 16972 6128 ne
rect 16972 5972 17128 6128
tri 17128 5972 17284 6128 sw
tri 17366 5972 17522 6128 ne
rect 17522 5972 17678 6128
tri 17678 5972 17834 6128 sw
tri 17916 5972 18072 6128 ne
rect 18072 5972 18228 6128
tri 18228 5972 18384 6128 sw
tri 18466 5972 18622 6128 ne
rect 18622 5972 18778 6128
tri 18778 5972 18934 6128 sw
tri 19016 5972 19172 6128 ne
rect 19172 5972 19328 6128
tri 19328 5972 19484 6128 sw
tri 19566 5972 19722 6128 ne
rect 19722 5972 21800 6128
rect -500 5835 234 5972
tri 234 5835 371 5972 sw
tri 472 5835 609 5972 ne
rect 609 5835 784 5972
tri 784 5835 921 5972 sw
tri 1022 5835 1159 5972 ne
rect 1159 5835 1334 5972
tri 1334 5835 1471 5972 sw
tri 1572 5835 1709 5972 ne
rect 1709 5835 1884 5972
tri 1884 5835 2021 5972 sw
tri 2122 5835 2259 5972 ne
rect 2259 5835 2434 5972
tri 2434 5835 2571 5972 sw
tri 2672 5835 2809 5972 ne
rect 2809 5835 2984 5972
tri 2984 5835 3121 5972 sw
tri 3222 5835 3359 5972 ne
rect 3359 5835 3534 5972
tri 3534 5835 3671 5972 sw
tri 3772 5835 3909 5972 ne
rect 3909 5835 4084 5972
tri 4084 5835 4221 5972 sw
tri 4322 5835 4459 5972 ne
rect 4459 5835 4634 5972
tri 4634 5835 4771 5972 sw
tri 4872 5835 5009 5972 ne
rect 5009 5835 5184 5972
tri 5184 5835 5321 5972 sw
tri 5422 5835 5559 5972 ne
rect 5559 5835 5734 5972
tri 5734 5835 5871 5972 sw
tri 5972 5835 6109 5972 ne
rect 6109 5835 6284 5972
tri 6284 5835 6421 5972 sw
tri 6522 5835 6659 5972 ne
rect 6659 5835 6834 5972
tri 6834 5835 6971 5972 sw
tri 7072 5835 7209 5972 ne
rect 7209 5835 7384 5972
tri 7384 5835 7521 5972 sw
tri 7622 5835 7759 5972 ne
rect 7759 5835 7934 5972
tri 7934 5835 8071 5972 sw
tri 8172 5835 8309 5972 ne
rect 8309 5835 8484 5972
tri 8484 5835 8621 5972 sw
tri 8722 5835 8859 5972 ne
rect 8859 5835 9034 5972
tri 9034 5835 9171 5972 sw
tri 9272 5835 9409 5972 ne
rect 9409 5835 9584 5972
tri 9584 5835 9721 5972 sw
tri 9822 5835 9959 5972 ne
rect 9959 5835 10134 5972
tri 10134 5835 10271 5972 sw
tri 10372 5835 10509 5972 ne
rect 10509 5835 10684 5972
tri 10684 5835 10821 5972 sw
tri 10922 5835 11059 5972 ne
rect 11059 5835 11234 5972
tri 11234 5835 11371 5972 sw
tri 11472 5835 11609 5972 ne
rect 11609 5835 11784 5972
tri 11784 5835 11921 5972 sw
tri 12022 5835 12159 5972 ne
rect 12159 5835 12334 5972
tri 12334 5835 12471 5972 sw
tri 12572 5835 12709 5972 ne
rect 12709 5835 12884 5972
tri 12884 5835 13021 5972 sw
tri 13122 5835 13259 5972 ne
rect 13259 5835 13434 5972
tri 13434 5835 13571 5972 sw
tri 13672 5835 13809 5972 ne
rect 13809 5835 13984 5972
tri 13984 5835 14121 5972 sw
tri 14222 5835 14359 5972 ne
rect 14359 5835 14534 5972
tri 14534 5835 14671 5972 sw
tri 14772 5835 14909 5972 ne
rect 14909 5835 15084 5972
tri 15084 5835 15221 5972 sw
tri 15322 5835 15459 5972 ne
rect 15459 5835 15634 5972
tri 15634 5835 15771 5972 sw
tri 15872 5835 16009 5972 ne
rect 16009 5835 16184 5972
tri 16184 5835 16321 5972 sw
tri 16422 5835 16559 5972 ne
rect 16559 5835 16734 5972
tri 16734 5835 16871 5972 sw
tri 16972 5835 17109 5972 ne
rect 17109 5835 17284 5972
tri 17284 5835 17421 5972 sw
tri 17522 5835 17659 5972 ne
rect 17659 5835 17834 5972
tri 17834 5835 17971 5972 sw
tri 18072 5835 18209 5972 ne
rect 18209 5835 18384 5972
tri 18384 5835 18521 5972 sw
tri 18622 5835 18759 5972 ne
rect 18759 5835 18934 5972
tri 18934 5835 19071 5972 sw
tri 19172 5835 19309 5972 ne
rect 19309 5835 19484 5972
tri 19484 5835 19621 5972 sw
rect -500 5817 215 5835
tri 77 5715 179 5817 ne
rect 179 5715 215 5817
rect 335 5715 371 5835
tri 179 5578 316 5715 ne
rect 316 5660 371 5715
tri 371 5660 546 5835 sw
tri 609 5715 729 5835 ne
rect 729 5715 765 5835
rect 885 5715 921 5835
rect 316 5578 546 5660
tri 546 5578 628 5660 sw
tri 729 5578 866 5715 ne
rect 866 5660 921 5715
tri 921 5660 1096 5835 sw
tri 1159 5715 1279 5835 ne
rect 1279 5715 1315 5835
rect 1435 5715 1471 5835
rect 866 5578 1096 5660
tri 1096 5578 1178 5660 sw
tri 1279 5578 1416 5715 ne
rect 1416 5660 1471 5715
tri 1471 5660 1646 5835 sw
tri 1709 5715 1829 5835 ne
rect 1829 5715 1865 5835
rect 1985 5715 2021 5835
rect 1416 5578 1646 5660
tri 1646 5578 1728 5660 sw
tri 1829 5578 1966 5715 ne
rect 1966 5660 2021 5715
tri 2021 5660 2196 5835 sw
tri 2259 5715 2379 5835 ne
rect 2379 5715 2415 5835
rect 2535 5715 2571 5835
rect 1966 5578 2196 5660
tri 2196 5578 2278 5660 sw
tri 2379 5578 2516 5715 ne
rect 2516 5660 2571 5715
tri 2571 5660 2746 5835 sw
tri 2809 5715 2929 5835 ne
rect 2929 5715 2965 5835
rect 3085 5715 3121 5835
rect 2516 5578 2746 5660
tri 2746 5578 2828 5660 sw
tri 2929 5578 3066 5715 ne
rect 3066 5660 3121 5715
tri 3121 5660 3296 5835 sw
tri 3359 5715 3479 5835 ne
rect 3479 5715 3515 5835
rect 3635 5715 3671 5835
rect 3066 5578 3296 5660
tri 3296 5578 3378 5660 sw
tri 3479 5578 3616 5715 ne
rect 3616 5660 3671 5715
tri 3671 5660 3846 5835 sw
tri 3909 5715 4029 5835 ne
rect 4029 5715 4065 5835
rect 4185 5715 4221 5835
rect 3616 5578 3846 5660
tri 3846 5578 3928 5660 sw
tri 4029 5578 4166 5715 ne
rect 4166 5660 4221 5715
tri 4221 5660 4396 5835 sw
tri 4459 5715 4579 5835 ne
rect 4579 5715 4615 5835
rect 4735 5715 4771 5835
rect 4166 5578 4396 5660
tri 4396 5578 4478 5660 sw
tri 4579 5578 4716 5715 ne
rect 4716 5660 4771 5715
tri 4771 5660 4946 5835 sw
tri 5009 5715 5129 5835 ne
rect 5129 5715 5165 5835
rect 5285 5715 5321 5835
rect 4716 5578 4946 5660
tri 4946 5578 5028 5660 sw
tri 5129 5578 5266 5715 ne
rect 5266 5660 5321 5715
tri 5321 5660 5496 5835 sw
tri 5559 5715 5679 5835 ne
rect 5679 5715 5715 5835
rect 5835 5715 5871 5835
rect 5266 5578 5496 5660
tri 5496 5578 5578 5660 sw
tri 5679 5578 5816 5715 ne
rect 5816 5660 5871 5715
tri 5871 5660 6046 5835 sw
tri 6109 5715 6229 5835 ne
rect 6229 5715 6265 5835
rect 6385 5715 6421 5835
rect 5816 5578 6046 5660
tri 6046 5578 6128 5660 sw
tri 6229 5578 6366 5715 ne
rect 6366 5660 6421 5715
tri 6421 5660 6596 5835 sw
tri 6659 5715 6779 5835 ne
rect 6779 5715 6815 5835
rect 6935 5715 6971 5835
rect 6366 5578 6596 5660
tri 6596 5578 6678 5660 sw
tri 6779 5578 6916 5715 ne
rect 6916 5660 6971 5715
tri 6971 5660 7146 5835 sw
tri 7209 5715 7329 5835 ne
rect 7329 5715 7365 5835
rect 7485 5715 7521 5835
rect 6916 5578 7146 5660
tri 7146 5578 7228 5660 sw
tri 7329 5578 7466 5715 ne
rect 7466 5660 7521 5715
tri 7521 5660 7696 5835 sw
tri 7759 5715 7879 5835 ne
rect 7879 5715 7915 5835
rect 8035 5715 8071 5835
rect 7466 5578 7696 5660
tri 7696 5578 7778 5660 sw
tri 7879 5578 8016 5715 ne
rect 8016 5660 8071 5715
tri 8071 5660 8246 5835 sw
tri 8309 5715 8429 5835 ne
rect 8429 5715 8465 5835
rect 8585 5715 8621 5835
rect 8016 5578 8246 5660
tri 8246 5578 8328 5660 sw
tri 8429 5578 8566 5715 ne
rect 8566 5660 8621 5715
tri 8621 5660 8796 5835 sw
tri 8859 5715 8979 5835 ne
rect 8979 5715 9015 5835
rect 9135 5715 9171 5835
rect 8566 5578 8796 5660
tri 8796 5578 8878 5660 sw
tri 8979 5578 9116 5715 ne
rect 9116 5660 9171 5715
tri 9171 5660 9346 5835 sw
tri 9409 5715 9529 5835 ne
rect 9529 5715 9565 5835
rect 9685 5715 9721 5835
rect 9116 5578 9346 5660
tri 9346 5578 9428 5660 sw
tri 9529 5578 9666 5715 ne
rect 9666 5660 9721 5715
tri 9721 5660 9896 5835 sw
tri 9959 5715 10079 5835 ne
rect 10079 5715 10115 5835
rect 10235 5715 10271 5835
rect 9666 5578 9896 5660
tri 9896 5578 9978 5660 sw
tri 10079 5578 10216 5715 ne
rect 10216 5660 10271 5715
tri 10271 5660 10446 5835 sw
tri 10509 5715 10629 5835 ne
rect 10629 5715 10665 5835
rect 10785 5715 10821 5835
rect 10216 5578 10446 5660
tri 10446 5578 10528 5660 sw
tri 10629 5578 10766 5715 ne
rect 10766 5660 10821 5715
tri 10821 5660 10996 5835 sw
tri 11059 5715 11179 5835 ne
rect 11179 5715 11215 5835
rect 11335 5715 11371 5835
rect 10766 5578 10996 5660
tri 10996 5578 11078 5660 sw
tri 11179 5578 11316 5715 ne
rect 11316 5660 11371 5715
tri 11371 5660 11546 5835 sw
tri 11609 5715 11729 5835 ne
rect 11729 5715 11765 5835
rect 11885 5715 11921 5835
rect 11316 5578 11546 5660
tri 11546 5578 11628 5660 sw
tri 11729 5578 11866 5715 ne
rect 11866 5660 11921 5715
tri 11921 5660 12096 5835 sw
tri 12159 5715 12279 5835 ne
rect 12279 5715 12315 5835
rect 12435 5715 12471 5835
rect 11866 5578 12096 5660
tri 12096 5578 12178 5660 sw
tri 12279 5578 12416 5715 ne
rect 12416 5660 12471 5715
tri 12471 5660 12646 5835 sw
tri 12709 5715 12829 5835 ne
rect 12829 5715 12865 5835
rect 12985 5715 13021 5835
rect 12416 5578 12646 5660
tri 12646 5578 12728 5660 sw
tri 12829 5578 12966 5715 ne
rect 12966 5660 13021 5715
tri 13021 5660 13196 5835 sw
tri 13259 5715 13379 5835 ne
rect 13379 5715 13415 5835
rect 13535 5715 13571 5835
rect 12966 5578 13196 5660
tri 13196 5578 13278 5660 sw
tri 13379 5578 13516 5715 ne
rect 13516 5660 13571 5715
tri 13571 5660 13746 5835 sw
tri 13809 5715 13929 5835 ne
rect 13929 5715 13965 5835
rect 14085 5715 14121 5835
rect 13516 5578 13746 5660
tri 13746 5578 13828 5660 sw
tri 13929 5578 14066 5715 ne
rect 14066 5660 14121 5715
tri 14121 5660 14296 5835 sw
tri 14359 5715 14479 5835 ne
rect 14479 5715 14515 5835
rect 14635 5715 14671 5835
rect 14066 5578 14296 5660
tri 14296 5578 14378 5660 sw
tri 14479 5578 14616 5715 ne
rect 14616 5660 14671 5715
tri 14671 5660 14846 5835 sw
tri 14909 5715 15029 5835 ne
rect 15029 5715 15065 5835
rect 15185 5715 15221 5835
rect 14616 5578 14846 5660
tri 14846 5578 14928 5660 sw
tri 15029 5578 15166 5715 ne
rect 15166 5660 15221 5715
tri 15221 5660 15396 5835 sw
tri 15459 5715 15579 5835 ne
rect 15579 5715 15615 5835
rect 15735 5715 15771 5835
rect 15166 5578 15396 5660
tri 15396 5578 15478 5660 sw
tri 15579 5578 15716 5715 ne
rect 15716 5660 15771 5715
tri 15771 5660 15946 5835 sw
tri 16009 5715 16129 5835 ne
rect 16129 5715 16165 5835
rect 16285 5715 16321 5835
rect 15716 5578 15946 5660
tri 15946 5578 16028 5660 sw
tri 16129 5578 16266 5715 ne
rect 16266 5660 16321 5715
tri 16321 5660 16496 5835 sw
tri 16559 5715 16679 5835 ne
rect 16679 5715 16715 5835
rect 16835 5715 16871 5835
rect 16266 5578 16496 5660
tri 16496 5578 16578 5660 sw
tri 16679 5578 16816 5715 ne
rect 16816 5660 16871 5715
tri 16871 5660 17046 5835 sw
tri 17109 5715 17229 5835 ne
rect 17229 5715 17265 5835
rect 17385 5715 17421 5835
rect 16816 5578 17046 5660
tri 17046 5578 17128 5660 sw
tri 17229 5578 17366 5715 ne
rect 17366 5660 17421 5715
tri 17421 5660 17596 5835 sw
tri 17659 5715 17779 5835 ne
rect 17779 5715 17815 5835
rect 17935 5715 17971 5835
rect 17366 5578 17596 5660
tri 17596 5578 17678 5660 sw
tri 17779 5578 17916 5715 ne
rect 17916 5660 17971 5715
tri 17971 5660 18146 5835 sw
tri 18209 5715 18329 5835 ne
rect 18329 5715 18365 5835
rect 18485 5715 18521 5835
rect 17916 5578 18146 5660
tri 18146 5578 18228 5660 sw
tri 18329 5578 18466 5715 ne
rect 18466 5660 18521 5715
tri 18521 5660 18696 5835 sw
tri 18759 5715 18879 5835 ne
rect 18879 5715 18915 5835
rect 19035 5715 19071 5835
rect 18466 5578 18696 5660
tri 18696 5578 18778 5660 sw
tri 18879 5578 19016 5715 ne
rect 19016 5660 19071 5715
tri 19071 5660 19246 5835 sw
tri 19309 5715 19429 5835 ne
rect 19429 5715 19465 5835
rect 19585 5733 19621 5835
tri 19621 5733 19723 5835 sw
rect 19585 5715 20300 5733
rect 19016 5578 19246 5660
tri 19246 5578 19328 5660 sw
tri 19429 5578 19566 5715 ne
rect 19566 5578 20300 5715
rect -2000 5422 78 5578
tri 78 5422 234 5578 sw
tri 316 5422 472 5578 ne
rect 472 5422 628 5578
tri 628 5422 784 5578 sw
tri 866 5422 1022 5578 ne
rect 1022 5422 1178 5578
tri 1178 5422 1334 5578 sw
tri 1416 5422 1572 5578 ne
rect 1572 5422 1728 5578
tri 1728 5422 1884 5578 sw
tri 1966 5422 2122 5578 ne
rect 2122 5422 2278 5578
tri 2278 5422 2434 5578 sw
tri 2516 5422 2672 5578 ne
rect 2672 5422 2828 5578
tri 2828 5422 2984 5578 sw
tri 3066 5422 3222 5578 ne
rect 3222 5422 3378 5578
tri 3378 5422 3534 5578 sw
tri 3616 5422 3772 5578 ne
rect 3772 5422 3928 5578
tri 3928 5422 4084 5578 sw
tri 4166 5422 4322 5578 ne
rect 4322 5422 4478 5578
tri 4478 5422 4634 5578 sw
tri 4716 5422 4872 5578 ne
rect 4872 5422 5028 5578
tri 5028 5422 5184 5578 sw
tri 5266 5422 5422 5578 ne
rect 5422 5422 5578 5578
tri 5578 5422 5734 5578 sw
tri 5816 5422 5972 5578 ne
rect 5972 5422 6128 5578
tri 6128 5422 6284 5578 sw
tri 6366 5422 6522 5578 ne
rect 6522 5422 6678 5578
tri 6678 5422 6834 5578 sw
tri 6916 5422 7072 5578 ne
rect 7072 5422 7228 5578
tri 7228 5422 7384 5578 sw
tri 7466 5422 7622 5578 ne
rect 7622 5422 7778 5578
tri 7778 5422 7934 5578 sw
tri 8016 5422 8172 5578 ne
rect 8172 5422 8328 5578
tri 8328 5422 8484 5578 sw
tri 8566 5422 8722 5578 ne
rect 8722 5422 8878 5578
tri 8878 5422 9034 5578 sw
tri 9116 5422 9272 5578 ne
rect 9272 5422 9428 5578
tri 9428 5422 9584 5578 sw
tri 9666 5422 9822 5578 ne
rect 9822 5422 9978 5578
tri 9978 5422 10134 5578 sw
tri 10216 5422 10372 5578 ne
rect 10372 5422 10528 5578
tri 10528 5422 10684 5578 sw
tri 10766 5422 10922 5578 ne
rect 10922 5422 11078 5578
tri 11078 5422 11234 5578 sw
tri 11316 5422 11472 5578 ne
rect 11472 5422 11628 5578
tri 11628 5422 11784 5578 sw
tri 11866 5422 12022 5578 ne
rect 12022 5422 12178 5578
tri 12178 5422 12334 5578 sw
tri 12416 5422 12572 5578 ne
rect 12572 5422 12728 5578
tri 12728 5422 12884 5578 sw
tri 12966 5422 13122 5578 ne
rect 13122 5422 13278 5578
tri 13278 5422 13434 5578 sw
tri 13516 5422 13672 5578 ne
rect 13672 5422 13828 5578
tri 13828 5422 13984 5578 sw
tri 14066 5422 14222 5578 ne
rect 14222 5422 14378 5578
tri 14378 5422 14534 5578 sw
tri 14616 5422 14772 5578 ne
rect 14772 5422 14928 5578
tri 14928 5422 15084 5578 sw
tri 15166 5422 15322 5578 ne
rect 15322 5422 15478 5578
tri 15478 5422 15634 5578 sw
tri 15716 5422 15872 5578 ne
rect 15872 5422 16028 5578
tri 16028 5422 16184 5578 sw
tri 16266 5422 16422 5578 ne
rect 16422 5422 16578 5578
tri 16578 5422 16734 5578 sw
tri 16816 5422 16972 5578 ne
rect 16972 5422 17128 5578
tri 17128 5422 17284 5578 sw
tri 17366 5422 17522 5578 ne
rect 17522 5422 17678 5578
tri 17678 5422 17834 5578 sw
tri 17916 5422 18072 5578 ne
rect 18072 5422 18228 5578
tri 18228 5422 18384 5578 sw
tri 18466 5422 18622 5578 ne
rect 18622 5422 18778 5578
tri 18778 5422 18934 5578 sw
tri 19016 5422 19172 5578 ne
rect 19172 5422 19328 5578
tri 19328 5422 19484 5578 sw
tri 19566 5422 19722 5578 ne
rect 19722 5422 20300 5578
rect -2000 5285 234 5422
tri 234 5285 371 5422 sw
tri 472 5285 609 5422 ne
rect 609 5285 784 5422
tri 784 5285 921 5422 sw
tri 1022 5285 1159 5422 ne
rect 1159 5285 1334 5422
tri 1334 5285 1471 5422 sw
tri 1572 5285 1709 5422 ne
rect 1709 5285 1884 5422
tri 1884 5285 2021 5422 sw
tri 2122 5285 2259 5422 ne
rect 2259 5285 2434 5422
tri 2434 5285 2571 5422 sw
tri 2672 5285 2809 5422 ne
rect 2809 5285 2984 5422
tri 2984 5285 3121 5422 sw
tri 3222 5285 3359 5422 ne
rect 3359 5285 3534 5422
tri 3534 5285 3671 5422 sw
tri 3772 5285 3909 5422 ne
rect 3909 5285 4084 5422
tri 4084 5285 4221 5422 sw
tri 4322 5285 4459 5422 ne
rect 4459 5285 4634 5422
tri 4634 5285 4771 5422 sw
tri 4872 5285 5009 5422 ne
rect 5009 5285 5184 5422
tri 5184 5285 5321 5422 sw
tri 5422 5285 5559 5422 ne
rect 5559 5285 5734 5422
tri 5734 5285 5871 5422 sw
tri 5972 5285 6109 5422 ne
rect 6109 5285 6284 5422
tri 6284 5285 6421 5422 sw
tri 6522 5285 6659 5422 ne
rect 6659 5285 6834 5422
tri 6834 5285 6971 5422 sw
tri 7072 5285 7209 5422 ne
rect 7209 5285 7384 5422
tri 7384 5285 7521 5422 sw
tri 7622 5285 7759 5422 ne
rect 7759 5285 7934 5422
tri 7934 5285 8071 5422 sw
tri 8172 5285 8309 5422 ne
rect 8309 5285 8484 5422
tri 8484 5285 8621 5422 sw
tri 8722 5285 8859 5422 ne
rect 8859 5285 9034 5422
tri 9034 5285 9171 5422 sw
tri 9272 5285 9409 5422 ne
rect 9409 5285 9584 5422
tri 9584 5285 9721 5422 sw
tri 9822 5285 9959 5422 ne
rect 9959 5285 10134 5422
tri 10134 5285 10271 5422 sw
tri 10372 5285 10509 5422 ne
rect 10509 5285 10684 5422
tri 10684 5285 10821 5422 sw
tri 10922 5285 11059 5422 ne
rect 11059 5285 11234 5422
tri 11234 5285 11371 5422 sw
tri 11472 5285 11609 5422 ne
rect 11609 5285 11784 5422
tri 11784 5285 11921 5422 sw
tri 12022 5285 12159 5422 ne
rect 12159 5285 12334 5422
tri 12334 5285 12471 5422 sw
tri 12572 5285 12709 5422 ne
rect 12709 5285 12884 5422
tri 12884 5285 13021 5422 sw
tri 13122 5285 13259 5422 ne
rect 13259 5285 13434 5422
tri 13434 5285 13571 5422 sw
tri 13672 5285 13809 5422 ne
rect 13809 5285 13984 5422
tri 13984 5285 14121 5422 sw
tri 14222 5285 14359 5422 ne
rect 14359 5285 14534 5422
tri 14534 5285 14671 5422 sw
tri 14772 5285 14909 5422 ne
rect 14909 5285 15084 5422
tri 15084 5285 15221 5422 sw
tri 15322 5285 15459 5422 ne
rect 15459 5285 15634 5422
tri 15634 5285 15771 5422 sw
tri 15872 5285 16009 5422 ne
rect 16009 5285 16184 5422
tri 16184 5285 16321 5422 sw
tri 16422 5285 16559 5422 ne
rect 16559 5285 16734 5422
tri 16734 5285 16871 5422 sw
tri 16972 5285 17109 5422 ne
rect 17109 5285 17284 5422
tri 17284 5285 17421 5422 sw
tri 17522 5285 17659 5422 ne
rect 17659 5285 17834 5422
tri 17834 5285 17971 5422 sw
tri 18072 5285 18209 5422 ne
rect 18209 5285 18384 5422
tri 18384 5285 18521 5422 sw
tri 18622 5285 18759 5422 ne
rect 18759 5285 18934 5422
tri 18934 5285 19071 5422 sw
tri 19172 5285 19309 5422 ne
rect 19309 5285 19484 5422
tri 19484 5285 19621 5422 sw
rect -2000 5267 215 5285
rect -2000 4478 -1000 5267
tri 77 5165 179 5267 ne
rect 179 5165 215 5267
rect 335 5165 371 5285
tri 179 5028 316 5165 ne
rect 316 5110 371 5165
tri 371 5110 546 5285 sw
tri 609 5165 729 5285 ne
rect 729 5165 765 5285
rect 885 5165 921 5285
rect 316 5028 546 5110
tri 546 5028 628 5110 sw
tri 729 5028 866 5165 ne
rect 866 5110 921 5165
tri 921 5110 1096 5285 sw
tri 1159 5165 1279 5285 ne
rect 1279 5165 1315 5285
rect 1435 5165 1471 5285
rect 866 5028 1096 5110
tri 1096 5028 1178 5110 sw
tri 1279 5028 1416 5165 ne
rect 1416 5110 1471 5165
tri 1471 5110 1646 5285 sw
tri 1709 5165 1829 5285 ne
rect 1829 5165 1865 5285
rect 1985 5165 2021 5285
rect 1416 5028 1646 5110
tri 1646 5028 1728 5110 sw
tri 1829 5028 1966 5165 ne
rect 1966 5110 2021 5165
tri 2021 5110 2196 5285 sw
tri 2259 5165 2379 5285 ne
rect 2379 5165 2415 5285
rect 2535 5165 2571 5285
rect 1966 5028 2196 5110
tri 2196 5028 2278 5110 sw
tri 2379 5028 2516 5165 ne
rect 2516 5110 2571 5165
tri 2571 5110 2746 5285 sw
tri 2809 5165 2929 5285 ne
rect 2929 5165 2965 5285
rect 3085 5165 3121 5285
rect 2516 5028 2746 5110
tri 2746 5028 2828 5110 sw
tri 2929 5028 3066 5165 ne
rect 3066 5110 3121 5165
tri 3121 5110 3296 5285 sw
tri 3359 5165 3479 5285 ne
rect 3479 5165 3515 5285
rect 3635 5165 3671 5285
rect 3066 5028 3296 5110
tri 3296 5028 3378 5110 sw
tri 3479 5028 3616 5165 ne
rect 3616 5110 3671 5165
tri 3671 5110 3846 5285 sw
tri 3909 5165 4029 5285 ne
rect 4029 5165 4065 5285
rect 4185 5165 4221 5285
rect 3616 5028 3846 5110
tri 3846 5028 3928 5110 sw
tri 4029 5028 4166 5165 ne
rect 4166 5110 4221 5165
tri 4221 5110 4396 5285 sw
tri 4459 5165 4579 5285 ne
rect 4579 5165 4615 5285
rect 4735 5165 4771 5285
rect 4166 5028 4396 5110
tri 4396 5028 4478 5110 sw
tri 4579 5028 4716 5165 ne
rect 4716 5110 4771 5165
tri 4771 5110 4946 5285 sw
tri 5009 5165 5129 5285 ne
rect 5129 5165 5165 5285
rect 5285 5165 5321 5285
rect 4716 5028 4946 5110
tri 4946 5028 5028 5110 sw
tri 5129 5028 5266 5165 ne
rect 5266 5110 5321 5165
tri 5321 5110 5496 5285 sw
tri 5559 5165 5679 5285 ne
rect 5679 5165 5715 5285
rect 5835 5165 5871 5285
rect 5266 5028 5496 5110
tri 5496 5028 5578 5110 sw
tri 5679 5028 5816 5165 ne
rect 5816 5110 5871 5165
tri 5871 5110 6046 5285 sw
tri 6109 5165 6229 5285 ne
rect 6229 5165 6265 5285
rect 6385 5165 6421 5285
rect 5816 5028 6046 5110
tri 6046 5028 6128 5110 sw
tri 6229 5028 6366 5165 ne
rect 6366 5110 6421 5165
tri 6421 5110 6596 5285 sw
tri 6659 5165 6779 5285 ne
rect 6779 5165 6815 5285
rect 6935 5165 6971 5285
rect 6366 5028 6596 5110
tri 6596 5028 6678 5110 sw
tri 6779 5028 6916 5165 ne
rect 6916 5110 6971 5165
tri 6971 5110 7146 5285 sw
tri 7209 5165 7329 5285 ne
rect 7329 5165 7365 5285
rect 7485 5165 7521 5285
rect 6916 5028 7146 5110
tri 7146 5028 7228 5110 sw
tri 7329 5028 7466 5165 ne
rect 7466 5110 7521 5165
tri 7521 5110 7696 5285 sw
tri 7759 5165 7879 5285 ne
rect 7879 5165 7915 5285
rect 8035 5165 8071 5285
rect 7466 5028 7696 5110
tri 7696 5028 7778 5110 sw
tri 7879 5028 8016 5165 ne
rect 8016 5110 8071 5165
tri 8071 5110 8246 5285 sw
tri 8309 5165 8429 5285 ne
rect 8429 5165 8465 5285
rect 8585 5165 8621 5285
rect 8016 5028 8246 5110
tri 8246 5028 8328 5110 sw
tri 8429 5028 8566 5165 ne
rect 8566 5110 8621 5165
tri 8621 5110 8796 5285 sw
tri 8859 5165 8979 5285 ne
rect 8979 5165 9015 5285
rect 9135 5165 9171 5285
rect 8566 5028 8796 5110
tri 8796 5028 8878 5110 sw
tri 8979 5028 9116 5165 ne
rect 9116 5110 9171 5165
tri 9171 5110 9346 5285 sw
tri 9409 5165 9529 5285 ne
rect 9529 5165 9565 5285
rect 9685 5165 9721 5285
rect 9116 5028 9346 5110
tri 9346 5028 9428 5110 sw
tri 9529 5028 9666 5165 ne
rect 9666 5110 9721 5165
tri 9721 5110 9896 5285 sw
tri 9959 5165 10079 5285 ne
rect 10079 5165 10115 5285
rect 10235 5165 10271 5285
rect 9666 5028 9896 5110
tri 9896 5028 9978 5110 sw
tri 10079 5028 10216 5165 ne
rect 10216 5110 10271 5165
tri 10271 5110 10446 5285 sw
tri 10509 5165 10629 5285 ne
rect 10629 5165 10665 5285
rect 10785 5165 10821 5285
rect 10216 5028 10446 5110
tri 10446 5028 10528 5110 sw
tri 10629 5028 10766 5165 ne
rect 10766 5110 10821 5165
tri 10821 5110 10996 5285 sw
tri 11059 5165 11179 5285 ne
rect 11179 5165 11215 5285
rect 11335 5165 11371 5285
rect 10766 5028 10996 5110
tri 10996 5028 11078 5110 sw
tri 11179 5028 11316 5165 ne
rect 11316 5110 11371 5165
tri 11371 5110 11546 5285 sw
tri 11609 5165 11729 5285 ne
rect 11729 5165 11765 5285
rect 11885 5165 11921 5285
rect 11316 5028 11546 5110
tri 11546 5028 11628 5110 sw
tri 11729 5028 11866 5165 ne
rect 11866 5110 11921 5165
tri 11921 5110 12096 5285 sw
tri 12159 5165 12279 5285 ne
rect 12279 5165 12315 5285
rect 12435 5165 12471 5285
rect 11866 5028 12096 5110
tri 12096 5028 12178 5110 sw
tri 12279 5028 12416 5165 ne
rect 12416 5110 12471 5165
tri 12471 5110 12646 5285 sw
tri 12709 5165 12829 5285 ne
rect 12829 5165 12865 5285
rect 12985 5165 13021 5285
rect 12416 5028 12646 5110
tri 12646 5028 12728 5110 sw
tri 12829 5028 12966 5165 ne
rect 12966 5110 13021 5165
tri 13021 5110 13196 5285 sw
tri 13259 5165 13379 5285 ne
rect 13379 5165 13415 5285
rect 13535 5165 13571 5285
rect 12966 5028 13196 5110
tri 13196 5028 13278 5110 sw
tri 13379 5028 13516 5165 ne
rect 13516 5110 13571 5165
tri 13571 5110 13746 5285 sw
tri 13809 5165 13929 5285 ne
rect 13929 5165 13965 5285
rect 14085 5165 14121 5285
rect 13516 5028 13746 5110
tri 13746 5028 13828 5110 sw
tri 13929 5028 14066 5165 ne
rect 14066 5110 14121 5165
tri 14121 5110 14296 5285 sw
tri 14359 5165 14479 5285 ne
rect 14479 5165 14515 5285
rect 14635 5165 14671 5285
rect 14066 5028 14296 5110
tri 14296 5028 14378 5110 sw
tri 14479 5028 14616 5165 ne
rect 14616 5110 14671 5165
tri 14671 5110 14846 5285 sw
tri 14909 5165 15029 5285 ne
rect 15029 5165 15065 5285
rect 15185 5165 15221 5285
rect 14616 5028 14846 5110
tri 14846 5028 14928 5110 sw
tri 15029 5028 15166 5165 ne
rect 15166 5110 15221 5165
tri 15221 5110 15396 5285 sw
tri 15459 5165 15579 5285 ne
rect 15579 5165 15615 5285
rect 15735 5165 15771 5285
rect 15166 5028 15396 5110
tri 15396 5028 15478 5110 sw
tri 15579 5028 15716 5165 ne
rect 15716 5110 15771 5165
tri 15771 5110 15946 5285 sw
tri 16009 5165 16129 5285 ne
rect 16129 5165 16165 5285
rect 16285 5165 16321 5285
rect 15716 5028 15946 5110
tri 15946 5028 16028 5110 sw
tri 16129 5028 16266 5165 ne
rect 16266 5110 16321 5165
tri 16321 5110 16496 5285 sw
tri 16559 5165 16679 5285 ne
rect 16679 5165 16715 5285
rect 16835 5165 16871 5285
rect 16266 5028 16496 5110
tri 16496 5028 16578 5110 sw
tri 16679 5028 16816 5165 ne
rect 16816 5110 16871 5165
tri 16871 5110 17046 5285 sw
tri 17109 5165 17229 5285 ne
rect 17229 5165 17265 5285
rect 17385 5165 17421 5285
rect 16816 5028 17046 5110
tri 17046 5028 17128 5110 sw
tri 17229 5028 17366 5165 ne
rect 17366 5110 17421 5165
tri 17421 5110 17596 5285 sw
tri 17659 5165 17779 5285 ne
rect 17779 5165 17815 5285
rect 17935 5165 17971 5285
rect 17366 5028 17596 5110
tri 17596 5028 17678 5110 sw
tri 17779 5028 17916 5165 ne
rect 17916 5110 17971 5165
tri 17971 5110 18146 5285 sw
tri 18209 5165 18329 5285 ne
rect 18329 5165 18365 5285
rect 18485 5165 18521 5285
rect 17916 5028 18146 5110
tri 18146 5028 18228 5110 sw
tri 18329 5028 18466 5165 ne
rect 18466 5110 18521 5165
tri 18521 5110 18696 5285 sw
tri 18759 5165 18879 5285 ne
rect 18879 5165 18915 5285
rect 19035 5165 19071 5285
rect 18466 5028 18696 5110
tri 18696 5028 18778 5110 sw
tri 18879 5028 19016 5165 ne
rect 19016 5110 19071 5165
tri 19071 5110 19246 5285 sw
tri 19309 5165 19429 5285 ne
rect 19429 5165 19465 5285
rect 19585 5183 19621 5285
tri 19621 5183 19723 5285 sw
rect 20800 5183 21800 5972
rect 19585 5165 21800 5183
rect 19016 5028 19246 5110
tri 19246 5028 19328 5110 sw
tri 19429 5028 19566 5165 ne
rect 19566 5028 21800 5165
rect -500 4872 78 5028
tri 78 4872 234 5028 sw
tri 316 4872 472 5028 ne
rect 472 4872 628 5028
tri 628 4872 784 5028 sw
tri 866 4872 1022 5028 ne
rect 1022 4872 1178 5028
tri 1178 4872 1334 5028 sw
tri 1416 4872 1572 5028 ne
rect 1572 4872 1728 5028
tri 1728 4872 1884 5028 sw
tri 1966 4872 2122 5028 ne
rect 2122 4872 2278 5028
tri 2278 4872 2434 5028 sw
tri 2516 4872 2672 5028 ne
rect 2672 4872 2828 5028
tri 2828 4872 2984 5028 sw
tri 3066 4872 3222 5028 ne
rect 3222 4872 3378 5028
tri 3378 4872 3534 5028 sw
tri 3616 4872 3772 5028 ne
rect 3772 4872 3928 5028
tri 3928 4872 4084 5028 sw
tri 4166 4872 4322 5028 ne
rect 4322 4872 4478 5028
tri 4478 4872 4634 5028 sw
tri 4716 4872 4872 5028 ne
rect 4872 4872 5028 5028
tri 5028 4872 5184 5028 sw
tri 5266 4872 5422 5028 ne
rect 5422 4872 5578 5028
tri 5578 4872 5734 5028 sw
tri 5816 4872 5972 5028 ne
rect 5972 4872 6128 5028
tri 6128 4872 6284 5028 sw
tri 6366 4872 6522 5028 ne
rect 6522 4872 6678 5028
tri 6678 4872 6834 5028 sw
tri 6916 4872 7072 5028 ne
rect 7072 4872 7228 5028
tri 7228 4872 7384 5028 sw
tri 7466 4872 7622 5028 ne
rect 7622 4872 7778 5028
tri 7778 4872 7934 5028 sw
tri 8016 4872 8172 5028 ne
rect 8172 4872 8328 5028
tri 8328 4872 8484 5028 sw
tri 8566 4872 8722 5028 ne
rect 8722 4872 8878 5028
tri 8878 4872 9034 5028 sw
tri 9116 4872 9272 5028 ne
rect 9272 4872 9428 5028
tri 9428 4872 9584 5028 sw
tri 9666 4872 9822 5028 ne
rect 9822 4872 9978 5028
tri 9978 4872 10134 5028 sw
tri 10216 4872 10372 5028 ne
rect 10372 4872 10528 5028
tri 10528 4872 10684 5028 sw
tri 10766 4872 10922 5028 ne
rect 10922 4872 11078 5028
tri 11078 4872 11234 5028 sw
tri 11316 4872 11472 5028 ne
rect 11472 4872 11628 5028
tri 11628 4872 11784 5028 sw
tri 11866 4872 12022 5028 ne
rect 12022 4872 12178 5028
tri 12178 4872 12334 5028 sw
tri 12416 4872 12572 5028 ne
rect 12572 4872 12728 5028
tri 12728 4872 12884 5028 sw
tri 12966 4872 13122 5028 ne
rect 13122 4872 13278 5028
tri 13278 4872 13434 5028 sw
tri 13516 4872 13672 5028 ne
rect 13672 4872 13828 5028
tri 13828 4872 13984 5028 sw
tri 14066 4872 14222 5028 ne
rect 14222 4872 14378 5028
tri 14378 4872 14534 5028 sw
tri 14616 4872 14772 5028 ne
rect 14772 4872 14928 5028
tri 14928 4872 15084 5028 sw
tri 15166 4872 15322 5028 ne
rect 15322 4872 15478 5028
tri 15478 4872 15634 5028 sw
tri 15716 4872 15872 5028 ne
rect 15872 4872 16028 5028
tri 16028 4872 16184 5028 sw
tri 16266 4872 16422 5028 ne
rect 16422 4872 16578 5028
tri 16578 4872 16734 5028 sw
tri 16816 4872 16972 5028 ne
rect 16972 4872 17128 5028
tri 17128 4872 17284 5028 sw
tri 17366 4872 17522 5028 ne
rect 17522 4872 17678 5028
tri 17678 4872 17834 5028 sw
tri 17916 4872 18072 5028 ne
rect 18072 4872 18228 5028
tri 18228 4872 18384 5028 sw
tri 18466 4872 18622 5028 ne
rect 18622 4872 18778 5028
tri 18778 4872 18934 5028 sw
tri 19016 4872 19172 5028 ne
rect 19172 4872 19328 5028
tri 19328 4872 19484 5028 sw
tri 19566 4872 19722 5028 ne
rect 19722 4872 21800 5028
rect -500 4735 234 4872
tri 234 4735 371 4872 sw
tri 472 4735 609 4872 ne
rect 609 4735 784 4872
tri 784 4735 921 4872 sw
tri 1022 4735 1159 4872 ne
rect 1159 4735 1334 4872
tri 1334 4735 1471 4872 sw
tri 1572 4735 1709 4872 ne
rect 1709 4735 1884 4872
tri 1884 4735 2021 4872 sw
tri 2122 4735 2259 4872 ne
rect 2259 4735 2434 4872
tri 2434 4735 2571 4872 sw
tri 2672 4735 2809 4872 ne
rect 2809 4735 2984 4872
tri 2984 4735 3121 4872 sw
tri 3222 4735 3359 4872 ne
rect 3359 4735 3534 4872
tri 3534 4735 3671 4872 sw
tri 3772 4735 3909 4872 ne
rect 3909 4735 4084 4872
tri 4084 4735 4221 4872 sw
tri 4322 4735 4459 4872 ne
rect 4459 4735 4634 4872
tri 4634 4735 4771 4872 sw
tri 4872 4735 5009 4872 ne
rect 5009 4735 5184 4872
tri 5184 4735 5321 4872 sw
tri 5422 4735 5559 4872 ne
rect 5559 4735 5734 4872
tri 5734 4735 5871 4872 sw
tri 5972 4735 6109 4872 ne
rect 6109 4735 6284 4872
tri 6284 4735 6421 4872 sw
tri 6522 4735 6659 4872 ne
rect 6659 4735 6834 4872
tri 6834 4735 6971 4872 sw
tri 7072 4735 7209 4872 ne
rect 7209 4735 7384 4872
tri 7384 4735 7521 4872 sw
tri 7622 4735 7759 4872 ne
rect 7759 4735 7934 4872
tri 7934 4735 8071 4872 sw
tri 8172 4735 8309 4872 ne
rect 8309 4735 8484 4872
tri 8484 4735 8621 4872 sw
tri 8722 4735 8859 4872 ne
rect 8859 4735 9034 4872
tri 9034 4735 9171 4872 sw
tri 9272 4735 9409 4872 ne
rect 9409 4735 9584 4872
tri 9584 4735 9721 4872 sw
tri 9822 4735 9959 4872 ne
rect 9959 4735 10134 4872
tri 10134 4735 10271 4872 sw
tri 10372 4735 10509 4872 ne
rect 10509 4735 10684 4872
tri 10684 4735 10821 4872 sw
tri 10922 4735 11059 4872 ne
rect 11059 4735 11234 4872
tri 11234 4735 11371 4872 sw
tri 11472 4735 11609 4872 ne
rect 11609 4735 11784 4872
tri 11784 4735 11921 4872 sw
tri 12022 4735 12159 4872 ne
rect 12159 4735 12334 4872
tri 12334 4735 12471 4872 sw
tri 12572 4735 12709 4872 ne
rect 12709 4735 12884 4872
tri 12884 4735 13021 4872 sw
tri 13122 4735 13259 4872 ne
rect 13259 4735 13434 4872
tri 13434 4735 13571 4872 sw
tri 13672 4735 13809 4872 ne
rect 13809 4735 13984 4872
tri 13984 4735 14121 4872 sw
tri 14222 4735 14359 4872 ne
rect 14359 4735 14534 4872
tri 14534 4735 14671 4872 sw
tri 14772 4735 14909 4872 ne
rect 14909 4735 15084 4872
tri 15084 4735 15221 4872 sw
tri 15322 4735 15459 4872 ne
rect 15459 4735 15634 4872
tri 15634 4735 15771 4872 sw
tri 15872 4735 16009 4872 ne
rect 16009 4735 16184 4872
tri 16184 4735 16321 4872 sw
tri 16422 4735 16559 4872 ne
rect 16559 4735 16734 4872
tri 16734 4735 16871 4872 sw
tri 16972 4735 17109 4872 ne
rect 17109 4735 17284 4872
tri 17284 4735 17421 4872 sw
tri 17522 4735 17659 4872 ne
rect 17659 4735 17834 4872
tri 17834 4735 17971 4872 sw
tri 18072 4735 18209 4872 ne
rect 18209 4735 18384 4872
tri 18384 4735 18521 4872 sw
tri 18622 4735 18759 4872 ne
rect 18759 4735 18934 4872
tri 18934 4735 19071 4872 sw
tri 19172 4735 19309 4872 ne
rect 19309 4735 19484 4872
tri 19484 4735 19621 4872 sw
rect -500 4717 215 4735
tri 77 4615 179 4717 ne
rect 179 4615 215 4717
rect 335 4615 371 4735
tri 179 4478 316 4615 ne
rect 316 4560 371 4615
tri 371 4560 546 4735 sw
tri 609 4615 729 4735 ne
rect 729 4615 765 4735
rect 885 4615 921 4735
rect 316 4478 546 4560
tri 546 4478 628 4560 sw
tri 729 4478 866 4615 ne
rect 866 4560 921 4615
tri 921 4560 1096 4735 sw
tri 1159 4615 1279 4735 ne
rect 1279 4615 1315 4735
rect 1435 4615 1471 4735
rect 866 4478 1096 4560
tri 1096 4478 1178 4560 sw
tri 1279 4478 1416 4615 ne
rect 1416 4560 1471 4615
tri 1471 4560 1646 4735 sw
tri 1709 4615 1829 4735 ne
rect 1829 4615 1865 4735
rect 1985 4615 2021 4735
rect 1416 4478 1646 4560
tri 1646 4478 1728 4560 sw
tri 1829 4478 1966 4615 ne
rect 1966 4560 2021 4615
tri 2021 4560 2196 4735 sw
tri 2259 4615 2379 4735 ne
rect 2379 4615 2415 4735
rect 2535 4615 2571 4735
rect 1966 4478 2196 4560
tri 2196 4478 2278 4560 sw
tri 2379 4478 2516 4615 ne
rect 2516 4560 2571 4615
tri 2571 4560 2746 4735 sw
tri 2809 4615 2929 4735 ne
rect 2929 4615 2965 4735
rect 3085 4615 3121 4735
rect 2516 4478 2746 4560
tri 2746 4478 2828 4560 sw
tri 2929 4478 3066 4615 ne
rect 3066 4560 3121 4615
tri 3121 4560 3296 4735 sw
tri 3359 4615 3479 4735 ne
rect 3479 4615 3515 4735
rect 3635 4615 3671 4735
rect 3066 4478 3296 4560
tri 3296 4478 3378 4560 sw
tri 3479 4478 3616 4615 ne
rect 3616 4560 3671 4615
tri 3671 4560 3846 4735 sw
tri 3909 4615 4029 4735 ne
rect 4029 4615 4065 4735
rect 4185 4615 4221 4735
rect 3616 4478 3846 4560
tri 3846 4478 3928 4560 sw
tri 4029 4478 4166 4615 ne
rect 4166 4560 4221 4615
tri 4221 4560 4396 4735 sw
tri 4459 4615 4579 4735 ne
rect 4579 4615 4615 4735
rect 4735 4615 4771 4735
rect 4166 4478 4396 4560
tri 4396 4478 4478 4560 sw
tri 4579 4478 4716 4615 ne
rect 4716 4560 4771 4615
tri 4771 4560 4946 4735 sw
tri 5009 4615 5129 4735 ne
rect 5129 4615 5165 4735
rect 5285 4615 5321 4735
rect 4716 4478 4946 4560
tri 4946 4478 5028 4560 sw
tri 5129 4478 5266 4615 ne
rect 5266 4560 5321 4615
tri 5321 4560 5496 4735 sw
tri 5559 4615 5679 4735 ne
rect 5679 4615 5715 4735
rect 5835 4615 5871 4735
rect 5266 4478 5496 4560
tri 5496 4478 5578 4560 sw
tri 5679 4478 5816 4615 ne
rect 5816 4560 5871 4615
tri 5871 4560 6046 4735 sw
tri 6109 4615 6229 4735 ne
rect 6229 4615 6265 4735
rect 6385 4615 6421 4735
rect 5816 4478 6046 4560
tri 6046 4478 6128 4560 sw
tri 6229 4478 6366 4615 ne
rect 6366 4560 6421 4615
tri 6421 4560 6596 4735 sw
tri 6659 4615 6779 4735 ne
rect 6779 4615 6815 4735
rect 6935 4615 6971 4735
rect 6366 4478 6596 4560
tri 6596 4478 6678 4560 sw
tri 6779 4478 6916 4615 ne
rect 6916 4560 6971 4615
tri 6971 4560 7146 4735 sw
tri 7209 4615 7329 4735 ne
rect 7329 4615 7365 4735
rect 7485 4615 7521 4735
rect 6916 4478 7146 4560
tri 7146 4478 7228 4560 sw
tri 7329 4478 7466 4615 ne
rect 7466 4560 7521 4615
tri 7521 4560 7696 4735 sw
tri 7759 4615 7879 4735 ne
rect 7879 4615 7915 4735
rect 8035 4615 8071 4735
rect 7466 4478 7696 4560
tri 7696 4478 7778 4560 sw
tri 7879 4478 8016 4615 ne
rect 8016 4560 8071 4615
tri 8071 4560 8246 4735 sw
tri 8309 4615 8429 4735 ne
rect 8429 4615 8465 4735
rect 8585 4615 8621 4735
rect 8016 4478 8246 4560
tri 8246 4478 8328 4560 sw
tri 8429 4478 8566 4615 ne
rect 8566 4560 8621 4615
tri 8621 4560 8796 4735 sw
tri 8859 4615 8979 4735 ne
rect 8979 4615 9015 4735
rect 9135 4615 9171 4735
rect 8566 4478 8796 4560
tri 8796 4478 8878 4560 sw
tri 8979 4478 9116 4615 ne
rect 9116 4560 9171 4615
tri 9171 4560 9346 4735 sw
tri 9409 4615 9529 4735 ne
rect 9529 4615 9565 4735
rect 9685 4615 9721 4735
rect 9116 4478 9346 4560
tri 9346 4478 9428 4560 sw
tri 9529 4478 9666 4615 ne
rect 9666 4560 9721 4615
tri 9721 4560 9896 4735 sw
tri 9959 4615 10079 4735 ne
rect 10079 4615 10115 4735
rect 10235 4615 10271 4735
rect 9666 4478 9896 4560
tri 9896 4478 9978 4560 sw
tri 10079 4478 10216 4615 ne
rect 10216 4560 10271 4615
tri 10271 4560 10446 4735 sw
tri 10509 4615 10629 4735 ne
rect 10629 4615 10665 4735
rect 10785 4615 10821 4735
rect 10216 4478 10446 4560
tri 10446 4478 10528 4560 sw
tri 10629 4478 10766 4615 ne
rect 10766 4560 10821 4615
tri 10821 4560 10996 4735 sw
tri 11059 4615 11179 4735 ne
rect 11179 4615 11215 4735
rect 11335 4615 11371 4735
rect 10766 4478 10996 4560
tri 10996 4478 11078 4560 sw
tri 11179 4478 11316 4615 ne
rect 11316 4560 11371 4615
tri 11371 4560 11546 4735 sw
tri 11609 4615 11729 4735 ne
rect 11729 4615 11765 4735
rect 11885 4615 11921 4735
rect 11316 4478 11546 4560
tri 11546 4478 11628 4560 sw
tri 11729 4478 11866 4615 ne
rect 11866 4560 11921 4615
tri 11921 4560 12096 4735 sw
tri 12159 4615 12279 4735 ne
rect 12279 4615 12315 4735
rect 12435 4615 12471 4735
rect 11866 4478 12096 4560
tri 12096 4478 12178 4560 sw
tri 12279 4478 12416 4615 ne
rect 12416 4560 12471 4615
tri 12471 4560 12646 4735 sw
tri 12709 4615 12829 4735 ne
rect 12829 4615 12865 4735
rect 12985 4615 13021 4735
rect 12416 4478 12646 4560
tri 12646 4478 12728 4560 sw
tri 12829 4478 12966 4615 ne
rect 12966 4560 13021 4615
tri 13021 4560 13196 4735 sw
tri 13259 4615 13379 4735 ne
rect 13379 4615 13415 4735
rect 13535 4615 13571 4735
rect 12966 4478 13196 4560
tri 13196 4478 13278 4560 sw
tri 13379 4478 13516 4615 ne
rect 13516 4560 13571 4615
tri 13571 4560 13746 4735 sw
tri 13809 4615 13929 4735 ne
rect 13929 4615 13965 4735
rect 14085 4615 14121 4735
rect 13516 4478 13746 4560
tri 13746 4478 13828 4560 sw
tri 13929 4478 14066 4615 ne
rect 14066 4560 14121 4615
tri 14121 4560 14296 4735 sw
tri 14359 4615 14479 4735 ne
rect 14479 4615 14515 4735
rect 14635 4615 14671 4735
rect 14066 4478 14296 4560
tri 14296 4478 14378 4560 sw
tri 14479 4478 14616 4615 ne
rect 14616 4560 14671 4615
tri 14671 4560 14846 4735 sw
tri 14909 4615 15029 4735 ne
rect 15029 4615 15065 4735
rect 15185 4615 15221 4735
rect 14616 4478 14846 4560
tri 14846 4478 14928 4560 sw
tri 15029 4478 15166 4615 ne
rect 15166 4560 15221 4615
tri 15221 4560 15396 4735 sw
tri 15459 4615 15579 4735 ne
rect 15579 4615 15615 4735
rect 15735 4615 15771 4735
rect 15166 4478 15396 4560
tri 15396 4478 15478 4560 sw
tri 15579 4478 15716 4615 ne
rect 15716 4560 15771 4615
tri 15771 4560 15946 4735 sw
tri 16009 4615 16129 4735 ne
rect 16129 4615 16165 4735
rect 16285 4615 16321 4735
rect 15716 4478 15946 4560
tri 15946 4478 16028 4560 sw
tri 16129 4478 16266 4615 ne
rect 16266 4560 16321 4615
tri 16321 4560 16496 4735 sw
tri 16559 4615 16679 4735 ne
rect 16679 4615 16715 4735
rect 16835 4615 16871 4735
rect 16266 4478 16496 4560
tri 16496 4478 16578 4560 sw
tri 16679 4478 16816 4615 ne
rect 16816 4560 16871 4615
tri 16871 4560 17046 4735 sw
tri 17109 4615 17229 4735 ne
rect 17229 4615 17265 4735
rect 17385 4615 17421 4735
rect 16816 4478 17046 4560
tri 17046 4478 17128 4560 sw
tri 17229 4478 17366 4615 ne
rect 17366 4560 17421 4615
tri 17421 4560 17596 4735 sw
tri 17659 4615 17779 4735 ne
rect 17779 4615 17815 4735
rect 17935 4615 17971 4735
rect 17366 4478 17596 4560
tri 17596 4478 17678 4560 sw
tri 17779 4478 17916 4615 ne
rect 17916 4560 17971 4615
tri 17971 4560 18146 4735 sw
tri 18209 4615 18329 4735 ne
rect 18329 4615 18365 4735
rect 18485 4615 18521 4735
rect 17916 4478 18146 4560
tri 18146 4478 18228 4560 sw
tri 18329 4478 18466 4615 ne
rect 18466 4560 18521 4615
tri 18521 4560 18696 4735 sw
tri 18759 4615 18879 4735 ne
rect 18879 4615 18915 4735
rect 19035 4615 19071 4735
rect 18466 4478 18696 4560
tri 18696 4478 18778 4560 sw
tri 18879 4478 19016 4615 ne
rect 19016 4560 19071 4615
tri 19071 4560 19246 4735 sw
tri 19309 4615 19429 4735 ne
rect 19429 4615 19465 4735
rect 19585 4633 19621 4735
tri 19621 4633 19723 4735 sw
rect 19585 4615 20300 4633
rect 19016 4478 19246 4560
tri 19246 4478 19328 4560 sw
tri 19429 4478 19566 4615 ne
rect 19566 4478 20300 4615
rect -2000 4322 78 4478
tri 78 4322 234 4478 sw
tri 316 4322 472 4478 ne
rect 472 4322 628 4478
tri 628 4322 784 4478 sw
tri 866 4322 1022 4478 ne
rect 1022 4322 1178 4478
tri 1178 4322 1334 4478 sw
tri 1416 4322 1572 4478 ne
rect 1572 4322 1728 4478
tri 1728 4322 1884 4478 sw
tri 1966 4322 2122 4478 ne
rect 2122 4322 2278 4478
tri 2278 4322 2434 4478 sw
tri 2516 4322 2672 4478 ne
rect 2672 4322 2828 4478
tri 2828 4322 2984 4478 sw
tri 3066 4322 3222 4478 ne
rect 3222 4322 3378 4478
tri 3378 4322 3534 4478 sw
tri 3616 4322 3772 4478 ne
rect 3772 4322 3928 4478
tri 3928 4322 4084 4478 sw
tri 4166 4322 4322 4478 ne
rect 4322 4322 4478 4478
tri 4478 4322 4634 4478 sw
tri 4716 4322 4872 4478 ne
rect 4872 4322 5028 4478
tri 5028 4322 5184 4478 sw
tri 5266 4322 5422 4478 ne
rect 5422 4322 5578 4478
tri 5578 4322 5734 4478 sw
tri 5816 4322 5972 4478 ne
rect 5972 4322 6128 4478
tri 6128 4322 6284 4478 sw
tri 6366 4322 6522 4478 ne
rect 6522 4322 6678 4478
tri 6678 4322 6834 4478 sw
tri 6916 4322 7072 4478 ne
rect 7072 4322 7228 4478
tri 7228 4322 7384 4478 sw
tri 7466 4322 7622 4478 ne
rect 7622 4322 7778 4478
tri 7778 4322 7934 4478 sw
tri 8016 4322 8172 4478 ne
rect 8172 4322 8328 4478
tri 8328 4322 8484 4478 sw
tri 8566 4322 8722 4478 ne
rect 8722 4322 8878 4478
tri 8878 4322 9034 4478 sw
tri 9116 4322 9272 4478 ne
rect 9272 4322 9428 4478
tri 9428 4322 9584 4478 sw
tri 9666 4322 9822 4478 ne
rect 9822 4322 9978 4478
tri 9978 4322 10134 4478 sw
tri 10216 4322 10372 4478 ne
rect 10372 4322 10528 4478
tri 10528 4322 10684 4478 sw
tri 10766 4322 10922 4478 ne
rect 10922 4322 11078 4478
tri 11078 4322 11234 4478 sw
tri 11316 4322 11472 4478 ne
rect 11472 4322 11628 4478
tri 11628 4322 11784 4478 sw
tri 11866 4322 12022 4478 ne
rect 12022 4322 12178 4478
tri 12178 4322 12334 4478 sw
tri 12416 4322 12572 4478 ne
rect 12572 4322 12728 4478
tri 12728 4322 12884 4478 sw
tri 12966 4322 13122 4478 ne
rect 13122 4322 13278 4478
tri 13278 4322 13434 4478 sw
tri 13516 4322 13672 4478 ne
rect 13672 4322 13828 4478
tri 13828 4322 13984 4478 sw
tri 14066 4322 14222 4478 ne
rect 14222 4322 14378 4478
tri 14378 4322 14534 4478 sw
tri 14616 4322 14772 4478 ne
rect 14772 4322 14928 4478
tri 14928 4322 15084 4478 sw
tri 15166 4322 15322 4478 ne
rect 15322 4322 15478 4478
tri 15478 4322 15634 4478 sw
tri 15716 4322 15872 4478 ne
rect 15872 4322 16028 4478
tri 16028 4322 16184 4478 sw
tri 16266 4322 16422 4478 ne
rect 16422 4322 16578 4478
tri 16578 4322 16734 4478 sw
tri 16816 4322 16972 4478 ne
rect 16972 4322 17128 4478
tri 17128 4322 17284 4478 sw
tri 17366 4322 17522 4478 ne
rect 17522 4322 17678 4478
tri 17678 4322 17834 4478 sw
tri 17916 4322 18072 4478 ne
rect 18072 4322 18228 4478
tri 18228 4322 18384 4478 sw
tri 18466 4322 18622 4478 ne
rect 18622 4322 18778 4478
tri 18778 4322 18934 4478 sw
tri 19016 4322 19172 4478 ne
rect 19172 4322 19328 4478
tri 19328 4322 19484 4478 sw
tri 19566 4322 19722 4478 ne
rect 19722 4322 20300 4478
rect -2000 4185 234 4322
tri 234 4185 371 4322 sw
tri 472 4185 609 4322 ne
rect 609 4185 784 4322
tri 784 4185 921 4322 sw
tri 1022 4185 1159 4322 ne
rect 1159 4185 1334 4322
tri 1334 4185 1471 4322 sw
tri 1572 4185 1709 4322 ne
rect 1709 4185 1884 4322
tri 1884 4185 2021 4322 sw
tri 2122 4185 2259 4322 ne
rect 2259 4185 2434 4322
tri 2434 4185 2571 4322 sw
tri 2672 4185 2809 4322 ne
rect 2809 4185 2984 4322
tri 2984 4185 3121 4322 sw
tri 3222 4185 3359 4322 ne
rect 3359 4185 3534 4322
tri 3534 4185 3671 4322 sw
tri 3772 4185 3909 4322 ne
rect 3909 4185 4084 4322
tri 4084 4185 4221 4322 sw
tri 4322 4185 4459 4322 ne
rect 4459 4185 4634 4322
tri 4634 4185 4771 4322 sw
tri 4872 4185 5009 4322 ne
rect 5009 4185 5184 4322
tri 5184 4185 5321 4322 sw
tri 5422 4185 5559 4322 ne
rect 5559 4185 5734 4322
tri 5734 4185 5871 4322 sw
tri 5972 4185 6109 4322 ne
rect 6109 4185 6284 4322
tri 6284 4185 6421 4322 sw
tri 6522 4185 6659 4322 ne
rect 6659 4185 6834 4322
tri 6834 4185 6971 4322 sw
tri 7072 4185 7209 4322 ne
rect 7209 4185 7384 4322
tri 7384 4185 7521 4322 sw
tri 7622 4185 7759 4322 ne
rect 7759 4185 7934 4322
tri 7934 4185 8071 4322 sw
tri 8172 4185 8309 4322 ne
rect 8309 4185 8484 4322
tri 8484 4185 8621 4322 sw
tri 8722 4185 8859 4322 ne
rect 8859 4185 9034 4322
tri 9034 4185 9171 4322 sw
tri 9272 4185 9409 4322 ne
rect 9409 4185 9584 4322
tri 9584 4185 9721 4322 sw
tri 9822 4185 9959 4322 ne
rect 9959 4185 10134 4322
tri 10134 4185 10271 4322 sw
tri 10372 4185 10509 4322 ne
rect 10509 4185 10684 4322
tri 10684 4185 10821 4322 sw
tri 10922 4185 11059 4322 ne
rect 11059 4185 11234 4322
tri 11234 4185 11371 4322 sw
tri 11472 4185 11609 4322 ne
rect 11609 4185 11784 4322
tri 11784 4185 11921 4322 sw
tri 12022 4185 12159 4322 ne
rect 12159 4185 12334 4322
tri 12334 4185 12471 4322 sw
tri 12572 4185 12709 4322 ne
rect 12709 4185 12884 4322
tri 12884 4185 13021 4322 sw
tri 13122 4185 13259 4322 ne
rect 13259 4185 13434 4322
tri 13434 4185 13571 4322 sw
tri 13672 4185 13809 4322 ne
rect 13809 4185 13984 4322
tri 13984 4185 14121 4322 sw
tri 14222 4185 14359 4322 ne
rect 14359 4185 14534 4322
tri 14534 4185 14671 4322 sw
tri 14772 4185 14909 4322 ne
rect 14909 4185 15084 4322
tri 15084 4185 15221 4322 sw
tri 15322 4185 15459 4322 ne
rect 15459 4185 15634 4322
tri 15634 4185 15771 4322 sw
tri 15872 4185 16009 4322 ne
rect 16009 4185 16184 4322
tri 16184 4185 16321 4322 sw
tri 16422 4185 16559 4322 ne
rect 16559 4185 16734 4322
tri 16734 4185 16871 4322 sw
tri 16972 4185 17109 4322 ne
rect 17109 4185 17284 4322
tri 17284 4185 17421 4322 sw
tri 17522 4185 17659 4322 ne
rect 17659 4185 17834 4322
tri 17834 4185 17971 4322 sw
tri 18072 4185 18209 4322 ne
rect 18209 4185 18384 4322
tri 18384 4185 18521 4322 sw
tri 18622 4185 18759 4322 ne
rect 18759 4185 18934 4322
tri 18934 4185 19071 4322 sw
tri 19172 4185 19309 4322 ne
rect 19309 4185 19484 4322
tri 19484 4185 19621 4322 sw
rect -2000 4167 215 4185
rect -2000 3378 -1000 4167
tri 77 4065 179 4167 ne
rect 179 4065 215 4167
rect 335 4065 371 4185
tri 179 3928 316 4065 ne
rect 316 4010 371 4065
tri 371 4010 546 4185 sw
tri 609 4065 729 4185 ne
rect 729 4065 765 4185
rect 885 4065 921 4185
rect 316 3928 546 4010
tri 546 3928 628 4010 sw
tri 729 3928 866 4065 ne
rect 866 4010 921 4065
tri 921 4010 1096 4185 sw
tri 1159 4065 1279 4185 ne
rect 1279 4065 1315 4185
rect 1435 4065 1471 4185
rect 866 3928 1096 4010
tri 1096 3928 1178 4010 sw
tri 1279 3928 1416 4065 ne
rect 1416 4010 1471 4065
tri 1471 4010 1646 4185 sw
tri 1709 4065 1829 4185 ne
rect 1829 4065 1865 4185
rect 1985 4065 2021 4185
rect 1416 3928 1646 4010
tri 1646 3928 1728 4010 sw
tri 1829 3928 1966 4065 ne
rect 1966 4010 2021 4065
tri 2021 4010 2196 4185 sw
tri 2259 4065 2379 4185 ne
rect 2379 4065 2415 4185
rect 2535 4065 2571 4185
rect 1966 3928 2196 4010
tri 2196 3928 2278 4010 sw
tri 2379 3928 2516 4065 ne
rect 2516 4010 2571 4065
tri 2571 4010 2746 4185 sw
tri 2809 4065 2929 4185 ne
rect 2929 4065 2965 4185
rect 3085 4065 3121 4185
rect 2516 3928 2746 4010
tri 2746 3928 2828 4010 sw
tri 2929 3928 3066 4065 ne
rect 3066 4010 3121 4065
tri 3121 4010 3296 4185 sw
tri 3359 4065 3479 4185 ne
rect 3479 4065 3515 4185
rect 3635 4065 3671 4185
rect 3066 3928 3296 4010
tri 3296 3928 3378 4010 sw
tri 3479 3928 3616 4065 ne
rect 3616 4010 3671 4065
tri 3671 4010 3846 4185 sw
tri 3909 4065 4029 4185 ne
rect 4029 4065 4065 4185
rect 4185 4065 4221 4185
rect 3616 3928 3846 4010
tri 3846 3928 3928 4010 sw
tri 4029 3928 4166 4065 ne
rect 4166 4010 4221 4065
tri 4221 4010 4396 4185 sw
tri 4459 4065 4579 4185 ne
rect 4579 4065 4615 4185
rect 4735 4065 4771 4185
rect 4166 3928 4396 4010
tri 4396 3928 4478 4010 sw
tri 4579 3928 4716 4065 ne
rect 4716 4010 4771 4065
tri 4771 4010 4946 4185 sw
tri 5009 4065 5129 4185 ne
rect 5129 4065 5165 4185
rect 5285 4065 5321 4185
rect 4716 3928 4946 4010
tri 4946 3928 5028 4010 sw
tri 5129 3928 5266 4065 ne
rect 5266 4010 5321 4065
tri 5321 4010 5496 4185 sw
tri 5559 4065 5679 4185 ne
rect 5679 4065 5715 4185
rect 5835 4065 5871 4185
rect 5266 3928 5496 4010
tri 5496 3928 5578 4010 sw
tri 5679 3928 5816 4065 ne
rect 5816 4010 5871 4065
tri 5871 4010 6046 4185 sw
tri 6109 4065 6229 4185 ne
rect 6229 4065 6265 4185
rect 6385 4065 6421 4185
rect 5816 3928 6046 4010
tri 6046 3928 6128 4010 sw
tri 6229 3928 6366 4065 ne
rect 6366 4010 6421 4065
tri 6421 4010 6596 4185 sw
tri 6659 4065 6779 4185 ne
rect 6779 4065 6815 4185
rect 6935 4065 6971 4185
rect 6366 3928 6596 4010
tri 6596 3928 6678 4010 sw
tri 6779 3928 6916 4065 ne
rect 6916 4010 6971 4065
tri 6971 4010 7146 4185 sw
tri 7209 4065 7329 4185 ne
rect 7329 4065 7365 4185
rect 7485 4065 7521 4185
rect 6916 3928 7146 4010
tri 7146 3928 7228 4010 sw
tri 7329 3928 7466 4065 ne
rect 7466 4010 7521 4065
tri 7521 4010 7696 4185 sw
tri 7759 4065 7879 4185 ne
rect 7879 4065 7915 4185
rect 8035 4065 8071 4185
rect 7466 3928 7696 4010
tri 7696 3928 7778 4010 sw
tri 7879 3928 8016 4065 ne
rect 8016 4010 8071 4065
tri 8071 4010 8246 4185 sw
tri 8309 4065 8429 4185 ne
rect 8429 4065 8465 4185
rect 8585 4065 8621 4185
rect 8016 3928 8246 4010
tri 8246 3928 8328 4010 sw
tri 8429 3928 8566 4065 ne
rect 8566 4010 8621 4065
tri 8621 4010 8796 4185 sw
tri 8859 4065 8979 4185 ne
rect 8979 4065 9015 4185
rect 9135 4065 9171 4185
rect 8566 3928 8796 4010
tri 8796 3928 8878 4010 sw
tri 8979 3928 9116 4065 ne
rect 9116 4010 9171 4065
tri 9171 4010 9346 4185 sw
tri 9409 4065 9529 4185 ne
rect 9529 4065 9565 4185
rect 9685 4065 9721 4185
rect 9116 3928 9346 4010
tri 9346 3928 9428 4010 sw
tri 9529 3928 9666 4065 ne
rect 9666 4010 9721 4065
tri 9721 4010 9896 4185 sw
tri 9959 4065 10079 4185 ne
rect 10079 4065 10115 4185
rect 10235 4065 10271 4185
rect 9666 3928 9896 4010
tri 9896 3928 9978 4010 sw
tri 10079 3928 10216 4065 ne
rect 10216 4010 10271 4065
tri 10271 4010 10446 4185 sw
tri 10509 4065 10629 4185 ne
rect 10629 4065 10665 4185
rect 10785 4065 10821 4185
rect 10216 3928 10446 4010
tri 10446 3928 10528 4010 sw
tri 10629 3928 10766 4065 ne
rect 10766 4010 10821 4065
tri 10821 4010 10996 4185 sw
tri 11059 4065 11179 4185 ne
rect 11179 4065 11215 4185
rect 11335 4065 11371 4185
rect 10766 3928 10996 4010
tri 10996 3928 11078 4010 sw
tri 11179 3928 11316 4065 ne
rect 11316 4010 11371 4065
tri 11371 4010 11546 4185 sw
tri 11609 4065 11729 4185 ne
rect 11729 4065 11765 4185
rect 11885 4065 11921 4185
rect 11316 3928 11546 4010
tri 11546 3928 11628 4010 sw
tri 11729 3928 11866 4065 ne
rect 11866 4010 11921 4065
tri 11921 4010 12096 4185 sw
tri 12159 4065 12279 4185 ne
rect 12279 4065 12315 4185
rect 12435 4065 12471 4185
rect 11866 3928 12096 4010
tri 12096 3928 12178 4010 sw
tri 12279 3928 12416 4065 ne
rect 12416 4010 12471 4065
tri 12471 4010 12646 4185 sw
tri 12709 4065 12829 4185 ne
rect 12829 4065 12865 4185
rect 12985 4065 13021 4185
rect 12416 3928 12646 4010
tri 12646 3928 12728 4010 sw
tri 12829 3928 12966 4065 ne
rect 12966 4010 13021 4065
tri 13021 4010 13196 4185 sw
tri 13259 4065 13379 4185 ne
rect 13379 4065 13415 4185
rect 13535 4065 13571 4185
rect 12966 3928 13196 4010
tri 13196 3928 13278 4010 sw
tri 13379 3928 13516 4065 ne
rect 13516 4010 13571 4065
tri 13571 4010 13746 4185 sw
tri 13809 4065 13929 4185 ne
rect 13929 4065 13965 4185
rect 14085 4065 14121 4185
rect 13516 3928 13746 4010
tri 13746 3928 13828 4010 sw
tri 13929 3928 14066 4065 ne
rect 14066 4010 14121 4065
tri 14121 4010 14296 4185 sw
tri 14359 4065 14479 4185 ne
rect 14479 4065 14515 4185
rect 14635 4065 14671 4185
rect 14066 3928 14296 4010
tri 14296 3928 14378 4010 sw
tri 14479 3928 14616 4065 ne
rect 14616 4010 14671 4065
tri 14671 4010 14846 4185 sw
tri 14909 4065 15029 4185 ne
rect 15029 4065 15065 4185
rect 15185 4065 15221 4185
rect 14616 3928 14846 4010
tri 14846 3928 14928 4010 sw
tri 15029 3928 15166 4065 ne
rect 15166 4010 15221 4065
tri 15221 4010 15396 4185 sw
tri 15459 4065 15579 4185 ne
rect 15579 4065 15615 4185
rect 15735 4065 15771 4185
rect 15166 3928 15396 4010
tri 15396 3928 15478 4010 sw
tri 15579 3928 15716 4065 ne
rect 15716 4010 15771 4065
tri 15771 4010 15946 4185 sw
tri 16009 4065 16129 4185 ne
rect 16129 4065 16165 4185
rect 16285 4065 16321 4185
rect 15716 3928 15946 4010
tri 15946 3928 16028 4010 sw
tri 16129 3928 16266 4065 ne
rect 16266 4010 16321 4065
tri 16321 4010 16496 4185 sw
tri 16559 4065 16679 4185 ne
rect 16679 4065 16715 4185
rect 16835 4065 16871 4185
rect 16266 3928 16496 4010
tri 16496 3928 16578 4010 sw
tri 16679 3928 16816 4065 ne
rect 16816 4010 16871 4065
tri 16871 4010 17046 4185 sw
tri 17109 4065 17229 4185 ne
rect 17229 4065 17265 4185
rect 17385 4065 17421 4185
rect 16816 3928 17046 4010
tri 17046 3928 17128 4010 sw
tri 17229 3928 17366 4065 ne
rect 17366 4010 17421 4065
tri 17421 4010 17596 4185 sw
tri 17659 4065 17779 4185 ne
rect 17779 4065 17815 4185
rect 17935 4065 17971 4185
rect 17366 3928 17596 4010
tri 17596 3928 17678 4010 sw
tri 17779 3928 17916 4065 ne
rect 17916 4010 17971 4065
tri 17971 4010 18146 4185 sw
tri 18209 4065 18329 4185 ne
rect 18329 4065 18365 4185
rect 18485 4065 18521 4185
rect 17916 3928 18146 4010
tri 18146 3928 18228 4010 sw
tri 18329 3928 18466 4065 ne
rect 18466 4010 18521 4065
tri 18521 4010 18696 4185 sw
tri 18759 4065 18879 4185 ne
rect 18879 4065 18915 4185
rect 19035 4065 19071 4185
rect 18466 3928 18696 4010
tri 18696 3928 18778 4010 sw
tri 18879 3928 19016 4065 ne
rect 19016 4010 19071 4065
tri 19071 4010 19246 4185 sw
tri 19309 4065 19429 4185 ne
rect 19429 4065 19465 4185
rect 19585 4083 19621 4185
tri 19621 4083 19723 4185 sw
rect 20800 4083 21800 4872
rect 19585 4065 21800 4083
rect 19016 3928 19246 4010
tri 19246 3928 19328 4010 sw
tri 19429 3928 19566 4065 ne
rect 19566 3928 21800 4065
rect -500 3772 78 3928
tri 78 3772 234 3928 sw
tri 316 3772 472 3928 ne
rect 472 3772 628 3928
tri 628 3772 784 3928 sw
tri 866 3772 1022 3928 ne
rect 1022 3772 1178 3928
tri 1178 3772 1334 3928 sw
tri 1416 3772 1572 3928 ne
rect 1572 3772 1728 3928
tri 1728 3772 1884 3928 sw
tri 1966 3772 2122 3928 ne
rect 2122 3772 2278 3928
tri 2278 3772 2434 3928 sw
tri 2516 3772 2672 3928 ne
rect 2672 3772 2828 3928
tri 2828 3772 2984 3928 sw
tri 3066 3772 3222 3928 ne
rect 3222 3772 3378 3928
tri 3378 3772 3534 3928 sw
tri 3616 3772 3772 3928 ne
rect 3772 3772 3928 3928
tri 3928 3772 4084 3928 sw
tri 4166 3772 4322 3928 ne
rect 4322 3772 4478 3928
tri 4478 3772 4634 3928 sw
tri 4716 3772 4872 3928 ne
rect 4872 3772 5028 3928
tri 5028 3772 5184 3928 sw
tri 5266 3772 5422 3928 ne
rect 5422 3772 5578 3928
tri 5578 3772 5734 3928 sw
tri 5816 3772 5972 3928 ne
rect 5972 3772 6128 3928
tri 6128 3772 6284 3928 sw
tri 6366 3772 6522 3928 ne
rect 6522 3772 6678 3928
tri 6678 3772 6834 3928 sw
tri 6916 3772 7072 3928 ne
rect 7072 3772 7228 3928
tri 7228 3772 7384 3928 sw
tri 7466 3772 7622 3928 ne
rect 7622 3772 7778 3928
tri 7778 3772 7934 3928 sw
tri 8016 3772 8172 3928 ne
rect 8172 3772 8328 3928
tri 8328 3772 8484 3928 sw
tri 8566 3772 8722 3928 ne
rect 8722 3772 8878 3928
tri 8878 3772 9034 3928 sw
tri 9116 3772 9272 3928 ne
rect 9272 3772 9428 3928
tri 9428 3772 9584 3928 sw
tri 9666 3772 9822 3928 ne
rect 9822 3772 9978 3928
tri 9978 3772 10134 3928 sw
tri 10216 3772 10372 3928 ne
rect 10372 3772 10528 3928
tri 10528 3772 10684 3928 sw
tri 10766 3772 10922 3928 ne
rect 10922 3772 11078 3928
tri 11078 3772 11234 3928 sw
tri 11316 3772 11472 3928 ne
rect 11472 3772 11628 3928
tri 11628 3772 11784 3928 sw
tri 11866 3772 12022 3928 ne
rect 12022 3772 12178 3928
tri 12178 3772 12334 3928 sw
tri 12416 3772 12572 3928 ne
rect 12572 3772 12728 3928
tri 12728 3772 12884 3928 sw
tri 12966 3772 13122 3928 ne
rect 13122 3772 13278 3928
tri 13278 3772 13434 3928 sw
tri 13516 3772 13672 3928 ne
rect 13672 3772 13828 3928
tri 13828 3772 13984 3928 sw
tri 14066 3772 14222 3928 ne
rect 14222 3772 14378 3928
tri 14378 3772 14534 3928 sw
tri 14616 3772 14772 3928 ne
rect 14772 3772 14928 3928
tri 14928 3772 15084 3928 sw
tri 15166 3772 15322 3928 ne
rect 15322 3772 15478 3928
tri 15478 3772 15634 3928 sw
tri 15716 3772 15872 3928 ne
rect 15872 3772 16028 3928
tri 16028 3772 16184 3928 sw
tri 16266 3772 16422 3928 ne
rect 16422 3772 16578 3928
tri 16578 3772 16734 3928 sw
tri 16816 3772 16972 3928 ne
rect 16972 3772 17128 3928
tri 17128 3772 17284 3928 sw
tri 17366 3772 17522 3928 ne
rect 17522 3772 17678 3928
tri 17678 3772 17834 3928 sw
tri 17916 3772 18072 3928 ne
rect 18072 3772 18228 3928
tri 18228 3772 18384 3928 sw
tri 18466 3772 18622 3928 ne
rect 18622 3772 18778 3928
tri 18778 3772 18934 3928 sw
tri 19016 3772 19172 3928 ne
rect 19172 3772 19328 3928
tri 19328 3772 19484 3928 sw
tri 19566 3772 19722 3928 ne
rect 19722 3772 21800 3928
rect -500 3635 234 3772
tri 234 3635 371 3772 sw
tri 472 3635 609 3772 ne
rect 609 3635 784 3772
tri 784 3635 921 3772 sw
tri 1022 3635 1159 3772 ne
rect 1159 3635 1334 3772
tri 1334 3635 1471 3772 sw
tri 1572 3635 1709 3772 ne
rect 1709 3635 1884 3772
tri 1884 3635 2021 3772 sw
tri 2122 3635 2259 3772 ne
rect 2259 3635 2434 3772
tri 2434 3635 2571 3772 sw
tri 2672 3635 2809 3772 ne
rect 2809 3635 2984 3772
tri 2984 3635 3121 3772 sw
tri 3222 3635 3359 3772 ne
rect 3359 3635 3534 3772
tri 3534 3635 3671 3772 sw
tri 3772 3635 3909 3772 ne
rect 3909 3635 4084 3772
tri 4084 3635 4221 3772 sw
tri 4322 3635 4459 3772 ne
rect 4459 3635 4634 3772
tri 4634 3635 4771 3772 sw
tri 4872 3635 5009 3772 ne
rect 5009 3635 5184 3772
tri 5184 3635 5321 3772 sw
tri 5422 3635 5559 3772 ne
rect 5559 3635 5734 3772
tri 5734 3635 5871 3772 sw
tri 5972 3635 6109 3772 ne
rect 6109 3635 6284 3772
tri 6284 3635 6421 3772 sw
tri 6522 3635 6659 3772 ne
rect 6659 3635 6834 3772
tri 6834 3635 6971 3772 sw
tri 7072 3635 7209 3772 ne
rect 7209 3635 7384 3772
tri 7384 3635 7521 3772 sw
tri 7622 3635 7759 3772 ne
rect 7759 3635 7934 3772
tri 7934 3635 8071 3772 sw
tri 8172 3635 8309 3772 ne
rect 8309 3635 8484 3772
tri 8484 3635 8621 3772 sw
tri 8722 3635 8859 3772 ne
rect 8859 3635 9034 3772
tri 9034 3635 9171 3772 sw
tri 9272 3635 9409 3772 ne
rect 9409 3635 9584 3772
tri 9584 3635 9721 3772 sw
tri 9822 3635 9959 3772 ne
rect 9959 3635 10134 3772
tri 10134 3635 10271 3772 sw
tri 10372 3635 10509 3772 ne
rect 10509 3635 10684 3772
tri 10684 3635 10821 3772 sw
tri 10922 3635 11059 3772 ne
rect 11059 3635 11234 3772
tri 11234 3635 11371 3772 sw
tri 11472 3635 11609 3772 ne
rect 11609 3635 11784 3772
tri 11784 3635 11921 3772 sw
tri 12022 3635 12159 3772 ne
rect 12159 3635 12334 3772
tri 12334 3635 12471 3772 sw
tri 12572 3635 12709 3772 ne
rect 12709 3635 12884 3772
tri 12884 3635 13021 3772 sw
tri 13122 3635 13259 3772 ne
rect 13259 3635 13434 3772
tri 13434 3635 13571 3772 sw
tri 13672 3635 13809 3772 ne
rect 13809 3635 13984 3772
tri 13984 3635 14121 3772 sw
tri 14222 3635 14359 3772 ne
rect 14359 3635 14534 3772
tri 14534 3635 14671 3772 sw
tri 14772 3635 14909 3772 ne
rect 14909 3635 15084 3772
tri 15084 3635 15221 3772 sw
tri 15322 3635 15459 3772 ne
rect 15459 3635 15634 3772
tri 15634 3635 15771 3772 sw
tri 15872 3635 16009 3772 ne
rect 16009 3635 16184 3772
tri 16184 3635 16321 3772 sw
tri 16422 3635 16559 3772 ne
rect 16559 3635 16734 3772
tri 16734 3635 16871 3772 sw
tri 16972 3635 17109 3772 ne
rect 17109 3635 17284 3772
tri 17284 3635 17421 3772 sw
tri 17522 3635 17659 3772 ne
rect 17659 3635 17834 3772
tri 17834 3635 17971 3772 sw
tri 18072 3635 18209 3772 ne
rect 18209 3635 18384 3772
tri 18384 3635 18521 3772 sw
tri 18622 3635 18759 3772 ne
rect 18759 3635 18934 3772
tri 18934 3635 19071 3772 sw
tri 19172 3635 19309 3772 ne
rect 19309 3635 19484 3772
tri 19484 3635 19621 3772 sw
rect -500 3617 215 3635
tri 77 3515 179 3617 ne
rect 179 3515 215 3617
rect 335 3515 371 3635
tri 179 3378 316 3515 ne
rect 316 3460 371 3515
tri 371 3460 546 3635 sw
tri 609 3515 729 3635 ne
rect 729 3515 765 3635
rect 885 3515 921 3635
rect 316 3378 546 3460
tri 546 3378 628 3460 sw
tri 729 3378 866 3515 ne
rect 866 3460 921 3515
tri 921 3460 1096 3635 sw
tri 1159 3515 1279 3635 ne
rect 1279 3515 1315 3635
rect 1435 3515 1471 3635
rect 866 3378 1096 3460
tri 1096 3378 1178 3460 sw
tri 1279 3378 1416 3515 ne
rect 1416 3460 1471 3515
tri 1471 3460 1646 3635 sw
tri 1709 3515 1829 3635 ne
rect 1829 3515 1865 3635
rect 1985 3515 2021 3635
rect 1416 3378 1646 3460
tri 1646 3378 1728 3460 sw
tri 1829 3378 1966 3515 ne
rect 1966 3460 2021 3515
tri 2021 3460 2196 3635 sw
tri 2259 3515 2379 3635 ne
rect 2379 3515 2415 3635
rect 2535 3515 2571 3635
rect 1966 3378 2196 3460
tri 2196 3378 2278 3460 sw
tri 2379 3378 2516 3515 ne
rect 2516 3460 2571 3515
tri 2571 3460 2746 3635 sw
tri 2809 3515 2929 3635 ne
rect 2929 3515 2965 3635
rect 3085 3515 3121 3635
rect 2516 3378 2746 3460
tri 2746 3378 2828 3460 sw
tri 2929 3378 3066 3515 ne
rect 3066 3460 3121 3515
tri 3121 3460 3296 3635 sw
tri 3359 3515 3479 3635 ne
rect 3479 3515 3515 3635
rect 3635 3515 3671 3635
rect 3066 3378 3296 3460
tri 3296 3378 3378 3460 sw
tri 3479 3378 3616 3515 ne
rect 3616 3460 3671 3515
tri 3671 3460 3846 3635 sw
tri 3909 3515 4029 3635 ne
rect 4029 3515 4065 3635
rect 4185 3515 4221 3635
rect 3616 3378 3846 3460
tri 3846 3378 3928 3460 sw
tri 4029 3378 4166 3515 ne
rect 4166 3460 4221 3515
tri 4221 3460 4396 3635 sw
tri 4459 3515 4579 3635 ne
rect 4579 3515 4615 3635
rect 4735 3515 4771 3635
rect 4166 3378 4396 3460
tri 4396 3378 4478 3460 sw
tri 4579 3378 4716 3515 ne
rect 4716 3460 4771 3515
tri 4771 3460 4946 3635 sw
tri 5009 3515 5129 3635 ne
rect 5129 3515 5165 3635
rect 5285 3515 5321 3635
rect 4716 3378 4946 3460
tri 4946 3378 5028 3460 sw
tri 5129 3378 5266 3515 ne
rect 5266 3460 5321 3515
tri 5321 3460 5496 3635 sw
tri 5559 3515 5679 3635 ne
rect 5679 3515 5715 3635
rect 5835 3515 5871 3635
rect 5266 3378 5496 3460
tri 5496 3378 5578 3460 sw
tri 5679 3378 5816 3515 ne
rect 5816 3460 5871 3515
tri 5871 3460 6046 3635 sw
tri 6109 3515 6229 3635 ne
rect 6229 3515 6265 3635
rect 6385 3515 6421 3635
rect 5816 3378 6046 3460
tri 6046 3378 6128 3460 sw
tri 6229 3378 6366 3515 ne
rect 6366 3460 6421 3515
tri 6421 3460 6596 3635 sw
tri 6659 3515 6779 3635 ne
rect 6779 3515 6815 3635
rect 6935 3515 6971 3635
rect 6366 3378 6596 3460
tri 6596 3378 6678 3460 sw
tri 6779 3378 6916 3515 ne
rect 6916 3460 6971 3515
tri 6971 3460 7146 3635 sw
tri 7209 3515 7329 3635 ne
rect 7329 3515 7365 3635
rect 7485 3515 7521 3635
rect 6916 3378 7146 3460
tri 7146 3378 7228 3460 sw
tri 7329 3378 7466 3515 ne
rect 7466 3460 7521 3515
tri 7521 3460 7696 3635 sw
tri 7759 3515 7879 3635 ne
rect 7879 3515 7915 3635
rect 8035 3515 8071 3635
rect 7466 3378 7696 3460
tri 7696 3378 7778 3460 sw
tri 7879 3378 8016 3515 ne
rect 8016 3460 8071 3515
tri 8071 3460 8246 3635 sw
tri 8309 3515 8429 3635 ne
rect 8429 3515 8465 3635
rect 8585 3515 8621 3635
rect 8016 3378 8246 3460
tri 8246 3378 8328 3460 sw
tri 8429 3378 8566 3515 ne
rect 8566 3460 8621 3515
tri 8621 3460 8796 3635 sw
tri 8859 3515 8979 3635 ne
rect 8979 3515 9015 3635
rect 9135 3515 9171 3635
rect 8566 3378 8796 3460
tri 8796 3378 8878 3460 sw
tri 8979 3378 9116 3515 ne
rect 9116 3460 9171 3515
tri 9171 3460 9346 3635 sw
tri 9409 3515 9529 3635 ne
rect 9529 3515 9565 3635
rect 9685 3515 9721 3635
rect 9116 3378 9346 3460
tri 9346 3378 9428 3460 sw
tri 9529 3378 9666 3515 ne
rect 9666 3460 9721 3515
tri 9721 3460 9896 3635 sw
tri 9959 3515 10079 3635 ne
rect 10079 3515 10115 3635
rect 10235 3515 10271 3635
rect 9666 3378 9896 3460
tri 9896 3378 9978 3460 sw
tri 10079 3378 10216 3515 ne
rect 10216 3460 10271 3515
tri 10271 3460 10446 3635 sw
tri 10509 3515 10629 3635 ne
rect 10629 3515 10665 3635
rect 10785 3515 10821 3635
rect 10216 3378 10446 3460
tri 10446 3378 10528 3460 sw
tri 10629 3378 10766 3515 ne
rect 10766 3460 10821 3515
tri 10821 3460 10996 3635 sw
tri 11059 3515 11179 3635 ne
rect 11179 3515 11215 3635
rect 11335 3515 11371 3635
rect 10766 3378 10996 3460
tri 10996 3378 11078 3460 sw
tri 11179 3378 11316 3515 ne
rect 11316 3460 11371 3515
tri 11371 3460 11546 3635 sw
tri 11609 3515 11729 3635 ne
rect 11729 3515 11765 3635
rect 11885 3515 11921 3635
rect 11316 3378 11546 3460
tri 11546 3378 11628 3460 sw
tri 11729 3378 11866 3515 ne
rect 11866 3460 11921 3515
tri 11921 3460 12096 3635 sw
tri 12159 3515 12279 3635 ne
rect 12279 3515 12315 3635
rect 12435 3515 12471 3635
rect 11866 3378 12096 3460
tri 12096 3378 12178 3460 sw
tri 12279 3378 12416 3515 ne
rect 12416 3460 12471 3515
tri 12471 3460 12646 3635 sw
tri 12709 3515 12829 3635 ne
rect 12829 3515 12865 3635
rect 12985 3515 13021 3635
rect 12416 3378 12646 3460
tri 12646 3378 12728 3460 sw
tri 12829 3378 12966 3515 ne
rect 12966 3460 13021 3515
tri 13021 3460 13196 3635 sw
tri 13259 3515 13379 3635 ne
rect 13379 3515 13415 3635
rect 13535 3515 13571 3635
rect 12966 3378 13196 3460
tri 13196 3378 13278 3460 sw
tri 13379 3378 13516 3515 ne
rect 13516 3460 13571 3515
tri 13571 3460 13746 3635 sw
tri 13809 3515 13929 3635 ne
rect 13929 3515 13965 3635
rect 14085 3515 14121 3635
rect 13516 3378 13746 3460
tri 13746 3378 13828 3460 sw
tri 13929 3378 14066 3515 ne
rect 14066 3460 14121 3515
tri 14121 3460 14296 3635 sw
tri 14359 3515 14479 3635 ne
rect 14479 3515 14515 3635
rect 14635 3515 14671 3635
rect 14066 3378 14296 3460
tri 14296 3378 14378 3460 sw
tri 14479 3378 14616 3515 ne
rect 14616 3460 14671 3515
tri 14671 3460 14846 3635 sw
tri 14909 3515 15029 3635 ne
rect 15029 3515 15065 3635
rect 15185 3515 15221 3635
rect 14616 3378 14846 3460
tri 14846 3378 14928 3460 sw
tri 15029 3378 15166 3515 ne
rect 15166 3460 15221 3515
tri 15221 3460 15396 3635 sw
tri 15459 3515 15579 3635 ne
rect 15579 3515 15615 3635
rect 15735 3515 15771 3635
rect 15166 3378 15396 3460
tri 15396 3378 15478 3460 sw
tri 15579 3378 15716 3515 ne
rect 15716 3460 15771 3515
tri 15771 3460 15946 3635 sw
tri 16009 3515 16129 3635 ne
rect 16129 3515 16165 3635
rect 16285 3515 16321 3635
rect 15716 3378 15946 3460
tri 15946 3378 16028 3460 sw
tri 16129 3378 16266 3515 ne
rect 16266 3460 16321 3515
tri 16321 3460 16496 3635 sw
tri 16559 3515 16679 3635 ne
rect 16679 3515 16715 3635
rect 16835 3515 16871 3635
rect 16266 3378 16496 3460
tri 16496 3378 16578 3460 sw
tri 16679 3378 16816 3515 ne
rect 16816 3460 16871 3515
tri 16871 3460 17046 3635 sw
tri 17109 3515 17229 3635 ne
rect 17229 3515 17265 3635
rect 17385 3515 17421 3635
rect 16816 3378 17046 3460
tri 17046 3378 17128 3460 sw
tri 17229 3378 17366 3515 ne
rect 17366 3460 17421 3515
tri 17421 3460 17596 3635 sw
tri 17659 3515 17779 3635 ne
rect 17779 3515 17815 3635
rect 17935 3515 17971 3635
rect 17366 3378 17596 3460
tri 17596 3378 17678 3460 sw
tri 17779 3378 17916 3515 ne
rect 17916 3460 17971 3515
tri 17971 3460 18146 3635 sw
tri 18209 3515 18329 3635 ne
rect 18329 3515 18365 3635
rect 18485 3515 18521 3635
rect 17916 3378 18146 3460
tri 18146 3378 18228 3460 sw
tri 18329 3378 18466 3515 ne
rect 18466 3460 18521 3515
tri 18521 3460 18696 3635 sw
tri 18759 3515 18879 3635 ne
rect 18879 3515 18915 3635
rect 19035 3515 19071 3635
rect 18466 3378 18696 3460
tri 18696 3378 18778 3460 sw
tri 18879 3378 19016 3515 ne
rect 19016 3460 19071 3515
tri 19071 3460 19246 3635 sw
tri 19309 3515 19429 3635 ne
rect 19429 3515 19465 3635
rect 19585 3533 19621 3635
tri 19621 3533 19723 3635 sw
rect 19585 3515 20300 3533
rect 19016 3378 19246 3460
tri 19246 3378 19328 3460 sw
tri 19429 3378 19566 3515 ne
rect 19566 3378 20300 3515
rect -2000 3222 78 3378
tri 78 3222 234 3378 sw
tri 316 3222 472 3378 ne
rect 472 3222 628 3378
tri 628 3222 784 3378 sw
tri 866 3222 1022 3378 ne
rect 1022 3222 1178 3378
tri 1178 3222 1334 3378 sw
tri 1416 3222 1572 3378 ne
rect 1572 3222 1728 3378
tri 1728 3222 1884 3378 sw
tri 1966 3222 2122 3378 ne
rect 2122 3222 2278 3378
tri 2278 3222 2434 3378 sw
tri 2516 3222 2672 3378 ne
rect 2672 3222 2828 3378
tri 2828 3222 2984 3378 sw
tri 3066 3222 3222 3378 ne
rect 3222 3222 3378 3378
tri 3378 3222 3534 3378 sw
tri 3616 3222 3772 3378 ne
rect 3772 3222 3928 3378
tri 3928 3222 4084 3378 sw
tri 4166 3222 4322 3378 ne
rect 4322 3222 4478 3378
tri 4478 3222 4634 3378 sw
tri 4716 3222 4872 3378 ne
rect 4872 3222 5028 3378
tri 5028 3222 5184 3378 sw
tri 5266 3222 5422 3378 ne
rect 5422 3222 5578 3378
tri 5578 3222 5734 3378 sw
tri 5816 3222 5972 3378 ne
rect 5972 3222 6128 3378
tri 6128 3222 6284 3378 sw
tri 6366 3222 6522 3378 ne
rect 6522 3222 6678 3378
tri 6678 3222 6834 3378 sw
tri 6916 3222 7072 3378 ne
rect 7072 3222 7228 3378
tri 7228 3222 7384 3378 sw
tri 7466 3222 7622 3378 ne
rect 7622 3222 7778 3378
tri 7778 3222 7934 3378 sw
tri 8016 3222 8172 3378 ne
rect 8172 3222 8328 3378
tri 8328 3222 8484 3378 sw
tri 8566 3222 8722 3378 ne
rect 8722 3222 8878 3378
tri 8878 3222 9034 3378 sw
tri 9116 3222 9272 3378 ne
rect 9272 3222 9428 3378
tri 9428 3222 9584 3378 sw
tri 9666 3222 9822 3378 ne
rect 9822 3222 9978 3378
tri 9978 3222 10134 3378 sw
tri 10216 3222 10372 3378 ne
rect 10372 3222 10528 3378
tri 10528 3222 10684 3378 sw
tri 10766 3222 10922 3378 ne
rect 10922 3222 11078 3378
tri 11078 3222 11234 3378 sw
tri 11316 3222 11472 3378 ne
rect 11472 3222 11628 3378
tri 11628 3222 11784 3378 sw
tri 11866 3222 12022 3378 ne
rect 12022 3222 12178 3378
tri 12178 3222 12334 3378 sw
tri 12416 3222 12572 3378 ne
rect 12572 3222 12728 3378
tri 12728 3222 12884 3378 sw
tri 12966 3222 13122 3378 ne
rect 13122 3222 13278 3378
tri 13278 3222 13434 3378 sw
tri 13516 3222 13672 3378 ne
rect 13672 3222 13828 3378
tri 13828 3222 13984 3378 sw
tri 14066 3222 14222 3378 ne
rect 14222 3222 14378 3378
tri 14378 3222 14534 3378 sw
tri 14616 3222 14772 3378 ne
rect 14772 3222 14928 3378
tri 14928 3222 15084 3378 sw
tri 15166 3222 15322 3378 ne
rect 15322 3222 15478 3378
tri 15478 3222 15634 3378 sw
tri 15716 3222 15872 3378 ne
rect 15872 3222 16028 3378
tri 16028 3222 16184 3378 sw
tri 16266 3222 16422 3378 ne
rect 16422 3222 16578 3378
tri 16578 3222 16734 3378 sw
tri 16816 3222 16972 3378 ne
rect 16972 3222 17128 3378
tri 17128 3222 17284 3378 sw
tri 17366 3222 17522 3378 ne
rect 17522 3222 17678 3378
tri 17678 3222 17834 3378 sw
tri 17916 3222 18072 3378 ne
rect 18072 3222 18228 3378
tri 18228 3222 18384 3378 sw
tri 18466 3222 18622 3378 ne
rect 18622 3222 18778 3378
tri 18778 3222 18934 3378 sw
tri 19016 3222 19172 3378 ne
rect 19172 3222 19328 3378
tri 19328 3222 19484 3378 sw
tri 19566 3222 19722 3378 ne
rect 19722 3222 20300 3378
rect -2000 3085 234 3222
tri 234 3085 371 3222 sw
tri 472 3085 609 3222 ne
rect 609 3085 784 3222
tri 784 3085 921 3222 sw
tri 1022 3085 1159 3222 ne
rect 1159 3085 1334 3222
tri 1334 3085 1471 3222 sw
tri 1572 3085 1709 3222 ne
rect 1709 3085 1884 3222
tri 1884 3085 2021 3222 sw
tri 2122 3085 2259 3222 ne
rect 2259 3085 2434 3222
tri 2434 3085 2571 3222 sw
tri 2672 3085 2809 3222 ne
rect 2809 3085 2984 3222
tri 2984 3085 3121 3222 sw
tri 3222 3085 3359 3222 ne
rect 3359 3085 3534 3222
tri 3534 3085 3671 3222 sw
tri 3772 3085 3909 3222 ne
rect 3909 3085 4084 3222
tri 4084 3085 4221 3222 sw
tri 4322 3085 4459 3222 ne
rect 4459 3085 4634 3222
tri 4634 3085 4771 3222 sw
tri 4872 3085 5009 3222 ne
rect 5009 3085 5184 3222
tri 5184 3085 5321 3222 sw
tri 5422 3085 5559 3222 ne
rect 5559 3085 5734 3222
tri 5734 3085 5871 3222 sw
tri 5972 3085 6109 3222 ne
rect 6109 3085 6284 3222
tri 6284 3085 6421 3222 sw
tri 6522 3085 6659 3222 ne
rect 6659 3085 6834 3222
tri 6834 3085 6971 3222 sw
tri 7072 3085 7209 3222 ne
rect 7209 3085 7384 3222
tri 7384 3085 7521 3222 sw
tri 7622 3085 7759 3222 ne
rect 7759 3085 7934 3222
tri 7934 3085 8071 3222 sw
tri 8172 3085 8309 3222 ne
rect 8309 3085 8484 3222
tri 8484 3085 8621 3222 sw
tri 8722 3085 8859 3222 ne
rect 8859 3085 9034 3222
tri 9034 3085 9171 3222 sw
tri 9272 3085 9409 3222 ne
rect 9409 3085 9584 3222
tri 9584 3085 9721 3222 sw
tri 9822 3085 9959 3222 ne
rect 9959 3085 10134 3222
tri 10134 3085 10271 3222 sw
tri 10372 3085 10509 3222 ne
rect 10509 3085 10684 3222
tri 10684 3085 10821 3222 sw
tri 10922 3085 11059 3222 ne
rect 11059 3085 11234 3222
tri 11234 3085 11371 3222 sw
tri 11472 3085 11609 3222 ne
rect 11609 3085 11784 3222
tri 11784 3085 11921 3222 sw
tri 12022 3085 12159 3222 ne
rect 12159 3085 12334 3222
tri 12334 3085 12471 3222 sw
tri 12572 3085 12709 3222 ne
rect 12709 3085 12884 3222
tri 12884 3085 13021 3222 sw
tri 13122 3085 13259 3222 ne
rect 13259 3085 13434 3222
tri 13434 3085 13571 3222 sw
tri 13672 3085 13809 3222 ne
rect 13809 3085 13984 3222
tri 13984 3085 14121 3222 sw
tri 14222 3085 14359 3222 ne
rect 14359 3085 14534 3222
tri 14534 3085 14671 3222 sw
tri 14772 3085 14909 3222 ne
rect 14909 3085 15084 3222
tri 15084 3085 15221 3222 sw
tri 15322 3085 15459 3222 ne
rect 15459 3085 15634 3222
tri 15634 3085 15771 3222 sw
tri 15872 3085 16009 3222 ne
rect 16009 3085 16184 3222
tri 16184 3085 16321 3222 sw
tri 16422 3085 16559 3222 ne
rect 16559 3085 16734 3222
tri 16734 3085 16871 3222 sw
tri 16972 3085 17109 3222 ne
rect 17109 3085 17284 3222
tri 17284 3085 17421 3222 sw
tri 17522 3085 17659 3222 ne
rect 17659 3085 17834 3222
tri 17834 3085 17971 3222 sw
tri 18072 3085 18209 3222 ne
rect 18209 3085 18384 3222
tri 18384 3085 18521 3222 sw
tri 18622 3085 18759 3222 ne
rect 18759 3085 18934 3222
tri 18934 3085 19071 3222 sw
tri 19172 3085 19309 3222 ne
rect 19309 3085 19484 3222
tri 19484 3085 19621 3222 sw
rect -2000 3067 215 3085
rect -2000 2278 -1000 3067
tri 77 2965 179 3067 ne
rect 179 2965 215 3067
rect 335 2965 371 3085
tri 179 2828 316 2965 ne
rect 316 2910 371 2965
tri 371 2910 546 3085 sw
tri 609 2965 729 3085 ne
rect 729 2965 765 3085
rect 885 2965 921 3085
rect 316 2828 546 2910
tri 546 2828 628 2910 sw
tri 729 2828 866 2965 ne
rect 866 2910 921 2965
tri 921 2910 1096 3085 sw
tri 1159 2965 1279 3085 ne
rect 1279 2965 1315 3085
rect 1435 2965 1471 3085
rect 866 2828 1096 2910
tri 1096 2828 1178 2910 sw
tri 1279 2828 1416 2965 ne
rect 1416 2910 1471 2965
tri 1471 2910 1646 3085 sw
tri 1709 2965 1829 3085 ne
rect 1829 2965 1865 3085
rect 1985 2965 2021 3085
rect 1416 2828 1646 2910
tri 1646 2828 1728 2910 sw
tri 1829 2828 1966 2965 ne
rect 1966 2910 2021 2965
tri 2021 2910 2196 3085 sw
tri 2259 2965 2379 3085 ne
rect 2379 2965 2415 3085
rect 2535 2965 2571 3085
rect 1966 2828 2196 2910
tri 2196 2828 2278 2910 sw
tri 2379 2828 2516 2965 ne
rect 2516 2910 2571 2965
tri 2571 2910 2746 3085 sw
tri 2809 2965 2929 3085 ne
rect 2929 2965 2965 3085
rect 3085 2965 3121 3085
rect 2516 2828 2746 2910
tri 2746 2828 2828 2910 sw
tri 2929 2828 3066 2965 ne
rect 3066 2910 3121 2965
tri 3121 2910 3296 3085 sw
tri 3359 2965 3479 3085 ne
rect 3479 2965 3515 3085
rect 3635 2965 3671 3085
rect 3066 2828 3296 2910
tri 3296 2828 3378 2910 sw
tri 3479 2828 3616 2965 ne
rect 3616 2910 3671 2965
tri 3671 2910 3846 3085 sw
tri 3909 2965 4029 3085 ne
rect 4029 2965 4065 3085
rect 4185 2965 4221 3085
rect 3616 2828 3846 2910
tri 3846 2828 3928 2910 sw
tri 4029 2828 4166 2965 ne
rect 4166 2910 4221 2965
tri 4221 2910 4396 3085 sw
tri 4459 2965 4579 3085 ne
rect 4579 2965 4615 3085
rect 4735 2965 4771 3085
rect 4166 2828 4396 2910
tri 4396 2828 4478 2910 sw
tri 4579 2828 4716 2965 ne
rect 4716 2910 4771 2965
tri 4771 2910 4946 3085 sw
tri 5009 2965 5129 3085 ne
rect 5129 2965 5165 3085
rect 5285 2965 5321 3085
rect 4716 2828 4946 2910
tri 4946 2828 5028 2910 sw
tri 5129 2828 5266 2965 ne
rect 5266 2910 5321 2965
tri 5321 2910 5496 3085 sw
tri 5559 2965 5679 3085 ne
rect 5679 2965 5715 3085
rect 5835 2965 5871 3085
rect 5266 2828 5496 2910
tri 5496 2828 5578 2910 sw
tri 5679 2828 5816 2965 ne
rect 5816 2910 5871 2965
tri 5871 2910 6046 3085 sw
tri 6109 2965 6229 3085 ne
rect 6229 2965 6265 3085
rect 6385 2965 6421 3085
rect 5816 2828 6046 2910
tri 6046 2828 6128 2910 sw
tri 6229 2828 6366 2965 ne
rect 6366 2910 6421 2965
tri 6421 2910 6596 3085 sw
tri 6659 2965 6779 3085 ne
rect 6779 2965 6815 3085
rect 6935 2965 6971 3085
rect 6366 2828 6596 2910
tri 6596 2828 6678 2910 sw
tri 6779 2828 6916 2965 ne
rect 6916 2910 6971 2965
tri 6971 2910 7146 3085 sw
tri 7209 2965 7329 3085 ne
rect 7329 2965 7365 3085
rect 7485 2965 7521 3085
rect 6916 2828 7146 2910
tri 7146 2828 7228 2910 sw
tri 7329 2828 7466 2965 ne
rect 7466 2910 7521 2965
tri 7521 2910 7696 3085 sw
tri 7759 2965 7879 3085 ne
rect 7879 2965 7915 3085
rect 8035 2965 8071 3085
rect 7466 2828 7696 2910
tri 7696 2828 7778 2910 sw
tri 7879 2828 8016 2965 ne
rect 8016 2910 8071 2965
tri 8071 2910 8246 3085 sw
tri 8309 2965 8429 3085 ne
rect 8429 2965 8465 3085
rect 8585 2965 8621 3085
rect 8016 2828 8246 2910
tri 8246 2828 8328 2910 sw
tri 8429 2828 8566 2965 ne
rect 8566 2910 8621 2965
tri 8621 2910 8796 3085 sw
tri 8859 2965 8979 3085 ne
rect 8979 2965 9015 3085
rect 9135 2965 9171 3085
rect 8566 2828 8796 2910
tri 8796 2828 8878 2910 sw
tri 8979 2828 9116 2965 ne
rect 9116 2910 9171 2965
tri 9171 2910 9346 3085 sw
tri 9409 2965 9529 3085 ne
rect 9529 2965 9565 3085
rect 9685 2965 9721 3085
rect 9116 2828 9346 2910
tri 9346 2828 9428 2910 sw
tri 9529 2828 9666 2965 ne
rect 9666 2910 9721 2965
tri 9721 2910 9896 3085 sw
tri 9959 2965 10079 3085 ne
rect 10079 2965 10115 3085
rect 10235 2965 10271 3085
rect 9666 2828 9896 2910
tri 9896 2828 9978 2910 sw
tri 10079 2828 10216 2965 ne
rect 10216 2910 10271 2965
tri 10271 2910 10446 3085 sw
tri 10509 2965 10629 3085 ne
rect 10629 2965 10665 3085
rect 10785 2965 10821 3085
rect 10216 2828 10446 2910
tri 10446 2828 10528 2910 sw
tri 10629 2828 10766 2965 ne
rect 10766 2910 10821 2965
tri 10821 2910 10996 3085 sw
tri 11059 2965 11179 3085 ne
rect 11179 2965 11215 3085
rect 11335 2965 11371 3085
rect 10766 2828 10996 2910
tri 10996 2828 11078 2910 sw
tri 11179 2828 11316 2965 ne
rect 11316 2910 11371 2965
tri 11371 2910 11546 3085 sw
tri 11609 2965 11729 3085 ne
rect 11729 2965 11765 3085
rect 11885 2965 11921 3085
rect 11316 2828 11546 2910
tri 11546 2828 11628 2910 sw
tri 11729 2828 11866 2965 ne
rect 11866 2910 11921 2965
tri 11921 2910 12096 3085 sw
tri 12159 2965 12279 3085 ne
rect 12279 2965 12315 3085
rect 12435 2965 12471 3085
rect 11866 2828 12096 2910
tri 12096 2828 12178 2910 sw
tri 12279 2828 12416 2965 ne
rect 12416 2910 12471 2965
tri 12471 2910 12646 3085 sw
tri 12709 2965 12829 3085 ne
rect 12829 2965 12865 3085
rect 12985 2965 13021 3085
rect 12416 2828 12646 2910
tri 12646 2828 12728 2910 sw
tri 12829 2828 12966 2965 ne
rect 12966 2910 13021 2965
tri 13021 2910 13196 3085 sw
tri 13259 2965 13379 3085 ne
rect 13379 2965 13415 3085
rect 13535 2965 13571 3085
rect 12966 2828 13196 2910
tri 13196 2828 13278 2910 sw
tri 13379 2828 13516 2965 ne
rect 13516 2910 13571 2965
tri 13571 2910 13746 3085 sw
tri 13809 2965 13929 3085 ne
rect 13929 2965 13965 3085
rect 14085 2965 14121 3085
rect 13516 2828 13746 2910
tri 13746 2828 13828 2910 sw
tri 13929 2828 14066 2965 ne
rect 14066 2910 14121 2965
tri 14121 2910 14296 3085 sw
tri 14359 2965 14479 3085 ne
rect 14479 2965 14515 3085
rect 14635 2965 14671 3085
rect 14066 2828 14296 2910
tri 14296 2828 14378 2910 sw
tri 14479 2828 14616 2965 ne
rect 14616 2910 14671 2965
tri 14671 2910 14846 3085 sw
tri 14909 2965 15029 3085 ne
rect 15029 2965 15065 3085
rect 15185 2965 15221 3085
rect 14616 2828 14846 2910
tri 14846 2828 14928 2910 sw
tri 15029 2828 15166 2965 ne
rect 15166 2910 15221 2965
tri 15221 2910 15396 3085 sw
tri 15459 2965 15579 3085 ne
rect 15579 2965 15615 3085
rect 15735 2965 15771 3085
rect 15166 2828 15396 2910
tri 15396 2828 15478 2910 sw
tri 15579 2828 15716 2965 ne
rect 15716 2910 15771 2965
tri 15771 2910 15946 3085 sw
tri 16009 2965 16129 3085 ne
rect 16129 2965 16165 3085
rect 16285 2965 16321 3085
rect 15716 2828 15946 2910
tri 15946 2828 16028 2910 sw
tri 16129 2828 16266 2965 ne
rect 16266 2910 16321 2965
tri 16321 2910 16496 3085 sw
tri 16559 2965 16679 3085 ne
rect 16679 2965 16715 3085
rect 16835 2965 16871 3085
rect 16266 2828 16496 2910
tri 16496 2828 16578 2910 sw
tri 16679 2828 16816 2965 ne
rect 16816 2910 16871 2965
tri 16871 2910 17046 3085 sw
tri 17109 2965 17229 3085 ne
rect 17229 2965 17265 3085
rect 17385 2965 17421 3085
rect 16816 2828 17046 2910
tri 17046 2828 17128 2910 sw
tri 17229 2828 17366 2965 ne
rect 17366 2910 17421 2965
tri 17421 2910 17596 3085 sw
tri 17659 2965 17779 3085 ne
rect 17779 2965 17815 3085
rect 17935 2965 17971 3085
rect 17366 2828 17596 2910
tri 17596 2828 17678 2910 sw
tri 17779 2828 17916 2965 ne
rect 17916 2910 17971 2965
tri 17971 2910 18146 3085 sw
tri 18209 2965 18329 3085 ne
rect 18329 2965 18365 3085
rect 18485 2965 18521 3085
rect 17916 2828 18146 2910
tri 18146 2828 18228 2910 sw
tri 18329 2828 18466 2965 ne
rect 18466 2910 18521 2965
tri 18521 2910 18696 3085 sw
tri 18759 2965 18879 3085 ne
rect 18879 2965 18915 3085
rect 19035 2965 19071 3085
rect 18466 2828 18696 2910
tri 18696 2828 18778 2910 sw
tri 18879 2828 19016 2965 ne
rect 19016 2910 19071 2965
tri 19071 2910 19246 3085 sw
tri 19309 2965 19429 3085 ne
rect 19429 2965 19465 3085
rect 19585 2983 19621 3085
tri 19621 2983 19723 3085 sw
rect 20800 2983 21800 3772
rect 19585 2965 21800 2983
rect 19016 2828 19246 2910
tri 19246 2828 19328 2910 sw
tri 19429 2828 19566 2965 ne
rect 19566 2828 21800 2965
rect -500 2672 78 2828
tri 78 2672 234 2828 sw
tri 316 2672 472 2828 ne
rect 472 2672 628 2828
tri 628 2672 784 2828 sw
tri 866 2672 1022 2828 ne
rect 1022 2672 1178 2828
tri 1178 2672 1334 2828 sw
tri 1416 2672 1572 2828 ne
rect 1572 2672 1728 2828
tri 1728 2672 1884 2828 sw
tri 1966 2672 2122 2828 ne
rect 2122 2672 2278 2828
tri 2278 2672 2434 2828 sw
tri 2516 2672 2672 2828 ne
rect 2672 2672 2828 2828
tri 2828 2672 2984 2828 sw
tri 3066 2672 3222 2828 ne
rect 3222 2672 3378 2828
tri 3378 2672 3534 2828 sw
tri 3616 2672 3772 2828 ne
rect 3772 2672 3928 2828
tri 3928 2672 4084 2828 sw
tri 4166 2672 4322 2828 ne
rect 4322 2672 4478 2828
tri 4478 2672 4634 2828 sw
tri 4716 2672 4872 2828 ne
rect 4872 2672 5028 2828
tri 5028 2672 5184 2828 sw
tri 5266 2672 5422 2828 ne
rect 5422 2672 5578 2828
tri 5578 2672 5734 2828 sw
tri 5816 2672 5972 2828 ne
rect 5972 2672 6128 2828
tri 6128 2672 6284 2828 sw
tri 6366 2672 6522 2828 ne
rect 6522 2672 6678 2828
tri 6678 2672 6834 2828 sw
tri 6916 2672 7072 2828 ne
rect 7072 2672 7228 2828
tri 7228 2672 7384 2828 sw
tri 7466 2672 7622 2828 ne
rect 7622 2672 7778 2828
tri 7778 2672 7934 2828 sw
tri 8016 2672 8172 2828 ne
rect 8172 2672 8328 2828
tri 8328 2672 8484 2828 sw
tri 8566 2672 8722 2828 ne
rect 8722 2672 8878 2828
tri 8878 2672 9034 2828 sw
tri 9116 2672 9272 2828 ne
rect 9272 2672 9428 2828
tri 9428 2672 9584 2828 sw
tri 9666 2672 9822 2828 ne
rect 9822 2672 9978 2828
tri 9978 2672 10134 2828 sw
tri 10216 2672 10372 2828 ne
rect 10372 2672 10528 2828
tri 10528 2672 10684 2828 sw
tri 10766 2672 10922 2828 ne
rect 10922 2672 11078 2828
tri 11078 2672 11234 2828 sw
tri 11316 2672 11472 2828 ne
rect 11472 2672 11628 2828
tri 11628 2672 11784 2828 sw
tri 11866 2672 12022 2828 ne
rect 12022 2672 12178 2828
tri 12178 2672 12334 2828 sw
tri 12416 2672 12572 2828 ne
rect 12572 2672 12728 2828
tri 12728 2672 12884 2828 sw
tri 12966 2672 13122 2828 ne
rect 13122 2672 13278 2828
tri 13278 2672 13434 2828 sw
tri 13516 2672 13672 2828 ne
rect 13672 2672 13828 2828
tri 13828 2672 13984 2828 sw
tri 14066 2672 14222 2828 ne
rect 14222 2672 14378 2828
tri 14378 2672 14534 2828 sw
tri 14616 2672 14772 2828 ne
rect 14772 2672 14928 2828
tri 14928 2672 15084 2828 sw
tri 15166 2672 15322 2828 ne
rect 15322 2672 15478 2828
tri 15478 2672 15634 2828 sw
tri 15716 2672 15872 2828 ne
rect 15872 2672 16028 2828
tri 16028 2672 16184 2828 sw
tri 16266 2672 16422 2828 ne
rect 16422 2672 16578 2828
tri 16578 2672 16734 2828 sw
tri 16816 2672 16972 2828 ne
rect 16972 2672 17128 2828
tri 17128 2672 17284 2828 sw
tri 17366 2672 17522 2828 ne
rect 17522 2672 17678 2828
tri 17678 2672 17834 2828 sw
tri 17916 2672 18072 2828 ne
rect 18072 2672 18228 2828
tri 18228 2672 18384 2828 sw
tri 18466 2672 18622 2828 ne
rect 18622 2672 18778 2828
tri 18778 2672 18934 2828 sw
tri 19016 2672 19172 2828 ne
rect 19172 2672 19328 2828
tri 19328 2672 19484 2828 sw
tri 19566 2672 19722 2828 ne
rect 19722 2672 21800 2828
rect -500 2535 234 2672
tri 234 2535 371 2672 sw
tri 472 2535 609 2672 ne
rect 609 2535 784 2672
tri 784 2535 921 2672 sw
tri 1022 2535 1159 2672 ne
rect 1159 2535 1334 2672
tri 1334 2535 1471 2672 sw
tri 1572 2535 1709 2672 ne
rect 1709 2535 1884 2672
tri 1884 2535 2021 2672 sw
tri 2122 2535 2259 2672 ne
rect 2259 2535 2434 2672
tri 2434 2535 2571 2672 sw
tri 2672 2535 2809 2672 ne
rect 2809 2535 2984 2672
tri 2984 2535 3121 2672 sw
tri 3222 2535 3359 2672 ne
rect 3359 2535 3534 2672
tri 3534 2535 3671 2672 sw
tri 3772 2535 3909 2672 ne
rect 3909 2535 4084 2672
tri 4084 2535 4221 2672 sw
tri 4322 2535 4459 2672 ne
rect 4459 2535 4634 2672
tri 4634 2535 4771 2672 sw
tri 4872 2535 5009 2672 ne
rect 5009 2535 5184 2672
tri 5184 2535 5321 2672 sw
tri 5422 2535 5559 2672 ne
rect 5559 2535 5734 2672
tri 5734 2535 5871 2672 sw
tri 5972 2535 6109 2672 ne
rect 6109 2535 6284 2672
tri 6284 2535 6421 2672 sw
tri 6522 2535 6659 2672 ne
rect 6659 2535 6834 2672
tri 6834 2535 6971 2672 sw
tri 7072 2535 7209 2672 ne
rect 7209 2535 7384 2672
tri 7384 2535 7521 2672 sw
tri 7622 2535 7759 2672 ne
rect 7759 2535 7934 2672
tri 7934 2535 8071 2672 sw
tri 8172 2535 8309 2672 ne
rect 8309 2535 8484 2672
tri 8484 2535 8621 2672 sw
tri 8722 2535 8859 2672 ne
rect 8859 2535 9034 2672
tri 9034 2535 9171 2672 sw
tri 9272 2535 9409 2672 ne
rect 9409 2535 9584 2672
tri 9584 2535 9721 2672 sw
tri 9822 2535 9959 2672 ne
rect 9959 2535 10134 2672
tri 10134 2535 10271 2672 sw
tri 10372 2535 10509 2672 ne
rect 10509 2535 10684 2672
tri 10684 2535 10821 2672 sw
tri 10922 2535 11059 2672 ne
rect 11059 2535 11234 2672
tri 11234 2535 11371 2672 sw
tri 11472 2535 11609 2672 ne
rect 11609 2535 11784 2672
tri 11784 2535 11921 2672 sw
tri 12022 2535 12159 2672 ne
rect 12159 2535 12334 2672
tri 12334 2535 12471 2672 sw
tri 12572 2535 12709 2672 ne
rect 12709 2535 12884 2672
tri 12884 2535 13021 2672 sw
tri 13122 2535 13259 2672 ne
rect 13259 2535 13434 2672
tri 13434 2535 13571 2672 sw
tri 13672 2535 13809 2672 ne
rect 13809 2535 13984 2672
tri 13984 2535 14121 2672 sw
tri 14222 2535 14359 2672 ne
rect 14359 2535 14534 2672
tri 14534 2535 14671 2672 sw
tri 14772 2535 14909 2672 ne
rect 14909 2535 15084 2672
tri 15084 2535 15221 2672 sw
tri 15322 2535 15459 2672 ne
rect 15459 2535 15634 2672
tri 15634 2535 15771 2672 sw
tri 15872 2535 16009 2672 ne
rect 16009 2535 16184 2672
tri 16184 2535 16321 2672 sw
tri 16422 2535 16559 2672 ne
rect 16559 2535 16734 2672
tri 16734 2535 16871 2672 sw
tri 16972 2535 17109 2672 ne
rect 17109 2535 17284 2672
tri 17284 2535 17421 2672 sw
tri 17522 2535 17659 2672 ne
rect 17659 2535 17834 2672
tri 17834 2535 17971 2672 sw
tri 18072 2535 18209 2672 ne
rect 18209 2535 18384 2672
tri 18384 2535 18521 2672 sw
tri 18622 2535 18759 2672 ne
rect 18759 2535 18934 2672
tri 18934 2535 19071 2672 sw
tri 19172 2535 19309 2672 ne
rect 19309 2535 19484 2672
tri 19484 2535 19621 2672 sw
rect -500 2517 215 2535
tri 77 2415 179 2517 ne
rect 179 2415 215 2517
rect 335 2415 371 2535
tri 179 2278 316 2415 ne
rect 316 2360 371 2415
tri 371 2360 546 2535 sw
tri 609 2415 729 2535 ne
rect 729 2415 765 2535
rect 885 2415 921 2535
rect 316 2278 546 2360
tri 546 2278 628 2360 sw
tri 729 2278 866 2415 ne
rect 866 2360 921 2415
tri 921 2360 1096 2535 sw
tri 1159 2415 1279 2535 ne
rect 1279 2415 1315 2535
rect 1435 2415 1471 2535
rect 866 2278 1096 2360
tri 1096 2278 1178 2360 sw
tri 1279 2278 1416 2415 ne
rect 1416 2360 1471 2415
tri 1471 2360 1646 2535 sw
tri 1709 2415 1829 2535 ne
rect 1829 2415 1865 2535
rect 1985 2415 2021 2535
rect 1416 2278 1646 2360
tri 1646 2278 1728 2360 sw
tri 1829 2278 1966 2415 ne
rect 1966 2360 2021 2415
tri 2021 2360 2196 2535 sw
tri 2259 2415 2379 2535 ne
rect 2379 2415 2415 2535
rect 2535 2415 2571 2535
rect 1966 2278 2196 2360
tri 2196 2278 2278 2360 sw
tri 2379 2278 2516 2415 ne
rect 2516 2360 2571 2415
tri 2571 2360 2746 2535 sw
tri 2809 2415 2929 2535 ne
rect 2929 2415 2965 2535
rect 3085 2415 3121 2535
rect 2516 2278 2746 2360
tri 2746 2278 2828 2360 sw
tri 2929 2278 3066 2415 ne
rect 3066 2360 3121 2415
tri 3121 2360 3296 2535 sw
tri 3359 2415 3479 2535 ne
rect 3479 2415 3515 2535
rect 3635 2415 3671 2535
rect 3066 2278 3296 2360
tri 3296 2278 3378 2360 sw
tri 3479 2278 3616 2415 ne
rect 3616 2360 3671 2415
tri 3671 2360 3846 2535 sw
tri 3909 2415 4029 2535 ne
rect 4029 2415 4065 2535
rect 4185 2415 4221 2535
rect 3616 2278 3846 2360
tri 3846 2278 3928 2360 sw
tri 4029 2278 4166 2415 ne
rect 4166 2360 4221 2415
tri 4221 2360 4396 2535 sw
tri 4459 2415 4579 2535 ne
rect 4579 2415 4615 2535
rect 4735 2415 4771 2535
rect 4166 2278 4396 2360
tri 4396 2278 4478 2360 sw
tri 4579 2278 4716 2415 ne
rect 4716 2360 4771 2415
tri 4771 2360 4946 2535 sw
tri 5009 2415 5129 2535 ne
rect 5129 2415 5165 2535
rect 5285 2415 5321 2535
rect 4716 2278 4946 2360
tri 4946 2278 5028 2360 sw
tri 5129 2278 5266 2415 ne
rect 5266 2360 5321 2415
tri 5321 2360 5496 2535 sw
tri 5559 2415 5679 2535 ne
rect 5679 2415 5715 2535
rect 5835 2415 5871 2535
rect 5266 2278 5496 2360
tri 5496 2278 5578 2360 sw
tri 5679 2278 5816 2415 ne
rect 5816 2360 5871 2415
tri 5871 2360 6046 2535 sw
tri 6109 2415 6229 2535 ne
rect 6229 2415 6265 2535
rect 6385 2415 6421 2535
rect 5816 2278 6046 2360
tri 6046 2278 6128 2360 sw
tri 6229 2278 6366 2415 ne
rect 6366 2360 6421 2415
tri 6421 2360 6596 2535 sw
tri 6659 2415 6779 2535 ne
rect 6779 2415 6815 2535
rect 6935 2415 6971 2535
rect 6366 2278 6596 2360
tri 6596 2278 6678 2360 sw
tri 6779 2278 6916 2415 ne
rect 6916 2360 6971 2415
tri 6971 2360 7146 2535 sw
tri 7209 2415 7329 2535 ne
rect 7329 2415 7365 2535
rect 7485 2415 7521 2535
rect 6916 2278 7146 2360
tri 7146 2278 7228 2360 sw
tri 7329 2278 7466 2415 ne
rect 7466 2360 7521 2415
tri 7521 2360 7696 2535 sw
tri 7759 2415 7879 2535 ne
rect 7879 2415 7915 2535
rect 8035 2415 8071 2535
rect 7466 2278 7696 2360
tri 7696 2278 7778 2360 sw
tri 7879 2278 8016 2415 ne
rect 8016 2360 8071 2415
tri 8071 2360 8246 2535 sw
tri 8309 2415 8429 2535 ne
rect 8429 2415 8465 2535
rect 8585 2415 8621 2535
rect 8016 2278 8246 2360
tri 8246 2278 8328 2360 sw
tri 8429 2278 8566 2415 ne
rect 8566 2360 8621 2415
tri 8621 2360 8796 2535 sw
tri 8859 2415 8979 2535 ne
rect 8979 2415 9015 2535
rect 9135 2415 9171 2535
rect 8566 2278 8796 2360
tri 8796 2278 8878 2360 sw
tri 8979 2278 9116 2415 ne
rect 9116 2360 9171 2415
tri 9171 2360 9346 2535 sw
tri 9409 2415 9529 2535 ne
rect 9529 2415 9565 2535
rect 9685 2415 9721 2535
rect 9116 2278 9346 2360
tri 9346 2278 9428 2360 sw
tri 9529 2278 9666 2415 ne
rect 9666 2360 9721 2415
tri 9721 2360 9896 2535 sw
tri 9959 2415 10079 2535 ne
rect 10079 2415 10115 2535
rect 10235 2415 10271 2535
rect 9666 2278 9896 2360
tri 9896 2278 9978 2360 sw
tri 10079 2278 10216 2415 ne
rect 10216 2360 10271 2415
tri 10271 2360 10446 2535 sw
tri 10509 2415 10629 2535 ne
rect 10629 2415 10665 2535
rect 10785 2415 10821 2535
rect 10216 2278 10446 2360
tri 10446 2278 10528 2360 sw
tri 10629 2278 10766 2415 ne
rect 10766 2360 10821 2415
tri 10821 2360 10996 2535 sw
tri 11059 2415 11179 2535 ne
rect 11179 2415 11215 2535
rect 11335 2415 11371 2535
rect 10766 2278 10996 2360
tri 10996 2278 11078 2360 sw
tri 11179 2278 11316 2415 ne
rect 11316 2360 11371 2415
tri 11371 2360 11546 2535 sw
tri 11609 2415 11729 2535 ne
rect 11729 2415 11765 2535
rect 11885 2415 11921 2535
rect 11316 2278 11546 2360
tri 11546 2278 11628 2360 sw
tri 11729 2278 11866 2415 ne
rect 11866 2360 11921 2415
tri 11921 2360 12096 2535 sw
tri 12159 2415 12279 2535 ne
rect 12279 2415 12315 2535
rect 12435 2415 12471 2535
rect 11866 2278 12096 2360
tri 12096 2278 12178 2360 sw
tri 12279 2278 12416 2415 ne
rect 12416 2360 12471 2415
tri 12471 2360 12646 2535 sw
tri 12709 2415 12829 2535 ne
rect 12829 2415 12865 2535
rect 12985 2415 13021 2535
rect 12416 2278 12646 2360
tri 12646 2278 12728 2360 sw
tri 12829 2278 12966 2415 ne
rect 12966 2360 13021 2415
tri 13021 2360 13196 2535 sw
tri 13259 2415 13379 2535 ne
rect 13379 2415 13415 2535
rect 13535 2415 13571 2535
rect 12966 2278 13196 2360
tri 13196 2278 13278 2360 sw
tri 13379 2278 13516 2415 ne
rect 13516 2360 13571 2415
tri 13571 2360 13746 2535 sw
tri 13809 2415 13929 2535 ne
rect 13929 2415 13965 2535
rect 14085 2415 14121 2535
rect 13516 2278 13746 2360
tri 13746 2278 13828 2360 sw
tri 13929 2278 14066 2415 ne
rect 14066 2360 14121 2415
tri 14121 2360 14296 2535 sw
tri 14359 2415 14479 2535 ne
rect 14479 2415 14515 2535
rect 14635 2415 14671 2535
rect 14066 2278 14296 2360
tri 14296 2278 14378 2360 sw
tri 14479 2278 14616 2415 ne
rect 14616 2360 14671 2415
tri 14671 2360 14846 2535 sw
tri 14909 2415 15029 2535 ne
rect 15029 2415 15065 2535
rect 15185 2415 15221 2535
rect 14616 2278 14846 2360
tri 14846 2278 14928 2360 sw
tri 15029 2278 15166 2415 ne
rect 15166 2360 15221 2415
tri 15221 2360 15396 2535 sw
tri 15459 2415 15579 2535 ne
rect 15579 2415 15615 2535
rect 15735 2415 15771 2535
rect 15166 2278 15396 2360
tri 15396 2278 15478 2360 sw
tri 15579 2278 15716 2415 ne
rect 15716 2360 15771 2415
tri 15771 2360 15946 2535 sw
tri 16009 2415 16129 2535 ne
rect 16129 2415 16165 2535
rect 16285 2415 16321 2535
rect 15716 2278 15946 2360
tri 15946 2278 16028 2360 sw
tri 16129 2278 16266 2415 ne
rect 16266 2360 16321 2415
tri 16321 2360 16496 2535 sw
tri 16559 2415 16679 2535 ne
rect 16679 2415 16715 2535
rect 16835 2415 16871 2535
rect 16266 2278 16496 2360
tri 16496 2278 16578 2360 sw
tri 16679 2278 16816 2415 ne
rect 16816 2360 16871 2415
tri 16871 2360 17046 2535 sw
tri 17109 2415 17229 2535 ne
rect 17229 2415 17265 2535
rect 17385 2415 17421 2535
rect 16816 2278 17046 2360
tri 17046 2278 17128 2360 sw
tri 17229 2278 17366 2415 ne
rect 17366 2360 17421 2415
tri 17421 2360 17596 2535 sw
tri 17659 2415 17779 2535 ne
rect 17779 2415 17815 2535
rect 17935 2415 17971 2535
rect 17366 2278 17596 2360
tri 17596 2278 17678 2360 sw
tri 17779 2278 17916 2415 ne
rect 17916 2360 17971 2415
tri 17971 2360 18146 2535 sw
tri 18209 2415 18329 2535 ne
rect 18329 2415 18365 2535
rect 18485 2415 18521 2535
rect 17916 2278 18146 2360
tri 18146 2278 18228 2360 sw
tri 18329 2278 18466 2415 ne
rect 18466 2360 18521 2415
tri 18521 2360 18696 2535 sw
tri 18759 2415 18879 2535 ne
rect 18879 2415 18915 2535
rect 19035 2415 19071 2535
rect 18466 2278 18696 2360
tri 18696 2278 18778 2360 sw
tri 18879 2278 19016 2415 ne
rect 19016 2360 19071 2415
tri 19071 2360 19246 2535 sw
tri 19309 2415 19429 2535 ne
rect 19429 2415 19465 2535
rect 19585 2433 19621 2535
tri 19621 2433 19723 2535 sw
rect 19585 2415 20300 2433
rect 19016 2278 19246 2360
tri 19246 2278 19328 2360 sw
tri 19429 2278 19566 2415 ne
rect 19566 2278 20300 2415
rect -2000 2122 78 2278
tri 78 2122 234 2278 sw
tri 316 2122 472 2278 ne
rect 472 2122 628 2278
tri 628 2122 784 2278 sw
tri 866 2122 1022 2278 ne
rect 1022 2122 1178 2278
tri 1178 2122 1334 2278 sw
tri 1416 2122 1572 2278 ne
rect 1572 2122 1728 2278
tri 1728 2122 1884 2278 sw
tri 1966 2122 2122 2278 ne
rect 2122 2122 2278 2278
tri 2278 2122 2434 2278 sw
tri 2516 2122 2672 2278 ne
rect 2672 2122 2828 2278
tri 2828 2122 2984 2278 sw
tri 3066 2122 3222 2278 ne
rect 3222 2122 3378 2278
tri 3378 2122 3534 2278 sw
tri 3616 2122 3772 2278 ne
rect 3772 2122 3928 2278
tri 3928 2122 4084 2278 sw
tri 4166 2122 4322 2278 ne
rect 4322 2122 4478 2278
tri 4478 2122 4634 2278 sw
tri 4716 2122 4872 2278 ne
rect 4872 2122 5028 2278
tri 5028 2122 5184 2278 sw
tri 5266 2122 5422 2278 ne
rect 5422 2122 5578 2278
tri 5578 2122 5734 2278 sw
tri 5816 2122 5972 2278 ne
rect 5972 2122 6128 2278
tri 6128 2122 6284 2278 sw
tri 6366 2122 6522 2278 ne
rect 6522 2122 6678 2278
tri 6678 2122 6834 2278 sw
tri 6916 2122 7072 2278 ne
rect 7072 2122 7228 2278
tri 7228 2122 7384 2278 sw
tri 7466 2122 7622 2278 ne
rect 7622 2122 7778 2278
tri 7778 2122 7934 2278 sw
tri 8016 2122 8172 2278 ne
rect 8172 2122 8328 2278
tri 8328 2122 8484 2278 sw
tri 8566 2122 8722 2278 ne
rect 8722 2122 8878 2278
tri 8878 2122 9034 2278 sw
tri 9116 2122 9272 2278 ne
rect 9272 2122 9428 2278
tri 9428 2122 9584 2278 sw
tri 9666 2122 9822 2278 ne
rect 9822 2122 9978 2278
tri 9978 2122 10134 2278 sw
tri 10216 2122 10372 2278 ne
rect 10372 2122 10528 2278
tri 10528 2122 10684 2278 sw
tri 10766 2122 10922 2278 ne
rect 10922 2122 11078 2278
tri 11078 2122 11234 2278 sw
tri 11316 2122 11472 2278 ne
rect 11472 2122 11628 2278
tri 11628 2122 11784 2278 sw
tri 11866 2122 12022 2278 ne
rect 12022 2122 12178 2278
tri 12178 2122 12334 2278 sw
tri 12416 2122 12572 2278 ne
rect 12572 2122 12728 2278
tri 12728 2122 12884 2278 sw
tri 12966 2122 13122 2278 ne
rect 13122 2122 13278 2278
tri 13278 2122 13434 2278 sw
tri 13516 2122 13672 2278 ne
rect 13672 2122 13828 2278
tri 13828 2122 13984 2278 sw
tri 14066 2122 14222 2278 ne
rect 14222 2122 14378 2278
tri 14378 2122 14534 2278 sw
tri 14616 2122 14772 2278 ne
rect 14772 2122 14928 2278
tri 14928 2122 15084 2278 sw
tri 15166 2122 15322 2278 ne
rect 15322 2122 15478 2278
tri 15478 2122 15634 2278 sw
tri 15716 2122 15872 2278 ne
rect 15872 2122 16028 2278
tri 16028 2122 16184 2278 sw
tri 16266 2122 16422 2278 ne
rect 16422 2122 16578 2278
tri 16578 2122 16734 2278 sw
tri 16816 2122 16972 2278 ne
rect 16972 2122 17128 2278
tri 17128 2122 17284 2278 sw
tri 17366 2122 17522 2278 ne
rect 17522 2122 17678 2278
tri 17678 2122 17834 2278 sw
tri 17916 2122 18072 2278 ne
rect 18072 2122 18228 2278
tri 18228 2122 18384 2278 sw
tri 18466 2122 18622 2278 ne
rect 18622 2122 18778 2278
tri 18778 2122 18934 2278 sw
tri 19016 2122 19172 2278 ne
rect 19172 2122 19328 2278
tri 19328 2122 19484 2278 sw
tri 19566 2122 19722 2278 ne
rect 19722 2122 20300 2278
rect -2000 1985 234 2122
tri 234 1985 371 2122 sw
tri 472 1985 609 2122 ne
rect 609 1985 784 2122
tri 784 1985 921 2122 sw
tri 1022 1985 1159 2122 ne
rect 1159 1985 1334 2122
tri 1334 1985 1471 2122 sw
tri 1572 1985 1709 2122 ne
rect 1709 1985 1884 2122
tri 1884 1985 2021 2122 sw
tri 2122 1985 2259 2122 ne
rect 2259 1985 2434 2122
tri 2434 1985 2571 2122 sw
tri 2672 1985 2809 2122 ne
rect 2809 1985 2984 2122
tri 2984 1985 3121 2122 sw
tri 3222 1985 3359 2122 ne
rect 3359 1985 3534 2122
tri 3534 1985 3671 2122 sw
tri 3772 1985 3909 2122 ne
rect 3909 1985 4084 2122
tri 4084 1985 4221 2122 sw
tri 4322 1985 4459 2122 ne
rect 4459 1985 4634 2122
tri 4634 1985 4771 2122 sw
tri 4872 1985 5009 2122 ne
rect 5009 1985 5184 2122
tri 5184 1985 5321 2122 sw
tri 5422 1985 5559 2122 ne
rect 5559 1985 5734 2122
tri 5734 1985 5871 2122 sw
tri 5972 1985 6109 2122 ne
rect 6109 1985 6284 2122
tri 6284 1985 6421 2122 sw
tri 6522 1985 6659 2122 ne
rect 6659 1985 6834 2122
tri 6834 1985 6971 2122 sw
tri 7072 1985 7209 2122 ne
rect 7209 1985 7384 2122
tri 7384 1985 7521 2122 sw
tri 7622 1985 7759 2122 ne
rect 7759 1985 7934 2122
tri 7934 1985 8071 2122 sw
tri 8172 1985 8309 2122 ne
rect 8309 1985 8484 2122
tri 8484 1985 8621 2122 sw
tri 8722 1985 8859 2122 ne
rect 8859 1985 9034 2122
tri 9034 1985 9171 2122 sw
tri 9272 1985 9409 2122 ne
rect 9409 1985 9584 2122
tri 9584 1985 9721 2122 sw
tri 9822 1985 9959 2122 ne
rect 9959 1985 10134 2122
tri 10134 1985 10271 2122 sw
tri 10372 1985 10509 2122 ne
rect 10509 1985 10684 2122
tri 10684 1985 10821 2122 sw
tri 10922 1985 11059 2122 ne
rect 11059 1985 11234 2122
tri 11234 1985 11371 2122 sw
tri 11472 1985 11609 2122 ne
rect 11609 1985 11784 2122
tri 11784 1985 11921 2122 sw
tri 12022 1985 12159 2122 ne
rect 12159 1985 12334 2122
tri 12334 1985 12471 2122 sw
tri 12572 1985 12709 2122 ne
rect 12709 1985 12884 2122
tri 12884 1985 13021 2122 sw
tri 13122 1985 13259 2122 ne
rect 13259 1985 13434 2122
tri 13434 1985 13571 2122 sw
tri 13672 1985 13809 2122 ne
rect 13809 1985 13984 2122
tri 13984 1985 14121 2122 sw
tri 14222 1985 14359 2122 ne
rect 14359 1985 14534 2122
tri 14534 1985 14671 2122 sw
tri 14772 1985 14909 2122 ne
rect 14909 1985 15084 2122
tri 15084 1985 15221 2122 sw
tri 15322 1985 15459 2122 ne
rect 15459 1985 15634 2122
tri 15634 1985 15771 2122 sw
tri 15872 1985 16009 2122 ne
rect 16009 1985 16184 2122
tri 16184 1985 16321 2122 sw
tri 16422 1985 16559 2122 ne
rect 16559 1985 16734 2122
tri 16734 1985 16871 2122 sw
tri 16972 1985 17109 2122 ne
rect 17109 1985 17284 2122
tri 17284 1985 17421 2122 sw
tri 17522 1985 17659 2122 ne
rect 17659 1985 17834 2122
tri 17834 1985 17971 2122 sw
tri 18072 1985 18209 2122 ne
rect 18209 1985 18384 2122
tri 18384 1985 18521 2122 sw
tri 18622 1985 18759 2122 ne
rect 18759 1985 18934 2122
tri 18934 1985 19071 2122 sw
tri 19172 1985 19309 2122 ne
rect 19309 1985 19484 2122
tri 19484 1985 19621 2122 sw
rect -2000 1967 215 1985
rect -2000 1650 -1000 1967
tri 77 1865 179 1967 ne
rect 179 1865 215 1967
rect 335 1865 371 1985
tri 179 1728 316 1865 ne
rect 316 1810 371 1865
tri 371 1810 546 1985 sw
tri 609 1865 729 1985 ne
rect 729 1865 765 1985
rect 885 1865 921 1985
rect 316 1728 546 1810
tri 546 1728 628 1810 sw
tri 729 1728 866 1865 ne
rect 866 1810 921 1865
tri 921 1810 1096 1985 sw
tri 1159 1865 1279 1985 ne
rect 1279 1865 1315 1985
rect 1435 1865 1471 1985
rect 866 1728 1096 1810
tri 1096 1728 1178 1810 sw
tri 1279 1728 1416 1865 ne
rect 1416 1810 1471 1865
tri 1471 1810 1646 1985 sw
tri 1709 1865 1829 1985 ne
rect 1829 1865 1865 1985
rect 1985 1865 2021 1985
rect 1416 1728 1646 1810
tri 1646 1728 1728 1810 sw
tri 1829 1728 1966 1865 ne
rect 1966 1810 2021 1865
tri 2021 1810 2196 1985 sw
tri 2259 1865 2379 1985 ne
rect 2379 1865 2415 1985
rect 2535 1865 2571 1985
rect 1966 1728 2196 1810
tri 2196 1728 2278 1810 sw
tri 2379 1728 2516 1865 ne
rect 2516 1810 2571 1865
tri 2571 1810 2746 1985 sw
tri 2809 1865 2929 1985 ne
rect 2929 1865 2965 1985
rect 3085 1865 3121 1985
rect 2516 1728 2746 1810
tri 2746 1728 2828 1810 sw
tri 2929 1728 3066 1865 ne
rect 3066 1810 3121 1865
tri 3121 1810 3296 1985 sw
tri 3359 1865 3479 1985 ne
rect 3479 1865 3515 1985
rect 3635 1865 3671 1985
rect 3066 1728 3296 1810
tri 3296 1728 3378 1810 sw
tri 3479 1728 3616 1865 ne
rect 3616 1810 3671 1865
tri 3671 1810 3846 1985 sw
tri 3909 1865 4029 1985 ne
rect 4029 1865 4065 1985
rect 4185 1865 4221 1985
rect 3616 1728 3846 1810
tri 3846 1728 3928 1810 sw
tri 4029 1728 4166 1865 ne
rect 4166 1810 4221 1865
tri 4221 1810 4396 1985 sw
tri 4459 1865 4579 1985 ne
rect 4579 1865 4615 1985
rect 4735 1865 4771 1985
rect 4166 1728 4396 1810
tri 4396 1728 4478 1810 sw
tri 4579 1728 4716 1865 ne
rect 4716 1810 4771 1865
tri 4771 1810 4946 1985 sw
tri 5009 1865 5129 1985 ne
rect 5129 1865 5165 1985
rect 5285 1865 5321 1985
rect 4716 1728 4946 1810
tri 4946 1728 5028 1810 sw
tri 5129 1728 5266 1865 ne
rect 5266 1810 5321 1865
tri 5321 1810 5496 1985 sw
tri 5559 1865 5679 1985 ne
rect 5679 1865 5715 1985
rect 5835 1865 5871 1985
rect 5266 1728 5496 1810
tri 5496 1728 5578 1810 sw
tri 5679 1728 5816 1865 ne
rect 5816 1810 5871 1865
tri 5871 1810 6046 1985 sw
tri 6109 1865 6229 1985 ne
rect 6229 1865 6265 1985
rect 6385 1865 6421 1985
rect 5816 1728 6046 1810
tri 6046 1728 6128 1810 sw
tri 6229 1728 6366 1865 ne
rect 6366 1810 6421 1865
tri 6421 1810 6596 1985 sw
tri 6659 1865 6779 1985 ne
rect 6779 1865 6815 1985
rect 6935 1865 6971 1985
rect 6366 1728 6596 1810
tri 6596 1728 6678 1810 sw
tri 6779 1728 6916 1865 ne
rect 6916 1810 6971 1865
tri 6971 1810 7146 1985 sw
tri 7209 1865 7329 1985 ne
rect 7329 1865 7365 1985
rect 7485 1865 7521 1985
rect 6916 1728 7146 1810
tri 7146 1728 7228 1810 sw
tri 7329 1728 7466 1865 ne
rect 7466 1810 7521 1865
tri 7521 1810 7696 1985 sw
tri 7759 1865 7879 1985 ne
rect 7879 1865 7915 1985
rect 8035 1865 8071 1985
rect 7466 1728 7696 1810
tri 7696 1728 7778 1810 sw
tri 7879 1728 8016 1865 ne
rect 8016 1810 8071 1865
tri 8071 1810 8246 1985 sw
tri 8309 1865 8429 1985 ne
rect 8429 1865 8465 1985
rect 8585 1865 8621 1985
rect 8016 1728 8246 1810
tri 8246 1728 8328 1810 sw
tri 8429 1728 8566 1865 ne
rect 8566 1810 8621 1865
tri 8621 1810 8796 1985 sw
tri 8859 1865 8979 1985 ne
rect 8979 1865 9015 1985
rect 9135 1865 9171 1985
rect 8566 1728 8796 1810
tri 8796 1728 8878 1810 sw
tri 8979 1728 9116 1865 ne
rect 9116 1810 9171 1865
tri 9171 1810 9346 1985 sw
tri 9409 1865 9529 1985 ne
rect 9529 1865 9565 1985
rect 9685 1865 9721 1985
rect 9116 1728 9346 1810
tri 9346 1728 9428 1810 sw
tri 9529 1728 9666 1865 ne
rect 9666 1810 9721 1865
tri 9721 1810 9896 1985 sw
tri 9959 1865 10079 1985 ne
rect 10079 1865 10115 1985
rect 10235 1865 10271 1985
rect 9666 1728 9896 1810
tri 9896 1728 9978 1810 sw
tri 10079 1728 10216 1865 ne
rect 10216 1810 10271 1865
tri 10271 1810 10446 1985 sw
tri 10509 1865 10629 1985 ne
rect 10629 1865 10665 1985
rect 10785 1865 10821 1985
rect 10216 1728 10446 1810
tri 10446 1728 10528 1810 sw
tri 10629 1728 10766 1865 ne
rect 10766 1810 10821 1865
tri 10821 1810 10996 1985 sw
tri 11059 1865 11179 1985 ne
rect 11179 1865 11215 1985
rect 11335 1865 11371 1985
rect 10766 1728 10996 1810
tri 10996 1728 11078 1810 sw
tri 11179 1728 11316 1865 ne
rect 11316 1810 11371 1865
tri 11371 1810 11546 1985 sw
tri 11609 1865 11729 1985 ne
rect 11729 1865 11765 1985
rect 11885 1865 11921 1985
rect 11316 1728 11546 1810
tri 11546 1728 11628 1810 sw
tri 11729 1728 11866 1865 ne
rect 11866 1810 11921 1865
tri 11921 1810 12096 1985 sw
tri 12159 1865 12279 1985 ne
rect 12279 1865 12315 1985
rect 12435 1865 12471 1985
rect 11866 1728 12096 1810
tri 12096 1728 12178 1810 sw
tri 12279 1728 12416 1865 ne
rect 12416 1810 12471 1865
tri 12471 1810 12646 1985 sw
tri 12709 1865 12829 1985 ne
rect 12829 1865 12865 1985
rect 12985 1865 13021 1985
rect 12416 1728 12646 1810
tri 12646 1728 12728 1810 sw
tri 12829 1728 12966 1865 ne
rect 12966 1810 13021 1865
tri 13021 1810 13196 1985 sw
tri 13259 1865 13379 1985 ne
rect 13379 1865 13415 1985
rect 13535 1865 13571 1985
rect 12966 1728 13196 1810
tri 13196 1728 13278 1810 sw
tri 13379 1728 13516 1865 ne
rect 13516 1810 13571 1865
tri 13571 1810 13746 1985 sw
tri 13809 1865 13929 1985 ne
rect 13929 1865 13965 1985
rect 14085 1865 14121 1985
rect 13516 1728 13746 1810
tri 13746 1728 13828 1810 sw
tri 13929 1728 14066 1865 ne
rect 14066 1810 14121 1865
tri 14121 1810 14296 1985 sw
tri 14359 1865 14479 1985 ne
rect 14479 1865 14515 1985
rect 14635 1865 14671 1985
rect 14066 1728 14296 1810
tri 14296 1728 14378 1810 sw
tri 14479 1728 14616 1865 ne
rect 14616 1810 14671 1865
tri 14671 1810 14846 1985 sw
tri 14909 1865 15029 1985 ne
rect 15029 1865 15065 1985
rect 15185 1865 15221 1985
rect 14616 1728 14846 1810
tri 14846 1728 14928 1810 sw
tri 15029 1728 15166 1865 ne
rect 15166 1810 15221 1865
tri 15221 1810 15396 1985 sw
tri 15459 1865 15579 1985 ne
rect 15579 1865 15615 1985
rect 15735 1865 15771 1985
rect 15166 1728 15396 1810
tri 15396 1728 15478 1810 sw
tri 15579 1728 15716 1865 ne
rect 15716 1810 15771 1865
tri 15771 1810 15946 1985 sw
tri 16009 1865 16129 1985 ne
rect 16129 1865 16165 1985
rect 16285 1865 16321 1985
rect 15716 1728 15946 1810
tri 15946 1728 16028 1810 sw
tri 16129 1728 16266 1865 ne
rect 16266 1810 16321 1865
tri 16321 1810 16496 1985 sw
tri 16559 1865 16679 1985 ne
rect 16679 1865 16715 1985
rect 16835 1865 16871 1985
rect 16266 1728 16496 1810
tri 16496 1728 16578 1810 sw
tri 16679 1728 16816 1865 ne
rect 16816 1810 16871 1865
tri 16871 1810 17046 1985 sw
tri 17109 1865 17229 1985 ne
rect 17229 1865 17265 1985
rect 17385 1865 17421 1985
rect 16816 1728 17046 1810
tri 17046 1728 17128 1810 sw
tri 17229 1728 17366 1865 ne
rect 17366 1810 17421 1865
tri 17421 1810 17596 1985 sw
tri 17659 1865 17779 1985 ne
rect 17779 1865 17815 1985
rect 17935 1865 17971 1985
rect 17366 1728 17596 1810
tri 17596 1728 17678 1810 sw
tri 17779 1728 17916 1865 ne
rect 17916 1810 17971 1865
tri 17971 1810 18146 1985 sw
tri 18209 1865 18329 1985 ne
rect 18329 1865 18365 1985
rect 18485 1865 18521 1985
rect 17916 1728 18146 1810
tri 18146 1728 18228 1810 sw
tri 18329 1728 18466 1865 ne
rect 18466 1810 18521 1865
tri 18521 1810 18696 1985 sw
tri 18759 1865 18879 1985 ne
rect 18879 1865 18915 1985
rect 19035 1865 19071 1985
rect 18466 1728 18696 1810
tri 18696 1728 18778 1810 sw
tri 18879 1728 19016 1865 ne
rect 19016 1810 19071 1865
tri 19071 1810 19246 1985 sw
tri 19309 1865 19429 1985 ne
rect 19429 1865 19465 1985
rect 19585 1883 19621 1985
tri 19621 1883 19723 1985 sw
rect 20800 1883 21800 2672
rect 19585 1865 21800 1883
rect 19016 1728 19246 1810
tri 19246 1728 19328 1810 sw
tri 19429 1728 19566 1865 ne
rect 19566 1728 21800 1865
rect -500 1572 78 1728
tri 78 1572 234 1728 sw
tri 316 1572 472 1728 ne
rect 472 1572 628 1728
tri 628 1572 784 1728 sw
tri 866 1572 1022 1728 ne
rect 1022 1572 1178 1728
tri 1178 1572 1334 1728 sw
tri 1416 1572 1572 1728 ne
rect 1572 1572 1728 1728
tri 1728 1572 1884 1728 sw
tri 1966 1572 2122 1728 ne
rect 2122 1572 2278 1728
tri 2278 1572 2434 1728 sw
tri 2516 1572 2672 1728 ne
rect 2672 1572 2828 1728
tri 2828 1572 2984 1728 sw
tri 3066 1572 3222 1728 ne
rect 3222 1572 3378 1728
tri 3378 1572 3534 1728 sw
tri 3616 1572 3772 1728 ne
rect 3772 1572 3928 1728
tri 3928 1572 4084 1728 sw
tri 4166 1572 4322 1728 ne
rect 4322 1572 4478 1728
tri 4478 1572 4634 1728 sw
tri 4716 1572 4872 1728 ne
rect 4872 1572 5028 1728
tri 5028 1572 5184 1728 sw
tri 5266 1572 5422 1728 ne
rect 5422 1572 5578 1728
tri 5578 1572 5734 1728 sw
tri 5816 1572 5972 1728 ne
rect 5972 1572 6128 1728
tri 6128 1572 6284 1728 sw
tri 6366 1572 6522 1728 ne
rect 6522 1572 6678 1728
tri 6678 1572 6834 1728 sw
tri 6916 1572 7072 1728 ne
rect 7072 1572 7228 1728
tri 7228 1572 7384 1728 sw
tri 7466 1572 7622 1728 ne
rect 7622 1572 7778 1728
tri 7778 1572 7934 1728 sw
tri 8016 1572 8172 1728 ne
rect 8172 1572 8328 1728
tri 8328 1572 8484 1728 sw
tri 8566 1572 8722 1728 ne
rect 8722 1572 8878 1728
tri 8878 1572 9034 1728 sw
tri 9116 1572 9272 1728 ne
rect 9272 1572 9428 1728
tri 9428 1572 9584 1728 sw
tri 9666 1572 9822 1728 ne
rect 9822 1572 9978 1728
tri 9978 1572 10134 1728 sw
tri 10216 1572 10372 1728 ne
rect 10372 1572 10528 1728
tri 10528 1572 10684 1728 sw
tri 10766 1572 10922 1728 ne
rect 10922 1572 11078 1728
tri 11078 1572 11234 1728 sw
tri 11316 1572 11472 1728 ne
rect 11472 1572 11628 1728
tri 11628 1572 11784 1728 sw
tri 11866 1572 12022 1728 ne
rect 12022 1572 12178 1728
tri 12178 1572 12334 1728 sw
tri 12416 1572 12572 1728 ne
rect 12572 1572 12728 1728
tri 12728 1572 12884 1728 sw
tri 12966 1572 13122 1728 ne
rect 13122 1572 13278 1728
tri 13278 1572 13434 1728 sw
tri 13516 1572 13672 1728 ne
rect 13672 1572 13828 1728
tri 13828 1572 13984 1728 sw
tri 14066 1572 14222 1728 ne
rect 14222 1572 14378 1728
tri 14378 1572 14534 1728 sw
tri 14616 1572 14772 1728 ne
rect 14772 1572 14928 1728
tri 14928 1572 15084 1728 sw
tri 15166 1572 15322 1728 ne
rect 15322 1572 15478 1728
tri 15478 1572 15634 1728 sw
tri 15716 1572 15872 1728 ne
rect 15872 1572 16028 1728
tri 16028 1572 16184 1728 sw
tri 16266 1572 16422 1728 ne
rect 16422 1572 16578 1728
tri 16578 1572 16734 1728 sw
tri 16816 1572 16972 1728 ne
rect 16972 1572 17128 1728
tri 17128 1572 17284 1728 sw
tri 17366 1572 17522 1728 ne
rect 17522 1572 17678 1728
tri 17678 1572 17834 1728 sw
tri 17916 1572 18072 1728 ne
rect 18072 1572 18228 1728
tri 18228 1572 18384 1728 sw
tri 18466 1572 18622 1728 ne
rect 18622 1572 18778 1728
tri 18778 1572 18934 1728 sw
tri 19016 1572 19172 1728 ne
rect 19172 1572 19328 1728
tri 19328 1572 19484 1728 sw
tri 19566 1572 19722 1728 ne
rect 19722 1572 21800 1728
rect -500 1435 234 1572
tri 234 1435 371 1572 sw
tri 472 1435 609 1572 ne
rect 609 1435 784 1572
tri 784 1435 921 1572 sw
tri 1022 1435 1159 1572 ne
rect 1159 1435 1334 1572
tri 1334 1435 1471 1572 sw
tri 1572 1435 1709 1572 ne
rect 1709 1435 1884 1572
tri 1884 1435 2021 1572 sw
tri 2122 1435 2259 1572 ne
rect 2259 1435 2434 1572
tri 2434 1435 2571 1572 sw
tri 2672 1435 2809 1572 ne
rect 2809 1435 2984 1572
tri 2984 1435 3121 1572 sw
tri 3222 1435 3359 1572 ne
rect 3359 1435 3534 1572
tri 3534 1435 3671 1572 sw
tri 3772 1435 3909 1572 ne
rect 3909 1435 4084 1572
tri 4084 1435 4221 1572 sw
tri 4322 1435 4459 1572 ne
rect 4459 1435 4634 1572
tri 4634 1435 4771 1572 sw
tri 4872 1435 5009 1572 ne
rect 5009 1435 5184 1572
tri 5184 1435 5321 1572 sw
tri 5422 1435 5559 1572 ne
rect 5559 1435 5734 1572
tri 5734 1435 5871 1572 sw
tri 5972 1435 6109 1572 ne
rect 6109 1435 6284 1572
tri 6284 1435 6421 1572 sw
tri 6522 1435 6659 1572 ne
rect 6659 1435 6834 1572
tri 6834 1435 6971 1572 sw
tri 7072 1435 7209 1572 ne
rect 7209 1435 7384 1572
tri 7384 1435 7521 1572 sw
tri 7622 1435 7759 1572 ne
rect 7759 1435 7934 1572
tri 7934 1435 8071 1572 sw
tri 8172 1435 8309 1572 ne
rect 8309 1435 8484 1572
tri 8484 1435 8621 1572 sw
tri 8722 1435 8859 1572 ne
rect 8859 1435 9034 1572
tri 9034 1435 9171 1572 sw
tri 9272 1435 9409 1572 ne
rect 9409 1435 9584 1572
tri 9584 1435 9721 1572 sw
tri 9822 1435 9959 1572 ne
rect 9959 1435 10134 1572
tri 10134 1435 10271 1572 sw
tri 10372 1435 10509 1572 ne
rect 10509 1435 10684 1572
tri 10684 1435 10821 1572 sw
tri 10922 1435 11059 1572 ne
rect 11059 1435 11234 1572
tri 11234 1435 11371 1572 sw
tri 11472 1435 11609 1572 ne
rect 11609 1435 11784 1572
tri 11784 1435 11921 1572 sw
tri 12022 1435 12159 1572 ne
rect 12159 1435 12334 1572
tri 12334 1435 12471 1572 sw
tri 12572 1435 12709 1572 ne
rect 12709 1435 12884 1572
tri 12884 1435 13021 1572 sw
tri 13122 1435 13259 1572 ne
rect 13259 1435 13434 1572
tri 13434 1435 13571 1572 sw
tri 13672 1435 13809 1572 ne
rect 13809 1435 13984 1572
tri 13984 1435 14121 1572 sw
tri 14222 1435 14359 1572 ne
rect 14359 1435 14534 1572
tri 14534 1435 14671 1572 sw
tri 14772 1435 14909 1572 ne
rect 14909 1435 15084 1572
tri 15084 1435 15221 1572 sw
tri 15322 1435 15459 1572 ne
rect 15459 1435 15634 1572
tri 15634 1435 15771 1572 sw
tri 15872 1435 16009 1572 ne
rect 16009 1435 16184 1572
tri 16184 1435 16321 1572 sw
tri 16422 1435 16559 1572 ne
rect 16559 1435 16734 1572
tri 16734 1435 16871 1572 sw
tri 16972 1435 17109 1572 ne
rect 17109 1435 17284 1572
tri 17284 1435 17421 1572 sw
tri 17522 1435 17659 1572 ne
rect 17659 1435 17834 1572
tri 17834 1435 17971 1572 sw
tri 18072 1435 18209 1572 ne
rect 18209 1435 18384 1572
tri 18384 1435 18521 1572 sw
tri 18622 1435 18759 1572 ne
rect 18759 1435 18934 1572
tri 18934 1435 19071 1572 sw
tri 19172 1435 19309 1572 ne
rect 19309 1435 19484 1572
tri 19484 1435 19621 1572 sw
rect -500 1417 215 1435
tri 77 1315 179 1417 ne
rect 179 1315 215 1417
rect 335 1315 371 1435
tri 179 1178 316 1315 ne
rect 316 1260 371 1315
tri 371 1260 546 1435 sw
tri 609 1315 729 1435 ne
rect 729 1315 765 1435
rect 885 1315 921 1435
rect 316 1178 546 1260
tri 546 1178 628 1260 sw
tri 729 1178 866 1315 ne
rect 866 1260 921 1315
tri 921 1260 1096 1435 sw
tri 1159 1315 1279 1435 ne
rect 1279 1315 1315 1435
rect 1435 1315 1471 1435
rect 866 1178 1096 1260
tri 1096 1178 1178 1260 sw
tri 1279 1178 1416 1315 ne
rect 1416 1260 1471 1315
tri 1471 1260 1646 1435 sw
tri 1709 1315 1829 1435 ne
rect 1829 1315 1865 1435
rect 1985 1315 2021 1435
rect 1416 1178 1646 1260
tri 1646 1178 1728 1260 sw
tri 1829 1178 1966 1315 ne
rect 1966 1260 2021 1315
tri 2021 1260 2196 1435 sw
tri 2259 1315 2379 1435 ne
rect 2379 1315 2415 1435
rect 2535 1315 2571 1435
rect 1966 1178 2196 1260
tri 2196 1178 2278 1260 sw
tri 2379 1178 2516 1315 ne
rect 2516 1260 2571 1315
tri 2571 1260 2746 1435 sw
tri 2809 1315 2929 1435 ne
rect 2929 1315 2965 1435
rect 3085 1315 3121 1435
rect 2516 1178 2746 1260
tri 2746 1178 2828 1260 sw
tri 2929 1178 3066 1315 ne
rect 3066 1260 3121 1315
tri 3121 1260 3296 1435 sw
tri 3359 1315 3479 1435 ne
rect 3479 1315 3515 1435
rect 3635 1315 3671 1435
rect 3066 1178 3296 1260
tri 3296 1178 3378 1260 sw
tri 3479 1178 3616 1315 ne
rect 3616 1260 3671 1315
tri 3671 1260 3846 1435 sw
tri 3909 1315 4029 1435 ne
rect 4029 1315 4065 1435
rect 4185 1315 4221 1435
rect 3616 1178 3846 1260
tri 3846 1178 3928 1260 sw
tri 4029 1178 4166 1315 ne
rect 4166 1260 4221 1315
tri 4221 1260 4396 1435 sw
tri 4459 1315 4579 1435 ne
rect 4579 1315 4615 1435
rect 4735 1315 4771 1435
rect 4166 1178 4396 1260
tri 4396 1178 4478 1260 sw
tri 4579 1178 4716 1315 ne
rect 4716 1260 4771 1315
tri 4771 1260 4946 1435 sw
tri 5009 1315 5129 1435 ne
rect 5129 1315 5165 1435
rect 5285 1315 5321 1435
rect 4716 1178 4946 1260
tri 4946 1178 5028 1260 sw
tri 5129 1178 5266 1315 ne
rect 5266 1260 5321 1315
tri 5321 1260 5496 1435 sw
tri 5559 1315 5679 1435 ne
rect 5679 1315 5715 1435
rect 5835 1315 5871 1435
rect 5266 1178 5496 1260
tri 5496 1178 5578 1260 sw
tri 5679 1178 5816 1315 ne
rect 5816 1260 5871 1315
tri 5871 1260 6046 1435 sw
tri 6109 1315 6229 1435 ne
rect 6229 1315 6265 1435
rect 6385 1315 6421 1435
rect 5816 1178 6046 1260
tri 6046 1178 6128 1260 sw
tri 6229 1178 6366 1315 ne
rect 6366 1260 6421 1315
tri 6421 1260 6596 1435 sw
tri 6659 1315 6779 1435 ne
rect 6779 1315 6815 1435
rect 6935 1315 6971 1435
rect 6366 1178 6596 1260
tri 6596 1178 6678 1260 sw
tri 6779 1178 6916 1315 ne
rect 6916 1260 6971 1315
tri 6971 1260 7146 1435 sw
tri 7209 1315 7329 1435 ne
rect 7329 1315 7365 1435
rect 7485 1315 7521 1435
rect 6916 1178 7146 1260
tri 7146 1178 7228 1260 sw
tri 7329 1178 7466 1315 ne
rect 7466 1260 7521 1315
tri 7521 1260 7696 1435 sw
tri 7759 1315 7879 1435 ne
rect 7879 1315 7915 1435
rect 8035 1315 8071 1435
rect 7466 1178 7696 1260
tri 7696 1178 7778 1260 sw
tri 7879 1178 8016 1315 ne
rect 8016 1260 8071 1315
tri 8071 1260 8246 1435 sw
tri 8309 1315 8429 1435 ne
rect 8429 1315 8465 1435
rect 8585 1315 8621 1435
rect 8016 1178 8246 1260
tri 8246 1178 8328 1260 sw
tri 8429 1178 8566 1315 ne
rect 8566 1260 8621 1315
tri 8621 1260 8796 1435 sw
tri 8859 1315 8979 1435 ne
rect 8979 1315 9015 1435
rect 9135 1315 9171 1435
rect 8566 1178 8796 1260
tri 8796 1178 8878 1260 sw
tri 8979 1178 9116 1315 ne
rect 9116 1260 9171 1315
tri 9171 1260 9346 1435 sw
tri 9409 1315 9529 1435 ne
rect 9529 1315 9565 1435
rect 9685 1315 9721 1435
rect 9116 1178 9346 1260
tri 9346 1178 9428 1260 sw
tri 9529 1178 9666 1315 ne
rect 9666 1260 9721 1315
tri 9721 1260 9896 1435 sw
tri 9959 1315 10079 1435 ne
rect 10079 1315 10115 1435
rect 10235 1315 10271 1435
rect 9666 1178 9896 1260
tri 9896 1178 9978 1260 sw
tri 10079 1178 10216 1315 ne
rect 10216 1260 10271 1315
tri 10271 1260 10446 1435 sw
tri 10509 1315 10629 1435 ne
rect 10629 1315 10665 1435
rect 10785 1315 10821 1435
rect 10216 1178 10446 1260
tri 10446 1178 10528 1260 sw
tri 10629 1178 10766 1315 ne
rect 10766 1260 10821 1315
tri 10821 1260 10996 1435 sw
tri 11059 1315 11179 1435 ne
rect 11179 1315 11215 1435
rect 11335 1315 11371 1435
rect 10766 1178 10996 1260
tri 10996 1178 11078 1260 sw
tri 11179 1178 11316 1315 ne
rect 11316 1260 11371 1315
tri 11371 1260 11546 1435 sw
tri 11609 1315 11729 1435 ne
rect 11729 1315 11765 1435
rect 11885 1315 11921 1435
rect 11316 1178 11546 1260
tri 11546 1178 11628 1260 sw
tri 11729 1178 11866 1315 ne
rect 11866 1260 11921 1315
tri 11921 1260 12096 1435 sw
tri 12159 1315 12279 1435 ne
rect 12279 1315 12315 1435
rect 12435 1315 12471 1435
rect 11866 1178 12096 1260
tri 12096 1178 12178 1260 sw
tri 12279 1178 12416 1315 ne
rect 12416 1260 12471 1315
tri 12471 1260 12646 1435 sw
tri 12709 1315 12829 1435 ne
rect 12829 1315 12865 1435
rect 12985 1315 13021 1435
rect 12416 1178 12646 1260
tri 12646 1178 12728 1260 sw
tri 12829 1178 12966 1315 ne
rect 12966 1260 13021 1315
tri 13021 1260 13196 1435 sw
tri 13259 1315 13379 1435 ne
rect 13379 1315 13415 1435
rect 13535 1315 13571 1435
rect 12966 1178 13196 1260
tri 13196 1178 13278 1260 sw
tri 13379 1178 13516 1315 ne
rect 13516 1260 13571 1315
tri 13571 1260 13746 1435 sw
tri 13809 1315 13929 1435 ne
rect 13929 1315 13965 1435
rect 14085 1315 14121 1435
rect 13516 1178 13746 1260
tri 13746 1178 13828 1260 sw
tri 13929 1178 14066 1315 ne
rect 14066 1260 14121 1315
tri 14121 1260 14296 1435 sw
tri 14359 1315 14479 1435 ne
rect 14479 1315 14515 1435
rect 14635 1315 14671 1435
rect 14066 1178 14296 1260
tri 14296 1178 14378 1260 sw
tri 14479 1178 14616 1315 ne
rect 14616 1260 14671 1315
tri 14671 1260 14846 1435 sw
tri 14909 1315 15029 1435 ne
rect 15029 1315 15065 1435
rect 15185 1315 15221 1435
rect 14616 1178 14846 1260
tri 14846 1178 14928 1260 sw
tri 15029 1178 15166 1315 ne
rect 15166 1260 15221 1315
tri 15221 1260 15396 1435 sw
tri 15459 1315 15579 1435 ne
rect 15579 1315 15615 1435
rect 15735 1315 15771 1435
rect 15166 1178 15396 1260
tri 15396 1178 15478 1260 sw
tri 15579 1178 15716 1315 ne
rect 15716 1260 15771 1315
tri 15771 1260 15946 1435 sw
tri 16009 1315 16129 1435 ne
rect 16129 1315 16165 1435
rect 16285 1315 16321 1435
rect 15716 1178 15946 1260
tri 15946 1178 16028 1260 sw
tri 16129 1178 16266 1315 ne
rect 16266 1260 16321 1315
tri 16321 1260 16496 1435 sw
tri 16559 1315 16679 1435 ne
rect 16679 1315 16715 1435
rect 16835 1315 16871 1435
rect 16266 1178 16496 1260
tri 16496 1178 16578 1260 sw
tri 16679 1178 16816 1315 ne
rect 16816 1260 16871 1315
tri 16871 1260 17046 1435 sw
tri 17109 1315 17229 1435 ne
rect 17229 1315 17265 1435
rect 17385 1315 17421 1435
rect 16816 1178 17046 1260
tri 17046 1178 17128 1260 sw
tri 17229 1178 17366 1315 ne
rect 17366 1260 17421 1315
tri 17421 1260 17596 1435 sw
tri 17659 1315 17779 1435 ne
rect 17779 1315 17815 1435
rect 17935 1315 17971 1435
rect 17366 1178 17596 1260
tri 17596 1178 17678 1260 sw
tri 17779 1178 17916 1315 ne
rect 17916 1260 17971 1315
tri 17971 1260 18146 1435 sw
tri 18209 1315 18329 1435 ne
rect 18329 1315 18365 1435
rect 18485 1315 18521 1435
rect 17916 1178 18146 1260
tri 18146 1178 18228 1260 sw
tri 18329 1178 18466 1315 ne
rect 18466 1260 18521 1315
tri 18521 1260 18696 1435 sw
tri 18759 1315 18879 1435 ne
rect 18879 1315 18915 1435
rect 19035 1315 19071 1435
rect 18466 1178 18696 1260
tri 18696 1178 18778 1260 sw
tri 18879 1178 19016 1315 ne
rect 19016 1260 19071 1315
tri 19071 1260 19246 1435 sw
tri 19309 1315 19429 1435 ne
rect 19429 1315 19465 1435
rect 19585 1333 19621 1435
tri 19621 1333 19723 1435 sw
rect 19585 1315 20300 1333
rect 19016 1178 19246 1260
tri 19246 1178 19328 1260 sw
tri 19429 1178 19566 1315 ne
rect 19566 1178 20300 1315
rect -1000 1022 78 1178
tri 78 1022 234 1178 sw
tri 316 1022 472 1178 ne
rect 472 1022 628 1178
tri 628 1022 784 1178 sw
tri 866 1022 1022 1178 ne
rect 1022 1022 1178 1178
tri 1178 1022 1334 1178 sw
tri 1416 1022 1572 1178 ne
rect 1572 1022 1728 1178
tri 1728 1022 1884 1178 sw
tri 1966 1022 2122 1178 ne
rect 2122 1022 2278 1178
tri 2278 1022 2434 1178 sw
tri 2516 1022 2672 1178 ne
rect 2672 1022 2828 1178
tri 2828 1022 2984 1178 sw
tri 3066 1022 3222 1178 ne
rect 3222 1022 3378 1178
tri 3378 1022 3534 1178 sw
tri 3616 1022 3772 1178 ne
rect 3772 1022 3928 1178
tri 3928 1022 4084 1178 sw
tri 4166 1022 4322 1178 ne
rect 4322 1022 4478 1178
tri 4478 1022 4634 1178 sw
tri 4716 1022 4872 1178 ne
rect 4872 1022 5028 1178
tri 5028 1022 5184 1178 sw
tri 5266 1022 5422 1178 ne
rect 5422 1022 5578 1178
tri 5578 1022 5734 1178 sw
tri 5816 1022 5972 1178 ne
rect 5972 1022 6128 1178
tri 6128 1022 6284 1178 sw
tri 6366 1022 6522 1178 ne
rect 6522 1022 6678 1178
tri 6678 1022 6834 1178 sw
tri 6916 1022 7072 1178 ne
rect 7072 1022 7228 1178
tri 7228 1022 7384 1178 sw
tri 7466 1022 7622 1178 ne
rect 7622 1022 7778 1178
tri 7778 1022 7934 1178 sw
tri 8016 1022 8172 1178 ne
rect 8172 1022 8328 1178
tri 8328 1022 8484 1178 sw
tri 8566 1022 8722 1178 ne
rect 8722 1022 8878 1178
tri 8878 1022 9034 1178 sw
tri 9116 1022 9272 1178 ne
rect 9272 1022 9428 1178
tri 9428 1022 9584 1178 sw
tri 9666 1022 9822 1178 ne
rect 9822 1022 9978 1178
tri 9978 1022 10134 1178 sw
tri 10216 1022 10372 1178 ne
rect 10372 1022 10528 1178
tri 10528 1022 10684 1178 sw
tri 10766 1022 10922 1178 ne
rect 10922 1022 11078 1178
tri 11078 1022 11234 1178 sw
tri 11316 1022 11472 1178 ne
rect 11472 1022 11628 1178
tri 11628 1022 11784 1178 sw
tri 11866 1022 12022 1178 ne
rect 12022 1022 12178 1178
tri 12178 1022 12334 1178 sw
tri 12416 1022 12572 1178 ne
rect 12572 1022 12728 1178
tri 12728 1022 12884 1178 sw
tri 12966 1022 13122 1178 ne
rect 13122 1022 13278 1178
tri 13278 1022 13434 1178 sw
tri 13516 1022 13672 1178 ne
rect 13672 1022 13828 1178
tri 13828 1022 13984 1178 sw
tri 14066 1022 14222 1178 ne
rect 14222 1022 14378 1178
tri 14378 1022 14534 1178 sw
tri 14616 1022 14772 1178 ne
rect 14772 1022 14928 1178
tri 14928 1022 15084 1178 sw
tri 15166 1022 15322 1178 ne
rect 15322 1022 15478 1178
tri 15478 1022 15634 1178 sw
tri 15716 1022 15872 1178 ne
rect 15872 1022 16028 1178
tri 16028 1022 16184 1178 sw
tri 16266 1022 16422 1178 ne
rect 16422 1022 16578 1178
tri 16578 1022 16734 1178 sw
tri 16816 1022 16972 1178 ne
rect 16972 1022 17128 1178
tri 17128 1022 17284 1178 sw
tri 17366 1022 17522 1178 ne
rect 17522 1022 17678 1178
tri 17678 1022 17834 1178 sw
tri 17916 1022 18072 1178 ne
rect 18072 1022 18228 1178
tri 18228 1022 18384 1178 sw
tri 18466 1022 18622 1178 ne
rect 18622 1022 18778 1178
tri 18778 1022 18934 1178 sw
tri 19016 1022 19172 1178 ne
rect 19172 1022 19328 1178
tri 19328 1022 19484 1178 sw
tri 19566 1022 19722 1178 ne
rect 19722 1022 20300 1178
rect -1000 885 234 1022
tri 234 885 371 1022 sw
tri 472 885 609 1022 ne
rect 609 885 784 1022
tri 784 885 921 1022 sw
tri 1022 885 1159 1022 ne
rect 1159 885 1334 1022
tri 1334 885 1471 1022 sw
tri 1572 885 1709 1022 ne
rect 1709 885 1884 1022
tri 1884 885 2021 1022 sw
tri 2122 885 2259 1022 ne
rect 2259 885 2434 1022
tri 2434 885 2571 1022 sw
tri 2672 885 2809 1022 ne
rect 2809 885 2984 1022
tri 2984 885 3121 1022 sw
tri 3222 885 3359 1022 ne
rect 3359 885 3534 1022
tri 3534 885 3671 1022 sw
tri 3772 885 3909 1022 ne
rect 3909 885 4084 1022
tri 4084 885 4221 1022 sw
tri 4322 885 4459 1022 ne
rect 4459 885 4634 1022
tri 4634 885 4771 1022 sw
tri 4872 885 5009 1022 ne
rect 5009 885 5184 1022
tri 5184 885 5321 1022 sw
tri 5422 885 5559 1022 ne
rect 5559 885 5734 1022
tri 5734 885 5871 1022 sw
tri 5972 885 6109 1022 ne
rect 6109 885 6284 1022
tri 6284 885 6421 1022 sw
tri 6522 885 6659 1022 ne
rect 6659 885 6834 1022
tri 6834 885 6971 1022 sw
tri 7072 885 7209 1022 ne
rect 7209 885 7384 1022
tri 7384 885 7521 1022 sw
tri 7622 885 7759 1022 ne
rect 7759 885 7934 1022
tri 7934 885 8071 1022 sw
tri 8172 885 8309 1022 ne
rect 8309 885 8484 1022
tri 8484 885 8621 1022 sw
tri 8722 885 8859 1022 ne
rect 8859 885 9034 1022
tri 9034 885 9171 1022 sw
tri 9272 885 9409 1022 ne
rect 9409 885 9584 1022
tri 9584 885 9721 1022 sw
tri 9822 885 9959 1022 ne
rect 9959 885 10134 1022
tri 10134 885 10271 1022 sw
tri 10372 885 10509 1022 ne
rect 10509 885 10684 1022
tri 10684 885 10821 1022 sw
tri 10922 885 11059 1022 ne
rect 11059 885 11234 1022
tri 11234 885 11371 1022 sw
tri 11472 885 11609 1022 ne
rect 11609 885 11784 1022
tri 11784 885 11921 1022 sw
tri 12022 885 12159 1022 ne
rect 12159 885 12334 1022
tri 12334 885 12471 1022 sw
tri 12572 885 12709 1022 ne
rect 12709 885 12884 1022
tri 12884 885 13021 1022 sw
tri 13122 885 13259 1022 ne
rect 13259 885 13434 1022
tri 13434 885 13571 1022 sw
tri 13672 885 13809 1022 ne
rect 13809 885 13984 1022
tri 13984 885 14121 1022 sw
tri 14222 885 14359 1022 ne
rect 14359 885 14534 1022
tri 14534 885 14671 1022 sw
tri 14772 885 14909 1022 ne
rect 14909 885 15084 1022
tri 15084 885 15221 1022 sw
tri 15322 885 15459 1022 ne
rect 15459 885 15634 1022
tri 15634 885 15771 1022 sw
tri 15872 885 16009 1022 ne
rect 16009 885 16184 1022
tri 16184 885 16321 1022 sw
tri 16422 885 16559 1022 ne
rect 16559 885 16734 1022
tri 16734 885 16871 1022 sw
tri 16972 885 17109 1022 ne
rect 17109 885 17284 1022
tri 17284 885 17421 1022 sw
tri 17522 885 17659 1022 ne
rect 17659 885 17834 1022
tri 17834 885 17971 1022 sw
tri 18072 885 18209 1022 ne
rect 18209 885 18384 1022
tri 18384 885 18521 1022 sw
tri 18622 885 18759 1022 ne
rect 18759 885 18934 1022
tri 18934 885 19071 1022 sw
tri 19172 885 19309 1022 ne
rect 19309 885 19484 1022
tri 19484 885 19621 1022 sw
rect -1000 867 215 885
tri 77 765 179 867 ne
rect 179 765 215 867
rect 335 765 371 885
tri 179 628 316 765 ne
rect 316 710 371 765
tri 371 710 546 885 sw
tri 609 765 729 885 ne
rect 729 765 765 885
rect 885 765 921 885
rect 316 628 546 710
tri 546 628 628 710 sw
tri 729 628 866 765 ne
rect 866 710 921 765
tri 921 710 1096 885 sw
tri 1159 765 1279 885 ne
rect 1279 765 1315 885
rect 1435 765 1471 885
rect 866 628 1096 710
tri 1096 628 1178 710 sw
tri 1279 628 1416 765 ne
rect 1416 710 1471 765
tri 1471 710 1646 885 sw
tri 1709 765 1829 885 ne
rect 1829 765 1865 885
rect 1985 765 2021 885
rect 1416 628 1646 710
tri 1646 628 1728 710 sw
tri 1829 628 1966 765 ne
rect 1966 710 2021 765
tri 2021 710 2196 885 sw
tri 2259 765 2379 885 ne
rect 2379 765 2415 885
rect 2535 765 2571 885
rect 1966 628 2196 710
tri 2196 628 2278 710 sw
tri 2379 628 2516 765 ne
rect 2516 710 2571 765
tri 2571 710 2746 885 sw
tri 2809 765 2929 885 ne
rect 2929 765 2965 885
rect 3085 765 3121 885
rect 2516 628 2746 710
tri 2746 628 2828 710 sw
tri 2929 628 3066 765 ne
rect 3066 710 3121 765
tri 3121 710 3296 885 sw
tri 3359 765 3479 885 ne
rect 3479 765 3515 885
rect 3635 765 3671 885
rect 3066 628 3296 710
tri 3296 628 3378 710 sw
tri 3479 628 3616 765 ne
rect 3616 710 3671 765
tri 3671 710 3846 885 sw
tri 3909 765 4029 885 ne
rect 4029 765 4065 885
rect 4185 765 4221 885
rect 3616 628 3846 710
tri 3846 628 3928 710 sw
tri 4029 628 4166 765 ne
rect 4166 710 4221 765
tri 4221 710 4396 885 sw
tri 4459 765 4579 885 ne
rect 4579 765 4615 885
rect 4735 765 4771 885
rect 4166 628 4396 710
tri 4396 628 4478 710 sw
tri 4579 628 4716 765 ne
rect 4716 710 4771 765
tri 4771 710 4946 885 sw
tri 5009 765 5129 885 ne
rect 5129 765 5165 885
rect 5285 765 5321 885
rect 4716 628 4946 710
tri 4946 628 5028 710 sw
tri 5129 628 5266 765 ne
rect 5266 710 5321 765
tri 5321 710 5496 885 sw
tri 5559 765 5679 885 ne
rect 5679 765 5715 885
rect 5835 765 5871 885
rect 5266 628 5496 710
tri 5496 628 5578 710 sw
tri 5679 628 5816 765 ne
rect 5816 710 5871 765
tri 5871 710 6046 885 sw
tri 6109 765 6229 885 ne
rect 6229 765 6265 885
rect 6385 765 6421 885
rect 5816 628 6046 710
tri 6046 628 6128 710 sw
tri 6229 628 6366 765 ne
rect 6366 710 6421 765
tri 6421 710 6596 885 sw
tri 6659 765 6779 885 ne
rect 6779 765 6815 885
rect 6935 765 6971 885
rect 6366 628 6596 710
tri 6596 628 6678 710 sw
tri 6779 628 6916 765 ne
rect 6916 710 6971 765
tri 6971 710 7146 885 sw
tri 7209 765 7329 885 ne
rect 7329 765 7365 885
rect 7485 765 7521 885
rect 6916 628 7146 710
tri 7146 628 7228 710 sw
tri 7329 628 7466 765 ne
rect 7466 710 7521 765
tri 7521 710 7696 885 sw
tri 7759 765 7879 885 ne
rect 7879 765 7915 885
rect 8035 765 8071 885
rect 7466 628 7696 710
tri 7696 628 7778 710 sw
tri 7879 628 8016 765 ne
rect 8016 710 8071 765
tri 8071 710 8246 885 sw
tri 8309 765 8429 885 ne
rect 8429 765 8465 885
rect 8585 765 8621 885
rect 8016 628 8246 710
tri 8246 628 8328 710 sw
tri 8429 628 8566 765 ne
rect 8566 710 8621 765
tri 8621 710 8796 885 sw
tri 8859 765 8979 885 ne
rect 8979 765 9015 885
rect 9135 765 9171 885
rect 8566 628 8796 710
tri 8796 628 8878 710 sw
tri 8979 628 9116 765 ne
rect 9116 710 9171 765
tri 9171 710 9346 885 sw
tri 9409 765 9529 885 ne
rect 9529 765 9565 885
rect 9685 765 9721 885
rect 9116 628 9346 710
tri 9346 628 9428 710 sw
tri 9529 628 9666 765 ne
rect 9666 710 9721 765
tri 9721 710 9896 885 sw
tri 9959 765 10079 885 ne
rect 10079 765 10115 885
rect 10235 765 10271 885
rect 9666 628 9896 710
tri 9896 628 9978 710 sw
tri 10079 628 10216 765 ne
rect 10216 710 10271 765
tri 10271 710 10446 885 sw
tri 10509 765 10629 885 ne
rect 10629 765 10665 885
rect 10785 765 10821 885
rect 10216 628 10446 710
tri 10446 628 10528 710 sw
tri 10629 628 10766 765 ne
rect 10766 710 10821 765
tri 10821 710 10996 885 sw
tri 11059 765 11179 885 ne
rect 11179 765 11215 885
rect 11335 765 11371 885
rect 10766 628 10996 710
tri 10996 628 11078 710 sw
tri 11179 628 11316 765 ne
rect 11316 710 11371 765
tri 11371 710 11546 885 sw
tri 11609 765 11729 885 ne
rect 11729 765 11765 885
rect 11885 765 11921 885
rect 11316 628 11546 710
tri 11546 628 11628 710 sw
tri 11729 628 11866 765 ne
rect 11866 710 11921 765
tri 11921 710 12096 885 sw
tri 12159 765 12279 885 ne
rect 12279 765 12315 885
rect 12435 765 12471 885
rect 11866 628 12096 710
tri 12096 628 12178 710 sw
tri 12279 628 12416 765 ne
rect 12416 710 12471 765
tri 12471 710 12646 885 sw
tri 12709 765 12829 885 ne
rect 12829 765 12865 885
rect 12985 765 13021 885
rect 12416 628 12646 710
tri 12646 628 12728 710 sw
tri 12829 628 12966 765 ne
rect 12966 710 13021 765
tri 13021 710 13196 885 sw
tri 13259 765 13379 885 ne
rect 13379 765 13415 885
rect 13535 765 13571 885
rect 12966 628 13196 710
tri 13196 628 13278 710 sw
tri 13379 628 13516 765 ne
rect 13516 710 13571 765
tri 13571 710 13746 885 sw
tri 13809 765 13929 885 ne
rect 13929 765 13965 885
rect 14085 765 14121 885
rect 13516 628 13746 710
tri 13746 628 13828 710 sw
tri 13929 628 14066 765 ne
rect 14066 710 14121 765
tri 14121 710 14296 885 sw
tri 14359 765 14479 885 ne
rect 14479 765 14515 885
rect 14635 765 14671 885
rect 14066 628 14296 710
tri 14296 628 14378 710 sw
tri 14479 628 14616 765 ne
rect 14616 710 14671 765
tri 14671 710 14846 885 sw
tri 14909 765 15029 885 ne
rect 15029 765 15065 885
rect 15185 765 15221 885
rect 14616 628 14846 710
tri 14846 628 14928 710 sw
tri 15029 628 15166 765 ne
rect 15166 710 15221 765
tri 15221 710 15396 885 sw
tri 15459 765 15579 885 ne
rect 15579 765 15615 885
rect 15735 765 15771 885
rect 15166 628 15396 710
tri 15396 628 15478 710 sw
tri 15579 628 15716 765 ne
rect 15716 710 15771 765
tri 15771 710 15946 885 sw
tri 16009 765 16129 885 ne
rect 16129 765 16165 885
rect 16285 765 16321 885
rect 15716 628 15946 710
tri 15946 628 16028 710 sw
tri 16129 628 16266 765 ne
rect 16266 710 16321 765
tri 16321 710 16496 885 sw
tri 16559 765 16679 885 ne
rect 16679 765 16715 885
rect 16835 765 16871 885
rect 16266 628 16496 710
tri 16496 628 16578 710 sw
tri 16679 628 16816 765 ne
rect 16816 710 16871 765
tri 16871 710 17046 885 sw
tri 17109 765 17229 885 ne
rect 17229 765 17265 885
rect 17385 765 17421 885
rect 16816 628 17046 710
tri 17046 628 17128 710 sw
tri 17229 628 17366 765 ne
rect 17366 710 17421 765
tri 17421 710 17596 885 sw
tri 17659 765 17779 885 ne
rect 17779 765 17815 885
rect 17935 765 17971 885
rect 17366 628 17596 710
tri 17596 628 17678 710 sw
tri 17779 628 17916 765 ne
rect 17916 710 17971 765
tri 17971 710 18146 885 sw
tri 18209 765 18329 885 ne
rect 18329 765 18365 885
rect 18485 765 18521 885
rect 17916 628 18146 710
tri 18146 628 18228 710 sw
tri 18329 628 18466 765 ne
rect 18466 710 18521 765
tri 18521 710 18696 885 sw
tri 18759 765 18879 885 ne
rect 18879 765 18915 885
rect 19035 765 19071 885
rect 18466 628 18696 710
tri 18696 628 18778 710 sw
tri 18879 628 19016 765 ne
rect 19016 710 19071 765
tri 19071 710 19246 885 sw
tri 19309 765 19429 885 ne
rect 19429 765 19465 885
rect 19585 783 19621 885
tri 19621 783 19723 885 sw
rect 20800 783 21800 1572
rect 19585 765 21800 783
rect 19016 628 19246 710
tri 19246 628 19328 710 sw
tri 19429 628 19566 765 ne
rect 19566 628 21800 765
rect -500 472 78 628
tri 78 472 234 628 sw
tri 316 472 472 628 ne
rect 472 472 628 628
tri 628 472 784 628 sw
tri 866 472 1022 628 ne
rect 1022 472 1178 628
tri 1178 472 1334 628 sw
tri 1416 472 1572 628 ne
rect 1572 472 1728 628
tri 1728 472 1884 628 sw
tri 1966 472 2122 628 ne
rect 2122 472 2278 628
tri 2278 472 2434 628 sw
tri 2516 472 2672 628 ne
rect 2672 472 2828 628
tri 2828 472 2984 628 sw
tri 3066 472 3222 628 ne
rect 3222 472 3378 628
tri 3378 472 3534 628 sw
tri 3616 472 3772 628 ne
rect 3772 472 3928 628
tri 3928 472 4084 628 sw
tri 4166 472 4322 628 ne
rect 4322 472 4478 628
tri 4478 472 4634 628 sw
tri 4716 472 4872 628 ne
rect 4872 472 5028 628
tri 5028 472 5184 628 sw
tri 5266 472 5422 628 ne
rect 5422 472 5578 628
tri 5578 472 5734 628 sw
tri 5816 472 5972 628 ne
rect 5972 472 6128 628
tri 6128 472 6284 628 sw
tri 6366 472 6522 628 ne
rect 6522 472 6678 628
tri 6678 472 6834 628 sw
tri 6916 472 7072 628 ne
rect 7072 472 7228 628
tri 7228 472 7384 628 sw
tri 7466 472 7622 628 ne
rect 7622 472 7778 628
tri 7778 472 7934 628 sw
tri 8016 472 8172 628 ne
rect 8172 472 8328 628
tri 8328 472 8484 628 sw
tri 8566 472 8722 628 ne
rect 8722 472 8878 628
tri 8878 472 9034 628 sw
tri 9116 472 9272 628 ne
rect 9272 472 9428 628
tri 9428 472 9584 628 sw
tri 9666 472 9822 628 ne
rect 9822 472 9978 628
tri 9978 472 10134 628 sw
tri 10216 472 10372 628 ne
rect 10372 472 10528 628
tri 10528 472 10684 628 sw
tri 10766 472 10922 628 ne
rect 10922 472 11078 628
tri 11078 472 11234 628 sw
tri 11316 472 11472 628 ne
rect 11472 472 11628 628
tri 11628 472 11784 628 sw
tri 11866 472 12022 628 ne
rect 12022 472 12178 628
tri 12178 472 12334 628 sw
tri 12416 472 12572 628 ne
rect 12572 472 12728 628
tri 12728 472 12884 628 sw
tri 12966 472 13122 628 ne
rect 13122 472 13278 628
tri 13278 472 13434 628 sw
tri 13516 472 13672 628 ne
rect 13672 472 13828 628
tri 13828 472 13984 628 sw
tri 14066 472 14222 628 ne
rect 14222 472 14378 628
tri 14378 472 14534 628 sw
tri 14616 472 14772 628 ne
rect 14772 472 14928 628
tri 14928 472 15084 628 sw
tri 15166 472 15322 628 ne
rect 15322 472 15478 628
tri 15478 472 15634 628 sw
tri 15716 472 15872 628 ne
rect 15872 472 16028 628
tri 16028 472 16184 628 sw
tri 16266 472 16422 628 ne
rect 16422 472 16578 628
tri 16578 472 16734 628 sw
tri 16816 472 16972 628 ne
rect 16972 472 17128 628
tri 17128 472 17284 628 sw
tri 17366 472 17522 628 ne
rect 17522 472 17678 628
tri 17678 472 17834 628 sw
tri 17916 472 18072 628 ne
rect 18072 472 18228 628
tri 18228 472 18384 628 sw
tri 18466 472 18622 628 ne
rect 18622 472 18778 628
tri 18778 472 18934 628 sw
tri 19016 472 19172 628 ne
rect 19172 472 19328 628
tri 19328 472 19484 628 sw
tri 19566 472 19722 628 ne
rect 19722 472 21800 628
rect -500 335 234 472
tri 234 335 371 472 sw
rect -500 317 215 335
tri 77 215 179 317 ne
rect 179 215 215 317
rect 335 234 371 335
tri 371 234 472 335 sw
tri 472 234 710 472 ne
rect 710 335 784 472
tri 784 335 921 472 sw
rect 710 234 765 335
rect 335 215 472 234
tri 179 77 317 215 ne
rect 317 78 472 215
tri 472 78 628 234 sw
tri 710 215 729 234 ne
rect 729 215 765 234
rect 885 234 921 335
tri 921 234 1022 335 sw
tri 1022 234 1260 472 ne
rect 1260 335 1334 472
tri 1334 335 1471 472 sw
rect 1260 234 1315 335
rect 885 215 1022 234
rect 317 -1000 628 78
tri 729 77 867 215 ne
rect 867 78 1022 215
tri 1022 78 1178 234 sw
tri 1260 215 1279 234 ne
rect 1279 215 1315 234
rect 1435 234 1471 335
tri 1471 234 1572 335 sw
tri 1572 234 1810 472 ne
rect 1810 335 1884 472
tri 1884 335 2021 472 sw
rect 1810 234 1865 335
rect 1435 215 1572 234
rect 867 -500 1178 78
tri 1279 77 1417 215 ne
rect 1417 78 1572 215
tri 1572 78 1728 234 sw
tri 1810 215 1829 234 ne
rect 1829 215 1865 234
rect 1985 234 2021 335
tri 2021 234 2122 335 sw
tri 2122 234 2360 472 ne
rect 2360 335 2434 472
tri 2434 335 2571 472 sw
rect 2360 234 2415 335
rect 1985 215 2122 234
rect 1417 -1000 1728 78
tri 1829 77 1967 215 ne
rect 1967 78 2122 215
tri 2122 78 2278 234 sw
tri 2360 215 2379 234 ne
rect 2379 215 2415 234
rect 2535 234 2571 335
tri 2571 234 2672 335 sw
tri 2672 234 2910 472 ne
rect 2910 335 2984 472
tri 2984 335 3121 472 sw
rect 2910 234 2965 335
rect 2535 215 2672 234
rect 1967 -500 2278 78
tri 2379 77 2517 215 ne
rect 2517 78 2672 215
tri 2672 78 2828 234 sw
tri 2910 215 2929 234 ne
rect 2929 215 2965 234
rect 3085 234 3121 335
tri 3121 234 3222 335 sw
tri 3222 234 3460 472 ne
rect 3460 335 3534 472
tri 3534 335 3671 472 sw
rect 3460 234 3515 335
rect 3085 215 3222 234
rect 2517 -1000 2828 78
tri 2929 77 3067 215 ne
rect 3067 78 3222 215
tri 3222 78 3378 234 sw
tri 3460 215 3479 234 ne
rect 3479 215 3515 234
rect 3635 234 3671 335
tri 3671 234 3772 335 sw
tri 3772 234 4010 472 ne
rect 4010 335 4084 472
tri 4084 335 4221 472 sw
rect 4010 234 4065 335
rect 3635 215 3772 234
rect 3067 -500 3378 78
tri 3479 77 3617 215 ne
rect 3617 78 3772 215
tri 3772 78 3928 234 sw
tri 4010 215 4029 234 ne
rect 4029 215 4065 234
rect 4185 234 4221 335
tri 4221 234 4322 335 sw
tri 4322 234 4560 472 ne
rect 4560 335 4634 472
tri 4634 335 4771 472 sw
rect 4560 234 4615 335
rect 4185 215 4322 234
rect 3617 -1000 3928 78
tri 4029 77 4167 215 ne
rect 4167 78 4322 215
tri 4322 78 4478 234 sw
tri 4560 215 4579 234 ne
rect 4579 215 4615 234
rect 4735 234 4771 335
tri 4771 234 4872 335 sw
tri 4872 234 5110 472 ne
rect 5110 335 5184 472
tri 5184 335 5321 472 sw
rect 5110 234 5165 335
rect 4735 215 4872 234
rect 4167 -500 4478 78
tri 4579 77 4717 215 ne
rect 4717 78 4872 215
tri 4872 78 5028 234 sw
tri 5110 215 5129 234 ne
rect 5129 215 5165 234
rect 5285 234 5321 335
tri 5321 234 5422 335 sw
tri 5422 234 5660 472 ne
rect 5660 335 5734 472
tri 5734 335 5871 472 sw
rect 5660 234 5715 335
rect 5285 215 5422 234
rect 4717 -1000 5028 78
tri 5129 77 5267 215 ne
rect 5267 78 5422 215
tri 5422 78 5578 234 sw
tri 5660 215 5679 234 ne
rect 5679 215 5715 234
rect 5835 234 5871 335
tri 5871 234 5972 335 sw
tri 5972 234 6210 472 ne
rect 6210 335 6284 472
tri 6284 335 6421 472 sw
rect 6210 234 6265 335
rect 5835 215 5972 234
rect 5267 -500 5578 78
tri 5679 77 5817 215 ne
rect 5817 78 5972 215
tri 5972 78 6128 234 sw
tri 6210 215 6229 234 ne
rect 6229 215 6265 234
rect 6385 234 6421 335
tri 6421 234 6522 335 sw
tri 6522 234 6760 472 ne
rect 6760 335 6834 472
tri 6834 335 6971 472 sw
rect 6760 234 6815 335
rect 6385 215 6522 234
rect 5817 -1000 6128 78
tri 6229 77 6367 215 ne
rect 6367 78 6522 215
tri 6522 78 6678 234 sw
tri 6760 215 6779 234 ne
rect 6779 215 6815 234
rect 6935 234 6971 335
tri 6971 234 7072 335 sw
tri 7072 234 7310 472 ne
rect 7310 335 7384 472
tri 7384 335 7521 472 sw
rect 7310 234 7365 335
rect 6935 215 7072 234
rect 6367 -500 6678 78
tri 6779 77 6917 215 ne
rect 6917 78 7072 215
tri 7072 78 7228 234 sw
tri 7310 215 7329 234 ne
rect 7329 215 7365 234
rect 7485 234 7521 335
tri 7521 234 7622 335 sw
tri 7622 234 7860 472 ne
rect 7860 335 7934 472
tri 7934 335 8071 472 sw
rect 7860 234 7915 335
rect 7485 215 7622 234
rect 6917 -1000 7228 78
tri 7329 77 7467 215 ne
rect 7467 78 7622 215
tri 7622 78 7778 234 sw
tri 7860 215 7879 234 ne
rect 7879 215 7915 234
rect 8035 234 8071 335
tri 8071 234 8172 335 sw
tri 8172 234 8410 472 ne
rect 8410 335 8484 472
tri 8484 335 8621 472 sw
rect 8410 234 8465 335
rect 8035 215 8172 234
rect 7467 -500 7778 78
tri 7879 77 8017 215 ne
rect 8017 78 8172 215
tri 8172 78 8328 234 sw
tri 8410 215 8429 234 ne
rect 8429 215 8465 234
rect 8585 234 8621 335
tri 8621 234 8722 335 sw
tri 8722 234 8960 472 ne
rect 8960 335 9034 472
tri 9034 335 9171 472 sw
rect 8960 234 9015 335
rect 8585 215 8722 234
rect 8017 -1000 8328 78
tri 8429 77 8567 215 ne
rect 8567 78 8722 215
tri 8722 78 8878 234 sw
tri 8960 215 8979 234 ne
rect 8979 215 9015 234
rect 9135 234 9171 335
tri 9171 234 9272 335 sw
tri 9272 234 9510 472 ne
rect 9510 335 9584 472
tri 9584 335 9721 472 sw
rect 9510 234 9565 335
rect 9135 215 9272 234
rect 8567 -500 8878 78
tri 8979 77 9117 215 ne
rect 9117 78 9272 215
tri 9272 78 9428 234 sw
tri 9510 215 9529 234 ne
rect 9529 215 9565 234
rect 9685 234 9721 335
tri 9721 234 9822 335 sw
tri 9822 234 10060 472 ne
rect 10060 335 10134 472
tri 10134 335 10271 472 sw
rect 10060 234 10115 335
rect 9685 215 9822 234
rect 9117 -1000 9428 78
tri 9529 77 9667 215 ne
rect 9667 78 9822 215
tri 9822 78 9978 234 sw
tri 10060 215 10079 234 ne
rect 10079 215 10115 234
rect 10235 234 10271 335
tri 10271 234 10372 335 sw
tri 10372 234 10610 472 ne
rect 10610 335 10684 472
tri 10684 335 10821 472 sw
rect 10610 234 10665 335
rect 10235 215 10372 234
rect 9667 -500 9978 78
tri 10079 77 10217 215 ne
rect 10217 78 10372 215
tri 10372 78 10528 234 sw
tri 10610 215 10629 234 ne
rect 10629 215 10665 234
rect 10785 234 10821 335
tri 10821 234 10922 335 sw
tri 10922 234 11160 472 ne
rect 11160 335 11234 472
tri 11234 335 11371 472 sw
rect 11160 234 11215 335
rect 10785 215 10922 234
rect 10217 -1000 10528 78
tri 10629 77 10767 215 ne
rect 10767 78 10922 215
tri 10922 78 11078 234 sw
tri 11160 215 11179 234 ne
rect 11179 215 11215 234
rect 11335 234 11371 335
tri 11371 234 11472 335 sw
tri 11472 234 11710 472 ne
rect 11710 335 11784 472
tri 11784 335 11921 472 sw
rect 11710 234 11765 335
rect 11335 215 11472 234
rect 10767 -500 11078 78
tri 11179 77 11317 215 ne
rect 11317 78 11472 215
tri 11472 78 11628 234 sw
tri 11710 215 11729 234 ne
rect 11729 215 11765 234
rect 11885 234 11921 335
tri 11921 234 12022 335 sw
tri 12022 234 12260 472 ne
rect 12260 335 12334 472
tri 12334 335 12471 472 sw
rect 12260 234 12315 335
rect 11885 215 12022 234
rect 11317 -1000 11628 78
tri 11729 77 11867 215 ne
rect 11867 78 12022 215
tri 12022 78 12178 234 sw
tri 12260 215 12279 234 ne
rect 12279 215 12315 234
rect 12435 234 12471 335
tri 12471 234 12572 335 sw
tri 12572 234 12810 472 ne
rect 12810 335 12884 472
tri 12884 335 13021 472 sw
rect 12810 234 12865 335
rect 12435 215 12572 234
rect 11867 -500 12178 78
tri 12279 77 12417 215 ne
rect 12417 78 12572 215
tri 12572 78 12728 234 sw
tri 12810 215 12829 234 ne
rect 12829 215 12865 234
rect 12985 234 13021 335
tri 13021 234 13122 335 sw
tri 13122 234 13360 472 ne
rect 13360 335 13434 472
tri 13434 335 13571 472 sw
rect 13360 234 13415 335
rect 12985 215 13122 234
rect 12417 -1000 12728 78
tri 12829 77 12967 215 ne
rect 12967 78 13122 215
tri 13122 78 13278 234 sw
tri 13360 215 13379 234 ne
rect 13379 215 13415 234
rect 13535 234 13571 335
tri 13571 234 13672 335 sw
tri 13672 234 13910 472 ne
rect 13910 335 13984 472
tri 13984 335 14121 472 sw
rect 13910 234 13965 335
rect 13535 215 13672 234
rect 12967 -500 13278 78
tri 13379 77 13517 215 ne
rect 13517 78 13672 215
tri 13672 78 13828 234 sw
tri 13910 215 13929 234 ne
rect 13929 215 13965 234
rect 14085 234 14121 335
tri 14121 234 14222 335 sw
tri 14222 234 14460 472 ne
rect 14460 335 14534 472
tri 14534 335 14671 472 sw
rect 14460 234 14515 335
rect 14085 215 14222 234
rect 13517 -1000 13828 78
tri 13929 77 14067 215 ne
rect 14067 78 14222 215
tri 14222 78 14378 234 sw
tri 14460 215 14479 234 ne
rect 14479 215 14515 234
rect 14635 234 14671 335
tri 14671 234 14772 335 sw
tri 14772 234 15010 472 ne
rect 15010 335 15084 472
tri 15084 335 15221 472 sw
rect 15010 234 15065 335
rect 14635 215 14772 234
rect 14067 -500 14378 78
tri 14479 77 14617 215 ne
rect 14617 78 14772 215
tri 14772 78 14928 234 sw
tri 15010 215 15029 234 ne
rect 15029 215 15065 234
rect 15185 234 15221 335
tri 15221 234 15322 335 sw
tri 15322 234 15560 472 ne
rect 15560 335 15634 472
tri 15634 335 15771 472 sw
rect 15560 234 15615 335
rect 15185 215 15322 234
rect 14617 -1000 14928 78
tri 15029 77 15167 215 ne
rect 15167 78 15322 215
tri 15322 78 15478 234 sw
tri 15560 215 15579 234 ne
rect 15579 215 15615 234
rect 15735 234 15771 335
tri 15771 234 15872 335 sw
tri 15872 234 16110 472 ne
rect 16110 335 16184 472
tri 16184 335 16321 472 sw
rect 16110 234 16165 335
rect 15735 215 15872 234
rect 15167 -500 15478 78
tri 15579 77 15717 215 ne
rect 15717 78 15872 215
tri 15872 78 16028 234 sw
tri 16110 215 16129 234 ne
rect 16129 215 16165 234
rect 16285 234 16321 335
tri 16321 234 16422 335 sw
tri 16422 234 16660 472 ne
rect 16660 335 16734 472
tri 16734 335 16871 472 sw
rect 16660 234 16715 335
rect 16285 215 16422 234
rect 15717 -1000 16028 78
tri 16129 77 16267 215 ne
rect 16267 78 16422 215
tri 16422 78 16578 234 sw
tri 16660 215 16679 234 ne
rect 16679 215 16715 234
rect 16835 234 16871 335
tri 16871 234 16972 335 sw
tri 16972 234 17210 472 ne
rect 17210 335 17284 472
tri 17284 335 17421 472 sw
rect 17210 234 17265 335
rect 16835 215 16972 234
rect 16267 -500 16578 78
tri 16679 77 16817 215 ne
rect 16817 78 16972 215
tri 16972 78 17128 234 sw
tri 17210 215 17229 234 ne
rect 17229 215 17265 234
rect 17385 234 17421 335
tri 17421 234 17522 335 sw
tri 17522 234 17760 472 ne
rect 17760 335 17834 472
tri 17834 335 17971 472 sw
rect 17760 234 17815 335
rect 17385 215 17522 234
rect 16817 -1000 17128 78
tri 17229 77 17367 215 ne
rect 17367 78 17522 215
tri 17522 78 17678 234 sw
tri 17760 215 17779 234 ne
rect 17779 215 17815 234
rect 17935 234 17971 335
tri 17971 234 18072 335 sw
tri 18072 234 18310 472 ne
rect 18310 335 18384 472
tri 18384 335 18521 472 sw
rect 18310 234 18365 335
rect 17935 215 18072 234
rect 17367 -500 17678 78
tri 17779 77 17917 215 ne
rect 17917 78 18072 215
tri 18072 78 18228 234 sw
tri 18310 215 18329 234 ne
rect 18329 215 18365 234
rect 18485 234 18521 335
tri 18521 234 18622 335 sw
tri 18622 234 18860 472 ne
rect 18860 335 18934 472
tri 18934 335 19071 472 sw
rect 18860 234 18915 335
rect 18485 215 18622 234
rect 17917 -1000 18228 78
tri 18329 77 18467 215 ne
rect 18467 78 18622 215
tri 18622 78 18778 234 sw
tri 18860 215 18879 234 ne
rect 18879 215 18915 234
rect 19035 234 19071 335
tri 19071 234 19172 335 sw
tri 19172 234 19410 472 ne
rect 19410 335 19484 472
tri 19484 335 19621 472 sw
rect 19410 234 19465 335
rect 19035 215 19172 234
rect 18467 -500 18778 78
tri 18879 77 19017 215 ne
rect 19017 78 19172 215
tri 19172 78 19328 234 sw
tri 19410 215 19429 234 ne
rect 19429 215 19465 234
rect 19585 233 19621 335
tri 19621 233 19723 335 sw
rect 19585 215 20300 233
rect 19017 -1000 19328 78
tri 19429 77 19567 215 ne
rect 19567 -78 20300 215
rect 19567 -500 19878 -78
rect 20800 -1000 21800 472
rect 0 -2000 21800 -1000
<< properties >>
string MASKHINTS_HVNTM 43 39417 39557 39557 43 43 39557 183 43 183 183 39417 39417 183 39557 39417
<< end >>
