magic
tech sky130A
timestamp 1666382007
<< metal1 >>
rect 1000 41045 136600 41050
rect 1000 40855 4897 41045
rect 4930 40855 56597 41045
rect 56630 40855 65597 41045
rect 65630 40855 130597 41045
rect 130630 40855 136600 41045
rect 1000 40850 136600 40855
rect 1000 40795 136900 40800
rect 1000 40605 5335 40795
rect 5425 40605 57035 40795
rect 57125 40605 66035 40795
rect 66125 40605 131035 40795
rect 131125 40605 136900 40795
rect 1000 40600 136900 40605
rect 1000 37995 1500 40600
rect 2000 40350 137200 40550
rect 1000 37505 1005 37995
rect 1495 37505 1500 37995
rect 1000 37500 1500 37505
rect 135500 37995 136000 40350
rect 135500 37505 135505 37995
rect 135995 37505 136000 37995
rect 135500 37500 136000 37505
<< via1 >>
rect 4897 40855 4930 41045
rect 56597 40855 56630 41045
rect 65597 40855 65630 41045
rect 130597 40855 130630 41045
rect 5335 40605 5425 40795
rect 57035 40605 57125 40795
rect 66035 40605 66125 40795
rect 131035 40605 131125 40795
rect 4897 39906 4930 40136
rect 5335 39806 5425 40096
rect 56597 39906 56630 40136
rect 57035 39806 57125 40096
rect 65597 39906 65630 40136
rect 66035 39806 66125 40096
rect 130597 39906 130630 40136
rect 131035 39806 131125 40096
rect 1005 37505 1495 37995
rect 135505 37505 135995 37995
<< metal2 >>
rect 5050 41550 136600 41650
rect 4892 41045 4935 41050
rect 4892 40855 4897 41045
rect 4930 40855 4935 41045
rect 4892 40136 4935 40855
rect 5050 40266 5150 41550
rect 56750 41400 136800 41500
rect 56592 41045 56635 41050
rect 56592 40855 56597 41045
rect 56630 40855 56635 41045
rect 5330 40795 5430 40800
rect 5330 40605 5335 40795
rect 5425 40605 5430 40795
rect 4892 39906 4897 40136
rect 4930 39906 4935 40136
rect 4892 39901 4935 39906
rect 5330 40096 5430 40605
rect 5330 39806 5335 40096
rect 5425 39806 5430 40096
rect 56592 40136 56635 40855
rect 56750 40266 56850 41400
rect 65750 41250 137000 41350
rect 65592 41045 65635 41050
rect 65592 40855 65597 41045
rect 65630 40855 65635 41045
rect 57030 40795 57130 40800
rect 57030 40605 57035 40795
rect 57125 40605 57130 40795
rect 56592 39906 56597 40136
rect 56630 39906 56635 40136
rect 56592 39901 56635 39906
rect 57030 40096 57130 40605
rect 5330 39801 5430 39806
rect 57030 39806 57035 40096
rect 57125 39806 57130 40096
rect 65592 40136 65635 40855
rect 65750 40266 65850 41250
rect 130750 41100 137200 41200
rect 130592 41045 130635 41050
rect 130592 40855 130597 41045
rect 130630 40855 130635 41045
rect 66030 40795 66130 40800
rect 66030 40605 66035 40795
rect 66125 40605 66130 40795
rect 65592 39906 65597 40136
rect 65630 39906 65635 40136
rect 65592 39901 65635 39906
rect 66030 40096 66130 40605
rect 57030 39801 57130 39806
rect 66030 39806 66035 40096
rect 66125 39806 66130 40096
rect 130592 40136 130635 40855
rect 130750 40266 130850 41100
rect 131030 40795 131130 40800
rect 131030 40605 131035 40795
rect 131125 40605 131130 40795
rect 130592 39906 130597 40136
rect 130630 39906 130635 40136
rect 130592 39901 130635 39906
rect 131030 40096 131130 40605
rect 66030 39801 66130 39806
rect 131030 39806 131035 40096
rect 131125 39806 131130 40096
rect 131030 39801 131130 39806
rect 1000 37995 1500 38000
rect 1000 37505 1005 37995
rect 1495 37505 1500 37995
rect 135500 37995 136000 38000
rect 1000 37500 1500 37505
rect 5409 34000 5519 37666
rect 57109 34000 57219 37666
rect 66109 34000 66219 37666
rect 131109 34000 131219 37666
rect 135500 37505 135505 37995
rect 135995 37505 136000 37995
rect 135500 37500 136000 37505
<< via2 >>
rect 1005 37505 1495 37995
rect 135505 37505 135995 37995
<< metal3 >>
rect 1000 37995 1500 38000
rect 1000 37505 1005 37995
rect 1495 37505 1500 37995
rect 1000 31000 1500 37505
rect 135500 37995 136000 38000
rect 135500 37505 135505 37995
rect 135995 37505 136000 37995
rect 135500 31000 136000 37505
use converter  converter_0
timestamp 1666362992
transform 1 0 0 0 1 0
box 0 0 137200 208000
use level_shifter  level_shifter_0
timestamp 1665425771
transform 0 1 129000 -1 0 39203
box -1223 0 1802 4468
use level_shifter  level_shifter_1
timestamp 1665425771
transform 0 1 64000 -1 0 39203
box -1223 0 1802 4468
use level_shifter  level_shifter_2
timestamp 1665425771
transform 0 1 55000 -1 0 39203
box -1223 0 1802 4468
use level_shifter  level_shifter_3
timestamp 1665425771
transform 0 1 3300 -1 0 39203
box -1223 0 1802 4468
<< labels >>
rlabel metal1 136400 40850 136600 41050 7 VDD
rlabel metal2 137100 41100 137200 41200 7 D1
rlabel metal2 136900 41250 137000 41350 7 D2
rlabel metal2 136700 41400 136800 41500 7 D3
rlabel metal2 136500 41550 136600 41650 7 D1
<< end >>
