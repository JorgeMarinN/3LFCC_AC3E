magic
tech sky130A
timestamp 1668091195
<< metal1 >>
rect -40 9920 29960 9960
rect -40 0 0 9920
rect 29920 0 29960 9920
rect -40 -40 29960 0
<< metal2 >>
rect -40 9920 29960 9960
rect -40 0 0 9920
rect 29920 0 29960 9920
rect -40 -40 29960 0
<< metal3 >>
rect -40 9920 29960 9960
rect -40 0 0 9920
rect 29920 0 29960 9920
rect -40 -40 29960 0
<< metal4 >>
rect -40 9920 29960 9960
rect -40 0 0 9920
rect 29920 0 29960 9920
rect -40 -40 29960 0
<< metal5 >>
rect -40 0 0 9960
rect -40 -40 29960 0
use unit_pad  unit_pad_0
timestamp 1668089732
transform 1 0 0 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_1
timestamp 1668089732
transform 1 0 0 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_2
timestamp 1668089732
transform 1 0 0 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_3
timestamp 1668089732
transform 1 0 0 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_4
timestamp 1668089732
transform 1 0 0 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_5
timestamp 1668089732
transform 1 0 0 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_6
timestamp 1668089732
transform 1 0 0 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_7
timestamp 1668089732
transform 1 0 0 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_8
timestamp 1668089732
transform 1 0 0 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_9
timestamp 1668089732
transform 1 0 0 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_10
timestamp 1668089732
transform 1 0 0 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_11
timestamp 1668089732
transform 1 0 0 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_12
timestamp 1668089732
transform 1 0 0 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_13
timestamp 1668089732
transform 1 0 0 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_14
timestamp 1668089732
transform 1 0 0 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_15
timestamp 1668089732
transform 1 0 0 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_16
timestamp 1668089732
transform 1 0 0 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_17
timestamp 1668089732
transform 1 0 0 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_18
timestamp 1668089732
transform 1 0 0 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_19
timestamp 1668089732
transform 1 0 0 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_20
timestamp 1668089732
transform 1 0 0 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_21
timestamp 1668089732
transform 1 0 0 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_22
timestamp 1668089732
transform 1 0 0 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_23
timestamp 1668089732
transform 1 0 0 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_24
timestamp 1668089732
transform 1 0 0 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_25
timestamp 1668089732
transform 1 0 0 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_26
timestamp 1668089732
transform 1 0 0 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_27
timestamp 1668089732
transform 1 0 0 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_28
timestamp 1668089732
transform 1 0 0 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_29
timestamp 1668089732
transform 1 0 0 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_30
timestamp 1668089732
transform 1 0 0 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_31
timestamp 1668089732
transform 1 0 0 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_32
timestamp 1668089732
transform 1 0 0 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_33
timestamp 1668089732
transform 1 0 0 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_34
timestamp 1668089732
transform 1 0 0 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_35
timestamp 1668089732
transform 1 0 0 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_36
timestamp 1668089732
transform 1 0 0 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_37
timestamp 1668089732
transform 1 0 0 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_38
timestamp 1668089732
transform 1 0 0 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_39
timestamp 1668089732
transform 1 0 0 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_40
timestamp 1668089732
transform 1 0 0 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_41
timestamp 1668089732
transform 1 0 0 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_42
timestamp 1668089732
transform 1 0 0 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_43
timestamp 1668089732
transform 1 0 0 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_44
timestamp 1668089732
transform 1 0 0 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_45
timestamp 1668089732
transform 1 0 0 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_46
timestamp 1668089732
transform 1 0 0 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_47
timestamp 1668089732
transform 1 0 0 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_48
timestamp 1668089732
transform 1 0 0 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_49
timestamp 1668089732
transform 1 0 0 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_50
timestamp 1668089732
transform 1 0 0 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_51
timestamp 1668089732
transform 1 0 0 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_52
timestamp 1668089732
transform 1 0 0 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_53
timestamp 1668089732
transform 1 0 0 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_54
timestamp 1668089732
transform 1 0 0 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_55
timestamp 1668089732
transform 1 0 0 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_56
timestamp 1668089732
transform 1 0 0 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_57
timestamp 1668089732
transform 1 0 0 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_58
timestamp 1668089732
transform 1 0 0 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_59
timestamp 1668089732
transform 1 0 0 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_60
timestamp 1668089732
transform 1 0 0 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_61
timestamp 1668089732
transform 1 0 0 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_62
timestamp 1668089732
transform 1 0 160 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_63
timestamp 1668089732
transform 1 0 160 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_64
timestamp 1668089732
transform 1 0 160 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_65
timestamp 1668089732
transform 1 0 160 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_66
timestamp 1668089732
transform 1 0 160 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_67
timestamp 1668089732
transform 1 0 160 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_68
timestamp 1668089732
transform 1 0 160 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_69
timestamp 1668089732
transform 1 0 160 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_70
timestamp 1668089732
transform 1 0 160 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_71
timestamp 1668089732
transform 1 0 160 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_72
timestamp 1668089732
transform 1 0 160 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_73
timestamp 1668089732
transform 1 0 160 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_74
timestamp 1668089732
transform 1 0 160 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_75
timestamp 1668089732
transform 1 0 160 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_76
timestamp 1668089732
transform 1 0 160 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_77
timestamp 1668089732
transform 1 0 160 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_78
timestamp 1668089732
transform 1 0 160 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_79
timestamp 1668089732
transform 1 0 160 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_80
timestamp 1668089732
transform 1 0 160 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_81
timestamp 1668089732
transform 1 0 160 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_82
timestamp 1668089732
transform 1 0 160 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_83
timestamp 1668089732
transform 1 0 160 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_84
timestamp 1668089732
transform 1 0 160 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_85
timestamp 1668089732
transform 1 0 160 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_86
timestamp 1668089732
transform 1 0 160 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_87
timestamp 1668089732
transform 1 0 160 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_88
timestamp 1668089732
transform 1 0 160 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_89
timestamp 1668089732
transform 1 0 160 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_90
timestamp 1668089732
transform 1 0 160 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_91
timestamp 1668089732
transform 1 0 160 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_92
timestamp 1668089732
transform 1 0 160 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_93
timestamp 1668089732
transform 1 0 160 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_94
timestamp 1668089732
transform 1 0 160 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_95
timestamp 1668089732
transform 1 0 160 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_96
timestamp 1668089732
transform 1 0 160 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_97
timestamp 1668089732
transform 1 0 160 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_98
timestamp 1668089732
transform 1 0 160 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_99
timestamp 1668089732
transform 1 0 160 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_100
timestamp 1668089732
transform 1 0 160 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_101
timestamp 1668089732
transform 1 0 160 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_102
timestamp 1668089732
transform 1 0 160 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_103
timestamp 1668089732
transform 1 0 160 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_104
timestamp 1668089732
transform 1 0 160 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_105
timestamp 1668089732
transform 1 0 160 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_106
timestamp 1668089732
transform 1 0 160 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_107
timestamp 1668089732
transform 1 0 160 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_108
timestamp 1668089732
transform 1 0 160 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_109
timestamp 1668089732
transform 1 0 160 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_110
timestamp 1668089732
transform 1 0 160 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_111
timestamp 1668089732
transform 1 0 160 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_112
timestamp 1668089732
transform 1 0 160 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_113
timestamp 1668089732
transform 1 0 160 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_114
timestamp 1668089732
transform 1 0 160 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_115
timestamp 1668089732
transform 1 0 160 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_116
timestamp 1668089732
transform 1 0 160 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_117
timestamp 1668089732
transform 1 0 160 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_118
timestamp 1668089732
transform 1 0 160 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_119
timestamp 1668089732
transform 1 0 160 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_120
timestamp 1668089732
transform 1 0 160 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_121
timestamp 1668089732
transform 1 0 160 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_122
timestamp 1668089732
transform 1 0 160 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_123
timestamp 1668089732
transform 1 0 160 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_124
timestamp 1668089732
transform 1 0 320 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_125
timestamp 1668089732
transform 1 0 320 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_126
timestamp 1668089732
transform 1 0 320 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_127
timestamp 1668089732
transform 1 0 320 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_128
timestamp 1668089732
transform 1 0 320 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_129
timestamp 1668089732
transform 1 0 320 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_130
timestamp 1668089732
transform 1 0 320 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_131
timestamp 1668089732
transform 1 0 320 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_132
timestamp 1668089732
transform 1 0 320 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_133
timestamp 1668089732
transform 1 0 320 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_134
timestamp 1668089732
transform 1 0 320 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_135
timestamp 1668089732
transform 1 0 320 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_136
timestamp 1668089732
transform 1 0 320 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_137
timestamp 1668089732
transform 1 0 320 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_138
timestamp 1668089732
transform 1 0 320 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_139
timestamp 1668089732
transform 1 0 320 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_140
timestamp 1668089732
transform 1 0 320 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_141
timestamp 1668089732
transform 1 0 320 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_142
timestamp 1668089732
transform 1 0 320 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_143
timestamp 1668089732
transform 1 0 320 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_144
timestamp 1668089732
transform 1 0 320 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_145
timestamp 1668089732
transform 1 0 320 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_146
timestamp 1668089732
transform 1 0 320 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_147
timestamp 1668089732
transform 1 0 320 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_148
timestamp 1668089732
transform 1 0 320 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_149
timestamp 1668089732
transform 1 0 320 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_150
timestamp 1668089732
transform 1 0 320 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_151
timestamp 1668089732
transform 1 0 320 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_152
timestamp 1668089732
transform 1 0 320 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_153
timestamp 1668089732
transform 1 0 320 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_154
timestamp 1668089732
transform 1 0 320 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_155
timestamp 1668089732
transform 1 0 320 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_156
timestamp 1668089732
transform 1 0 320 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_157
timestamp 1668089732
transform 1 0 320 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_158
timestamp 1668089732
transform 1 0 320 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_159
timestamp 1668089732
transform 1 0 320 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_160
timestamp 1668089732
transform 1 0 320 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_161
timestamp 1668089732
transform 1 0 320 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_162
timestamp 1668089732
transform 1 0 320 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_163
timestamp 1668089732
transform 1 0 320 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_164
timestamp 1668089732
transform 1 0 320 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_165
timestamp 1668089732
transform 1 0 320 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_166
timestamp 1668089732
transform 1 0 320 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_167
timestamp 1668089732
transform 1 0 320 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_168
timestamp 1668089732
transform 1 0 320 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_169
timestamp 1668089732
transform 1 0 320 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_170
timestamp 1668089732
transform 1 0 320 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_171
timestamp 1668089732
transform 1 0 320 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_172
timestamp 1668089732
transform 1 0 320 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_173
timestamp 1668089732
transform 1 0 320 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_174
timestamp 1668089732
transform 1 0 320 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_175
timestamp 1668089732
transform 1 0 320 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_176
timestamp 1668089732
transform 1 0 320 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_177
timestamp 1668089732
transform 1 0 320 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_178
timestamp 1668089732
transform 1 0 320 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_179
timestamp 1668089732
transform 1 0 320 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_180
timestamp 1668089732
transform 1 0 320 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_181
timestamp 1668089732
transform 1 0 320 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_182
timestamp 1668089732
transform 1 0 320 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_183
timestamp 1668089732
transform 1 0 320 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_184
timestamp 1668089732
transform 1 0 320 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_185
timestamp 1668089732
transform 1 0 320 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_186
timestamp 1668089732
transform 1 0 480 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_187
timestamp 1668089732
transform 1 0 480 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_188
timestamp 1668089732
transform 1 0 480 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_189
timestamp 1668089732
transform 1 0 480 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_190
timestamp 1668089732
transform 1 0 480 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_191
timestamp 1668089732
transform 1 0 480 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_192
timestamp 1668089732
transform 1 0 480 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_193
timestamp 1668089732
transform 1 0 480 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_194
timestamp 1668089732
transform 1 0 480 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_195
timestamp 1668089732
transform 1 0 480 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_196
timestamp 1668089732
transform 1 0 480 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_197
timestamp 1668089732
transform 1 0 480 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_198
timestamp 1668089732
transform 1 0 480 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_199
timestamp 1668089732
transform 1 0 480 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_200
timestamp 1668089732
transform 1 0 480 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_201
timestamp 1668089732
transform 1 0 480 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_202
timestamp 1668089732
transform 1 0 480 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_203
timestamp 1668089732
transform 1 0 480 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_204
timestamp 1668089732
transform 1 0 480 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_205
timestamp 1668089732
transform 1 0 480 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_206
timestamp 1668089732
transform 1 0 480 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_207
timestamp 1668089732
transform 1 0 480 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_208
timestamp 1668089732
transform 1 0 480 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_209
timestamp 1668089732
transform 1 0 480 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_210
timestamp 1668089732
transform 1 0 480 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_211
timestamp 1668089732
transform 1 0 480 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_212
timestamp 1668089732
transform 1 0 480 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_213
timestamp 1668089732
transform 1 0 480 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_214
timestamp 1668089732
transform 1 0 480 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_215
timestamp 1668089732
transform 1 0 480 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_216
timestamp 1668089732
transform 1 0 480 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_217
timestamp 1668089732
transform 1 0 480 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_218
timestamp 1668089732
transform 1 0 480 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_219
timestamp 1668089732
transform 1 0 480 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_220
timestamp 1668089732
transform 1 0 480 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_221
timestamp 1668089732
transform 1 0 480 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_222
timestamp 1668089732
transform 1 0 480 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_223
timestamp 1668089732
transform 1 0 480 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_224
timestamp 1668089732
transform 1 0 480 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_225
timestamp 1668089732
transform 1 0 480 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_226
timestamp 1668089732
transform 1 0 480 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_227
timestamp 1668089732
transform 1 0 480 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_228
timestamp 1668089732
transform 1 0 480 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_229
timestamp 1668089732
transform 1 0 480 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_230
timestamp 1668089732
transform 1 0 480 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_231
timestamp 1668089732
transform 1 0 480 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_232
timestamp 1668089732
transform 1 0 480 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_233
timestamp 1668089732
transform 1 0 480 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_234
timestamp 1668089732
transform 1 0 480 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_235
timestamp 1668089732
transform 1 0 480 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_236
timestamp 1668089732
transform 1 0 480 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_237
timestamp 1668089732
transform 1 0 480 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_238
timestamp 1668089732
transform 1 0 480 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_239
timestamp 1668089732
transform 1 0 480 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_240
timestamp 1668089732
transform 1 0 480 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_241
timestamp 1668089732
transform 1 0 480 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_242
timestamp 1668089732
transform 1 0 480 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_243
timestamp 1668089732
transform 1 0 480 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_244
timestamp 1668089732
transform 1 0 480 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_245
timestamp 1668089732
transform 1 0 480 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_246
timestamp 1668089732
transform 1 0 480 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_247
timestamp 1668089732
transform 1 0 480 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_248
timestamp 1668089732
transform 1 0 640 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_249
timestamp 1668089732
transform 1 0 640 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_250
timestamp 1668089732
transform 1 0 640 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_251
timestamp 1668089732
transform 1 0 640 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_252
timestamp 1668089732
transform 1 0 640 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_253
timestamp 1668089732
transform 1 0 640 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_254
timestamp 1668089732
transform 1 0 640 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_255
timestamp 1668089732
transform 1 0 640 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_256
timestamp 1668089732
transform 1 0 640 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_257
timestamp 1668089732
transform 1 0 640 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_258
timestamp 1668089732
transform 1 0 640 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_259
timestamp 1668089732
transform 1 0 640 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_260
timestamp 1668089732
transform 1 0 640 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_261
timestamp 1668089732
transform 1 0 640 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_262
timestamp 1668089732
transform 1 0 640 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_263
timestamp 1668089732
transform 1 0 640 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_264
timestamp 1668089732
transform 1 0 640 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_265
timestamp 1668089732
transform 1 0 640 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_266
timestamp 1668089732
transform 1 0 640 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_267
timestamp 1668089732
transform 1 0 640 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_268
timestamp 1668089732
transform 1 0 640 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_269
timestamp 1668089732
transform 1 0 640 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_270
timestamp 1668089732
transform 1 0 640 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_271
timestamp 1668089732
transform 1 0 640 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_272
timestamp 1668089732
transform 1 0 640 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_273
timestamp 1668089732
transform 1 0 640 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_274
timestamp 1668089732
transform 1 0 640 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_275
timestamp 1668089732
transform 1 0 640 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_276
timestamp 1668089732
transform 1 0 640 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_277
timestamp 1668089732
transform 1 0 640 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_278
timestamp 1668089732
transform 1 0 640 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_279
timestamp 1668089732
transform 1 0 640 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_280
timestamp 1668089732
transform 1 0 640 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_281
timestamp 1668089732
transform 1 0 640 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_282
timestamp 1668089732
transform 1 0 640 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_283
timestamp 1668089732
transform 1 0 640 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_284
timestamp 1668089732
transform 1 0 640 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_285
timestamp 1668089732
transform 1 0 640 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_286
timestamp 1668089732
transform 1 0 640 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_287
timestamp 1668089732
transform 1 0 640 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_288
timestamp 1668089732
transform 1 0 640 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_289
timestamp 1668089732
transform 1 0 640 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_290
timestamp 1668089732
transform 1 0 640 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_291
timestamp 1668089732
transform 1 0 640 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_292
timestamp 1668089732
transform 1 0 640 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_293
timestamp 1668089732
transform 1 0 640 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_294
timestamp 1668089732
transform 1 0 640 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_295
timestamp 1668089732
transform 1 0 640 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_296
timestamp 1668089732
transform 1 0 640 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_297
timestamp 1668089732
transform 1 0 640 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_298
timestamp 1668089732
transform 1 0 640 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_299
timestamp 1668089732
transform 1 0 640 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_300
timestamp 1668089732
transform 1 0 640 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_301
timestamp 1668089732
transform 1 0 640 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_302
timestamp 1668089732
transform 1 0 640 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_303
timestamp 1668089732
transform 1 0 640 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_304
timestamp 1668089732
transform 1 0 640 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_305
timestamp 1668089732
transform 1 0 640 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_306
timestamp 1668089732
transform 1 0 640 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_307
timestamp 1668089732
transform 1 0 640 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_308
timestamp 1668089732
transform 1 0 640 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_309
timestamp 1668089732
transform 1 0 640 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_310
timestamp 1668089732
transform 1 0 800 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_311
timestamp 1668089732
transform 1 0 800 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_312
timestamp 1668089732
transform 1 0 800 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_313
timestamp 1668089732
transform 1 0 800 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_314
timestamp 1668089732
transform 1 0 800 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_315
timestamp 1668089732
transform 1 0 800 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_316
timestamp 1668089732
transform 1 0 800 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_317
timestamp 1668089732
transform 1 0 800 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_318
timestamp 1668089732
transform 1 0 800 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_319
timestamp 1668089732
transform 1 0 800 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_320
timestamp 1668089732
transform 1 0 800 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_321
timestamp 1668089732
transform 1 0 800 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_322
timestamp 1668089732
transform 1 0 800 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_323
timestamp 1668089732
transform 1 0 800 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_324
timestamp 1668089732
transform 1 0 800 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_325
timestamp 1668089732
transform 1 0 800 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_326
timestamp 1668089732
transform 1 0 800 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_327
timestamp 1668089732
transform 1 0 800 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_328
timestamp 1668089732
transform 1 0 800 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_329
timestamp 1668089732
transform 1 0 800 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_330
timestamp 1668089732
transform 1 0 800 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_331
timestamp 1668089732
transform 1 0 800 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_332
timestamp 1668089732
transform 1 0 800 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_333
timestamp 1668089732
transform 1 0 800 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_334
timestamp 1668089732
transform 1 0 800 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_335
timestamp 1668089732
transform 1 0 800 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_336
timestamp 1668089732
transform 1 0 800 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_337
timestamp 1668089732
transform 1 0 800 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_338
timestamp 1668089732
transform 1 0 800 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_339
timestamp 1668089732
transform 1 0 800 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_340
timestamp 1668089732
transform 1 0 800 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_341
timestamp 1668089732
transform 1 0 800 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_342
timestamp 1668089732
transform 1 0 800 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_343
timestamp 1668089732
transform 1 0 800 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_344
timestamp 1668089732
transform 1 0 800 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_345
timestamp 1668089732
transform 1 0 800 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_346
timestamp 1668089732
transform 1 0 800 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_347
timestamp 1668089732
transform 1 0 800 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_348
timestamp 1668089732
transform 1 0 800 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_349
timestamp 1668089732
transform 1 0 800 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_350
timestamp 1668089732
transform 1 0 800 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_351
timestamp 1668089732
transform 1 0 800 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_352
timestamp 1668089732
transform 1 0 800 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_353
timestamp 1668089732
transform 1 0 800 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_354
timestamp 1668089732
transform 1 0 800 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_355
timestamp 1668089732
transform 1 0 800 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_356
timestamp 1668089732
transform 1 0 800 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_357
timestamp 1668089732
transform 1 0 800 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_358
timestamp 1668089732
transform 1 0 800 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_359
timestamp 1668089732
transform 1 0 800 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_360
timestamp 1668089732
transform 1 0 800 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_361
timestamp 1668089732
transform 1 0 800 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_362
timestamp 1668089732
transform 1 0 800 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_363
timestamp 1668089732
transform 1 0 800 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_364
timestamp 1668089732
transform 1 0 800 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_365
timestamp 1668089732
transform 1 0 800 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_366
timestamp 1668089732
transform 1 0 800 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_367
timestamp 1668089732
transform 1 0 800 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_368
timestamp 1668089732
transform 1 0 800 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_369
timestamp 1668089732
transform 1 0 800 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_370
timestamp 1668089732
transform 1 0 800 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_371
timestamp 1668089732
transform 1 0 800 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_372
timestamp 1668089732
transform 1 0 960 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_373
timestamp 1668089732
transform 1 0 960 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_374
timestamp 1668089732
transform 1 0 960 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_375
timestamp 1668089732
transform 1 0 960 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_376
timestamp 1668089732
transform 1 0 960 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_377
timestamp 1668089732
transform 1 0 960 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_378
timestamp 1668089732
transform 1 0 960 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_379
timestamp 1668089732
transform 1 0 960 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_380
timestamp 1668089732
transform 1 0 960 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_381
timestamp 1668089732
transform 1 0 960 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_382
timestamp 1668089732
transform 1 0 960 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_383
timestamp 1668089732
transform 1 0 960 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_384
timestamp 1668089732
transform 1 0 960 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_385
timestamp 1668089732
transform 1 0 960 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_386
timestamp 1668089732
transform 1 0 960 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_387
timestamp 1668089732
transform 1 0 960 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_388
timestamp 1668089732
transform 1 0 960 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_389
timestamp 1668089732
transform 1 0 960 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_390
timestamp 1668089732
transform 1 0 960 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_391
timestamp 1668089732
transform 1 0 960 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_392
timestamp 1668089732
transform 1 0 960 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_393
timestamp 1668089732
transform 1 0 960 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_394
timestamp 1668089732
transform 1 0 960 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_395
timestamp 1668089732
transform 1 0 960 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_396
timestamp 1668089732
transform 1 0 960 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_397
timestamp 1668089732
transform 1 0 960 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_398
timestamp 1668089732
transform 1 0 960 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_399
timestamp 1668089732
transform 1 0 960 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_400
timestamp 1668089732
transform 1 0 960 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_401
timestamp 1668089732
transform 1 0 960 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_402
timestamp 1668089732
transform 1 0 960 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_403
timestamp 1668089732
transform 1 0 960 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_404
timestamp 1668089732
transform 1 0 960 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_405
timestamp 1668089732
transform 1 0 960 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_406
timestamp 1668089732
transform 1 0 960 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_407
timestamp 1668089732
transform 1 0 960 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_408
timestamp 1668089732
transform 1 0 960 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_409
timestamp 1668089732
transform 1 0 960 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_410
timestamp 1668089732
transform 1 0 960 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_411
timestamp 1668089732
transform 1 0 960 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_412
timestamp 1668089732
transform 1 0 960 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_413
timestamp 1668089732
transform 1 0 960 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_414
timestamp 1668089732
transform 1 0 960 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_415
timestamp 1668089732
transform 1 0 960 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_416
timestamp 1668089732
transform 1 0 960 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_417
timestamp 1668089732
transform 1 0 960 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_418
timestamp 1668089732
transform 1 0 960 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_419
timestamp 1668089732
transform 1 0 960 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_420
timestamp 1668089732
transform 1 0 960 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_421
timestamp 1668089732
transform 1 0 960 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_422
timestamp 1668089732
transform 1 0 960 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_423
timestamp 1668089732
transform 1 0 960 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_424
timestamp 1668089732
transform 1 0 960 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_425
timestamp 1668089732
transform 1 0 960 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_426
timestamp 1668089732
transform 1 0 960 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_427
timestamp 1668089732
transform 1 0 960 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_428
timestamp 1668089732
transform 1 0 960 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_429
timestamp 1668089732
transform 1 0 960 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_430
timestamp 1668089732
transform 1 0 960 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_431
timestamp 1668089732
transform 1 0 960 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_432
timestamp 1668089732
transform 1 0 960 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_433
timestamp 1668089732
transform 1 0 960 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_434
timestamp 1668089732
transform 1 0 1120 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_435
timestamp 1668089732
transform 1 0 1120 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_436
timestamp 1668089732
transform 1 0 1120 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_437
timestamp 1668089732
transform 1 0 1120 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_438
timestamp 1668089732
transform 1 0 1120 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_439
timestamp 1668089732
transform 1 0 1120 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_440
timestamp 1668089732
transform 1 0 1120 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_441
timestamp 1668089732
transform 1 0 1120 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_442
timestamp 1668089732
transform 1 0 1120 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_443
timestamp 1668089732
transform 1 0 1120 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_444
timestamp 1668089732
transform 1 0 1120 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_445
timestamp 1668089732
transform 1 0 1120 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_446
timestamp 1668089732
transform 1 0 1120 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_447
timestamp 1668089732
transform 1 0 1120 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_448
timestamp 1668089732
transform 1 0 1120 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_449
timestamp 1668089732
transform 1 0 1120 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_450
timestamp 1668089732
transform 1 0 1120 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_451
timestamp 1668089732
transform 1 0 1120 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_452
timestamp 1668089732
transform 1 0 1120 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_453
timestamp 1668089732
transform 1 0 1120 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_454
timestamp 1668089732
transform 1 0 1120 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_455
timestamp 1668089732
transform 1 0 1120 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_456
timestamp 1668089732
transform 1 0 1120 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_457
timestamp 1668089732
transform 1 0 1120 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_458
timestamp 1668089732
transform 1 0 1120 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_459
timestamp 1668089732
transform 1 0 1120 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_460
timestamp 1668089732
transform 1 0 1120 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_461
timestamp 1668089732
transform 1 0 1120 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_462
timestamp 1668089732
transform 1 0 1120 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_463
timestamp 1668089732
transform 1 0 1120 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_464
timestamp 1668089732
transform 1 0 1120 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_465
timestamp 1668089732
transform 1 0 1120 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_466
timestamp 1668089732
transform 1 0 1120 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_467
timestamp 1668089732
transform 1 0 1120 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_468
timestamp 1668089732
transform 1 0 1120 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_469
timestamp 1668089732
transform 1 0 1120 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_470
timestamp 1668089732
transform 1 0 1120 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_471
timestamp 1668089732
transform 1 0 1120 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_472
timestamp 1668089732
transform 1 0 1120 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_473
timestamp 1668089732
transform 1 0 1120 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_474
timestamp 1668089732
transform 1 0 1120 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_475
timestamp 1668089732
transform 1 0 1120 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_476
timestamp 1668089732
transform 1 0 1120 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_477
timestamp 1668089732
transform 1 0 1120 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_478
timestamp 1668089732
transform 1 0 1120 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_479
timestamp 1668089732
transform 1 0 1120 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_480
timestamp 1668089732
transform 1 0 1120 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_481
timestamp 1668089732
transform 1 0 1120 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_482
timestamp 1668089732
transform 1 0 1120 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_483
timestamp 1668089732
transform 1 0 1120 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_484
timestamp 1668089732
transform 1 0 1120 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_485
timestamp 1668089732
transform 1 0 1120 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_486
timestamp 1668089732
transform 1 0 1120 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_487
timestamp 1668089732
transform 1 0 1120 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_488
timestamp 1668089732
transform 1 0 1120 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_489
timestamp 1668089732
transform 1 0 1120 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_490
timestamp 1668089732
transform 1 0 1120 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_491
timestamp 1668089732
transform 1 0 1120 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_492
timestamp 1668089732
transform 1 0 1120 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_493
timestamp 1668089732
transform 1 0 1120 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_494
timestamp 1668089732
transform 1 0 1120 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_495
timestamp 1668089732
transform 1 0 1120 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_496
timestamp 1668089732
transform 1 0 1280 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_497
timestamp 1668089732
transform 1 0 1280 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_498
timestamp 1668089732
transform 1 0 1280 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_499
timestamp 1668089732
transform 1 0 1280 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_500
timestamp 1668089732
transform 1 0 1280 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_501
timestamp 1668089732
transform 1 0 1280 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_502
timestamp 1668089732
transform 1 0 1280 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_503
timestamp 1668089732
transform 1 0 1280 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_504
timestamp 1668089732
transform 1 0 1280 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_505
timestamp 1668089732
transform 1 0 1280 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_506
timestamp 1668089732
transform 1 0 1280 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_507
timestamp 1668089732
transform 1 0 1280 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_508
timestamp 1668089732
transform 1 0 1280 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_509
timestamp 1668089732
transform 1 0 1280 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_510
timestamp 1668089732
transform 1 0 1280 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_511
timestamp 1668089732
transform 1 0 1280 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_512
timestamp 1668089732
transform 1 0 1280 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_513
timestamp 1668089732
transform 1 0 1280 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_514
timestamp 1668089732
transform 1 0 1280 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_515
timestamp 1668089732
transform 1 0 1280 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_516
timestamp 1668089732
transform 1 0 1280 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_517
timestamp 1668089732
transform 1 0 1280 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_518
timestamp 1668089732
transform 1 0 1280 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_519
timestamp 1668089732
transform 1 0 1280 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_520
timestamp 1668089732
transform 1 0 1280 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_521
timestamp 1668089732
transform 1 0 1280 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_522
timestamp 1668089732
transform 1 0 1280 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_523
timestamp 1668089732
transform 1 0 1280 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_524
timestamp 1668089732
transform 1 0 1280 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_525
timestamp 1668089732
transform 1 0 1280 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_526
timestamp 1668089732
transform 1 0 1280 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_527
timestamp 1668089732
transform 1 0 1280 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_528
timestamp 1668089732
transform 1 0 1280 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_529
timestamp 1668089732
transform 1 0 1280 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_530
timestamp 1668089732
transform 1 0 1280 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_531
timestamp 1668089732
transform 1 0 1280 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_532
timestamp 1668089732
transform 1 0 1280 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_533
timestamp 1668089732
transform 1 0 1280 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_534
timestamp 1668089732
transform 1 0 1280 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_535
timestamp 1668089732
transform 1 0 1280 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_536
timestamp 1668089732
transform 1 0 1280 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_537
timestamp 1668089732
transform 1 0 1280 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_538
timestamp 1668089732
transform 1 0 1280 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_539
timestamp 1668089732
transform 1 0 1280 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_540
timestamp 1668089732
transform 1 0 1280 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_541
timestamp 1668089732
transform 1 0 1280 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_542
timestamp 1668089732
transform 1 0 1280 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_543
timestamp 1668089732
transform 1 0 1280 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_544
timestamp 1668089732
transform 1 0 1280 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_545
timestamp 1668089732
transform 1 0 1280 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_546
timestamp 1668089732
transform 1 0 1280 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_547
timestamp 1668089732
transform 1 0 1280 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_548
timestamp 1668089732
transform 1 0 1280 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_549
timestamp 1668089732
transform 1 0 1280 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_550
timestamp 1668089732
transform 1 0 1280 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_551
timestamp 1668089732
transform 1 0 1280 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_552
timestamp 1668089732
transform 1 0 1280 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_553
timestamp 1668089732
transform 1 0 1280 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_554
timestamp 1668089732
transform 1 0 1280 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_555
timestamp 1668089732
transform 1 0 1280 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_556
timestamp 1668089732
transform 1 0 1280 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_557
timestamp 1668089732
transform 1 0 1280 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_558
timestamp 1668089732
transform 1 0 1440 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_559
timestamp 1668089732
transform 1 0 1440 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_560
timestamp 1668089732
transform 1 0 1440 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_561
timestamp 1668089732
transform 1 0 1440 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_562
timestamp 1668089732
transform 1 0 1440 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_563
timestamp 1668089732
transform 1 0 1440 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_564
timestamp 1668089732
transform 1 0 1440 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_565
timestamp 1668089732
transform 1 0 1440 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_566
timestamp 1668089732
transform 1 0 1440 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_567
timestamp 1668089732
transform 1 0 1440 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_568
timestamp 1668089732
transform 1 0 1440 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_569
timestamp 1668089732
transform 1 0 1440 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_570
timestamp 1668089732
transform 1 0 1440 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_571
timestamp 1668089732
transform 1 0 1440 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_572
timestamp 1668089732
transform 1 0 1440 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_573
timestamp 1668089732
transform 1 0 1440 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_574
timestamp 1668089732
transform 1 0 1440 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_575
timestamp 1668089732
transform 1 0 1440 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_576
timestamp 1668089732
transform 1 0 1440 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_577
timestamp 1668089732
transform 1 0 1440 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_578
timestamp 1668089732
transform 1 0 1440 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_579
timestamp 1668089732
transform 1 0 1440 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_580
timestamp 1668089732
transform 1 0 1440 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_581
timestamp 1668089732
transform 1 0 1440 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_582
timestamp 1668089732
transform 1 0 1440 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_583
timestamp 1668089732
transform 1 0 1440 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_584
timestamp 1668089732
transform 1 0 1440 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_585
timestamp 1668089732
transform 1 0 1440 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_586
timestamp 1668089732
transform 1 0 1440 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_587
timestamp 1668089732
transform 1 0 1440 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_588
timestamp 1668089732
transform 1 0 1440 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_589
timestamp 1668089732
transform 1 0 1440 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_590
timestamp 1668089732
transform 1 0 1440 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_591
timestamp 1668089732
transform 1 0 1440 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_592
timestamp 1668089732
transform 1 0 1440 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_593
timestamp 1668089732
transform 1 0 1440 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_594
timestamp 1668089732
transform 1 0 1440 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_595
timestamp 1668089732
transform 1 0 1440 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_596
timestamp 1668089732
transform 1 0 1440 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_597
timestamp 1668089732
transform 1 0 1440 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_598
timestamp 1668089732
transform 1 0 1440 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_599
timestamp 1668089732
transform 1 0 1440 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_600
timestamp 1668089732
transform 1 0 1440 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_601
timestamp 1668089732
transform 1 0 1440 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_602
timestamp 1668089732
transform 1 0 1440 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_603
timestamp 1668089732
transform 1 0 1440 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_604
timestamp 1668089732
transform 1 0 1440 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_605
timestamp 1668089732
transform 1 0 1440 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_606
timestamp 1668089732
transform 1 0 1440 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_607
timestamp 1668089732
transform 1 0 1440 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_608
timestamp 1668089732
transform 1 0 1440 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_609
timestamp 1668089732
transform 1 0 1440 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_610
timestamp 1668089732
transform 1 0 1440 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_611
timestamp 1668089732
transform 1 0 1440 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_612
timestamp 1668089732
transform 1 0 1440 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_613
timestamp 1668089732
transform 1 0 1440 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_614
timestamp 1668089732
transform 1 0 1440 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_615
timestamp 1668089732
transform 1 0 1440 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_616
timestamp 1668089732
transform 1 0 1440 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_617
timestamp 1668089732
transform 1 0 1440 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_618
timestamp 1668089732
transform 1 0 1440 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_619
timestamp 1668089732
transform 1 0 1440 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_620
timestamp 1668089732
transform 1 0 1600 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_621
timestamp 1668089732
transform 1 0 1600 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_622
timestamp 1668089732
transform 1 0 1600 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_623
timestamp 1668089732
transform 1 0 1600 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_624
timestamp 1668089732
transform 1 0 1600 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_625
timestamp 1668089732
transform 1 0 1600 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_626
timestamp 1668089732
transform 1 0 1600 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_627
timestamp 1668089732
transform 1 0 1600 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_628
timestamp 1668089732
transform 1 0 1600 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_629
timestamp 1668089732
transform 1 0 1600 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_630
timestamp 1668089732
transform 1 0 1600 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_631
timestamp 1668089732
transform 1 0 1600 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_632
timestamp 1668089732
transform 1 0 1600 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_633
timestamp 1668089732
transform 1 0 1600 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_634
timestamp 1668089732
transform 1 0 1600 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_635
timestamp 1668089732
transform 1 0 1600 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_636
timestamp 1668089732
transform 1 0 1600 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_637
timestamp 1668089732
transform 1 0 1600 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_638
timestamp 1668089732
transform 1 0 1600 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_639
timestamp 1668089732
transform 1 0 1600 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_640
timestamp 1668089732
transform 1 0 1600 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_641
timestamp 1668089732
transform 1 0 1600 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_642
timestamp 1668089732
transform 1 0 1600 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_643
timestamp 1668089732
transform 1 0 1600 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_644
timestamp 1668089732
transform 1 0 1600 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_645
timestamp 1668089732
transform 1 0 1600 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_646
timestamp 1668089732
transform 1 0 1600 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_647
timestamp 1668089732
transform 1 0 1600 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_648
timestamp 1668089732
transform 1 0 1600 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_649
timestamp 1668089732
transform 1 0 1600 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_650
timestamp 1668089732
transform 1 0 1600 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_651
timestamp 1668089732
transform 1 0 1600 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_652
timestamp 1668089732
transform 1 0 1600 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_653
timestamp 1668089732
transform 1 0 1600 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_654
timestamp 1668089732
transform 1 0 1600 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_655
timestamp 1668089732
transform 1 0 1600 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_656
timestamp 1668089732
transform 1 0 1600 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_657
timestamp 1668089732
transform 1 0 1600 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_658
timestamp 1668089732
transform 1 0 1600 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_659
timestamp 1668089732
transform 1 0 1600 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_660
timestamp 1668089732
transform 1 0 1600 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_661
timestamp 1668089732
transform 1 0 1600 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_662
timestamp 1668089732
transform 1 0 1600 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_663
timestamp 1668089732
transform 1 0 1600 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_664
timestamp 1668089732
transform 1 0 1600 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_665
timestamp 1668089732
transform 1 0 1600 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_666
timestamp 1668089732
transform 1 0 1600 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_667
timestamp 1668089732
transform 1 0 1600 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_668
timestamp 1668089732
transform 1 0 1600 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_669
timestamp 1668089732
transform 1 0 1600 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_670
timestamp 1668089732
transform 1 0 1600 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_671
timestamp 1668089732
transform 1 0 1600 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_672
timestamp 1668089732
transform 1 0 1600 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_673
timestamp 1668089732
transform 1 0 1600 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_674
timestamp 1668089732
transform 1 0 1600 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_675
timestamp 1668089732
transform 1 0 1600 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_676
timestamp 1668089732
transform 1 0 1600 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_677
timestamp 1668089732
transform 1 0 1600 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_678
timestamp 1668089732
transform 1 0 1600 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_679
timestamp 1668089732
transform 1 0 1600 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_680
timestamp 1668089732
transform 1 0 1600 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_681
timestamp 1668089732
transform 1 0 1600 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_682
timestamp 1668089732
transform 1 0 1760 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_683
timestamp 1668089732
transform 1 0 1760 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_684
timestamp 1668089732
transform 1 0 1760 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_685
timestamp 1668089732
transform 1 0 1760 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_686
timestamp 1668089732
transform 1 0 1760 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_687
timestamp 1668089732
transform 1 0 1760 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_688
timestamp 1668089732
transform 1 0 1760 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_689
timestamp 1668089732
transform 1 0 1760 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_690
timestamp 1668089732
transform 1 0 1760 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_691
timestamp 1668089732
transform 1 0 1760 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_692
timestamp 1668089732
transform 1 0 1760 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_693
timestamp 1668089732
transform 1 0 1760 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_694
timestamp 1668089732
transform 1 0 1760 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_695
timestamp 1668089732
transform 1 0 1760 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_696
timestamp 1668089732
transform 1 0 1760 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_697
timestamp 1668089732
transform 1 0 1760 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_698
timestamp 1668089732
transform 1 0 1760 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_699
timestamp 1668089732
transform 1 0 1760 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_700
timestamp 1668089732
transform 1 0 1760 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_701
timestamp 1668089732
transform 1 0 1760 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_702
timestamp 1668089732
transform 1 0 1760 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_703
timestamp 1668089732
transform 1 0 1760 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_704
timestamp 1668089732
transform 1 0 1760 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_705
timestamp 1668089732
transform 1 0 1760 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_706
timestamp 1668089732
transform 1 0 1760 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_707
timestamp 1668089732
transform 1 0 1760 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_708
timestamp 1668089732
transform 1 0 1760 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_709
timestamp 1668089732
transform 1 0 1760 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_710
timestamp 1668089732
transform 1 0 1760 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_711
timestamp 1668089732
transform 1 0 1760 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_712
timestamp 1668089732
transform 1 0 1760 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_713
timestamp 1668089732
transform 1 0 1760 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_714
timestamp 1668089732
transform 1 0 1760 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_715
timestamp 1668089732
transform 1 0 1760 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_716
timestamp 1668089732
transform 1 0 1760 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_717
timestamp 1668089732
transform 1 0 1760 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_718
timestamp 1668089732
transform 1 0 1760 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_719
timestamp 1668089732
transform 1 0 1760 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_720
timestamp 1668089732
transform 1 0 1760 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_721
timestamp 1668089732
transform 1 0 1760 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_722
timestamp 1668089732
transform 1 0 1760 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_723
timestamp 1668089732
transform 1 0 1760 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_724
timestamp 1668089732
transform 1 0 1760 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_725
timestamp 1668089732
transform 1 0 1760 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_726
timestamp 1668089732
transform 1 0 1760 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_727
timestamp 1668089732
transform 1 0 1760 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_728
timestamp 1668089732
transform 1 0 1760 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_729
timestamp 1668089732
transform 1 0 1760 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_730
timestamp 1668089732
transform 1 0 1760 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_731
timestamp 1668089732
transform 1 0 1760 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_732
timestamp 1668089732
transform 1 0 1760 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_733
timestamp 1668089732
transform 1 0 1760 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_734
timestamp 1668089732
transform 1 0 1760 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_735
timestamp 1668089732
transform 1 0 1760 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_736
timestamp 1668089732
transform 1 0 1760 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_737
timestamp 1668089732
transform 1 0 1760 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_738
timestamp 1668089732
transform 1 0 1760 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_739
timestamp 1668089732
transform 1 0 1760 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_740
timestamp 1668089732
transform 1 0 1760 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_741
timestamp 1668089732
transform 1 0 1760 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_742
timestamp 1668089732
transform 1 0 1760 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_743
timestamp 1668089732
transform 1 0 1760 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_744
timestamp 1668089732
transform 1 0 1920 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_745
timestamp 1668089732
transform 1 0 1920 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_746
timestamp 1668089732
transform 1 0 1920 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_747
timestamp 1668089732
transform 1 0 1920 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_748
timestamp 1668089732
transform 1 0 1920 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_749
timestamp 1668089732
transform 1 0 1920 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_750
timestamp 1668089732
transform 1 0 1920 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_751
timestamp 1668089732
transform 1 0 1920 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_752
timestamp 1668089732
transform 1 0 1920 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_753
timestamp 1668089732
transform 1 0 1920 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_754
timestamp 1668089732
transform 1 0 1920 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_755
timestamp 1668089732
transform 1 0 1920 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_756
timestamp 1668089732
transform 1 0 1920 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_757
timestamp 1668089732
transform 1 0 1920 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_758
timestamp 1668089732
transform 1 0 1920 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_759
timestamp 1668089732
transform 1 0 1920 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_760
timestamp 1668089732
transform 1 0 1920 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_761
timestamp 1668089732
transform 1 0 1920 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_762
timestamp 1668089732
transform 1 0 1920 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_763
timestamp 1668089732
transform 1 0 1920 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_764
timestamp 1668089732
transform 1 0 1920 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_765
timestamp 1668089732
transform 1 0 1920 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_766
timestamp 1668089732
transform 1 0 1920 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_767
timestamp 1668089732
transform 1 0 1920 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_768
timestamp 1668089732
transform 1 0 1920 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_769
timestamp 1668089732
transform 1 0 1920 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_770
timestamp 1668089732
transform 1 0 1920 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_771
timestamp 1668089732
transform 1 0 1920 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_772
timestamp 1668089732
transform 1 0 1920 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_773
timestamp 1668089732
transform 1 0 1920 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_774
timestamp 1668089732
transform 1 0 1920 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_775
timestamp 1668089732
transform 1 0 1920 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_776
timestamp 1668089732
transform 1 0 1920 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_777
timestamp 1668089732
transform 1 0 1920 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_778
timestamp 1668089732
transform 1 0 1920 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_779
timestamp 1668089732
transform 1 0 1920 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_780
timestamp 1668089732
transform 1 0 1920 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_781
timestamp 1668089732
transform 1 0 1920 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_782
timestamp 1668089732
transform 1 0 1920 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_783
timestamp 1668089732
transform 1 0 1920 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_784
timestamp 1668089732
transform 1 0 1920 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_785
timestamp 1668089732
transform 1 0 1920 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_786
timestamp 1668089732
transform 1 0 1920 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_787
timestamp 1668089732
transform 1 0 1920 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_788
timestamp 1668089732
transform 1 0 1920 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_789
timestamp 1668089732
transform 1 0 1920 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_790
timestamp 1668089732
transform 1 0 1920 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_791
timestamp 1668089732
transform 1 0 1920 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_792
timestamp 1668089732
transform 1 0 1920 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_793
timestamp 1668089732
transform 1 0 1920 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_794
timestamp 1668089732
transform 1 0 1920 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_795
timestamp 1668089732
transform 1 0 1920 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_796
timestamp 1668089732
transform 1 0 1920 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_797
timestamp 1668089732
transform 1 0 1920 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_798
timestamp 1668089732
transform 1 0 1920 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_799
timestamp 1668089732
transform 1 0 1920 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_800
timestamp 1668089732
transform 1 0 1920 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_801
timestamp 1668089732
transform 1 0 1920 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_802
timestamp 1668089732
transform 1 0 1920 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_803
timestamp 1668089732
transform 1 0 1920 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_804
timestamp 1668089732
transform 1 0 1920 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_805
timestamp 1668089732
transform 1 0 1920 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_806
timestamp 1668089732
transform 1 0 2080 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_807
timestamp 1668089732
transform 1 0 2080 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_808
timestamp 1668089732
transform 1 0 2080 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_809
timestamp 1668089732
transform 1 0 2080 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_810
timestamp 1668089732
transform 1 0 2080 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_811
timestamp 1668089732
transform 1 0 2080 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_812
timestamp 1668089732
transform 1 0 2080 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_813
timestamp 1668089732
transform 1 0 2080 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_814
timestamp 1668089732
transform 1 0 2080 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_815
timestamp 1668089732
transform 1 0 2080 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_816
timestamp 1668089732
transform 1 0 2080 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_817
timestamp 1668089732
transform 1 0 2080 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_818
timestamp 1668089732
transform 1 0 2080 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_819
timestamp 1668089732
transform 1 0 2080 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_820
timestamp 1668089732
transform 1 0 2080 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_821
timestamp 1668089732
transform 1 0 2080 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_822
timestamp 1668089732
transform 1 0 2080 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_823
timestamp 1668089732
transform 1 0 2080 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_824
timestamp 1668089732
transform 1 0 2080 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_825
timestamp 1668089732
transform 1 0 2080 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_826
timestamp 1668089732
transform 1 0 2080 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_827
timestamp 1668089732
transform 1 0 2080 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_828
timestamp 1668089732
transform 1 0 2080 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_829
timestamp 1668089732
transform 1 0 2080 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_830
timestamp 1668089732
transform 1 0 2080 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_831
timestamp 1668089732
transform 1 0 2080 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_832
timestamp 1668089732
transform 1 0 2080 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_833
timestamp 1668089732
transform 1 0 2080 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_834
timestamp 1668089732
transform 1 0 2080 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_835
timestamp 1668089732
transform 1 0 2080 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_836
timestamp 1668089732
transform 1 0 2080 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_837
timestamp 1668089732
transform 1 0 2080 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_838
timestamp 1668089732
transform 1 0 2080 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_839
timestamp 1668089732
transform 1 0 2080 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_840
timestamp 1668089732
transform 1 0 2080 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_841
timestamp 1668089732
transform 1 0 2080 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_842
timestamp 1668089732
transform 1 0 2080 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_843
timestamp 1668089732
transform 1 0 2080 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_844
timestamp 1668089732
transform 1 0 2080 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_845
timestamp 1668089732
transform 1 0 2080 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_846
timestamp 1668089732
transform 1 0 2080 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_847
timestamp 1668089732
transform 1 0 2080 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_848
timestamp 1668089732
transform 1 0 2080 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_849
timestamp 1668089732
transform 1 0 2080 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_850
timestamp 1668089732
transform 1 0 2080 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_851
timestamp 1668089732
transform 1 0 2080 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_852
timestamp 1668089732
transform 1 0 2080 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_853
timestamp 1668089732
transform 1 0 2080 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_854
timestamp 1668089732
transform 1 0 2080 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_855
timestamp 1668089732
transform 1 0 2080 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_856
timestamp 1668089732
transform 1 0 2080 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_857
timestamp 1668089732
transform 1 0 2080 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_858
timestamp 1668089732
transform 1 0 2080 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_859
timestamp 1668089732
transform 1 0 2080 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_860
timestamp 1668089732
transform 1 0 2080 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_861
timestamp 1668089732
transform 1 0 2080 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_862
timestamp 1668089732
transform 1 0 2080 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_863
timestamp 1668089732
transform 1 0 2080 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_864
timestamp 1668089732
transform 1 0 2080 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_865
timestamp 1668089732
transform 1 0 2080 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_866
timestamp 1668089732
transform 1 0 2080 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_867
timestamp 1668089732
transform 1 0 2080 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_868
timestamp 1668089732
transform 1 0 2240 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_869
timestamp 1668089732
transform 1 0 2240 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_870
timestamp 1668089732
transform 1 0 2240 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_871
timestamp 1668089732
transform 1 0 2240 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_872
timestamp 1668089732
transform 1 0 2240 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_873
timestamp 1668089732
transform 1 0 2240 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_874
timestamp 1668089732
transform 1 0 2240 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_875
timestamp 1668089732
transform 1 0 2240 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_876
timestamp 1668089732
transform 1 0 2240 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_877
timestamp 1668089732
transform 1 0 2240 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_878
timestamp 1668089732
transform 1 0 2240 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_879
timestamp 1668089732
transform 1 0 2240 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_880
timestamp 1668089732
transform 1 0 2240 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_881
timestamp 1668089732
transform 1 0 2240 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_882
timestamp 1668089732
transform 1 0 2240 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_883
timestamp 1668089732
transform 1 0 2240 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_884
timestamp 1668089732
transform 1 0 2240 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_885
timestamp 1668089732
transform 1 0 2240 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_886
timestamp 1668089732
transform 1 0 2240 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_887
timestamp 1668089732
transform 1 0 2240 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_888
timestamp 1668089732
transform 1 0 2240 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_889
timestamp 1668089732
transform 1 0 2240 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_890
timestamp 1668089732
transform 1 0 2240 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_891
timestamp 1668089732
transform 1 0 2240 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_892
timestamp 1668089732
transform 1 0 2240 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_893
timestamp 1668089732
transform 1 0 2240 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_894
timestamp 1668089732
transform 1 0 2240 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_895
timestamp 1668089732
transform 1 0 2240 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_896
timestamp 1668089732
transform 1 0 2240 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_897
timestamp 1668089732
transform 1 0 2240 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_898
timestamp 1668089732
transform 1 0 2240 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_899
timestamp 1668089732
transform 1 0 2240 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_900
timestamp 1668089732
transform 1 0 2240 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_901
timestamp 1668089732
transform 1 0 2240 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_902
timestamp 1668089732
transform 1 0 2240 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_903
timestamp 1668089732
transform 1 0 2240 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_904
timestamp 1668089732
transform 1 0 2240 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_905
timestamp 1668089732
transform 1 0 2240 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_906
timestamp 1668089732
transform 1 0 2240 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_907
timestamp 1668089732
transform 1 0 2240 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_908
timestamp 1668089732
transform 1 0 2240 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_909
timestamp 1668089732
transform 1 0 2240 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_910
timestamp 1668089732
transform 1 0 2240 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_911
timestamp 1668089732
transform 1 0 2240 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_912
timestamp 1668089732
transform 1 0 2240 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_913
timestamp 1668089732
transform 1 0 2240 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_914
timestamp 1668089732
transform 1 0 2240 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_915
timestamp 1668089732
transform 1 0 2240 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_916
timestamp 1668089732
transform 1 0 2240 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_917
timestamp 1668089732
transform 1 0 2240 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_918
timestamp 1668089732
transform 1 0 2240 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_919
timestamp 1668089732
transform 1 0 2240 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_920
timestamp 1668089732
transform 1 0 2240 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_921
timestamp 1668089732
transform 1 0 2240 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_922
timestamp 1668089732
transform 1 0 2240 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_923
timestamp 1668089732
transform 1 0 2240 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_924
timestamp 1668089732
transform 1 0 2240 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_925
timestamp 1668089732
transform 1 0 2240 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_926
timestamp 1668089732
transform 1 0 2240 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_927
timestamp 1668089732
transform 1 0 2240 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_928
timestamp 1668089732
transform 1 0 2240 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_929
timestamp 1668089732
transform 1 0 2240 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_930
timestamp 1668089732
transform 1 0 2400 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_931
timestamp 1668089732
transform 1 0 2400 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_932
timestamp 1668089732
transform 1 0 2400 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_933
timestamp 1668089732
transform 1 0 2400 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_934
timestamp 1668089732
transform 1 0 2400 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_935
timestamp 1668089732
transform 1 0 2400 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_936
timestamp 1668089732
transform 1 0 2400 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_937
timestamp 1668089732
transform 1 0 2400 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_938
timestamp 1668089732
transform 1 0 2400 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_939
timestamp 1668089732
transform 1 0 2400 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_940
timestamp 1668089732
transform 1 0 2400 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_941
timestamp 1668089732
transform 1 0 2400 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_942
timestamp 1668089732
transform 1 0 2400 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_943
timestamp 1668089732
transform 1 0 2400 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_944
timestamp 1668089732
transform 1 0 2400 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_945
timestamp 1668089732
transform 1 0 2400 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_946
timestamp 1668089732
transform 1 0 2400 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_947
timestamp 1668089732
transform 1 0 2400 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_948
timestamp 1668089732
transform 1 0 2400 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_949
timestamp 1668089732
transform 1 0 2400 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_950
timestamp 1668089732
transform 1 0 2400 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_951
timestamp 1668089732
transform 1 0 2400 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_952
timestamp 1668089732
transform 1 0 2400 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_953
timestamp 1668089732
transform 1 0 2400 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_954
timestamp 1668089732
transform 1 0 2400 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_955
timestamp 1668089732
transform 1 0 2400 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_956
timestamp 1668089732
transform 1 0 2400 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_957
timestamp 1668089732
transform 1 0 2400 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_958
timestamp 1668089732
transform 1 0 2400 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_959
timestamp 1668089732
transform 1 0 2400 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_960
timestamp 1668089732
transform 1 0 2400 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_961
timestamp 1668089732
transform 1 0 2400 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_962
timestamp 1668089732
transform 1 0 2400 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_963
timestamp 1668089732
transform 1 0 2400 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_964
timestamp 1668089732
transform 1 0 2400 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_965
timestamp 1668089732
transform 1 0 2400 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_966
timestamp 1668089732
transform 1 0 2400 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_967
timestamp 1668089732
transform 1 0 2400 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_968
timestamp 1668089732
transform 1 0 2400 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_969
timestamp 1668089732
transform 1 0 2400 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_970
timestamp 1668089732
transform 1 0 2400 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_971
timestamp 1668089732
transform 1 0 2400 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_972
timestamp 1668089732
transform 1 0 2400 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_973
timestamp 1668089732
transform 1 0 2400 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_974
timestamp 1668089732
transform 1 0 2400 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_975
timestamp 1668089732
transform 1 0 2400 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_976
timestamp 1668089732
transform 1 0 2400 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_977
timestamp 1668089732
transform 1 0 2400 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_978
timestamp 1668089732
transform 1 0 2400 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_979
timestamp 1668089732
transform 1 0 2400 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_980
timestamp 1668089732
transform 1 0 2400 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_981
timestamp 1668089732
transform 1 0 2400 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_982
timestamp 1668089732
transform 1 0 2400 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_983
timestamp 1668089732
transform 1 0 2400 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_984
timestamp 1668089732
transform 1 0 2400 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_985
timestamp 1668089732
transform 1 0 2400 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_986
timestamp 1668089732
transform 1 0 2400 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_987
timestamp 1668089732
transform 1 0 2400 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_988
timestamp 1668089732
transform 1 0 2400 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_989
timestamp 1668089732
transform 1 0 2400 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_990
timestamp 1668089732
transform 1 0 2400 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_991
timestamp 1668089732
transform 1 0 2400 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_992
timestamp 1668089732
transform 1 0 2560 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_993
timestamp 1668089732
transform 1 0 2560 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_994
timestamp 1668089732
transform 1 0 2560 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_995
timestamp 1668089732
transform 1 0 2560 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_996
timestamp 1668089732
transform 1 0 2560 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_997
timestamp 1668089732
transform 1 0 2560 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_998
timestamp 1668089732
transform 1 0 2560 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_999
timestamp 1668089732
transform 1 0 2560 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_1000
timestamp 1668089732
transform 1 0 2560 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_1001
timestamp 1668089732
transform 1 0 2560 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_1002
timestamp 1668089732
transform 1 0 2560 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_1003
timestamp 1668089732
transform 1 0 2560 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_1004
timestamp 1668089732
transform 1 0 2560 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_1005
timestamp 1668089732
transform 1 0 2560 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_1006
timestamp 1668089732
transform 1 0 2560 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_1007
timestamp 1668089732
transform 1 0 2560 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_1008
timestamp 1668089732
transform 1 0 2560 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_1009
timestamp 1668089732
transform 1 0 2560 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_1010
timestamp 1668089732
transform 1 0 2560 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_1011
timestamp 1668089732
transform 1 0 2560 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_1012
timestamp 1668089732
transform 1 0 2560 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_1013
timestamp 1668089732
transform 1 0 2560 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_1014
timestamp 1668089732
transform 1 0 2560 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_1015
timestamp 1668089732
transform 1 0 2560 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_1016
timestamp 1668089732
transform 1 0 2560 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_1017
timestamp 1668089732
transform 1 0 2560 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_1018
timestamp 1668089732
transform 1 0 2560 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_1019
timestamp 1668089732
transform 1 0 2560 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_1020
timestamp 1668089732
transform 1 0 2560 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_1021
timestamp 1668089732
transform 1 0 2560 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_1022
timestamp 1668089732
transform 1 0 2560 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_1023
timestamp 1668089732
transform 1 0 2560 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_1024
timestamp 1668089732
transform 1 0 2560 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_1025
timestamp 1668089732
transform 1 0 2560 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_1026
timestamp 1668089732
transform 1 0 2560 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_1027
timestamp 1668089732
transform 1 0 2560 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_1028
timestamp 1668089732
transform 1 0 2560 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_1029
timestamp 1668089732
transform 1 0 2560 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_1030
timestamp 1668089732
transform 1 0 2560 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_1031
timestamp 1668089732
transform 1 0 2560 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_1032
timestamp 1668089732
transform 1 0 2560 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_1033
timestamp 1668089732
transform 1 0 2560 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_1034
timestamp 1668089732
transform 1 0 2560 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_1035
timestamp 1668089732
transform 1 0 2560 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_1036
timestamp 1668089732
transform 1 0 2560 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_1037
timestamp 1668089732
transform 1 0 2560 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_1038
timestamp 1668089732
transform 1 0 2560 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_1039
timestamp 1668089732
transform 1 0 2560 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_1040
timestamp 1668089732
transform 1 0 2560 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_1041
timestamp 1668089732
transform 1 0 2560 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_1042
timestamp 1668089732
transform 1 0 2560 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_1043
timestamp 1668089732
transform 1 0 2560 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_1044
timestamp 1668089732
transform 1 0 2560 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_1045
timestamp 1668089732
transform 1 0 2560 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_1046
timestamp 1668089732
transform 1 0 2560 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_1047
timestamp 1668089732
transform 1 0 2560 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_1048
timestamp 1668089732
transform 1 0 2560 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_1049
timestamp 1668089732
transform 1 0 2560 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_1050
timestamp 1668089732
transform 1 0 2560 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_1051
timestamp 1668089732
transform 1 0 2560 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_1052
timestamp 1668089732
transform 1 0 2560 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_1053
timestamp 1668089732
transform 1 0 2560 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_1054
timestamp 1668089732
transform 1 0 2720 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_1055
timestamp 1668089732
transform 1 0 2720 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_1056
timestamp 1668089732
transform 1 0 2720 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_1057
timestamp 1668089732
transform 1 0 2720 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_1058
timestamp 1668089732
transform 1 0 2720 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_1059
timestamp 1668089732
transform 1 0 2720 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_1060
timestamp 1668089732
transform 1 0 2720 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_1061
timestamp 1668089732
transform 1 0 2720 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_1062
timestamp 1668089732
transform 1 0 2720 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_1063
timestamp 1668089732
transform 1 0 2720 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_1064
timestamp 1668089732
transform 1 0 2720 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_1065
timestamp 1668089732
transform 1 0 2720 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_1066
timestamp 1668089732
transform 1 0 2720 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_1067
timestamp 1668089732
transform 1 0 2720 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_1068
timestamp 1668089732
transform 1 0 2720 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_1069
timestamp 1668089732
transform 1 0 2720 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_1070
timestamp 1668089732
transform 1 0 2720 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_1071
timestamp 1668089732
transform 1 0 2720 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_1072
timestamp 1668089732
transform 1 0 2720 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_1073
timestamp 1668089732
transform 1 0 2720 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_1074
timestamp 1668089732
transform 1 0 2720 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_1075
timestamp 1668089732
transform 1 0 2720 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_1076
timestamp 1668089732
transform 1 0 2720 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_1077
timestamp 1668089732
transform 1 0 2720 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_1078
timestamp 1668089732
transform 1 0 2720 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_1079
timestamp 1668089732
transform 1 0 2720 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_1080
timestamp 1668089732
transform 1 0 2720 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_1081
timestamp 1668089732
transform 1 0 2720 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_1082
timestamp 1668089732
transform 1 0 2720 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_1083
timestamp 1668089732
transform 1 0 2720 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_1084
timestamp 1668089732
transform 1 0 2720 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_1085
timestamp 1668089732
transform 1 0 2720 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_1086
timestamp 1668089732
transform 1 0 2720 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_1087
timestamp 1668089732
transform 1 0 2720 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_1088
timestamp 1668089732
transform 1 0 2720 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_1089
timestamp 1668089732
transform 1 0 2720 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_1090
timestamp 1668089732
transform 1 0 2720 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_1091
timestamp 1668089732
transform 1 0 2720 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_1092
timestamp 1668089732
transform 1 0 2720 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_1093
timestamp 1668089732
transform 1 0 2720 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_1094
timestamp 1668089732
transform 1 0 2720 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_1095
timestamp 1668089732
transform 1 0 2720 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_1096
timestamp 1668089732
transform 1 0 2720 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_1097
timestamp 1668089732
transform 1 0 2720 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_1098
timestamp 1668089732
transform 1 0 2720 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_1099
timestamp 1668089732
transform 1 0 2720 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_1100
timestamp 1668089732
transform 1 0 2720 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_1101
timestamp 1668089732
transform 1 0 2720 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_1102
timestamp 1668089732
transform 1 0 2720 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_1103
timestamp 1668089732
transform 1 0 2720 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_1104
timestamp 1668089732
transform 1 0 2720 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_1105
timestamp 1668089732
transform 1 0 2720 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_1106
timestamp 1668089732
transform 1 0 2720 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_1107
timestamp 1668089732
transform 1 0 2720 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_1108
timestamp 1668089732
transform 1 0 2720 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_1109
timestamp 1668089732
transform 1 0 2720 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_1110
timestamp 1668089732
transform 1 0 2720 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_1111
timestamp 1668089732
transform 1 0 2720 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_1112
timestamp 1668089732
transform 1 0 2720 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_1113
timestamp 1668089732
transform 1 0 2720 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_1114
timestamp 1668089732
transform 1 0 2720 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_1115
timestamp 1668089732
transform 1 0 2720 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_1116
timestamp 1668089732
transform 1 0 2880 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_1117
timestamp 1668089732
transform 1 0 2880 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_1118
timestamp 1668089732
transform 1 0 2880 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_1119
timestamp 1668089732
transform 1 0 2880 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_1120
timestamp 1668089732
transform 1 0 2880 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_1121
timestamp 1668089732
transform 1 0 2880 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_1122
timestamp 1668089732
transform 1 0 2880 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_1123
timestamp 1668089732
transform 1 0 2880 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_1124
timestamp 1668089732
transform 1 0 2880 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_1125
timestamp 1668089732
transform 1 0 2880 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_1126
timestamp 1668089732
transform 1 0 2880 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_1127
timestamp 1668089732
transform 1 0 2880 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_1128
timestamp 1668089732
transform 1 0 2880 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_1129
timestamp 1668089732
transform 1 0 2880 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_1130
timestamp 1668089732
transform 1 0 2880 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_1131
timestamp 1668089732
transform 1 0 2880 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_1132
timestamp 1668089732
transform 1 0 2880 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_1133
timestamp 1668089732
transform 1 0 2880 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_1134
timestamp 1668089732
transform 1 0 2880 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_1135
timestamp 1668089732
transform 1 0 2880 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_1136
timestamp 1668089732
transform 1 0 2880 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_1137
timestamp 1668089732
transform 1 0 2880 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_1138
timestamp 1668089732
transform 1 0 2880 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_1139
timestamp 1668089732
transform 1 0 2880 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_1140
timestamp 1668089732
transform 1 0 2880 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_1141
timestamp 1668089732
transform 1 0 2880 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_1142
timestamp 1668089732
transform 1 0 2880 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_1143
timestamp 1668089732
transform 1 0 2880 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_1144
timestamp 1668089732
transform 1 0 2880 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_1145
timestamp 1668089732
transform 1 0 2880 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_1146
timestamp 1668089732
transform 1 0 2880 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_1147
timestamp 1668089732
transform 1 0 2880 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_1148
timestamp 1668089732
transform 1 0 2880 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_1149
timestamp 1668089732
transform 1 0 2880 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_1150
timestamp 1668089732
transform 1 0 2880 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_1151
timestamp 1668089732
transform 1 0 2880 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_1152
timestamp 1668089732
transform 1 0 2880 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_1153
timestamp 1668089732
transform 1 0 2880 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_1154
timestamp 1668089732
transform 1 0 2880 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_1155
timestamp 1668089732
transform 1 0 2880 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_1156
timestamp 1668089732
transform 1 0 2880 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_1157
timestamp 1668089732
transform 1 0 2880 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_1158
timestamp 1668089732
transform 1 0 2880 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_1159
timestamp 1668089732
transform 1 0 2880 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_1160
timestamp 1668089732
transform 1 0 2880 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_1161
timestamp 1668089732
transform 1 0 2880 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_1162
timestamp 1668089732
transform 1 0 2880 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_1163
timestamp 1668089732
transform 1 0 2880 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_1164
timestamp 1668089732
transform 1 0 2880 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_1165
timestamp 1668089732
transform 1 0 2880 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_1166
timestamp 1668089732
transform 1 0 2880 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_1167
timestamp 1668089732
transform 1 0 2880 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_1168
timestamp 1668089732
transform 1 0 2880 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_1169
timestamp 1668089732
transform 1 0 2880 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_1170
timestamp 1668089732
transform 1 0 2880 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_1171
timestamp 1668089732
transform 1 0 2880 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_1172
timestamp 1668089732
transform 1 0 2880 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_1173
timestamp 1668089732
transform 1 0 2880 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_1174
timestamp 1668089732
transform 1 0 2880 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_1175
timestamp 1668089732
transform 1 0 2880 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_1176
timestamp 1668089732
transform 1 0 2880 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_1177
timestamp 1668089732
transform 1 0 2880 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_1178
timestamp 1668089732
transform 1 0 3040 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_1179
timestamp 1668089732
transform 1 0 3040 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_1180
timestamp 1668089732
transform 1 0 3040 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_1181
timestamp 1668089732
transform 1 0 3040 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_1182
timestamp 1668089732
transform 1 0 3040 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_1183
timestamp 1668089732
transform 1 0 3040 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_1184
timestamp 1668089732
transform 1 0 3040 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_1185
timestamp 1668089732
transform 1 0 3040 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_1186
timestamp 1668089732
transform 1 0 3040 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_1187
timestamp 1668089732
transform 1 0 3040 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_1188
timestamp 1668089732
transform 1 0 3040 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_1189
timestamp 1668089732
transform 1 0 3040 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_1190
timestamp 1668089732
transform 1 0 3040 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_1191
timestamp 1668089732
transform 1 0 3040 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_1192
timestamp 1668089732
transform 1 0 3040 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_1193
timestamp 1668089732
transform 1 0 3040 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_1194
timestamp 1668089732
transform 1 0 3040 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_1195
timestamp 1668089732
transform 1 0 3040 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_1196
timestamp 1668089732
transform 1 0 3040 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_1197
timestamp 1668089732
transform 1 0 3040 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_1198
timestamp 1668089732
transform 1 0 3040 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_1199
timestamp 1668089732
transform 1 0 3040 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_1200
timestamp 1668089732
transform 1 0 3040 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_1201
timestamp 1668089732
transform 1 0 3040 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_1202
timestamp 1668089732
transform 1 0 3040 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_1203
timestamp 1668089732
transform 1 0 3040 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_1204
timestamp 1668089732
transform 1 0 3040 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_1205
timestamp 1668089732
transform 1 0 3040 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_1206
timestamp 1668089732
transform 1 0 3040 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_1207
timestamp 1668089732
transform 1 0 3040 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_1208
timestamp 1668089732
transform 1 0 3040 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_1209
timestamp 1668089732
transform 1 0 3040 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_1210
timestamp 1668089732
transform 1 0 3040 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_1211
timestamp 1668089732
transform 1 0 3040 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_1212
timestamp 1668089732
transform 1 0 3040 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_1213
timestamp 1668089732
transform 1 0 3040 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_1214
timestamp 1668089732
transform 1 0 3040 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_1215
timestamp 1668089732
transform 1 0 3040 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_1216
timestamp 1668089732
transform 1 0 3040 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_1217
timestamp 1668089732
transform 1 0 3040 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_1218
timestamp 1668089732
transform 1 0 3040 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_1219
timestamp 1668089732
transform 1 0 3040 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_1220
timestamp 1668089732
transform 1 0 3040 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_1221
timestamp 1668089732
transform 1 0 3040 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_1222
timestamp 1668089732
transform 1 0 3040 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_1223
timestamp 1668089732
transform 1 0 3040 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_1224
timestamp 1668089732
transform 1 0 3040 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_1225
timestamp 1668089732
transform 1 0 3040 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_1226
timestamp 1668089732
transform 1 0 3040 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_1227
timestamp 1668089732
transform 1 0 3040 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_1228
timestamp 1668089732
transform 1 0 3040 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_1229
timestamp 1668089732
transform 1 0 3040 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_1230
timestamp 1668089732
transform 1 0 3040 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_1231
timestamp 1668089732
transform 1 0 3040 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_1232
timestamp 1668089732
transform 1 0 3040 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_1233
timestamp 1668089732
transform 1 0 3040 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_1234
timestamp 1668089732
transform 1 0 3040 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_1235
timestamp 1668089732
transform 1 0 3040 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_1236
timestamp 1668089732
transform 1 0 3040 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_1237
timestamp 1668089732
transform 1 0 3040 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_1238
timestamp 1668089732
transform 1 0 3040 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_1239
timestamp 1668089732
transform 1 0 3040 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_1240
timestamp 1668089732
transform 1 0 3200 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_1241
timestamp 1668089732
transform 1 0 3200 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_1242
timestamp 1668089732
transform 1 0 3200 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_1243
timestamp 1668089732
transform 1 0 3200 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_1244
timestamp 1668089732
transform 1 0 3200 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_1245
timestamp 1668089732
transform 1 0 3200 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_1246
timestamp 1668089732
transform 1 0 3200 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_1247
timestamp 1668089732
transform 1 0 3200 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_1248
timestamp 1668089732
transform 1 0 3200 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_1249
timestamp 1668089732
transform 1 0 3200 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_1250
timestamp 1668089732
transform 1 0 3200 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_1251
timestamp 1668089732
transform 1 0 3200 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_1252
timestamp 1668089732
transform 1 0 3200 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_1253
timestamp 1668089732
transform 1 0 3200 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_1254
timestamp 1668089732
transform 1 0 3200 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_1255
timestamp 1668089732
transform 1 0 3200 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_1256
timestamp 1668089732
transform 1 0 3200 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_1257
timestamp 1668089732
transform 1 0 3200 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_1258
timestamp 1668089732
transform 1 0 3200 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_1259
timestamp 1668089732
transform 1 0 3200 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_1260
timestamp 1668089732
transform 1 0 3200 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_1261
timestamp 1668089732
transform 1 0 3200 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_1262
timestamp 1668089732
transform 1 0 3200 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_1263
timestamp 1668089732
transform 1 0 3200 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_1264
timestamp 1668089732
transform 1 0 3200 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_1265
timestamp 1668089732
transform 1 0 3200 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_1266
timestamp 1668089732
transform 1 0 3200 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_1267
timestamp 1668089732
transform 1 0 3200 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_1268
timestamp 1668089732
transform 1 0 3200 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_1269
timestamp 1668089732
transform 1 0 3200 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_1270
timestamp 1668089732
transform 1 0 3200 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_1271
timestamp 1668089732
transform 1 0 3200 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_1272
timestamp 1668089732
transform 1 0 3200 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_1273
timestamp 1668089732
transform 1 0 3200 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_1274
timestamp 1668089732
transform 1 0 3200 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_1275
timestamp 1668089732
transform 1 0 3200 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_1276
timestamp 1668089732
transform 1 0 3200 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_1277
timestamp 1668089732
transform 1 0 3200 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_1278
timestamp 1668089732
transform 1 0 3200 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_1279
timestamp 1668089732
transform 1 0 3200 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_1280
timestamp 1668089732
transform 1 0 3200 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_1281
timestamp 1668089732
transform 1 0 3200 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_1282
timestamp 1668089732
transform 1 0 3200 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_1283
timestamp 1668089732
transform 1 0 3200 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_1284
timestamp 1668089732
transform 1 0 3200 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_1285
timestamp 1668089732
transform 1 0 3200 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_1286
timestamp 1668089732
transform 1 0 3200 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_1287
timestamp 1668089732
transform 1 0 3200 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_1288
timestamp 1668089732
transform 1 0 3200 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_1289
timestamp 1668089732
transform 1 0 3200 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_1290
timestamp 1668089732
transform 1 0 3200 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_1291
timestamp 1668089732
transform 1 0 3200 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_1292
timestamp 1668089732
transform 1 0 3200 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_1293
timestamp 1668089732
transform 1 0 3200 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_1294
timestamp 1668089732
transform 1 0 3200 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_1295
timestamp 1668089732
transform 1 0 3200 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_1296
timestamp 1668089732
transform 1 0 3200 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_1297
timestamp 1668089732
transform 1 0 3200 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_1298
timestamp 1668089732
transform 1 0 3200 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_1299
timestamp 1668089732
transform 1 0 3200 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_1300
timestamp 1668089732
transform 1 0 3200 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_1301
timestamp 1668089732
transform 1 0 3200 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_1302
timestamp 1668089732
transform 1 0 3360 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_1303
timestamp 1668089732
transform 1 0 3360 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_1304
timestamp 1668089732
transform 1 0 3360 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_1305
timestamp 1668089732
transform 1 0 3360 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_1306
timestamp 1668089732
transform 1 0 3360 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_1307
timestamp 1668089732
transform 1 0 3360 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_1308
timestamp 1668089732
transform 1 0 3360 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_1309
timestamp 1668089732
transform 1 0 3360 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_1310
timestamp 1668089732
transform 1 0 3360 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_1311
timestamp 1668089732
transform 1 0 3360 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_1312
timestamp 1668089732
transform 1 0 3360 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_1313
timestamp 1668089732
transform 1 0 3360 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_1314
timestamp 1668089732
transform 1 0 3360 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_1315
timestamp 1668089732
transform 1 0 3360 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_1316
timestamp 1668089732
transform 1 0 3360 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_1317
timestamp 1668089732
transform 1 0 3360 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_1318
timestamp 1668089732
transform 1 0 3360 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_1319
timestamp 1668089732
transform 1 0 3360 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_1320
timestamp 1668089732
transform 1 0 3360 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_1321
timestamp 1668089732
transform 1 0 3360 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_1322
timestamp 1668089732
transform 1 0 3360 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_1323
timestamp 1668089732
transform 1 0 3360 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_1324
timestamp 1668089732
transform 1 0 3360 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_1325
timestamp 1668089732
transform 1 0 3360 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_1326
timestamp 1668089732
transform 1 0 3360 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_1327
timestamp 1668089732
transform 1 0 3360 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_1328
timestamp 1668089732
transform 1 0 3360 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_1329
timestamp 1668089732
transform 1 0 3360 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_1330
timestamp 1668089732
transform 1 0 3360 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_1331
timestamp 1668089732
transform 1 0 3360 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_1332
timestamp 1668089732
transform 1 0 3360 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_1333
timestamp 1668089732
transform 1 0 3360 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_1334
timestamp 1668089732
transform 1 0 3360 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_1335
timestamp 1668089732
transform 1 0 3360 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_1336
timestamp 1668089732
transform 1 0 3360 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_1337
timestamp 1668089732
transform 1 0 3360 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_1338
timestamp 1668089732
transform 1 0 3360 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_1339
timestamp 1668089732
transform 1 0 3360 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_1340
timestamp 1668089732
transform 1 0 3360 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_1341
timestamp 1668089732
transform 1 0 3360 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_1342
timestamp 1668089732
transform 1 0 3360 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_1343
timestamp 1668089732
transform 1 0 3360 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_1344
timestamp 1668089732
transform 1 0 3360 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_1345
timestamp 1668089732
transform 1 0 3360 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_1346
timestamp 1668089732
transform 1 0 3360 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_1347
timestamp 1668089732
transform 1 0 3360 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_1348
timestamp 1668089732
transform 1 0 3360 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_1349
timestamp 1668089732
transform 1 0 3360 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_1350
timestamp 1668089732
transform 1 0 3360 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_1351
timestamp 1668089732
transform 1 0 3360 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_1352
timestamp 1668089732
transform 1 0 3360 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_1353
timestamp 1668089732
transform 1 0 3360 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_1354
timestamp 1668089732
transform 1 0 3360 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_1355
timestamp 1668089732
transform 1 0 3360 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_1356
timestamp 1668089732
transform 1 0 3360 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_1357
timestamp 1668089732
transform 1 0 3360 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_1358
timestamp 1668089732
transform 1 0 3360 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_1359
timestamp 1668089732
transform 1 0 3360 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_1360
timestamp 1668089732
transform 1 0 3360 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_1361
timestamp 1668089732
transform 1 0 3360 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_1362
timestamp 1668089732
transform 1 0 3360 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_1363
timestamp 1668089732
transform 1 0 3360 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_1364
timestamp 1668089732
transform 1 0 3520 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_1365
timestamp 1668089732
transform 1 0 3520 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_1366
timestamp 1668089732
transform 1 0 3520 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_1367
timestamp 1668089732
transform 1 0 3520 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_1368
timestamp 1668089732
transform 1 0 3520 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_1369
timestamp 1668089732
transform 1 0 3520 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_1370
timestamp 1668089732
transform 1 0 3520 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_1371
timestamp 1668089732
transform 1 0 3520 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_1372
timestamp 1668089732
transform 1 0 3520 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_1373
timestamp 1668089732
transform 1 0 3520 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_1374
timestamp 1668089732
transform 1 0 3520 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_1375
timestamp 1668089732
transform 1 0 3520 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_1376
timestamp 1668089732
transform 1 0 3520 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_1377
timestamp 1668089732
transform 1 0 3520 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_1378
timestamp 1668089732
transform 1 0 3520 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_1379
timestamp 1668089732
transform 1 0 3520 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_1380
timestamp 1668089732
transform 1 0 3520 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_1381
timestamp 1668089732
transform 1 0 3520 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_1382
timestamp 1668089732
transform 1 0 3520 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_1383
timestamp 1668089732
transform 1 0 3520 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_1384
timestamp 1668089732
transform 1 0 3520 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_1385
timestamp 1668089732
transform 1 0 3520 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_1386
timestamp 1668089732
transform 1 0 3520 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_1387
timestamp 1668089732
transform 1 0 3520 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_1388
timestamp 1668089732
transform 1 0 3520 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_1389
timestamp 1668089732
transform 1 0 3520 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_1390
timestamp 1668089732
transform 1 0 3520 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_1391
timestamp 1668089732
transform 1 0 3520 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_1392
timestamp 1668089732
transform 1 0 3520 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_1393
timestamp 1668089732
transform 1 0 3520 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_1394
timestamp 1668089732
transform 1 0 3520 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_1395
timestamp 1668089732
transform 1 0 3520 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_1396
timestamp 1668089732
transform 1 0 3520 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_1397
timestamp 1668089732
transform 1 0 3520 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_1398
timestamp 1668089732
transform 1 0 3520 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_1399
timestamp 1668089732
transform 1 0 3520 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_1400
timestamp 1668089732
transform 1 0 3520 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_1401
timestamp 1668089732
transform 1 0 3520 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_1402
timestamp 1668089732
transform 1 0 3520 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_1403
timestamp 1668089732
transform 1 0 3520 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_1404
timestamp 1668089732
transform 1 0 3520 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_1405
timestamp 1668089732
transform 1 0 3520 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_1406
timestamp 1668089732
transform 1 0 3520 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_1407
timestamp 1668089732
transform 1 0 3520 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_1408
timestamp 1668089732
transform 1 0 3520 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_1409
timestamp 1668089732
transform 1 0 3520 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_1410
timestamp 1668089732
transform 1 0 3520 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_1411
timestamp 1668089732
transform 1 0 3520 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_1412
timestamp 1668089732
transform 1 0 3520 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_1413
timestamp 1668089732
transform 1 0 3520 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_1414
timestamp 1668089732
transform 1 0 3520 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_1415
timestamp 1668089732
transform 1 0 3520 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_1416
timestamp 1668089732
transform 1 0 3520 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_1417
timestamp 1668089732
transform 1 0 3520 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_1418
timestamp 1668089732
transform 1 0 3520 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_1419
timestamp 1668089732
transform 1 0 3520 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_1420
timestamp 1668089732
transform 1 0 3520 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_1421
timestamp 1668089732
transform 1 0 3520 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_1422
timestamp 1668089732
transform 1 0 3520 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_1423
timestamp 1668089732
transform 1 0 3520 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_1424
timestamp 1668089732
transform 1 0 3520 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_1425
timestamp 1668089732
transform 1 0 3520 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_1426
timestamp 1668089732
transform 1 0 3680 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_1427
timestamp 1668089732
transform 1 0 3680 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_1428
timestamp 1668089732
transform 1 0 3680 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_1429
timestamp 1668089732
transform 1 0 3680 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_1430
timestamp 1668089732
transform 1 0 3680 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_1431
timestamp 1668089732
transform 1 0 3680 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_1432
timestamp 1668089732
transform 1 0 3680 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_1433
timestamp 1668089732
transform 1 0 3680 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_1434
timestamp 1668089732
transform 1 0 3680 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_1435
timestamp 1668089732
transform 1 0 3680 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_1436
timestamp 1668089732
transform 1 0 3680 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_1437
timestamp 1668089732
transform 1 0 3680 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_1438
timestamp 1668089732
transform 1 0 3680 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_1439
timestamp 1668089732
transform 1 0 3680 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_1440
timestamp 1668089732
transform 1 0 3680 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_1441
timestamp 1668089732
transform 1 0 3680 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_1442
timestamp 1668089732
transform 1 0 3680 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_1443
timestamp 1668089732
transform 1 0 3680 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_1444
timestamp 1668089732
transform 1 0 3680 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_1445
timestamp 1668089732
transform 1 0 3680 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_1446
timestamp 1668089732
transform 1 0 3680 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_1447
timestamp 1668089732
transform 1 0 3680 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_1448
timestamp 1668089732
transform 1 0 3680 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_1449
timestamp 1668089732
transform 1 0 3680 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_1450
timestamp 1668089732
transform 1 0 3680 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_1451
timestamp 1668089732
transform 1 0 3680 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_1452
timestamp 1668089732
transform 1 0 3680 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_1453
timestamp 1668089732
transform 1 0 3680 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_1454
timestamp 1668089732
transform 1 0 3680 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_1455
timestamp 1668089732
transform 1 0 3680 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_1456
timestamp 1668089732
transform 1 0 3680 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_1457
timestamp 1668089732
transform 1 0 3680 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_1458
timestamp 1668089732
transform 1 0 3680 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_1459
timestamp 1668089732
transform 1 0 3680 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_1460
timestamp 1668089732
transform 1 0 3680 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_1461
timestamp 1668089732
transform 1 0 3680 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_1462
timestamp 1668089732
transform 1 0 3680 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_1463
timestamp 1668089732
transform 1 0 3680 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_1464
timestamp 1668089732
transform 1 0 3680 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_1465
timestamp 1668089732
transform 1 0 3680 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_1466
timestamp 1668089732
transform 1 0 3680 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_1467
timestamp 1668089732
transform 1 0 3680 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_1468
timestamp 1668089732
transform 1 0 3680 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_1469
timestamp 1668089732
transform 1 0 3680 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_1470
timestamp 1668089732
transform 1 0 3680 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_1471
timestamp 1668089732
transform 1 0 3680 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_1472
timestamp 1668089732
transform 1 0 3680 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_1473
timestamp 1668089732
transform 1 0 3680 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_1474
timestamp 1668089732
transform 1 0 3680 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_1475
timestamp 1668089732
transform 1 0 3680 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_1476
timestamp 1668089732
transform 1 0 3680 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_1477
timestamp 1668089732
transform 1 0 3680 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_1478
timestamp 1668089732
transform 1 0 3680 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_1479
timestamp 1668089732
transform 1 0 3680 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_1480
timestamp 1668089732
transform 1 0 3680 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_1481
timestamp 1668089732
transform 1 0 3680 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_1482
timestamp 1668089732
transform 1 0 3680 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_1483
timestamp 1668089732
transform 1 0 3680 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_1484
timestamp 1668089732
transform 1 0 3680 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_1485
timestamp 1668089732
transform 1 0 3680 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_1486
timestamp 1668089732
transform 1 0 3680 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_1487
timestamp 1668089732
transform 1 0 3680 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_1488
timestamp 1668089732
transform 1 0 3840 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_1489
timestamp 1668089732
transform 1 0 3840 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_1490
timestamp 1668089732
transform 1 0 3840 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_1491
timestamp 1668089732
transform 1 0 3840 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_1492
timestamp 1668089732
transform 1 0 3840 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_1493
timestamp 1668089732
transform 1 0 3840 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_1494
timestamp 1668089732
transform 1 0 3840 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_1495
timestamp 1668089732
transform 1 0 3840 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_1496
timestamp 1668089732
transform 1 0 3840 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_1497
timestamp 1668089732
transform 1 0 3840 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_1498
timestamp 1668089732
transform 1 0 3840 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_1499
timestamp 1668089732
transform 1 0 3840 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_1500
timestamp 1668089732
transform 1 0 3840 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_1501
timestamp 1668089732
transform 1 0 3840 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_1502
timestamp 1668089732
transform 1 0 3840 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_1503
timestamp 1668089732
transform 1 0 3840 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_1504
timestamp 1668089732
transform 1 0 3840 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_1505
timestamp 1668089732
transform 1 0 3840 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_1506
timestamp 1668089732
transform 1 0 3840 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_1507
timestamp 1668089732
transform 1 0 3840 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_1508
timestamp 1668089732
transform 1 0 3840 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_1509
timestamp 1668089732
transform 1 0 3840 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_1510
timestamp 1668089732
transform 1 0 3840 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_1511
timestamp 1668089732
transform 1 0 3840 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_1512
timestamp 1668089732
transform 1 0 3840 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_1513
timestamp 1668089732
transform 1 0 3840 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_1514
timestamp 1668089732
transform 1 0 3840 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_1515
timestamp 1668089732
transform 1 0 3840 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_1516
timestamp 1668089732
transform 1 0 3840 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_1517
timestamp 1668089732
transform 1 0 3840 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_1518
timestamp 1668089732
transform 1 0 3840 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_1519
timestamp 1668089732
transform 1 0 3840 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_1520
timestamp 1668089732
transform 1 0 3840 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_1521
timestamp 1668089732
transform 1 0 3840 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_1522
timestamp 1668089732
transform 1 0 3840 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_1523
timestamp 1668089732
transform 1 0 3840 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_1524
timestamp 1668089732
transform 1 0 3840 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_1525
timestamp 1668089732
transform 1 0 3840 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_1526
timestamp 1668089732
transform 1 0 3840 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_1527
timestamp 1668089732
transform 1 0 3840 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_1528
timestamp 1668089732
transform 1 0 3840 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_1529
timestamp 1668089732
transform 1 0 3840 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_1530
timestamp 1668089732
transform 1 0 3840 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_1531
timestamp 1668089732
transform 1 0 3840 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_1532
timestamp 1668089732
transform 1 0 3840 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_1533
timestamp 1668089732
transform 1 0 3840 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_1534
timestamp 1668089732
transform 1 0 3840 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_1535
timestamp 1668089732
transform 1 0 3840 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_1536
timestamp 1668089732
transform 1 0 3840 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_1537
timestamp 1668089732
transform 1 0 3840 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_1538
timestamp 1668089732
transform 1 0 3840 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_1539
timestamp 1668089732
transform 1 0 3840 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_1540
timestamp 1668089732
transform 1 0 3840 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_1541
timestamp 1668089732
transform 1 0 3840 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_1542
timestamp 1668089732
transform 1 0 3840 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_1543
timestamp 1668089732
transform 1 0 3840 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_1544
timestamp 1668089732
transform 1 0 3840 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_1545
timestamp 1668089732
transform 1 0 3840 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_1546
timestamp 1668089732
transform 1 0 3840 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_1547
timestamp 1668089732
transform 1 0 3840 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_1548
timestamp 1668089732
transform 1 0 3840 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_1549
timestamp 1668089732
transform 1 0 3840 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_1550
timestamp 1668089732
transform 1 0 4000 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_1551
timestamp 1668089732
transform 1 0 4000 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_1552
timestamp 1668089732
transform 1 0 4000 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_1553
timestamp 1668089732
transform 1 0 4000 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_1554
timestamp 1668089732
transform 1 0 4000 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_1555
timestamp 1668089732
transform 1 0 4000 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_1556
timestamp 1668089732
transform 1 0 4000 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_1557
timestamp 1668089732
transform 1 0 4000 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_1558
timestamp 1668089732
transform 1 0 4000 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_1559
timestamp 1668089732
transform 1 0 4000 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_1560
timestamp 1668089732
transform 1 0 4000 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_1561
timestamp 1668089732
transform 1 0 4000 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_1562
timestamp 1668089732
transform 1 0 4000 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_1563
timestamp 1668089732
transform 1 0 4000 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_1564
timestamp 1668089732
transform 1 0 4000 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_1565
timestamp 1668089732
transform 1 0 4000 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_1566
timestamp 1668089732
transform 1 0 4000 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_1567
timestamp 1668089732
transform 1 0 4000 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_1568
timestamp 1668089732
transform 1 0 4000 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_1569
timestamp 1668089732
transform 1 0 4000 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_1570
timestamp 1668089732
transform 1 0 4000 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_1571
timestamp 1668089732
transform 1 0 4000 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_1572
timestamp 1668089732
transform 1 0 4000 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_1573
timestamp 1668089732
transform 1 0 4000 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_1574
timestamp 1668089732
transform 1 0 4000 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_1575
timestamp 1668089732
transform 1 0 4000 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_1576
timestamp 1668089732
transform 1 0 4000 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_1577
timestamp 1668089732
transform 1 0 4000 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_1578
timestamp 1668089732
transform 1 0 4000 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_1579
timestamp 1668089732
transform 1 0 4000 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_1580
timestamp 1668089732
transform 1 0 4000 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_1581
timestamp 1668089732
transform 1 0 4000 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_1582
timestamp 1668089732
transform 1 0 4000 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_1583
timestamp 1668089732
transform 1 0 4000 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_1584
timestamp 1668089732
transform 1 0 4000 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_1585
timestamp 1668089732
transform 1 0 4000 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_1586
timestamp 1668089732
transform 1 0 4000 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_1587
timestamp 1668089732
transform 1 0 4000 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_1588
timestamp 1668089732
transform 1 0 4000 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_1589
timestamp 1668089732
transform 1 0 4000 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_1590
timestamp 1668089732
transform 1 0 4000 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_1591
timestamp 1668089732
transform 1 0 4000 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_1592
timestamp 1668089732
transform 1 0 4000 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_1593
timestamp 1668089732
transform 1 0 4000 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_1594
timestamp 1668089732
transform 1 0 4000 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_1595
timestamp 1668089732
transform 1 0 4000 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_1596
timestamp 1668089732
transform 1 0 4000 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_1597
timestamp 1668089732
transform 1 0 4000 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_1598
timestamp 1668089732
transform 1 0 4000 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_1599
timestamp 1668089732
transform 1 0 4000 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_1600
timestamp 1668089732
transform 1 0 4000 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_1601
timestamp 1668089732
transform 1 0 4000 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_1602
timestamp 1668089732
transform 1 0 4000 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_1603
timestamp 1668089732
transform 1 0 4000 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_1604
timestamp 1668089732
transform 1 0 4000 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_1605
timestamp 1668089732
transform 1 0 4000 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_1606
timestamp 1668089732
transform 1 0 4000 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_1607
timestamp 1668089732
transform 1 0 4000 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_1608
timestamp 1668089732
transform 1 0 4000 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_1609
timestamp 1668089732
transform 1 0 4000 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_1610
timestamp 1668089732
transform 1 0 4000 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_1611
timestamp 1668089732
transform 1 0 4000 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_1612
timestamp 1668089732
transform 1 0 4160 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_1613
timestamp 1668089732
transform 1 0 4160 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_1614
timestamp 1668089732
transform 1 0 4160 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_1615
timestamp 1668089732
transform 1 0 4160 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_1616
timestamp 1668089732
transform 1 0 4160 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_1617
timestamp 1668089732
transform 1 0 4160 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_1618
timestamp 1668089732
transform 1 0 4160 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_1619
timestamp 1668089732
transform 1 0 4160 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_1620
timestamp 1668089732
transform 1 0 4160 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_1621
timestamp 1668089732
transform 1 0 4160 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_1622
timestamp 1668089732
transform 1 0 4160 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_1623
timestamp 1668089732
transform 1 0 4160 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_1624
timestamp 1668089732
transform 1 0 4160 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_1625
timestamp 1668089732
transform 1 0 4160 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_1626
timestamp 1668089732
transform 1 0 4160 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_1627
timestamp 1668089732
transform 1 0 4160 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_1628
timestamp 1668089732
transform 1 0 4160 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_1629
timestamp 1668089732
transform 1 0 4160 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_1630
timestamp 1668089732
transform 1 0 4160 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_1631
timestamp 1668089732
transform 1 0 4160 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_1632
timestamp 1668089732
transform 1 0 4160 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_1633
timestamp 1668089732
transform 1 0 4160 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_1634
timestamp 1668089732
transform 1 0 4160 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_1635
timestamp 1668089732
transform 1 0 4160 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_1636
timestamp 1668089732
transform 1 0 4160 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_1637
timestamp 1668089732
transform 1 0 4160 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_1638
timestamp 1668089732
transform 1 0 4160 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_1639
timestamp 1668089732
transform 1 0 4160 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_1640
timestamp 1668089732
transform 1 0 4160 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_1641
timestamp 1668089732
transform 1 0 4160 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_1642
timestamp 1668089732
transform 1 0 4160 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_1643
timestamp 1668089732
transform 1 0 4160 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_1644
timestamp 1668089732
transform 1 0 4160 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_1645
timestamp 1668089732
transform 1 0 4160 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_1646
timestamp 1668089732
transform 1 0 4160 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_1647
timestamp 1668089732
transform 1 0 4160 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_1648
timestamp 1668089732
transform 1 0 4160 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_1649
timestamp 1668089732
transform 1 0 4160 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_1650
timestamp 1668089732
transform 1 0 4160 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_1651
timestamp 1668089732
transform 1 0 4160 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_1652
timestamp 1668089732
transform 1 0 4160 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_1653
timestamp 1668089732
transform 1 0 4160 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_1654
timestamp 1668089732
transform 1 0 4160 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_1655
timestamp 1668089732
transform 1 0 4160 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_1656
timestamp 1668089732
transform 1 0 4160 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_1657
timestamp 1668089732
transform 1 0 4160 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_1658
timestamp 1668089732
transform 1 0 4160 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_1659
timestamp 1668089732
transform 1 0 4160 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_1660
timestamp 1668089732
transform 1 0 4160 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_1661
timestamp 1668089732
transform 1 0 4160 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_1662
timestamp 1668089732
transform 1 0 4160 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_1663
timestamp 1668089732
transform 1 0 4160 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_1664
timestamp 1668089732
transform 1 0 4160 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_1665
timestamp 1668089732
transform 1 0 4160 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_1666
timestamp 1668089732
transform 1 0 4160 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_1667
timestamp 1668089732
transform 1 0 4160 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_1668
timestamp 1668089732
transform 1 0 4160 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_1669
timestamp 1668089732
transform 1 0 4160 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_1670
timestamp 1668089732
transform 1 0 4160 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_1671
timestamp 1668089732
transform 1 0 4160 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_1672
timestamp 1668089732
transform 1 0 4160 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_1673
timestamp 1668089732
transform 1 0 4160 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_1674
timestamp 1668089732
transform 1 0 4320 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_1675
timestamp 1668089732
transform 1 0 4320 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_1676
timestamp 1668089732
transform 1 0 4320 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_1677
timestamp 1668089732
transform 1 0 4320 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_1678
timestamp 1668089732
transform 1 0 4320 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_1679
timestamp 1668089732
transform 1 0 4320 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_1680
timestamp 1668089732
transform 1 0 4320 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_1681
timestamp 1668089732
transform 1 0 4320 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_1682
timestamp 1668089732
transform 1 0 4320 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_1683
timestamp 1668089732
transform 1 0 4320 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_1684
timestamp 1668089732
transform 1 0 4320 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_1685
timestamp 1668089732
transform 1 0 4320 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_1686
timestamp 1668089732
transform 1 0 4320 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_1687
timestamp 1668089732
transform 1 0 4320 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_1688
timestamp 1668089732
transform 1 0 4320 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_1689
timestamp 1668089732
transform 1 0 4320 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_1690
timestamp 1668089732
transform 1 0 4320 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_1691
timestamp 1668089732
transform 1 0 4320 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_1692
timestamp 1668089732
transform 1 0 4320 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_1693
timestamp 1668089732
transform 1 0 4320 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_1694
timestamp 1668089732
transform 1 0 4320 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_1695
timestamp 1668089732
transform 1 0 4320 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_1696
timestamp 1668089732
transform 1 0 4320 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_1697
timestamp 1668089732
transform 1 0 4320 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_1698
timestamp 1668089732
transform 1 0 4320 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_1699
timestamp 1668089732
transform 1 0 4320 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_1700
timestamp 1668089732
transform 1 0 4320 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_1701
timestamp 1668089732
transform 1 0 4320 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_1702
timestamp 1668089732
transform 1 0 4320 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_1703
timestamp 1668089732
transform 1 0 4320 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_1704
timestamp 1668089732
transform 1 0 4320 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_1705
timestamp 1668089732
transform 1 0 4320 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_1706
timestamp 1668089732
transform 1 0 4320 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_1707
timestamp 1668089732
transform 1 0 4320 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_1708
timestamp 1668089732
transform 1 0 4320 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_1709
timestamp 1668089732
transform 1 0 4320 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_1710
timestamp 1668089732
transform 1 0 4320 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_1711
timestamp 1668089732
transform 1 0 4320 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_1712
timestamp 1668089732
transform 1 0 4320 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_1713
timestamp 1668089732
transform 1 0 4320 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_1714
timestamp 1668089732
transform 1 0 4320 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_1715
timestamp 1668089732
transform 1 0 4320 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_1716
timestamp 1668089732
transform 1 0 4320 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_1717
timestamp 1668089732
transform 1 0 4320 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_1718
timestamp 1668089732
transform 1 0 4320 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_1719
timestamp 1668089732
transform 1 0 4320 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_1720
timestamp 1668089732
transform 1 0 4320 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_1721
timestamp 1668089732
transform 1 0 4320 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_1722
timestamp 1668089732
transform 1 0 4320 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_1723
timestamp 1668089732
transform 1 0 4320 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_1724
timestamp 1668089732
transform 1 0 4320 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_1725
timestamp 1668089732
transform 1 0 4320 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_1726
timestamp 1668089732
transform 1 0 4320 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_1727
timestamp 1668089732
transform 1 0 4320 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_1728
timestamp 1668089732
transform 1 0 4320 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_1729
timestamp 1668089732
transform 1 0 4320 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_1730
timestamp 1668089732
transform 1 0 4320 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_1731
timestamp 1668089732
transform 1 0 4320 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_1732
timestamp 1668089732
transform 1 0 4320 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_1733
timestamp 1668089732
transform 1 0 4320 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_1734
timestamp 1668089732
transform 1 0 4320 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_1735
timestamp 1668089732
transform 1 0 4320 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_1736
timestamp 1668089732
transform 1 0 4480 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_1737
timestamp 1668089732
transform 1 0 4480 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_1738
timestamp 1668089732
transform 1 0 4480 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_1739
timestamp 1668089732
transform 1 0 4480 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_1740
timestamp 1668089732
transform 1 0 4480 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_1741
timestamp 1668089732
transform 1 0 4480 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_1742
timestamp 1668089732
transform 1 0 4480 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_1743
timestamp 1668089732
transform 1 0 4480 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_1744
timestamp 1668089732
transform 1 0 4480 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_1745
timestamp 1668089732
transform 1 0 4480 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_1746
timestamp 1668089732
transform 1 0 4480 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_1747
timestamp 1668089732
transform 1 0 4480 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_1748
timestamp 1668089732
transform 1 0 4480 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_1749
timestamp 1668089732
transform 1 0 4480 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_1750
timestamp 1668089732
transform 1 0 4480 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_1751
timestamp 1668089732
transform 1 0 4480 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_1752
timestamp 1668089732
transform 1 0 4480 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_1753
timestamp 1668089732
transform 1 0 4480 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_1754
timestamp 1668089732
transform 1 0 4480 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_1755
timestamp 1668089732
transform 1 0 4480 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_1756
timestamp 1668089732
transform 1 0 4480 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_1757
timestamp 1668089732
transform 1 0 4480 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_1758
timestamp 1668089732
transform 1 0 4480 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_1759
timestamp 1668089732
transform 1 0 4480 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_1760
timestamp 1668089732
transform 1 0 4480 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_1761
timestamp 1668089732
transform 1 0 4480 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_1762
timestamp 1668089732
transform 1 0 4480 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_1763
timestamp 1668089732
transform 1 0 4480 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_1764
timestamp 1668089732
transform 1 0 4480 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_1765
timestamp 1668089732
transform 1 0 4480 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_1766
timestamp 1668089732
transform 1 0 4480 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_1767
timestamp 1668089732
transform 1 0 4480 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_1768
timestamp 1668089732
transform 1 0 4480 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_1769
timestamp 1668089732
transform 1 0 4480 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_1770
timestamp 1668089732
transform 1 0 4480 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_1771
timestamp 1668089732
transform 1 0 4480 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_1772
timestamp 1668089732
transform 1 0 4480 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_1773
timestamp 1668089732
transform 1 0 4480 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_1774
timestamp 1668089732
transform 1 0 4480 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_1775
timestamp 1668089732
transform 1 0 4480 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_1776
timestamp 1668089732
transform 1 0 4480 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_1777
timestamp 1668089732
transform 1 0 4480 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_1778
timestamp 1668089732
transform 1 0 4480 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_1779
timestamp 1668089732
transform 1 0 4480 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_1780
timestamp 1668089732
transform 1 0 4480 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_1781
timestamp 1668089732
transform 1 0 4480 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_1782
timestamp 1668089732
transform 1 0 4480 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_1783
timestamp 1668089732
transform 1 0 4480 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_1784
timestamp 1668089732
transform 1 0 4480 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_1785
timestamp 1668089732
transform 1 0 4480 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_1786
timestamp 1668089732
transform 1 0 4480 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_1787
timestamp 1668089732
transform 1 0 4480 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_1788
timestamp 1668089732
transform 1 0 4480 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_1789
timestamp 1668089732
transform 1 0 4480 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_1790
timestamp 1668089732
transform 1 0 4480 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_1791
timestamp 1668089732
transform 1 0 4480 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_1792
timestamp 1668089732
transform 1 0 4480 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_1793
timestamp 1668089732
transform 1 0 4480 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_1794
timestamp 1668089732
transform 1 0 4480 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_1795
timestamp 1668089732
transform 1 0 4480 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_1796
timestamp 1668089732
transform 1 0 4480 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_1797
timestamp 1668089732
transform 1 0 4480 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_1798
timestamp 1668089732
transform 1 0 4640 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_1799
timestamp 1668089732
transform 1 0 4640 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_1800
timestamp 1668089732
transform 1 0 4640 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_1801
timestamp 1668089732
transform 1 0 4640 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_1802
timestamp 1668089732
transform 1 0 4640 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_1803
timestamp 1668089732
transform 1 0 4640 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_1804
timestamp 1668089732
transform 1 0 4640 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_1805
timestamp 1668089732
transform 1 0 4640 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_1806
timestamp 1668089732
transform 1 0 4640 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_1807
timestamp 1668089732
transform 1 0 4640 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_1808
timestamp 1668089732
transform 1 0 4640 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_1809
timestamp 1668089732
transform 1 0 4640 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_1810
timestamp 1668089732
transform 1 0 4640 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_1811
timestamp 1668089732
transform 1 0 4640 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_1812
timestamp 1668089732
transform 1 0 4640 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_1813
timestamp 1668089732
transform 1 0 4640 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_1814
timestamp 1668089732
transform 1 0 4640 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_1815
timestamp 1668089732
transform 1 0 4640 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_1816
timestamp 1668089732
transform 1 0 4640 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_1817
timestamp 1668089732
transform 1 0 4640 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_1818
timestamp 1668089732
transform 1 0 4640 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_1819
timestamp 1668089732
transform 1 0 4640 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_1820
timestamp 1668089732
transform 1 0 4640 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_1821
timestamp 1668089732
transform 1 0 4640 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_1822
timestamp 1668089732
transform 1 0 4640 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_1823
timestamp 1668089732
transform 1 0 4640 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_1824
timestamp 1668089732
transform 1 0 4640 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_1825
timestamp 1668089732
transform 1 0 4640 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_1826
timestamp 1668089732
transform 1 0 4640 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_1827
timestamp 1668089732
transform 1 0 4640 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_1828
timestamp 1668089732
transform 1 0 4640 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_1829
timestamp 1668089732
transform 1 0 4640 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_1830
timestamp 1668089732
transform 1 0 4640 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_1831
timestamp 1668089732
transform 1 0 4640 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_1832
timestamp 1668089732
transform 1 0 4640 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_1833
timestamp 1668089732
transform 1 0 4640 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_1834
timestamp 1668089732
transform 1 0 4640 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_1835
timestamp 1668089732
transform 1 0 4640 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_1836
timestamp 1668089732
transform 1 0 4640 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_1837
timestamp 1668089732
transform 1 0 4640 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_1838
timestamp 1668089732
transform 1 0 4640 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_1839
timestamp 1668089732
transform 1 0 4640 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_1840
timestamp 1668089732
transform 1 0 4640 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_1841
timestamp 1668089732
transform 1 0 4640 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_1842
timestamp 1668089732
transform 1 0 4640 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_1843
timestamp 1668089732
transform 1 0 4640 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_1844
timestamp 1668089732
transform 1 0 4640 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_1845
timestamp 1668089732
transform 1 0 4640 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_1846
timestamp 1668089732
transform 1 0 4640 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_1847
timestamp 1668089732
transform 1 0 4640 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_1848
timestamp 1668089732
transform 1 0 4640 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_1849
timestamp 1668089732
transform 1 0 4640 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_1850
timestamp 1668089732
transform 1 0 4640 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_1851
timestamp 1668089732
transform 1 0 4640 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_1852
timestamp 1668089732
transform 1 0 4640 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_1853
timestamp 1668089732
transform 1 0 4640 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_1854
timestamp 1668089732
transform 1 0 4640 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_1855
timestamp 1668089732
transform 1 0 4640 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_1856
timestamp 1668089732
transform 1 0 4640 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_1857
timestamp 1668089732
transform 1 0 4640 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_1858
timestamp 1668089732
transform 1 0 4640 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_1859
timestamp 1668089732
transform 1 0 4640 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_1860
timestamp 1668089732
transform 1 0 4800 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_1861
timestamp 1668089732
transform 1 0 4800 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_1862
timestamp 1668089732
transform 1 0 4800 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_1863
timestamp 1668089732
transform 1 0 4800 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_1864
timestamp 1668089732
transform 1 0 4800 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_1865
timestamp 1668089732
transform 1 0 4800 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_1866
timestamp 1668089732
transform 1 0 4800 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_1867
timestamp 1668089732
transform 1 0 4800 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_1868
timestamp 1668089732
transform 1 0 4800 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_1869
timestamp 1668089732
transform 1 0 4800 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_1870
timestamp 1668089732
transform 1 0 4800 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_1871
timestamp 1668089732
transform 1 0 4800 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_1872
timestamp 1668089732
transform 1 0 4800 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_1873
timestamp 1668089732
transform 1 0 4800 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_1874
timestamp 1668089732
transform 1 0 4800 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_1875
timestamp 1668089732
transform 1 0 4800 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_1876
timestamp 1668089732
transform 1 0 4800 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_1877
timestamp 1668089732
transform 1 0 4800 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_1878
timestamp 1668089732
transform 1 0 4800 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_1879
timestamp 1668089732
transform 1 0 4800 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_1880
timestamp 1668089732
transform 1 0 4800 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_1881
timestamp 1668089732
transform 1 0 4800 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_1882
timestamp 1668089732
transform 1 0 4800 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_1883
timestamp 1668089732
transform 1 0 4800 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_1884
timestamp 1668089732
transform 1 0 4800 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_1885
timestamp 1668089732
transform 1 0 4800 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_1886
timestamp 1668089732
transform 1 0 4800 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_1887
timestamp 1668089732
transform 1 0 4800 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_1888
timestamp 1668089732
transform 1 0 4800 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_1889
timestamp 1668089732
transform 1 0 4800 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_1890
timestamp 1668089732
transform 1 0 4800 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_1891
timestamp 1668089732
transform 1 0 4800 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_1892
timestamp 1668089732
transform 1 0 4800 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_1893
timestamp 1668089732
transform 1 0 4800 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_1894
timestamp 1668089732
transform 1 0 4800 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_1895
timestamp 1668089732
transform 1 0 4800 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_1896
timestamp 1668089732
transform 1 0 4800 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_1897
timestamp 1668089732
transform 1 0 4800 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_1898
timestamp 1668089732
transform 1 0 4800 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_1899
timestamp 1668089732
transform 1 0 4800 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_1900
timestamp 1668089732
transform 1 0 4800 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_1901
timestamp 1668089732
transform 1 0 4800 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_1902
timestamp 1668089732
transform 1 0 4800 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_1903
timestamp 1668089732
transform 1 0 4800 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_1904
timestamp 1668089732
transform 1 0 4800 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_1905
timestamp 1668089732
transform 1 0 4800 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_1906
timestamp 1668089732
transform 1 0 4800 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_1907
timestamp 1668089732
transform 1 0 4800 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_1908
timestamp 1668089732
transform 1 0 4800 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_1909
timestamp 1668089732
transform 1 0 4800 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_1910
timestamp 1668089732
transform 1 0 4800 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_1911
timestamp 1668089732
transform 1 0 4800 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_1912
timestamp 1668089732
transform 1 0 4800 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_1913
timestamp 1668089732
transform 1 0 4800 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_1914
timestamp 1668089732
transform 1 0 4800 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_1915
timestamp 1668089732
transform 1 0 4800 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_1916
timestamp 1668089732
transform 1 0 4800 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_1917
timestamp 1668089732
transform 1 0 4800 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_1918
timestamp 1668089732
transform 1 0 4800 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_1919
timestamp 1668089732
transform 1 0 4800 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_1920
timestamp 1668089732
transform 1 0 4800 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_1921
timestamp 1668089732
transform 1 0 4800 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_1922
timestamp 1668089732
transform 1 0 4960 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_1923
timestamp 1668089732
transform 1 0 4960 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_1924
timestamp 1668089732
transform 1 0 4960 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_1925
timestamp 1668089732
transform 1 0 4960 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_1926
timestamp 1668089732
transform 1 0 4960 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_1927
timestamp 1668089732
transform 1 0 4960 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_1928
timestamp 1668089732
transform 1 0 4960 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_1929
timestamp 1668089732
transform 1 0 4960 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_1930
timestamp 1668089732
transform 1 0 4960 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_1931
timestamp 1668089732
transform 1 0 4960 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_1932
timestamp 1668089732
transform 1 0 4960 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_1933
timestamp 1668089732
transform 1 0 4960 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_1934
timestamp 1668089732
transform 1 0 4960 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_1935
timestamp 1668089732
transform 1 0 4960 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_1936
timestamp 1668089732
transform 1 0 4960 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_1937
timestamp 1668089732
transform 1 0 4960 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_1938
timestamp 1668089732
transform 1 0 4960 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_1939
timestamp 1668089732
transform 1 0 4960 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_1940
timestamp 1668089732
transform 1 0 4960 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_1941
timestamp 1668089732
transform 1 0 4960 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_1942
timestamp 1668089732
transform 1 0 4960 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_1943
timestamp 1668089732
transform 1 0 4960 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_1944
timestamp 1668089732
transform 1 0 4960 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_1945
timestamp 1668089732
transform 1 0 4960 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_1946
timestamp 1668089732
transform 1 0 4960 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_1947
timestamp 1668089732
transform 1 0 4960 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_1948
timestamp 1668089732
transform 1 0 4960 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_1949
timestamp 1668089732
transform 1 0 4960 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_1950
timestamp 1668089732
transform 1 0 4960 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_1951
timestamp 1668089732
transform 1 0 4960 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_1952
timestamp 1668089732
transform 1 0 4960 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_1953
timestamp 1668089732
transform 1 0 4960 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_1954
timestamp 1668089732
transform 1 0 4960 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_1955
timestamp 1668089732
transform 1 0 4960 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_1956
timestamp 1668089732
transform 1 0 4960 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_1957
timestamp 1668089732
transform 1 0 4960 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_1958
timestamp 1668089732
transform 1 0 4960 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_1959
timestamp 1668089732
transform 1 0 4960 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_1960
timestamp 1668089732
transform 1 0 4960 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_1961
timestamp 1668089732
transform 1 0 4960 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_1962
timestamp 1668089732
transform 1 0 4960 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_1963
timestamp 1668089732
transform 1 0 4960 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_1964
timestamp 1668089732
transform 1 0 4960 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_1965
timestamp 1668089732
transform 1 0 4960 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_1966
timestamp 1668089732
transform 1 0 4960 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_1967
timestamp 1668089732
transform 1 0 4960 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_1968
timestamp 1668089732
transform 1 0 4960 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_1969
timestamp 1668089732
transform 1 0 4960 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_1970
timestamp 1668089732
transform 1 0 4960 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_1971
timestamp 1668089732
transform 1 0 4960 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_1972
timestamp 1668089732
transform 1 0 4960 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_1973
timestamp 1668089732
transform 1 0 4960 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_1974
timestamp 1668089732
transform 1 0 4960 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_1975
timestamp 1668089732
transform 1 0 4960 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_1976
timestamp 1668089732
transform 1 0 4960 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_1977
timestamp 1668089732
transform 1 0 4960 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_1978
timestamp 1668089732
transform 1 0 4960 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_1979
timestamp 1668089732
transform 1 0 4960 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_1980
timestamp 1668089732
transform 1 0 4960 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_1981
timestamp 1668089732
transform 1 0 4960 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_1982
timestamp 1668089732
transform 1 0 4960 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_1983
timestamp 1668089732
transform 1 0 4960 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_1984
timestamp 1668089732
transform 1 0 5120 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_1985
timestamp 1668089732
transform 1 0 5120 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_1986
timestamp 1668089732
transform 1 0 5120 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_1987
timestamp 1668089732
transform 1 0 5120 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_1988
timestamp 1668089732
transform 1 0 5120 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_1989
timestamp 1668089732
transform 1 0 5120 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_1990
timestamp 1668089732
transform 1 0 5120 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_1991
timestamp 1668089732
transform 1 0 5120 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_1992
timestamp 1668089732
transform 1 0 5120 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_1993
timestamp 1668089732
transform 1 0 5120 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_1994
timestamp 1668089732
transform 1 0 5120 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_1995
timestamp 1668089732
transform 1 0 5120 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_1996
timestamp 1668089732
transform 1 0 5120 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_1997
timestamp 1668089732
transform 1 0 5120 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_1998
timestamp 1668089732
transform 1 0 5120 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_1999
timestamp 1668089732
transform 1 0 5120 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_2000
timestamp 1668089732
transform 1 0 5120 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_2001
timestamp 1668089732
transform 1 0 5120 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_2002
timestamp 1668089732
transform 1 0 5120 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_2003
timestamp 1668089732
transform 1 0 5120 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_2004
timestamp 1668089732
transform 1 0 5120 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_2005
timestamp 1668089732
transform 1 0 5120 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_2006
timestamp 1668089732
transform 1 0 5120 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_2007
timestamp 1668089732
transform 1 0 5120 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_2008
timestamp 1668089732
transform 1 0 5120 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_2009
timestamp 1668089732
transform 1 0 5120 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_2010
timestamp 1668089732
transform 1 0 5120 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_2011
timestamp 1668089732
transform 1 0 5120 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_2012
timestamp 1668089732
transform 1 0 5120 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_2013
timestamp 1668089732
transform 1 0 5120 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_2014
timestamp 1668089732
transform 1 0 5120 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_2015
timestamp 1668089732
transform 1 0 5120 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_2016
timestamp 1668089732
transform 1 0 5120 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_2017
timestamp 1668089732
transform 1 0 5120 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_2018
timestamp 1668089732
transform 1 0 5120 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_2019
timestamp 1668089732
transform 1 0 5120 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_2020
timestamp 1668089732
transform 1 0 5120 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_2021
timestamp 1668089732
transform 1 0 5120 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_2022
timestamp 1668089732
transform 1 0 5120 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_2023
timestamp 1668089732
transform 1 0 5120 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_2024
timestamp 1668089732
transform 1 0 5120 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_2025
timestamp 1668089732
transform 1 0 5120 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_2026
timestamp 1668089732
transform 1 0 5120 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_2027
timestamp 1668089732
transform 1 0 5120 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_2028
timestamp 1668089732
transform 1 0 5120 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_2029
timestamp 1668089732
transform 1 0 5120 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_2030
timestamp 1668089732
transform 1 0 5120 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_2031
timestamp 1668089732
transform 1 0 5120 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_2032
timestamp 1668089732
transform 1 0 5120 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_2033
timestamp 1668089732
transform 1 0 5120 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_2034
timestamp 1668089732
transform 1 0 5120 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_2035
timestamp 1668089732
transform 1 0 5120 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_2036
timestamp 1668089732
transform 1 0 5120 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_2037
timestamp 1668089732
transform 1 0 5120 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_2038
timestamp 1668089732
transform 1 0 5120 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_2039
timestamp 1668089732
transform 1 0 5120 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_2040
timestamp 1668089732
transform 1 0 5120 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_2041
timestamp 1668089732
transform 1 0 5120 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_2042
timestamp 1668089732
transform 1 0 5120 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_2043
timestamp 1668089732
transform 1 0 5120 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_2044
timestamp 1668089732
transform 1 0 5120 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_2045
timestamp 1668089732
transform 1 0 5120 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_2046
timestamp 1668089732
transform 1 0 5280 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_2047
timestamp 1668089732
transform 1 0 5280 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_2048
timestamp 1668089732
transform 1 0 5280 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_2049
timestamp 1668089732
transform 1 0 5280 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_2050
timestamp 1668089732
transform 1 0 5280 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_2051
timestamp 1668089732
transform 1 0 5280 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_2052
timestamp 1668089732
transform 1 0 5280 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_2053
timestamp 1668089732
transform 1 0 5280 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_2054
timestamp 1668089732
transform 1 0 5280 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_2055
timestamp 1668089732
transform 1 0 5280 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_2056
timestamp 1668089732
transform 1 0 5280 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_2057
timestamp 1668089732
transform 1 0 5280 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_2058
timestamp 1668089732
transform 1 0 5280 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_2059
timestamp 1668089732
transform 1 0 5280 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_2060
timestamp 1668089732
transform 1 0 5280 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_2061
timestamp 1668089732
transform 1 0 5280 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_2062
timestamp 1668089732
transform 1 0 5280 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_2063
timestamp 1668089732
transform 1 0 5280 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_2064
timestamp 1668089732
transform 1 0 5280 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_2065
timestamp 1668089732
transform 1 0 5280 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_2066
timestamp 1668089732
transform 1 0 5280 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_2067
timestamp 1668089732
transform 1 0 5280 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_2068
timestamp 1668089732
transform 1 0 5280 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_2069
timestamp 1668089732
transform 1 0 5280 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_2070
timestamp 1668089732
transform 1 0 5280 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_2071
timestamp 1668089732
transform 1 0 5280 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_2072
timestamp 1668089732
transform 1 0 5280 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_2073
timestamp 1668089732
transform 1 0 5280 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_2074
timestamp 1668089732
transform 1 0 5280 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_2075
timestamp 1668089732
transform 1 0 5280 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_2076
timestamp 1668089732
transform 1 0 5280 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_2077
timestamp 1668089732
transform 1 0 5280 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_2078
timestamp 1668089732
transform 1 0 5280 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_2079
timestamp 1668089732
transform 1 0 5280 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_2080
timestamp 1668089732
transform 1 0 5280 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_2081
timestamp 1668089732
transform 1 0 5280 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_2082
timestamp 1668089732
transform 1 0 5280 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_2083
timestamp 1668089732
transform 1 0 5280 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_2084
timestamp 1668089732
transform 1 0 5280 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_2085
timestamp 1668089732
transform 1 0 5280 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_2086
timestamp 1668089732
transform 1 0 5280 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_2087
timestamp 1668089732
transform 1 0 5280 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_2088
timestamp 1668089732
transform 1 0 5280 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_2089
timestamp 1668089732
transform 1 0 5280 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_2090
timestamp 1668089732
transform 1 0 5280 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_2091
timestamp 1668089732
transform 1 0 5280 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_2092
timestamp 1668089732
transform 1 0 5280 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_2093
timestamp 1668089732
transform 1 0 5280 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_2094
timestamp 1668089732
transform 1 0 5280 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_2095
timestamp 1668089732
transform 1 0 5280 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_2096
timestamp 1668089732
transform 1 0 5280 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_2097
timestamp 1668089732
transform 1 0 5280 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_2098
timestamp 1668089732
transform 1 0 5280 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_2099
timestamp 1668089732
transform 1 0 5280 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_2100
timestamp 1668089732
transform 1 0 5280 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_2101
timestamp 1668089732
transform 1 0 5280 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_2102
timestamp 1668089732
transform 1 0 5280 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_2103
timestamp 1668089732
transform 1 0 5280 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_2104
timestamp 1668089732
transform 1 0 5280 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_2105
timestamp 1668089732
transform 1 0 5280 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_2106
timestamp 1668089732
transform 1 0 5280 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_2107
timestamp 1668089732
transform 1 0 5280 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_2108
timestamp 1668089732
transform 1 0 5440 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_2109
timestamp 1668089732
transform 1 0 5440 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_2110
timestamp 1668089732
transform 1 0 5440 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_2111
timestamp 1668089732
transform 1 0 5440 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_2112
timestamp 1668089732
transform 1 0 5440 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_2113
timestamp 1668089732
transform 1 0 5440 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_2114
timestamp 1668089732
transform 1 0 5440 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_2115
timestamp 1668089732
transform 1 0 5440 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_2116
timestamp 1668089732
transform 1 0 5440 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_2117
timestamp 1668089732
transform 1 0 5440 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_2118
timestamp 1668089732
transform 1 0 5440 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_2119
timestamp 1668089732
transform 1 0 5440 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_2120
timestamp 1668089732
transform 1 0 5440 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_2121
timestamp 1668089732
transform 1 0 5440 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_2122
timestamp 1668089732
transform 1 0 5440 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_2123
timestamp 1668089732
transform 1 0 5440 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_2124
timestamp 1668089732
transform 1 0 5440 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_2125
timestamp 1668089732
transform 1 0 5440 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_2126
timestamp 1668089732
transform 1 0 5440 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_2127
timestamp 1668089732
transform 1 0 5440 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_2128
timestamp 1668089732
transform 1 0 5440 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_2129
timestamp 1668089732
transform 1 0 5440 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_2130
timestamp 1668089732
transform 1 0 5440 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_2131
timestamp 1668089732
transform 1 0 5440 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_2132
timestamp 1668089732
transform 1 0 5440 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_2133
timestamp 1668089732
transform 1 0 5440 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_2134
timestamp 1668089732
transform 1 0 5440 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_2135
timestamp 1668089732
transform 1 0 5440 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_2136
timestamp 1668089732
transform 1 0 5440 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_2137
timestamp 1668089732
transform 1 0 5440 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_2138
timestamp 1668089732
transform 1 0 5440 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_2139
timestamp 1668089732
transform 1 0 5440 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_2140
timestamp 1668089732
transform 1 0 5440 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_2141
timestamp 1668089732
transform 1 0 5440 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_2142
timestamp 1668089732
transform 1 0 5440 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_2143
timestamp 1668089732
transform 1 0 5440 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_2144
timestamp 1668089732
transform 1 0 5440 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_2145
timestamp 1668089732
transform 1 0 5440 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_2146
timestamp 1668089732
transform 1 0 5440 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_2147
timestamp 1668089732
transform 1 0 5440 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_2148
timestamp 1668089732
transform 1 0 5440 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_2149
timestamp 1668089732
transform 1 0 5440 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_2150
timestamp 1668089732
transform 1 0 5440 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_2151
timestamp 1668089732
transform 1 0 5440 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_2152
timestamp 1668089732
transform 1 0 5440 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_2153
timestamp 1668089732
transform 1 0 5440 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_2154
timestamp 1668089732
transform 1 0 5440 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_2155
timestamp 1668089732
transform 1 0 5440 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_2156
timestamp 1668089732
transform 1 0 5440 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_2157
timestamp 1668089732
transform 1 0 5440 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_2158
timestamp 1668089732
transform 1 0 5440 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_2159
timestamp 1668089732
transform 1 0 5440 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_2160
timestamp 1668089732
transform 1 0 5440 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_2161
timestamp 1668089732
transform 1 0 5440 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_2162
timestamp 1668089732
transform 1 0 5440 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_2163
timestamp 1668089732
transform 1 0 5440 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_2164
timestamp 1668089732
transform 1 0 5440 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_2165
timestamp 1668089732
transform 1 0 5440 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_2166
timestamp 1668089732
transform 1 0 5440 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_2167
timestamp 1668089732
transform 1 0 5440 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_2168
timestamp 1668089732
transform 1 0 5440 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_2169
timestamp 1668089732
transform 1 0 5440 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_2170
timestamp 1668089732
transform 1 0 5600 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_2171
timestamp 1668089732
transform 1 0 5600 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_2172
timestamp 1668089732
transform 1 0 5600 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_2173
timestamp 1668089732
transform 1 0 5600 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_2174
timestamp 1668089732
transform 1 0 5600 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_2175
timestamp 1668089732
transform 1 0 5600 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_2176
timestamp 1668089732
transform 1 0 5600 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_2177
timestamp 1668089732
transform 1 0 5600 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_2178
timestamp 1668089732
transform 1 0 5600 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_2179
timestamp 1668089732
transform 1 0 5600 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_2180
timestamp 1668089732
transform 1 0 5600 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_2181
timestamp 1668089732
transform 1 0 5600 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_2182
timestamp 1668089732
transform 1 0 5600 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_2183
timestamp 1668089732
transform 1 0 5600 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_2184
timestamp 1668089732
transform 1 0 5600 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_2185
timestamp 1668089732
transform 1 0 5600 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_2186
timestamp 1668089732
transform 1 0 5600 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_2187
timestamp 1668089732
transform 1 0 5600 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_2188
timestamp 1668089732
transform 1 0 5600 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_2189
timestamp 1668089732
transform 1 0 5600 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_2190
timestamp 1668089732
transform 1 0 5600 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_2191
timestamp 1668089732
transform 1 0 5600 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_2192
timestamp 1668089732
transform 1 0 5600 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_2193
timestamp 1668089732
transform 1 0 5600 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_2194
timestamp 1668089732
transform 1 0 5600 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_2195
timestamp 1668089732
transform 1 0 5600 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_2196
timestamp 1668089732
transform 1 0 5600 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_2197
timestamp 1668089732
transform 1 0 5600 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_2198
timestamp 1668089732
transform 1 0 5600 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_2199
timestamp 1668089732
transform 1 0 5600 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_2200
timestamp 1668089732
transform 1 0 5600 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_2201
timestamp 1668089732
transform 1 0 5600 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_2202
timestamp 1668089732
transform 1 0 5600 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_2203
timestamp 1668089732
transform 1 0 5600 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_2204
timestamp 1668089732
transform 1 0 5600 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_2205
timestamp 1668089732
transform 1 0 5600 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_2206
timestamp 1668089732
transform 1 0 5600 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_2207
timestamp 1668089732
transform 1 0 5600 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_2208
timestamp 1668089732
transform 1 0 5600 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_2209
timestamp 1668089732
transform 1 0 5600 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_2210
timestamp 1668089732
transform 1 0 5600 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_2211
timestamp 1668089732
transform 1 0 5600 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_2212
timestamp 1668089732
transform 1 0 5600 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_2213
timestamp 1668089732
transform 1 0 5600 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_2214
timestamp 1668089732
transform 1 0 5600 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_2215
timestamp 1668089732
transform 1 0 5600 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_2216
timestamp 1668089732
transform 1 0 5600 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_2217
timestamp 1668089732
transform 1 0 5600 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_2218
timestamp 1668089732
transform 1 0 5600 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_2219
timestamp 1668089732
transform 1 0 5600 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_2220
timestamp 1668089732
transform 1 0 5600 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_2221
timestamp 1668089732
transform 1 0 5600 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_2222
timestamp 1668089732
transform 1 0 5600 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_2223
timestamp 1668089732
transform 1 0 5600 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_2224
timestamp 1668089732
transform 1 0 5600 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_2225
timestamp 1668089732
transform 1 0 5600 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_2226
timestamp 1668089732
transform 1 0 5600 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_2227
timestamp 1668089732
transform 1 0 5600 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_2228
timestamp 1668089732
transform 1 0 5600 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_2229
timestamp 1668089732
transform 1 0 5600 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_2230
timestamp 1668089732
transform 1 0 5600 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_2231
timestamp 1668089732
transform 1 0 5600 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_2232
timestamp 1668089732
transform 1 0 5760 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_2233
timestamp 1668089732
transform 1 0 5760 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_2234
timestamp 1668089732
transform 1 0 5760 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_2235
timestamp 1668089732
transform 1 0 5760 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_2236
timestamp 1668089732
transform 1 0 5760 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_2237
timestamp 1668089732
transform 1 0 5760 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_2238
timestamp 1668089732
transform 1 0 5760 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_2239
timestamp 1668089732
transform 1 0 5760 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_2240
timestamp 1668089732
transform 1 0 5760 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_2241
timestamp 1668089732
transform 1 0 5760 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_2242
timestamp 1668089732
transform 1 0 5760 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_2243
timestamp 1668089732
transform 1 0 5760 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_2244
timestamp 1668089732
transform 1 0 5760 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_2245
timestamp 1668089732
transform 1 0 5760 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_2246
timestamp 1668089732
transform 1 0 5760 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_2247
timestamp 1668089732
transform 1 0 5760 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_2248
timestamp 1668089732
transform 1 0 5760 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_2249
timestamp 1668089732
transform 1 0 5760 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_2250
timestamp 1668089732
transform 1 0 5760 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_2251
timestamp 1668089732
transform 1 0 5760 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_2252
timestamp 1668089732
transform 1 0 5760 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_2253
timestamp 1668089732
transform 1 0 5760 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_2254
timestamp 1668089732
transform 1 0 5760 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_2255
timestamp 1668089732
transform 1 0 5760 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_2256
timestamp 1668089732
transform 1 0 5760 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_2257
timestamp 1668089732
transform 1 0 5760 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_2258
timestamp 1668089732
transform 1 0 5760 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_2259
timestamp 1668089732
transform 1 0 5760 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_2260
timestamp 1668089732
transform 1 0 5760 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_2261
timestamp 1668089732
transform 1 0 5760 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_2262
timestamp 1668089732
transform 1 0 5760 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_2263
timestamp 1668089732
transform 1 0 5760 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_2264
timestamp 1668089732
transform 1 0 5760 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_2265
timestamp 1668089732
transform 1 0 5760 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_2266
timestamp 1668089732
transform 1 0 5760 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_2267
timestamp 1668089732
transform 1 0 5760 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_2268
timestamp 1668089732
transform 1 0 5760 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_2269
timestamp 1668089732
transform 1 0 5760 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_2270
timestamp 1668089732
transform 1 0 5760 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_2271
timestamp 1668089732
transform 1 0 5760 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_2272
timestamp 1668089732
transform 1 0 5760 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_2273
timestamp 1668089732
transform 1 0 5760 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_2274
timestamp 1668089732
transform 1 0 5760 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_2275
timestamp 1668089732
transform 1 0 5760 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_2276
timestamp 1668089732
transform 1 0 5760 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_2277
timestamp 1668089732
transform 1 0 5760 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_2278
timestamp 1668089732
transform 1 0 5760 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_2279
timestamp 1668089732
transform 1 0 5760 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_2280
timestamp 1668089732
transform 1 0 5760 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_2281
timestamp 1668089732
transform 1 0 5760 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_2282
timestamp 1668089732
transform 1 0 5760 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_2283
timestamp 1668089732
transform 1 0 5760 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_2284
timestamp 1668089732
transform 1 0 5760 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_2285
timestamp 1668089732
transform 1 0 5760 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_2286
timestamp 1668089732
transform 1 0 5760 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_2287
timestamp 1668089732
transform 1 0 5760 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_2288
timestamp 1668089732
transform 1 0 5760 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_2289
timestamp 1668089732
transform 1 0 5760 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_2290
timestamp 1668089732
transform 1 0 5760 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_2291
timestamp 1668089732
transform 1 0 5760 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_2292
timestamp 1668089732
transform 1 0 5760 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_2293
timestamp 1668089732
transform 1 0 5760 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_2294
timestamp 1668089732
transform 1 0 5920 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_2295
timestamp 1668089732
transform 1 0 5920 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_2296
timestamp 1668089732
transform 1 0 5920 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_2297
timestamp 1668089732
transform 1 0 5920 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_2298
timestamp 1668089732
transform 1 0 5920 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_2299
timestamp 1668089732
transform 1 0 5920 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_2300
timestamp 1668089732
transform 1 0 5920 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_2301
timestamp 1668089732
transform 1 0 5920 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_2302
timestamp 1668089732
transform 1 0 5920 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_2303
timestamp 1668089732
transform 1 0 5920 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_2304
timestamp 1668089732
transform 1 0 5920 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_2305
timestamp 1668089732
transform 1 0 5920 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_2306
timestamp 1668089732
transform 1 0 5920 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_2307
timestamp 1668089732
transform 1 0 5920 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_2308
timestamp 1668089732
transform 1 0 5920 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_2309
timestamp 1668089732
transform 1 0 5920 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_2310
timestamp 1668089732
transform 1 0 5920 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_2311
timestamp 1668089732
transform 1 0 5920 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_2312
timestamp 1668089732
transform 1 0 5920 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_2313
timestamp 1668089732
transform 1 0 5920 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_2314
timestamp 1668089732
transform 1 0 5920 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_2315
timestamp 1668089732
transform 1 0 5920 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_2316
timestamp 1668089732
transform 1 0 5920 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_2317
timestamp 1668089732
transform 1 0 5920 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_2318
timestamp 1668089732
transform 1 0 5920 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_2319
timestamp 1668089732
transform 1 0 5920 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_2320
timestamp 1668089732
transform 1 0 5920 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_2321
timestamp 1668089732
transform 1 0 5920 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_2322
timestamp 1668089732
transform 1 0 5920 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_2323
timestamp 1668089732
transform 1 0 5920 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_2324
timestamp 1668089732
transform 1 0 5920 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_2325
timestamp 1668089732
transform 1 0 5920 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_2326
timestamp 1668089732
transform 1 0 5920 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_2327
timestamp 1668089732
transform 1 0 5920 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_2328
timestamp 1668089732
transform 1 0 5920 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_2329
timestamp 1668089732
transform 1 0 5920 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_2330
timestamp 1668089732
transform 1 0 5920 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_2331
timestamp 1668089732
transform 1 0 5920 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_2332
timestamp 1668089732
transform 1 0 5920 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_2333
timestamp 1668089732
transform 1 0 5920 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_2334
timestamp 1668089732
transform 1 0 5920 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_2335
timestamp 1668089732
transform 1 0 5920 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_2336
timestamp 1668089732
transform 1 0 5920 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_2337
timestamp 1668089732
transform 1 0 5920 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_2338
timestamp 1668089732
transform 1 0 5920 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_2339
timestamp 1668089732
transform 1 0 5920 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_2340
timestamp 1668089732
transform 1 0 5920 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_2341
timestamp 1668089732
transform 1 0 5920 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_2342
timestamp 1668089732
transform 1 0 5920 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_2343
timestamp 1668089732
transform 1 0 5920 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_2344
timestamp 1668089732
transform 1 0 5920 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_2345
timestamp 1668089732
transform 1 0 5920 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_2346
timestamp 1668089732
transform 1 0 5920 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_2347
timestamp 1668089732
transform 1 0 5920 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_2348
timestamp 1668089732
transform 1 0 5920 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_2349
timestamp 1668089732
transform 1 0 5920 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_2350
timestamp 1668089732
transform 1 0 5920 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_2351
timestamp 1668089732
transform 1 0 5920 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_2352
timestamp 1668089732
transform 1 0 5920 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_2353
timestamp 1668089732
transform 1 0 5920 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_2354
timestamp 1668089732
transform 1 0 5920 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_2355
timestamp 1668089732
transform 1 0 5920 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_2356
timestamp 1668089732
transform 1 0 6080 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_2357
timestamp 1668089732
transform 1 0 6080 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_2358
timestamp 1668089732
transform 1 0 6080 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_2359
timestamp 1668089732
transform 1 0 6080 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_2360
timestamp 1668089732
transform 1 0 6080 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_2361
timestamp 1668089732
transform 1 0 6080 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_2362
timestamp 1668089732
transform 1 0 6080 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_2363
timestamp 1668089732
transform 1 0 6080 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_2364
timestamp 1668089732
transform 1 0 6080 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_2365
timestamp 1668089732
transform 1 0 6080 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_2366
timestamp 1668089732
transform 1 0 6080 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_2367
timestamp 1668089732
transform 1 0 6080 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_2368
timestamp 1668089732
transform 1 0 6080 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_2369
timestamp 1668089732
transform 1 0 6080 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_2370
timestamp 1668089732
transform 1 0 6080 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_2371
timestamp 1668089732
transform 1 0 6080 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_2372
timestamp 1668089732
transform 1 0 6080 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_2373
timestamp 1668089732
transform 1 0 6080 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_2374
timestamp 1668089732
transform 1 0 6080 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_2375
timestamp 1668089732
transform 1 0 6080 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_2376
timestamp 1668089732
transform 1 0 6080 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_2377
timestamp 1668089732
transform 1 0 6080 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_2378
timestamp 1668089732
transform 1 0 6080 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_2379
timestamp 1668089732
transform 1 0 6080 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_2380
timestamp 1668089732
transform 1 0 6080 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_2381
timestamp 1668089732
transform 1 0 6080 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_2382
timestamp 1668089732
transform 1 0 6080 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_2383
timestamp 1668089732
transform 1 0 6080 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_2384
timestamp 1668089732
transform 1 0 6080 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_2385
timestamp 1668089732
transform 1 0 6080 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_2386
timestamp 1668089732
transform 1 0 6080 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_2387
timestamp 1668089732
transform 1 0 6080 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_2388
timestamp 1668089732
transform 1 0 6080 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_2389
timestamp 1668089732
transform 1 0 6080 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_2390
timestamp 1668089732
transform 1 0 6080 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_2391
timestamp 1668089732
transform 1 0 6080 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_2392
timestamp 1668089732
transform 1 0 6080 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_2393
timestamp 1668089732
transform 1 0 6080 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_2394
timestamp 1668089732
transform 1 0 6080 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_2395
timestamp 1668089732
transform 1 0 6080 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_2396
timestamp 1668089732
transform 1 0 6080 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_2397
timestamp 1668089732
transform 1 0 6080 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_2398
timestamp 1668089732
transform 1 0 6080 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_2399
timestamp 1668089732
transform 1 0 6080 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_2400
timestamp 1668089732
transform 1 0 6080 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_2401
timestamp 1668089732
transform 1 0 6080 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_2402
timestamp 1668089732
transform 1 0 6080 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_2403
timestamp 1668089732
transform 1 0 6080 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_2404
timestamp 1668089732
transform 1 0 6080 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_2405
timestamp 1668089732
transform 1 0 6080 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_2406
timestamp 1668089732
transform 1 0 6080 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_2407
timestamp 1668089732
transform 1 0 6080 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_2408
timestamp 1668089732
transform 1 0 6080 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_2409
timestamp 1668089732
transform 1 0 6080 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_2410
timestamp 1668089732
transform 1 0 6080 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_2411
timestamp 1668089732
transform 1 0 6080 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_2412
timestamp 1668089732
transform 1 0 6080 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_2413
timestamp 1668089732
transform 1 0 6080 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_2414
timestamp 1668089732
transform 1 0 6080 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_2415
timestamp 1668089732
transform 1 0 6080 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_2416
timestamp 1668089732
transform 1 0 6080 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_2417
timestamp 1668089732
transform 1 0 6080 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_2418
timestamp 1668089732
transform 1 0 6240 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_2419
timestamp 1668089732
transform 1 0 6240 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_2420
timestamp 1668089732
transform 1 0 6240 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_2421
timestamp 1668089732
transform 1 0 6240 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_2422
timestamp 1668089732
transform 1 0 6240 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_2423
timestamp 1668089732
transform 1 0 6240 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_2424
timestamp 1668089732
transform 1 0 6240 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_2425
timestamp 1668089732
transform 1 0 6240 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_2426
timestamp 1668089732
transform 1 0 6240 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_2427
timestamp 1668089732
transform 1 0 6240 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_2428
timestamp 1668089732
transform 1 0 6240 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_2429
timestamp 1668089732
transform 1 0 6240 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_2430
timestamp 1668089732
transform 1 0 6240 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_2431
timestamp 1668089732
transform 1 0 6240 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_2432
timestamp 1668089732
transform 1 0 6240 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_2433
timestamp 1668089732
transform 1 0 6240 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_2434
timestamp 1668089732
transform 1 0 6240 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_2435
timestamp 1668089732
transform 1 0 6240 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_2436
timestamp 1668089732
transform 1 0 6240 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_2437
timestamp 1668089732
transform 1 0 6240 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_2438
timestamp 1668089732
transform 1 0 6240 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_2439
timestamp 1668089732
transform 1 0 6240 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_2440
timestamp 1668089732
transform 1 0 6240 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_2441
timestamp 1668089732
transform 1 0 6240 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_2442
timestamp 1668089732
transform 1 0 6240 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_2443
timestamp 1668089732
transform 1 0 6240 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_2444
timestamp 1668089732
transform 1 0 6240 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_2445
timestamp 1668089732
transform 1 0 6240 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_2446
timestamp 1668089732
transform 1 0 6240 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_2447
timestamp 1668089732
transform 1 0 6240 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_2448
timestamp 1668089732
transform 1 0 6240 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_2449
timestamp 1668089732
transform 1 0 6240 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_2450
timestamp 1668089732
transform 1 0 6240 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_2451
timestamp 1668089732
transform 1 0 6240 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_2452
timestamp 1668089732
transform 1 0 6240 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_2453
timestamp 1668089732
transform 1 0 6240 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_2454
timestamp 1668089732
transform 1 0 6240 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_2455
timestamp 1668089732
transform 1 0 6240 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_2456
timestamp 1668089732
transform 1 0 6240 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_2457
timestamp 1668089732
transform 1 0 6240 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_2458
timestamp 1668089732
transform 1 0 6240 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_2459
timestamp 1668089732
transform 1 0 6240 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_2460
timestamp 1668089732
transform 1 0 6240 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_2461
timestamp 1668089732
transform 1 0 6240 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_2462
timestamp 1668089732
transform 1 0 6240 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_2463
timestamp 1668089732
transform 1 0 6240 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_2464
timestamp 1668089732
transform 1 0 6240 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_2465
timestamp 1668089732
transform 1 0 6240 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_2466
timestamp 1668089732
transform 1 0 6240 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_2467
timestamp 1668089732
transform 1 0 6240 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_2468
timestamp 1668089732
transform 1 0 6240 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_2469
timestamp 1668089732
transform 1 0 6240 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_2470
timestamp 1668089732
transform 1 0 6240 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_2471
timestamp 1668089732
transform 1 0 6240 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_2472
timestamp 1668089732
transform 1 0 6240 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_2473
timestamp 1668089732
transform 1 0 6240 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_2474
timestamp 1668089732
transform 1 0 6240 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_2475
timestamp 1668089732
transform 1 0 6240 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_2476
timestamp 1668089732
transform 1 0 6240 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_2477
timestamp 1668089732
transform 1 0 6240 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_2478
timestamp 1668089732
transform 1 0 6240 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_2479
timestamp 1668089732
transform 1 0 6240 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_2480
timestamp 1668089732
transform 1 0 6400 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_2481
timestamp 1668089732
transform 1 0 6400 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_2482
timestamp 1668089732
transform 1 0 6400 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_2483
timestamp 1668089732
transform 1 0 6400 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_2484
timestamp 1668089732
transform 1 0 6400 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_2485
timestamp 1668089732
transform 1 0 6400 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_2486
timestamp 1668089732
transform 1 0 6400 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_2487
timestamp 1668089732
transform 1 0 6400 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_2488
timestamp 1668089732
transform 1 0 6400 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_2489
timestamp 1668089732
transform 1 0 6400 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_2490
timestamp 1668089732
transform 1 0 6400 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_2491
timestamp 1668089732
transform 1 0 6400 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_2492
timestamp 1668089732
transform 1 0 6400 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_2493
timestamp 1668089732
transform 1 0 6400 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_2494
timestamp 1668089732
transform 1 0 6400 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_2495
timestamp 1668089732
transform 1 0 6400 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_2496
timestamp 1668089732
transform 1 0 6400 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_2497
timestamp 1668089732
transform 1 0 6400 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_2498
timestamp 1668089732
transform 1 0 6400 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_2499
timestamp 1668089732
transform 1 0 6400 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_2500
timestamp 1668089732
transform 1 0 6400 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_2501
timestamp 1668089732
transform 1 0 6400 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_2502
timestamp 1668089732
transform 1 0 6400 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_2503
timestamp 1668089732
transform 1 0 6400 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_2504
timestamp 1668089732
transform 1 0 6400 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_2505
timestamp 1668089732
transform 1 0 6400 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_2506
timestamp 1668089732
transform 1 0 6400 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_2507
timestamp 1668089732
transform 1 0 6400 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_2508
timestamp 1668089732
transform 1 0 6400 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_2509
timestamp 1668089732
transform 1 0 6400 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_2510
timestamp 1668089732
transform 1 0 6400 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_2511
timestamp 1668089732
transform 1 0 6400 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_2512
timestamp 1668089732
transform 1 0 6400 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_2513
timestamp 1668089732
transform 1 0 6400 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_2514
timestamp 1668089732
transform 1 0 6400 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_2515
timestamp 1668089732
transform 1 0 6400 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_2516
timestamp 1668089732
transform 1 0 6400 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_2517
timestamp 1668089732
transform 1 0 6400 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_2518
timestamp 1668089732
transform 1 0 6400 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_2519
timestamp 1668089732
transform 1 0 6400 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_2520
timestamp 1668089732
transform 1 0 6400 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_2521
timestamp 1668089732
transform 1 0 6400 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_2522
timestamp 1668089732
transform 1 0 6400 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_2523
timestamp 1668089732
transform 1 0 6400 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_2524
timestamp 1668089732
transform 1 0 6400 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_2525
timestamp 1668089732
transform 1 0 6400 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_2526
timestamp 1668089732
transform 1 0 6400 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_2527
timestamp 1668089732
transform 1 0 6400 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_2528
timestamp 1668089732
transform 1 0 6400 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_2529
timestamp 1668089732
transform 1 0 6400 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_2530
timestamp 1668089732
transform 1 0 6400 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_2531
timestamp 1668089732
transform 1 0 6400 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_2532
timestamp 1668089732
transform 1 0 6400 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_2533
timestamp 1668089732
transform 1 0 6400 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_2534
timestamp 1668089732
transform 1 0 6400 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_2535
timestamp 1668089732
transform 1 0 6400 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_2536
timestamp 1668089732
transform 1 0 6400 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_2537
timestamp 1668089732
transform 1 0 6400 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_2538
timestamp 1668089732
transform 1 0 6400 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_2539
timestamp 1668089732
transform 1 0 6400 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_2540
timestamp 1668089732
transform 1 0 6400 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_2541
timestamp 1668089732
transform 1 0 6400 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_2542
timestamp 1668089732
transform 1 0 6560 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_2543
timestamp 1668089732
transform 1 0 6560 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_2544
timestamp 1668089732
transform 1 0 6560 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_2545
timestamp 1668089732
transform 1 0 6560 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_2546
timestamp 1668089732
transform 1 0 6560 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_2547
timestamp 1668089732
transform 1 0 6560 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_2548
timestamp 1668089732
transform 1 0 6560 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_2549
timestamp 1668089732
transform 1 0 6560 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_2550
timestamp 1668089732
transform 1 0 6560 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_2551
timestamp 1668089732
transform 1 0 6560 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_2552
timestamp 1668089732
transform 1 0 6560 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_2553
timestamp 1668089732
transform 1 0 6560 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_2554
timestamp 1668089732
transform 1 0 6560 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_2555
timestamp 1668089732
transform 1 0 6560 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_2556
timestamp 1668089732
transform 1 0 6560 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_2557
timestamp 1668089732
transform 1 0 6560 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_2558
timestamp 1668089732
transform 1 0 6560 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_2559
timestamp 1668089732
transform 1 0 6560 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_2560
timestamp 1668089732
transform 1 0 6560 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_2561
timestamp 1668089732
transform 1 0 6560 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_2562
timestamp 1668089732
transform 1 0 6560 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_2563
timestamp 1668089732
transform 1 0 6560 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_2564
timestamp 1668089732
transform 1 0 6560 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_2565
timestamp 1668089732
transform 1 0 6560 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_2566
timestamp 1668089732
transform 1 0 6560 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_2567
timestamp 1668089732
transform 1 0 6560 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_2568
timestamp 1668089732
transform 1 0 6560 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_2569
timestamp 1668089732
transform 1 0 6560 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_2570
timestamp 1668089732
transform 1 0 6560 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_2571
timestamp 1668089732
transform 1 0 6560 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_2572
timestamp 1668089732
transform 1 0 6560 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_2573
timestamp 1668089732
transform 1 0 6560 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_2574
timestamp 1668089732
transform 1 0 6560 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_2575
timestamp 1668089732
transform 1 0 6560 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_2576
timestamp 1668089732
transform 1 0 6560 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_2577
timestamp 1668089732
transform 1 0 6560 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_2578
timestamp 1668089732
transform 1 0 6560 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_2579
timestamp 1668089732
transform 1 0 6560 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_2580
timestamp 1668089732
transform 1 0 6560 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_2581
timestamp 1668089732
transform 1 0 6560 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_2582
timestamp 1668089732
transform 1 0 6560 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_2583
timestamp 1668089732
transform 1 0 6560 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_2584
timestamp 1668089732
transform 1 0 6560 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_2585
timestamp 1668089732
transform 1 0 6560 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_2586
timestamp 1668089732
transform 1 0 6560 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_2587
timestamp 1668089732
transform 1 0 6560 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_2588
timestamp 1668089732
transform 1 0 6560 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_2589
timestamp 1668089732
transform 1 0 6560 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_2590
timestamp 1668089732
transform 1 0 6560 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_2591
timestamp 1668089732
transform 1 0 6560 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_2592
timestamp 1668089732
transform 1 0 6560 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_2593
timestamp 1668089732
transform 1 0 6560 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_2594
timestamp 1668089732
transform 1 0 6560 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_2595
timestamp 1668089732
transform 1 0 6560 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_2596
timestamp 1668089732
transform 1 0 6560 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_2597
timestamp 1668089732
transform 1 0 6560 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_2598
timestamp 1668089732
transform 1 0 6560 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_2599
timestamp 1668089732
transform 1 0 6560 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_2600
timestamp 1668089732
transform 1 0 6560 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_2601
timestamp 1668089732
transform 1 0 6560 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_2602
timestamp 1668089732
transform 1 0 6560 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_2603
timestamp 1668089732
transform 1 0 6560 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_2604
timestamp 1668089732
transform 1 0 6720 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_2605
timestamp 1668089732
transform 1 0 6720 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_2606
timestamp 1668089732
transform 1 0 6720 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_2607
timestamp 1668089732
transform 1 0 6720 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_2608
timestamp 1668089732
transform 1 0 6720 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_2609
timestamp 1668089732
transform 1 0 6720 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_2610
timestamp 1668089732
transform 1 0 6720 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_2611
timestamp 1668089732
transform 1 0 6720 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_2612
timestamp 1668089732
transform 1 0 6720 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_2613
timestamp 1668089732
transform 1 0 6720 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_2614
timestamp 1668089732
transform 1 0 6720 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_2615
timestamp 1668089732
transform 1 0 6720 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_2616
timestamp 1668089732
transform 1 0 6720 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_2617
timestamp 1668089732
transform 1 0 6720 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_2618
timestamp 1668089732
transform 1 0 6720 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_2619
timestamp 1668089732
transform 1 0 6720 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_2620
timestamp 1668089732
transform 1 0 6720 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_2621
timestamp 1668089732
transform 1 0 6720 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_2622
timestamp 1668089732
transform 1 0 6720 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_2623
timestamp 1668089732
transform 1 0 6720 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_2624
timestamp 1668089732
transform 1 0 6720 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_2625
timestamp 1668089732
transform 1 0 6720 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_2626
timestamp 1668089732
transform 1 0 6720 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_2627
timestamp 1668089732
transform 1 0 6720 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_2628
timestamp 1668089732
transform 1 0 6720 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_2629
timestamp 1668089732
transform 1 0 6720 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_2630
timestamp 1668089732
transform 1 0 6720 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_2631
timestamp 1668089732
transform 1 0 6720 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_2632
timestamp 1668089732
transform 1 0 6720 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_2633
timestamp 1668089732
transform 1 0 6720 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_2634
timestamp 1668089732
transform 1 0 6720 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_2635
timestamp 1668089732
transform 1 0 6720 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_2636
timestamp 1668089732
transform 1 0 6720 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_2637
timestamp 1668089732
transform 1 0 6720 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_2638
timestamp 1668089732
transform 1 0 6720 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_2639
timestamp 1668089732
transform 1 0 6720 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_2640
timestamp 1668089732
transform 1 0 6720 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_2641
timestamp 1668089732
transform 1 0 6720 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_2642
timestamp 1668089732
transform 1 0 6720 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_2643
timestamp 1668089732
transform 1 0 6720 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_2644
timestamp 1668089732
transform 1 0 6720 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_2645
timestamp 1668089732
transform 1 0 6720 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_2646
timestamp 1668089732
transform 1 0 6720 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_2647
timestamp 1668089732
transform 1 0 6720 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_2648
timestamp 1668089732
transform 1 0 6720 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_2649
timestamp 1668089732
transform 1 0 6720 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_2650
timestamp 1668089732
transform 1 0 6720 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_2651
timestamp 1668089732
transform 1 0 6720 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_2652
timestamp 1668089732
transform 1 0 6720 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_2653
timestamp 1668089732
transform 1 0 6720 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_2654
timestamp 1668089732
transform 1 0 6720 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_2655
timestamp 1668089732
transform 1 0 6720 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_2656
timestamp 1668089732
transform 1 0 6720 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_2657
timestamp 1668089732
transform 1 0 6720 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_2658
timestamp 1668089732
transform 1 0 6720 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_2659
timestamp 1668089732
transform 1 0 6720 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_2660
timestamp 1668089732
transform 1 0 6720 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_2661
timestamp 1668089732
transform 1 0 6720 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_2662
timestamp 1668089732
transform 1 0 6720 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_2663
timestamp 1668089732
transform 1 0 6720 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_2664
timestamp 1668089732
transform 1 0 6720 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_2665
timestamp 1668089732
transform 1 0 6720 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_2666
timestamp 1668089732
transform 1 0 6880 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_2667
timestamp 1668089732
transform 1 0 6880 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_2668
timestamp 1668089732
transform 1 0 6880 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_2669
timestamp 1668089732
transform 1 0 6880 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_2670
timestamp 1668089732
transform 1 0 6880 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_2671
timestamp 1668089732
transform 1 0 6880 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_2672
timestamp 1668089732
transform 1 0 6880 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_2673
timestamp 1668089732
transform 1 0 6880 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_2674
timestamp 1668089732
transform 1 0 6880 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_2675
timestamp 1668089732
transform 1 0 6880 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_2676
timestamp 1668089732
transform 1 0 6880 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_2677
timestamp 1668089732
transform 1 0 6880 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_2678
timestamp 1668089732
transform 1 0 6880 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_2679
timestamp 1668089732
transform 1 0 6880 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_2680
timestamp 1668089732
transform 1 0 6880 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_2681
timestamp 1668089732
transform 1 0 6880 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_2682
timestamp 1668089732
transform 1 0 6880 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_2683
timestamp 1668089732
transform 1 0 6880 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_2684
timestamp 1668089732
transform 1 0 6880 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_2685
timestamp 1668089732
transform 1 0 6880 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_2686
timestamp 1668089732
transform 1 0 6880 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_2687
timestamp 1668089732
transform 1 0 6880 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_2688
timestamp 1668089732
transform 1 0 6880 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_2689
timestamp 1668089732
transform 1 0 6880 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_2690
timestamp 1668089732
transform 1 0 6880 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_2691
timestamp 1668089732
transform 1 0 6880 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_2692
timestamp 1668089732
transform 1 0 6880 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_2693
timestamp 1668089732
transform 1 0 6880 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_2694
timestamp 1668089732
transform 1 0 6880 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_2695
timestamp 1668089732
transform 1 0 6880 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_2696
timestamp 1668089732
transform 1 0 6880 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_2697
timestamp 1668089732
transform 1 0 6880 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_2698
timestamp 1668089732
transform 1 0 6880 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_2699
timestamp 1668089732
transform 1 0 6880 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_2700
timestamp 1668089732
transform 1 0 6880 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_2701
timestamp 1668089732
transform 1 0 6880 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_2702
timestamp 1668089732
transform 1 0 6880 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_2703
timestamp 1668089732
transform 1 0 6880 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_2704
timestamp 1668089732
transform 1 0 6880 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_2705
timestamp 1668089732
transform 1 0 6880 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_2706
timestamp 1668089732
transform 1 0 6880 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_2707
timestamp 1668089732
transform 1 0 6880 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_2708
timestamp 1668089732
transform 1 0 6880 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_2709
timestamp 1668089732
transform 1 0 6880 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_2710
timestamp 1668089732
transform 1 0 6880 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_2711
timestamp 1668089732
transform 1 0 6880 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_2712
timestamp 1668089732
transform 1 0 6880 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_2713
timestamp 1668089732
transform 1 0 6880 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_2714
timestamp 1668089732
transform 1 0 6880 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_2715
timestamp 1668089732
transform 1 0 6880 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_2716
timestamp 1668089732
transform 1 0 6880 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_2717
timestamp 1668089732
transform 1 0 6880 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_2718
timestamp 1668089732
transform 1 0 6880 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_2719
timestamp 1668089732
transform 1 0 6880 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_2720
timestamp 1668089732
transform 1 0 6880 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_2721
timestamp 1668089732
transform 1 0 6880 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_2722
timestamp 1668089732
transform 1 0 6880 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_2723
timestamp 1668089732
transform 1 0 6880 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_2724
timestamp 1668089732
transform 1 0 6880 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_2725
timestamp 1668089732
transform 1 0 6880 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_2726
timestamp 1668089732
transform 1 0 6880 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_2727
timestamp 1668089732
transform 1 0 6880 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_2728
timestamp 1668089732
transform 1 0 7040 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_2729
timestamp 1668089732
transform 1 0 7040 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_2730
timestamp 1668089732
transform 1 0 7040 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_2731
timestamp 1668089732
transform 1 0 7040 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_2732
timestamp 1668089732
transform 1 0 7040 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_2733
timestamp 1668089732
transform 1 0 7040 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_2734
timestamp 1668089732
transform 1 0 7040 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_2735
timestamp 1668089732
transform 1 0 7040 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_2736
timestamp 1668089732
transform 1 0 7040 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_2737
timestamp 1668089732
transform 1 0 7040 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_2738
timestamp 1668089732
transform 1 0 7040 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_2739
timestamp 1668089732
transform 1 0 7040 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_2740
timestamp 1668089732
transform 1 0 7040 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_2741
timestamp 1668089732
transform 1 0 7040 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_2742
timestamp 1668089732
transform 1 0 7040 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_2743
timestamp 1668089732
transform 1 0 7040 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_2744
timestamp 1668089732
transform 1 0 7040 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_2745
timestamp 1668089732
transform 1 0 7040 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_2746
timestamp 1668089732
transform 1 0 7040 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_2747
timestamp 1668089732
transform 1 0 7040 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_2748
timestamp 1668089732
transform 1 0 7040 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_2749
timestamp 1668089732
transform 1 0 7040 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_2750
timestamp 1668089732
transform 1 0 7040 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_2751
timestamp 1668089732
transform 1 0 7040 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_2752
timestamp 1668089732
transform 1 0 7040 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_2753
timestamp 1668089732
transform 1 0 7040 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_2754
timestamp 1668089732
transform 1 0 7040 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_2755
timestamp 1668089732
transform 1 0 7040 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_2756
timestamp 1668089732
transform 1 0 7040 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_2757
timestamp 1668089732
transform 1 0 7040 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_2758
timestamp 1668089732
transform 1 0 7040 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_2759
timestamp 1668089732
transform 1 0 7040 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_2760
timestamp 1668089732
transform 1 0 7040 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_2761
timestamp 1668089732
transform 1 0 7040 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_2762
timestamp 1668089732
transform 1 0 7040 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_2763
timestamp 1668089732
transform 1 0 7040 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_2764
timestamp 1668089732
transform 1 0 7040 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_2765
timestamp 1668089732
transform 1 0 7040 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_2766
timestamp 1668089732
transform 1 0 7040 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_2767
timestamp 1668089732
transform 1 0 7040 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_2768
timestamp 1668089732
transform 1 0 7040 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_2769
timestamp 1668089732
transform 1 0 7040 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_2770
timestamp 1668089732
transform 1 0 7040 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_2771
timestamp 1668089732
transform 1 0 7040 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_2772
timestamp 1668089732
transform 1 0 7040 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_2773
timestamp 1668089732
transform 1 0 7040 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_2774
timestamp 1668089732
transform 1 0 7040 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_2775
timestamp 1668089732
transform 1 0 7040 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_2776
timestamp 1668089732
transform 1 0 7040 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_2777
timestamp 1668089732
transform 1 0 7040 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_2778
timestamp 1668089732
transform 1 0 7040 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_2779
timestamp 1668089732
transform 1 0 7040 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_2780
timestamp 1668089732
transform 1 0 7040 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_2781
timestamp 1668089732
transform 1 0 7040 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_2782
timestamp 1668089732
transform 1 0 7040 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_2783
timestamp 1668089732
transform 1 0 7040 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_2784
timestamp 1668089732
transform 1 0 7040 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_2785
timestamp 1668089732
transform 1 0 7040 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_2786
timestamp 1668089732
transform 1 0 7040 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_2787
timestamp 1668089732
transform 1 0 7040 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_2788
timestamp 1668089732
transform 1 0 7040 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_2789
timestamp 1668089732
transform 1 0 7040 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_2790
timestamp 1668089732
transform 1 0 7200 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_2791
timestamp 1668089732
transform 1 0 7200 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_2792
timestamp 1668089732
transform 1 0 7200 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_2793
timestamp 1668089732
transform 1 0 7200 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_2794
timestamp 1668089732
transform 1 0 7200 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_2795
timestamp 1668089732
transform 1 0 7200 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_2796
timestamp 1668089732
transform 1 0 7200 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_2797
timestamp 1668089732
transform 1 0 7200 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_2798
timestamp 1668089732
transform 1 0 7200 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_2799
timestamp 1668089732
transform 1 0 7200 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_2800
timestamp 1668089732
transform 1 0 7200 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_2801
timestamp 1668089732
transform 1 0 7200 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_2802
timestamp 1668089732
transform 1 0 7200 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_2803
timestamp 1668089732
transform 1 0 7200 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_2804
timestamp 1668089732
transform 1 0 7200 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_2805
timestamp 1668089732
transform 1 0 7200 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_2806
timestamp 1668089732
transform 1 0 7200 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_2807
timestamp 1668089732
transform 1 0 7200 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_2808
timestamp 1668089732
transform 1 0 7200 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_2809
timestamp 1668089732
transform 1 0 7200 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_2810
timestamp 1668089732
transform 1 0 7200 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_2811
timestamp 1668089732
transform 1 0 7200 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_2812
timestamp 1668089732
transform 1 0 7200 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_2813
timestamp 1668089732
transform 1 0 7200 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_2814
timestamp 1668089732
transform 1 0 7200 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_2815
timestamp 1668089732
transform 1 0 7200 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_2816
timestamp 1668089732
transform 1 0 7200 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_2817
timestamp 1668089732
transform 1 0 7200 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_2818
timestamp 1668089732
transform 1 0 7200 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_2819
timestamp 1668089732
transform 1 0 7200 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_2820
timestamp 1668089732
transform 1 0 7200 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_2821
timestamp 1668089732
transform 1 0 7200 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_2822
timestamp 1668089732
transform 1 0 7200 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_2823
timestamp 1668089732
transform 1 0 7200 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_2824
timestamp 1668089732
transform 1 0 7200 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_2825
timestamp 1668089732
transform 1 0 7200 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_2826
timestamp 1668089732
transform 1 0 7200 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_2827
timestamp 1668089732
transform 1 0 7200 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_2828
timestamp 1668089732
transform 1 0 7200 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_2829
timestamp 1668089732
transform 1 0 7200 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_2830
timestamp 1668089732
transform 1 0 7200 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_2831
timestamp 1668089732
transform 1 0 7200 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_2832
timestamp 1668089732
transform 1 0 7200 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_2833
timestamp 1668089732
transform 1 0 7200 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_2834
timestamp 1668089732
transform 1 0 7200 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_2835
timestamp 1668089732
transform 1 0 7200 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_2836
timestamp 1668089732
transform 1 0 7200 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_2837
timestamp 1668089732
transform 1 0 7200 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_2838
timestamp 1668089732
transform 1 0 7200 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_2839
timestamp 1668089732
transform 1 0 7200 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_2840
timestamp 1668089732
transform 1 0 7200 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_2841
timestamp 1668089732
transform 1 0 7200 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_2842
timestamp 1668089732
transform 1 0 7200 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_2843
timestamp 1668089732
transform 1 0 7200 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_2844
timestamp 1668089732
transform 1 0 7200 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_2845
timestamp 1668089732
transform 1 0 7200 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_2846
timestamp 1668089732
transform 1 0 7200 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_2847
timestamp 1668089732
transform 1 0 7200 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_2848
timestamp 1668089732
transform 1 0 7200 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_2849
timestamp 1668089732
transform 1 0 7200 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_2850
timestamp 1668089732
transform 1 0 7200 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_2851
timestamp 1668089732
transform 1 0 7200 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_2852
timestamp 1668089732
transform 1 0 7360 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_2853
timestamp 1668089732
transform 1 0 7360 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_2854
timestamp 1668089732
transform 1 0 7360 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_2855
timestamp 1668089732
transform 1 0 7360 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_2856
timestamp 1668089732
transform 1 0 7360 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_2857
timestamp 1668089732
transform 1 0 7360 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_2858
timestamp 1668089732
transform 1 0 7360 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_2859
timestamp 1668089732
transform 1 0 7360 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_2860
timestamp 1668089732
transform 1 0 7360 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_2861
timestamp 1668089732
transform 1 0 7360 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_2862
timestamp 1668089732
transform 1 0 7360 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_2863
timestamp 1668089732
transform 1 0 7360 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_2864
timestamp 1668089732
transform 1 0 7360 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_2865
timestamp 1668089732
transform 1 0 7360 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_2866
timestamp 1668089732
transform 1 0 7360 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_2867
timestamp 1668089732
transform 1 0 7360 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_2868
timestamp 1668089732
transform 1 0 7360 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_2869
timestamp 1668089732
transform 1 0 7360 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_2870
timestamp 1668089732
transform 1 0 7360 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_2871
timestamp 1668089732
transform 1 0 7360 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_2872
timestamp 1668089732
transform 1 0 7360 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_2873
timestamp 1668089732
transform 1 0 7360 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_2874
timestamp 1668089732
transform 1 0 7360 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_2875
timestamp 1668089732
transform 1 0 7360 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_2876
timestamp 1668089732
transform 1 0 7360 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_2877
timestamp 1668089732
transform 1 0 7360 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_2878
timestamp 1668089732
transform 1 0 7360 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_2879
timestamp 1668089732
transform 1 0 7360 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_2880
timestamp 1668089732
transform 1 0 7360 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_2881
timestamp 1668089732
transform 1 0 7360 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_2882
timestamp 1668089732
transform 1 0 7360 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_2883
timestamp 1668089732
transform 1 0 7360 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_2884
timestamp 1668089732
transform 1 0 7360 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_2885
timestamp 1668089732
transform 1 0 7360 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_2886
timestamp 1668089732
transform 1 0 7360 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_2887
timestamp 1668089732
transform 1 0 7360 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_2888
timestamp 1668089732
transform 1 0 7360 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_2889
timestamp 1668089732
transform 1 0 7360 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_2890
timestamp 1668089732
transform 1 0 7360 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_2891
timestamp 1668089732
transform 1 0 7360 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_2892
timestamp 1668089732
transform 1 0 7360 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_2893
timestamp 1668089732
transform 1 0 7360 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_2894
timestamp 1668089732
transform 1 0 7360 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_2895
timestamp 1668089732
transform 1 0 7360 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_2896
timestamp 1668089732
transform 1 0 7360 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_2897
timestamp 1668089732
transform 1 0 7360 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_2898
timestamp 1668089732
transform 1 0 7360 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_2899
timestamp 1668089732
transform 1 0 7360 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_2900
timestamp 1668089732
transform 1 0 7360 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_2901
timestamp 1668089732
transform 1 0 7360 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_2902
timestamp 1668089732
transform 1 0 7360 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_2903
timestamp 1668089732
transform 1 0 7360 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_2904
timestamp 1668089732
transform 1 0 7360 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_2905
timestamp 1668089732
transform 1 0 7360 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_2906
timestamp 1668089732
transform 1 0 7360 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_2907
timestamp 1668089732
transform 1 0 7360 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_2908
timestamp 1668089732
transform 1 0 7360 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_2909
timestamp 1668089732
transform 1 0 7360 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_2910
timestamp 1668089732
transform 1 0 7360 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_2911
timestamp 1668089732
transform 1 0 7360 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_2912
timestamp 1668089732
transform 1 0 7360 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_2913
timestamp 1668089732
transform 1 0 7360 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_2914
timestamp 1668089732
transform 1 0 7520 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_2915
timestamp 1668089732
transform 1 0 7520 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_2916
timestamp 1668089732
transform 1 0 7520 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_2917
timestamp 1668089732
transform 1 0 7520 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_2918
timestamp 1668089732
transform 1 0 7520 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_2919
timestamp 1668089732
transform 1 0 7520 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_2920
timestamp 1668089732
transform 1 0 7520 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_2921
timestamp 1668089732
transform 1 0 7520 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_2922
timestamp 1668089732
transform 1 0 7520 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_2923
timestamp 1668089732
transform 1 0 7520 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_2924
timestamp 1668089732
transform 1 0 7520 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_2925
timestamp 1668089732
transform 1 0 7520 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_2926
timestamp 1668089732
transform 1 0 7520 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_2927
timestamp 1668089732
transform 1 0 7520 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_2928
timestamp 1668089732
transform 1 0 7520 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_2929
timestamp 1668089732
transform 1 0 7520 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_2930
timestamp 1668089732
transform 1 0 7520 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_2931
timestamp 1668089732
transform 1 0 7520 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_2932
timestamp 1668089732
transform 1 0 7520 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_2933
timestamp 1668089732
transform 1 0 7520 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_2934
timestamp 1668089732
transform 1 0 7520 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_2935
timestamp 1668089732
transform 1 0 7520 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_2936
timestamp 1668089732
transform 1 0 7520 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_2937
timestamp 1668089732
transform 1 0 7520 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_2938
timestamp 1668089732
transform 1 0 7520 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_2939
timestamp 1668089732
transform 1 0 7520 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_2940
timestamp 1668089732
transform 1 0 7520 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_2941
timestamp 1668089732
transform 1 0 7520 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_2942
timestamp 1668089732
transform 1 0 7520 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_2943
timestamp 1668089732
transform 1 0 7520 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_2944
timestamp 1668089732
transform 1 0 7520 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_2945
timestamp 1668089732
transform 1 0 7520 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_2946
timestamp 1668089732
transform 1 0 7520 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_2947
timestamp 1668089732
transform 1 0 7520 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_2948
timestamp 1668089732
transform 1 0 7520 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_2949
timestamp 1668089732
transform 1 0 7520 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_2950
timestamp 1668089732
transform 1 0 7520 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_2951
timestamp 1668089732
transform 1 0 7520 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_2952
timestamp 1668089732
transform 1 0 7520 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_2953
timestamp 1668089732
transform 1 0 7520 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_2954
timestamp 1668089732
transform 1 0 7520 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_2955
timestamp 1668089732
transform 1 0 7520 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_2956
timestamp 1668089732
transform 1 0 7520 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_2957
timestamp 1668089732
transform 1 0 7520 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_2958
timestamp 1668089732
transform 1 0 7520 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_2959
timestamp 1668089732
transform 1 0 7520 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_2960
timestamp 1668089732
transform 1 0 7520 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_2961
timestamp 1668089732
transform 1 0 7520 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_2962
timestamp 1668089732
transform 1 0 7520 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_2963
timestamp 1668089732
transform 1 0 7520 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_2964
timestamp 1668089732
transform 1 0 7520 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_2965
timestamp 1668089732
transform 1 0 7520 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_2966
timestamp 1668089732
transform 1 0 7520 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_2967
timestamp 1668089732
transform 1 0 7520 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_2968
timestamp 1668089732
transform 1 0 7520 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_2969
timestamp 1668089732
transform 1 0 7520 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_2970
timestamp 1668089732
transform 1 0 7520 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_2971
timestamp 1668089732
transform 1 0 7520 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_2972
timestamp 1668089732
transform 1 0 7520 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_2973
timestamp 1668089732
transform 1 0 7520 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_2974
timestamp 1668089732
transform 1 0 7520 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_2975
timestamp 1668089732
transform 1 0 7520 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_2976
timestamp 1668089732
transform 1 0 7680 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_2977
timestamp 1668089732
transform 1 0 7680 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_2978
timestamp 1668089732
transform 1 0 7680 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_2979
timestamp 1668089732
transform 1 0 7680 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_2980
timestamp 1668089732
transform 1 0 7680 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_2981
timestamp 1668089732
transform 1 0 7680 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_2982
timestamp 1668089732
transform 1 0 7680 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_2983
timestamp 1668089732
transform 1 0 7680 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_2984
timestamp 1668089732
transform 1 0 7680 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_2985
timestamp 1668089732
transform 1 0 7680 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_2986
timestamp 1668089732
transform 1 0 7680 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_2987
timestamp 1668089732
transform 1 0 7680 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_2988
timestamp 1668089732
transform 1 0 7680 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_2989
timestamp 1668089732
transform 1 0 7680 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_2990
timestamp 1668089732
transform 1 0 7680 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_2991
timestamp 1668089732
transform 1 0 7680 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_2992
timestamp 1668089732
transform 1 0 7680 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_2993
timestamp 1668089732
transform 1 0 7680 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_2994
timestamp 1668089732
transform 1 0 7680 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_2995
timestamp 1668089732
transform 1 0 7680 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_2996
timestamp 1668089732
transform 1 0 7680 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_2997
timestamp 1668089732
transform 1 0 7680 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_2998
timestamp 1668089732
transform 1 0 7680 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_2999
timestamp 1668089732
transform 1 0 7680 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_3000
timestamp 1668089732
transform 1 0 7680 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_3001
timestamp 1668089732
transform 1 0 7680 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_3002
timestamp 1668089732
transform 1 0 7680 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_3003
timestamp 1668089732
transform 1 0 7680 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_3004
timestamp 1668089732
transform 1 0 7680 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_3005
timestamp 1668089732
transform 1 0 7680 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_3006
timestamp 1668089732
transform 1 0 7680 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_3007
timestamp 1668089732
transform 1 0 7680 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_3008
timestamp 1668089732
transform 1 0 7680 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_3009
timestamp 1668089732
transform 1 0 7680 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_3010
timestamp 1668089732
transform 1 0 7680 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_3011
timestamp 1668089732
transform 1 0 7680 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_3012
timestamp 1668089732
transform 1 0 7680 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_3013
timestamp 1668089732
transform 1 0 7680 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_3014
timestamp 1668089732
transform 1 0 7680 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_3015
timestamp 1668089732
transform 1 0 7680 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_3016
timestamp 1668089732
transform 1 0 7680 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_3017
timestamp 1668089732
transform 1 0 7680 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_3018
timestamp 1668089732
transform 1 0 7680 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_3019
timestamp 1668089732
transform 1 0 7680 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_3020
timestamp 1668089732
transform 1 0 7680 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_3021
timestamp 1668089732
transform 1 0 7680 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_3022
timestamp 1668089732
transform 1 0 7680 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_3023
timestamp 1668089732
transform 1 0 7680 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_3024
timestamp 1668089732
transform 1 0 7680 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_3025
timestamp 1668089732
transform 1 0 7680 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_3026
timestamp 1668089732
transform 1 0 7680 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_3027
timestamp 1668089732
transform 1 0 7680 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_3028
timestamp 1668089732
transform 1 0 7680 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_3029
timestamp 1668089732
transform 1 0 7680 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_3030
timestamp 1668089732
transform 1 0 7680 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_3031
timestamp 1668089732
transform 1 0 7680 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_3032
timestamp 1668089732
transform 1 0 7680 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_3033
timestamp 1668089732
transform 1 0 7680 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_3034
timestamp 1668089732
transform 1 0 7680 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_3035
timestamp 1668089732
transform 1 0 7680 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_3036
timestamp 1668089732
transform 1 0 7680 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_3037
timestamp 1668089732
transform 1 0 7680 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_3038
timestamp 1668089732
transform 1 0 7840 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_3039
timestamp 1668089732
transform 1 0 7840 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_3040
timestamp 1668089732
transform 1 0 7840 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_3041
timestamp 1668089732
transform 1 0 7840 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_3042
timestamp 1668089732
transform 1 0 7840 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_3043
timestamp 1668089732
transform 1 0 7840 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_3044
timestamp 1668089732
transform 1 0 7840 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_3045
timestamp 1668089732
transform 1 0 7840 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_3046
timestamp 1668089732
transform 1 0 7840 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_3047
timestamp 1668089732
transform 1 0 7840 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_3048
timestamp 1668089732
transform 1 0 7840 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_3049
timestamp 1668089732
transform 1 0 7840 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_3050
timestamp 1668089732
transform 1 0 7840 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_3051
timestamp 1668089732
transform 1 0 7840 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_3052
timestamp 1668089732
transform 1 0 7840 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_3053
timestamp 1668089732
transform 1 0 7840 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_3054
timestamp 1668089732
transform 1 0 7840 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_3055
timestamp 1668089732
transform 1 0 7840 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_3056
timestamp 1668089732
transform 1 0 7840 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_3057
timestamp 1668089732
transform 1 0 7840 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_3058
timestamp 1668089732
transform 1 0 7840 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_3059
timestamp 1668089732
transform 1 0 7840 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_3060
timestamp 1668089732
transform 1 0 7840 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_3061
timestamp 1668089732
transform 1 0 7840 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_3062
timestamp 1668089732
transform 1 0 7840 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_3063
timestamp 1668089732
transform 1 0 7840 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_3064
timestamp 1668089732
transform 1 0 7840 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_3065
timestamp 1668089732
transform 1 0 7840 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_3066
timestamp 1668089732
transform 1 0 7840 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_3067
timestamp 1668089732
transform 1 0 7840 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_3068
timestamp 1668089732
transform 1 0 7840 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_3069
timestamp 1668089732
transform 1 0 7840 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_3070
timestamp 1668089732
transform 1 0 7840 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_3071
timestamp 1668089732
transform 1 0 7840 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_3072
timestamp 1668089732
transform 1 0 7840 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_3073
timestamp 1668089732
transform 1 0 7840 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_3074
timestamp 1668089732
transform 1 0 7840 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_3075
timestamp 1668089732
transform 1 0 7840 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_3076
timestamp 1668089732
transform 1 0 7840 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_3077
timestamp 1668089732
transform 1 0 7840 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_3078
timestamp 1668089732
transform 1 0 7840 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_3079
timestamp 1668089732
transform 1 0 7840 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_3080
timestamp 1668089732
transform 1 0 7840 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_3081
timestamp 1668089732
transform 1 0 7840 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_3082
timestamp 1668089732
transform 1 0 7840 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_3083
timestamp 1668089732
transform 1 0 7840 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_3084
timestamp 1668089732
transform 1 0 7840 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_3085
timestamp 1668089732
transform 1 0 7840 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_3086
timestamp 1668089732
transform 1 0 7840 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_3087
timestamp 1668089732
transform 1 0 7840 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_3088
timestamp 1668089732
transform 1 0 7840 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_3089
timestamp 1668089732
transform 1 0 7840 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_3090
timestamp 1668089732
transform 1 0 7840 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_3091
timestamp 1668089732
transform 1 0 7840 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_3092
timestamp 1668089732
transform 1 0 7840 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_3093
timestamp 1668089732
transform 1 0 7840 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_3094
timestamp 1668089732
transform 1 0 7840 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_3095
timestamp 1668089732
transform 1 0 7840 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_3096
timestamp 1668089732
transform 1 0 7840 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_3097
timestamp 1668089732
transform 1 0 7840 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_3098
timestamp 1668089732
transform 1 0 7840 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_3099
timestamp 1668089732
transform 1 0 7840 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_3100
timestamp 1668089732
transform 1 0 8000 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_3101
timestamp 1668089732
transform 1 0 8000 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_3102
timestamp 1668089732
transform 1 0 8000 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_3103
timestamp 1668089732
transform 1 0 8000 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_3104
timestamp 1668089732
transform 1 0 8000 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_3105
timestamp 1668089732
transform 1 0 8000 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_3106
timestamp 1668089732
transform 1 0 8000 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_3107
timestamp 1668089732
transform 1 0 8000 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_3108
timestamp 1668089732
transform 1 0 8000 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_3109
timestamp 1668089732
transform 1 0 8000 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_3110
timestamp 1668089732
transform 1 0 8000 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_3111
timestamp 1668089732
transform 1 0 8000 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_3112
timestamp 1668089732
transform 1 0 8000 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_3113
timestamp 1668089732
transform 1 0 8000 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_3114
timestamp 1668089732
transform 1 0 8000 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_3115
timestamp 1668089732
transform 1 0 8000 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_3116
timestamp 1668089732
transform 1 0 8000 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_3117
timestamp 1668089732
transform 1 0 8000 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_3118
timestamp 1668089732
transform 1 0 8000 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_3119
timestamp 1668089732
transform 1 0 8000 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_3120
timestamp 1668089732
transform 1 0 8000 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_3121
timestamp 1668089732
transform 1 0 8000 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_3122
timestamp 1668089732
transform 1 0 8000 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_3123
timestamp 1668089732
transform 1 0 8000 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_3124
timestamp 1668089732
transform 1 0 8000 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_3125
timestamp 1668089732
transform 1 0 8000 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_3126
timestamp 1668089732
transform 1 0 8000 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_3127
timestamp 1668089732
transform 1 0 8000 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_3128
timestamp 1668089732
transform 1 0 8000 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_3129
timestamp 1668089732
transform 1 0 8000 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_3130
timestamp 1668089732
transform 1 0 8000 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_3131
timestamp 1668089732
transform 1 0 8000 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_3132
timestamp 1668089732
transform 1 0 8000 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_3133
timestamp 1668089732
transform 1 0 8000 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_3134
timestamp 1668089732
transform 1 0 8000 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_3135
timestamp 1668089732
transform 1 0 8000 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_3136
timestamp 1668089732
transform 1 0 8000 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_3137
timestamp 1668089732
transform 1 0 8000 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_3138
timestamp 1668089732
transform 1 0 8000 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_3139
timestamp 1668089732
transform 1 0 8000 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_3140
timestamp 1668089732
transform 1 0 8000 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_3141
timestamp 1668089732
transform 1 0 8000 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_3142
timestamp 1668089732
transform 1 0 8000 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_3143
timestamp 1668089732
transform 1 0 8000 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_3144
timestamp 1668089732
transform 1 0 8000 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_3145
timestamp 1668089732
transform 1 0 8000 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_3146
timestamp 1668089732
transform 1 0 8000 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_3147
timestamp 1668089732
transform 1 0 8000 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_3148
timestamp 1668089732
transform 1 0 8000 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_3149
timestamp 1668089732
transform 1 0 8000 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_3150
timestamp 1668089732
transform 1 0 8000 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_3151
timestamp 1668089732
transform 1 0 8000 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_3152
timestamp 1668089732
transform 1 0 8000 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_3153
timestamp 1668089732
transform 1 0 8000 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_3154
timestamp 1668089732
transform 1 0 8000 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_3155
timestamp 1668089732
transform 1 0 8000 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_3156
timestamp 1668089732
transform 1 0 8000 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_3157
timestamp 1668089732
transform 1 0 8000 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_3158
timestamp 1668089732
transform 1 0 8000 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_3159
timestamp 1668089732
transform 1 0 8000 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_3160
timestamp 1668089732
transform 1 0 8000 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_3161
timestamp 1668089732
transform 1 0 8000 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_3162
timestamp 1668089732
transform 1 0 8160 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_3163
timestamp 1668089732
transform 1 0 8160 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_3164
timestamp 1668089732
transform 1 0 8160 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_3165
timestamp 1668089732
transform 1 0 8160 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_3166
timestamp 1668089732
transform 1 0 8160 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_3167
timestamp 1668089732
transform 1 0 8160 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_3168
timestamp 1668089732
transform 1 0 8160 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_3169
timestamp 1668089732
transform 1 0 8160 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_3170
timestamp 1668089732
transform 1 0 8160 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_3171
timestamp 1668089732
transform 1 0 8160 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_3172
timestamp 1668089732
transform 1 0 8160 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_3173
timestamp 1668089732
transform 1 0 8160 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_3174
timestamp 1668089732
transform 1 0 8160 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_3175
timestamp 1668089732
transform 1 0 8160 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_3176
timestamp 1668089732
transform 1 0 8160 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_3177
timestamp 1668089732
transform 1 0 8160 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_3178
timestamp 1668089732
transform 1 0 8160 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_3179
timestamp 1668089732
transform 1 0 8160 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_3180
timestamp 1668089732
transform 1 0 8160 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_3181
timestamp 1668089732
transform 1 0 8160 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_3182
timestamp 1668089732
transform 1 0 8160 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_3183
timestamp 1668089732
transform 1 0 8160 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_3184
timestamp 1668089732
transform 1 0 8160 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_3185
timestamp 1668089732
transform 1 0 8160 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_3186
timestamp 1668089732
transform 1 0 8160 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_3187
timestamp 1668089732
transform 1 0 8160 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_3188
timestamp 1668089732
transform 1 0 8160 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_3189
timestamp 1668089732
transform 1 0 8160 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_3190
timestamp 1668089732
transform 1 0 8160 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_3191
timestamp 1668089732
transform 1 0 8160 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_3192
timestamp 1668089732
transform 1 0 8160 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_3193
timestamp 1668089732
transform 1 0 8160 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_3194
timestamp 1668089732
transform 1 0 8160 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_3195
timestamp 1668089732
transform 1 0 8160 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_3196
timestamp 1668089732
transform 1 0 8160 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_3197
timestamp 1668089732
transform 1 0 8160 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_3198
timestamp 1668089732
transform 1 0 8160 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_3199
timestamp 1668089732
transform 1 0 8160 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_3200
timestamp 1668089732
transform 1 0 8160 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_3201
timestamp 1668089732
transform 1 0 8160 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_3202
timestamp 1668089732
transform 1 0 8160 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_3203
timestamp 1668089732
transform 1 0 8160 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_3204
timestamp 1668089732
transform 1 0 8160 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_3205
timestamp 1668089732
transform 1 0 8160 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_3206
timestamp 1668089732
transform 1 0 8160 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_3207
timestamp 1668089732
transform 1 0 8160 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_3208
timestamp 1668089732
transform 1 0 8160 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_3209
timestamp 1668089732
transform 1 0 8160 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_3210
timestamp 1668089732
transform 1 0 8160 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_3211
timestamp 1668089732
transform 1 0 8160 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_3212
timestamp 1668089732
transform 1 0 8160 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_3213
timestamp 1668089732
transform 1 0 8160 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_3214
timestamp 1668089732
transform 1 0 8160 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_3215
timestamp 1668089732
transform 1 0 8160 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_3216
timestamp 1668089732
transform 1 0 8160 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_3217
timestamp 1668089732
transform 1 0 8160 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_3218
timestamp 1668089732
transform 1 0 8160 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_3219
timestamp 1668089732
transform 1 0 8160 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_3220
timestamp 1668089732
transform 1 0 8160 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_3221
timestamp 1668089732
transform 1 0 8160 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_3222
timestamp 1668089732
transform 1 0 8160 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_3223
timestamp 1668089732
transform 1 0 8160 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_3224
timestamp 1668089732
transform 1 0 8320 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_3225
timestamp 1668089732
transform 1 0 8320 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_3226
timestamp 1668089732
transform 1 0 8320 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_3227
timestamp 1668089732
transform 1 0 8320 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_3228
timestamp 1668089732
transform 1 0 8320 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_3229
timestamp 1668089732
transform 1 0 8320 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_3230
timestamp 1668089732
transform 1 0 8320 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_3231
timestamp 1668089732
transform 1 0 8320 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_3232
timestamp 1668089732
transform 1 0 8320 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_3233
timestamp 1668089732
transform 1 0 8320 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_3234
timestamp 1668089732
transform 1 0 8320 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_3235
timestamp 1668089732
transform 1 0 8320 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_3236
timestamp 1668089732
transform 1 0 8320 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_3237
timestamp 1668089732
transform 1 0 8320 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_3238
timestamp 1668089732
transform 1 0 8320 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_3239
timestamp 1668089732
transform 1 0 8320 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_3240
timestamp 1668089732
transform 1 0 8320 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_3241
timestamp 1668089732
transform 1 0 8320 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_3242
timestamp 1668089732
transform 1 0 8320 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_3243
timestamp 1668089732
transform 1 0 8320 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_3244
timestamp 1668089732
transform 1 0 8320 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_3245
timestamp 1668089732
transform 1 0 8320 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_3246
timestamp 1668089732
transform 1 0 8320 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_3247
timestamp 1668089732
transform 1 0 8320 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_3248
timestamp 1668089732
transform 1 0 8320 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_3249
timestamp 1668089732
transform 1 0 8320 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_3250
timestamp 1668089732
transform 1 0 8320 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_3251
timestamp 1668089732
transform 1 0 8320 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_3252
timestamp 1668089732
transform 1 0 8320 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_3253
timestamp 1668089732
transform 1 0 8320 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_3254
timestamp 1668089732
transform 1 0 8320 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_3255
timestamp 1668089732
transform 1 0 8320 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_3256
timestamp 1668089732
transform 1 0 8320 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_3257
timestamp 1668089732
transform 1 0 8320 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_3258
timestamp 1668089732
transform 1 0 8320 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_3259
timestamp 1668089732
transform 1 0 8320 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_3260
timestamp 1668089732
transform 1 0 8320 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_3261
timestamp 1668089732
transform 1 0 8320 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_3262
timestamp 1668089732
transform 1 0 8320 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_3263
timestamp 1668089732
transform 1 0 8320 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_3264
timestamp 1668089732
transform 1 0 8320 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_3265
timestamp 1668089732
transform 1 0 8320 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_3266
timestamp 1668089732
transform 1 0 8320 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_3267
timestamp 1668089732
transform 1 0 8320 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_3268
timestamp 1668089732
transform 1 0 8320 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_3269
timestamp 1668089732
transform 1 0 8320 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_3270
timestamp 1668089732
transform 1 0 8320 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_3271
timestamp 1668089732
transform 1 0 8320 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_3272
timestamp 1668089732
transform 1 0 8320 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_3273
timestamp 1668089732
transform 1 0 8320 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_3274
timestamp 1668089732
transform 1 0 8320 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_3275
timestamp 1668089732
transform 1 0 8320 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_3276
timestamp 1668089732
transform 1 0 8320 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_3277
timestamp 1668089732
transform 1 0 8320 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_3278
timestamp 1668089732
transform 1 0 8320 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_3279
timestamp 1668089732
transform 1 0 8320 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_3280
timestamp 1668089732
transform 1 0 8320 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_3281
timestamp 1668089732
transform 1 0 8320 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_3282
timestamp 1668089732
transform 1 0 8320 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_3283
timestamp 1668089732
transform 1 0 8320 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_3284
timestamp 1668089732
transform 1 0 8320 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_3285
timestamp 1668089732
transform 1 0 8320 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_3286
timestamp 1668089732
transform 1 0 8480 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_3287
timestamp 1668089732
transform 1 0 8480 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_3288
timestamp 1668089732
transform 1 0 8480 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_3289
timestamp 1668089732
transform 1 0 8480 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_3290
timestamp 1668089732
transform 1 0 8480 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_3291
timestamp 1668089732
transform 1 0 8480 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_3292
timestamp 1668089732
transform 1 0 8480 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_3293
timestamp 1668089732
transform 1 0 8480 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_3294
timestamp 1668089732
transform 1 0 8480 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_3295
timestamp 1668089732
transform 1 0 8480 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_3296
timestamp 1668089732
transform 1 0 8480 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_3297
timestamp 1668089732
transform 1 0 8480 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_3298
timestamp 1668089732
transform 1 0 8480 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_3299
timestamp 1668089732
transform 1 0 8480 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_3300
timestamp 1668089732
transform 1 0 8480 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_3301
timestamp 1668089732
transform 1 0 8480 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_3302
timestamp 1668089732
transform 1 0 8480 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_3303
timestamp 1668089732
transform 1 0 8480 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_3304
timestamp 1668089732
transform 1 0 8480 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_3305
timestamp 1668089732
transform 1 0 8480 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_3306
timestamp 1668089732
transform 1 0 8480 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_3307
timestamp 1668089732
transform 1 0 8480 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_3308
timestamp 1668089732
transform 1 0 8480 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_3309
timestamp 1668089732
transform 1 0 8480 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_3310
timestamp 1668089732
transform 1 0 8480 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_3311
timestamp 1668089732
transform 1 0 8480 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_3312
timestamp 1668089732
transform 1 0 8480 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_3313
timestamp 1668089732
transform 1 0 8480 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_3314
timestamp 1668089732
transform 1 0 8480 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_3315
timestamp 1668089732
transform 1 0 8480 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_3316
timestamp 1668089732
transform 1 0 8480 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_3317
timestamp 1668089732
transform 1 0 8480 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_3318
timestamp 1668089732
transform 1 0 8480 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_3319
timestamp 1668089732
transform 1 0 8480 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_3320
timestamp 1668089732
transform 1 0 8480 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_3321
timestamp 1668089732
transform 1 0 8480 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_3322
timestamp 1668089732
transform 1 0 8480 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_3323
timestamp 1668089732
transform 1 0 8480 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_3324
timestamp 1668089732
transform 1 0 8480 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_3325
timestamp 1668089732
transform 1 0 8480 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_3326
timestamp 1668089732
transform 1 0 8480 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_3327
timestamp 1668089732
transform 1 0 8480 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_3328
timestamp 1668089732
transform 1 0 8480 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_3329
timestamp 1668089732
transform 1 0 8480 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_3330
timestamp 1668089732
transform 1 0 8480 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_3331
timestamp 1668089732
transform 1 0 8480 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_3332
timestamp 1668089732
transform 1 0 8480 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_3333
timestamp 1668089732
transform 1 0 8480 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_3334
timestamp 1668089732
transform 1 0 8480 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_3335
timestamp 1668089732
transform 1 0 8480 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_3336
timestamp 1668089732
transform 1 0 8480 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_3337
timestamp 1668089732
transform 1 0 8480 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_3338
timestamp 1668089732
transform 1 0 8480 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_3339
timestamp 1668089732
transform 1 0 8480 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_3340
timestamp 1668089732
transform 1 0 8480 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_3341
timestamp 1668089732
transform 1 0 8480 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_3342
timestamp 1668089732
transform 1 0 8480 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_3343
timestamp 1668089732
transform 1 0 8480 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_3344
timestamp 1668089732
transform 1 0 8480 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_3345
timestamp 1668089732
transform 1 0 8480 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_3346
timestamp 1668089732
transform 1 0 8480 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_3347
timestamp 1668089732
transform 1 0 8480 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_3348
timestamp 1668089732
transform 1 0 8640 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_3349
timestamp 1668089732
transform 1 0 8640 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_3350
timestamp 1668089732
transform 1 0 8640 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_3351
timestamp 1668089732
transform 1 0 8640 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_3352
timestamp 1668089732
transform 1 0 8640 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_3353
timestamp 1668089732
transform 1 0 8640 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_3354
timestamp 1668089732
transform 1 0 8640 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_3355
timestamp 1668089732
transform 1 0 8640 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_3356
timestamp 1668089732
transform 1 0 8640 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_3357
timestamp 1668089732
transform 1 0 8640 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_3358
timestamp 1668089732
transform 1 0 8640 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_3359
timestamp 1668089732
transform 1 0 8640 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_3360
timestamp 1668089732
transform 1 0 8640 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_3361
timestamp 1668089732
transform 1 0 8640 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_3362
timestamp 1668089732
transform 1 0 8640 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_3363
timestamp 1668089732
transform 1 0 8640 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_3364
timestamp 1668089732
transform 1 0 8640 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_3365
timestamp 1668089732
transform 1 0 8640 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_3366
timestamp 1668089732
transform 1 0 8640 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_3367
timestamp 1668089732
transform 1 0 8640 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_3368
timestamp 1668089732
transform 1 0 8640 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_3369
timestamp 1668089732
transform 1 0 8640 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_3370
timestamp 1668089732
transform 1 0 8640 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_3371
timestamp 1668089732
transform 1 0 8640 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_3372
timestamp 1668089732
transform 1 0 8640 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_3373
timestamp 1668089732
transform 1 0 8640 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_3374
timestamp 1668089732
transform 1 0 8640 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_3375
timestamp 1668089732
transform 1 0 8640 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_3376
timestamp 1668089732
transform 1 0 8640 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_3377
timestamp 1668089732
transform 1 0 8640 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_3378
timestamp 1668089732
transform 1 0 8640 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_3379
timestamp 1668089732
transform 1 0 8640 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_3380
timestamp 1668089732
transform 1 0 8640 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_3381
timestamp 1668089732
transform 1 0 8640 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_3382
timestamp 1668089732
transform 1 0 8640 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_3383
timestamp 1668089732
transform 1 0 8640 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_3384
timestamp 1668089732
transform 1 0 8640 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_3385
timestamp 1668089732
transform 1 0 8640 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_3386
timestamp 1668089732
transform 1 0 8640 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_3387
timestamp 1668089732
transform 1 0 8640 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_3388
timestamp 1668089732
transform 1 0 8640 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_3389
timestamp 1668089732
transform 1 0 8640 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_3390
timestamp 1668089732
transform 1 0 8640 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_3391
timestamp 1668089732
transform 1 0 8640 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_3392
timestamp 1668089732
transform 1 0 8640 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_3393
timestamp 1668089732
transform 1 0 8640 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_3394
timestamp 1668089732
transform 1 0 8640 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_3395
timestamp 1668089732
transform 1 0 8640 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_3396
timestamp 1668089732
transform 1 0 8640 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_3397
timestamp 1668089732
transform 1 0 8640 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_3398
timestamp 1668089732
transform 1 0 8640 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_3399
timestamp 1668089732
transform 1 0 8640 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_3400
timestamp 1668089732
transform 1 0 8640 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_3401
timestamp 1668089732
transform 1 0 8640 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_3402
timestamp 1668089732
transform 1 0 8640 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_3403
timestamp 1668089732
transform 1 0 8640 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_3404
timestamp 1668089732
transform 1 0 8640 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_3405
timestamp 1668089732
transform 1 0 8640 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_3406
timestamp 1668089732
transform 1 0 8640 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_3407
timestamp 1668089732
transform 1 0 8640 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_3408
timestamp 1668089732
transform 1 0 8640 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_3409
timestamp 1668089732
transform 1 0 8640 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_3410
timestamp 1668089732
transform 1 0 8800 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_3411
timestamp 1668089732
transform 1 0 8800 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_3412
timestamp 1668089732
transform 1 0 8800 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_3413
timestamp 1668089732
transform 1 0 8800 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_3414
timestamp 1668089732
transform 1 0 8800 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_3415
timestamp 1668089732
transform 1 0 8800 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_3416
timestamp 1668089732
transform 1 0 8800 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_3417
timestamp 1668089732
transform 1 0 8800 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_3418
timestamp 1668089732
transform 1 0 8800 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_3419
timestamp 1668089732
transform 1 0 8800 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_3420
timestamp 1668089732
transform 1 0 8800 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_3421
timestamp 1668089732
transform 1 0 8800 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_3422
timestamp 1668089732
transform 1 0 8800 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_3423
timestamp 1668089732
transform 1 0 8800 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_3424
timestamp 1668089732
transform 1 0 8800 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_3425
timestamp 1668089732
transform 1 0 8800 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_3426
timestamp 1668089732
transform 1 0 8800 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_3427
timestamp 1668089732
transform 1 0 8800 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_3428
timestamp 1668089732
transform 1 0 8800 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_3429
timestamp 1668089732
transform 1 0 8800 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_3430
timestamp 1668089732
transform 1 0 8800 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_3431
timestamp 1668089732
transform 1 0 8800 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_3432
timestamp 1668089732
transform 1 0 8800 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_3433
timestamp 1668089732
transform 1 0 8800 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_3434
timestamp 1668089732
transform 1 0 8800 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_3435
timestamp 1668089732
transform 1 0 8800 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_3436
timestamp 1668089732
transform 1 0 8800 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_3437
timestamp 1668089732
transform 1 0 8800 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_3438
timestamp 1668089732
transform 1 0 8800 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_3439
timestamp 1668089732
transform 1 0 8800 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_3440
timestamp 1668089732
transform 1 0 8800 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_3441
timestamp 1668089732
transform 1 0 8800 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_3442
timestamp 1668089732
transform 1 0 8800 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_3443
timestamp 1668089732
transform 1 0 8800 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_3444
timestamp 1668089732
transform 1 0 8800 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_3445
timestamp 1668089732
transform 1 0 8800 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_3446
timestamp 1668089732
transform 1 0 8800 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_3447
timestamp 1668089732
transform 1 0 8800 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_3448
timestamp 1668089732
transform 1 0 8800 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_3449
timestamp 1668089732
transform 1 0 8800 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_3450
timestamp 1668089732
transform 1 0 8800 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_3451
timestamp 1668089732
transform 1 0 8800 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_3452
timestamp 1668089732
transform 1 0 8800 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_3453
timestamp 1668089732
transform 1 0 8800 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_3454
timestamp 1668089732
transform 1 0 8800 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_3455
timestamp 1668089732
transform 1 0 8800 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_3456
timestamp 1668089732
transform 1 0 8800 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_3457
timestamp 1668089732
transform 1 0 8800 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_3458
timestamp 1668089732
transform 1 0 8800 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_3459
timestamp 1668089732
transform 1 0 8800 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_3460
timestamp 1668089732
transform 1 0 8800 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_3461
timestamp 1668089732
transform 1 0 8800 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_3462
timestamp 1668089732
transform 1 0 8800 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_3463
timestamp 1668089732
transform 1 0 8800 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_3464
timestamp 1668089732
transform 1 0 8800 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_3465
timestamp 1668089732
transform 1 0 8800 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_3466
timestamp 1668089732
transform 1 0 8800 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_3467
timestamp 1668089732
transform 1 0 8800 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_3468
timestamp 1668089732
transform 1 0 8800 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_3469
timestamp 1668089732
transform 1 0 8800 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_3470
timestamp 1668089732
transform 1 0 8800 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_3471
timestamp 1668089732
transform 1 0 8800 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_3472
timestamp 1668089732
transform 1 0 8960 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_3473
timestamp 1668089732
transform 1 0 8960 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_3474
timestamp 1668089732
transform 1 0 8960 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_3475
timestamp 1668089732
transform 1 0 8960 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_3476
timestamp 1668089732
transform 1 0 8960 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_3477
timestamp 1668089732
transform 1 0 8960 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_3478
timestamp 1668089732
transform 1 0 8960 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_3479
timestamp 1668089732
transform 1 0 8960 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_3480
timestamp 1668089732
transform 1 0 8960 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_3481
timestamp 1668089732
transform 1 0 8960 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_3482
timestamp 1668089732
transform 1 0 8960 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_3483
timestamp 1668089732
transform 1 0 8960 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_3484
timestamp 1668089732
transform 1 0 8960 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_3485
timestamp 1668089732
transform 1 0 8960 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_3486
timestamp 1668089732
transform 1 0 8960 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_3487
timestamp 1668089732
transform 1 0 8960 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_3488
timestamp 1668089732
transform 1 0 8960 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_3489
timestamp 1668089732
transform 1 0 8960 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_3490
timestamp 1668089732
transform 1 0 8960 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_3491
timestamp 1668089732
transform 1 0 8960 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_3492
timestamp 1668089732
transform 1 0 8960 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_3493
timestamp 1668089732
transform 1 0 8960 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_3494
timestamp 1668089732
transform 1 0 8960 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_3495
timestamp 1668089732
transform 1 0 8960 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_3496
timestamp 1668089732
transform 1 0 8960 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_3497
timestamp 1668089732
transform 1 0 8960 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_3498
timestamp 1668089732
transform 1 0 8960 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_3499
timestamp 1668089732
transform 1 0 8960 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_3500
timestamp 1668089732
transform 1 0 8960 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_3501
timestamp 1668089732
transform 1 0 8960 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_3502
timestamp 1668089732
transform 1 0 8960 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_3503
timestamp 1668089732
transform 1 0 8960 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_3504
timestamp 1668089732
transform 1 0 8960 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_3505
timestamp 1668089732
transform 1 0 8960 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_3506
timestamp 1668089732
transform 1 0 8960 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_3507
timestamp 1668089732
transform 1 0 8960 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_3508
timestamp 1668089732
transform 1 0 8960 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_3509
timestamp 1668089732
transform 1 0 8960 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_3510
timestamp 1668089732
transform 1 0 8960 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_3511
timestamp 1668089732
transform 1 0 8960 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_3512
timestamp 1668089732
transform 1 0 8960 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_3513
timestamp 1668089732
transform 1 0 8960 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_3514
timestamp 1668089732
transform 1 0 8960 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_3515
timestamp 1668089732
transform 1 0 8960 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_3516
timestamp 1668089732
transform 1 0 8960 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_3517
timestamp 1668089732
transform 1 0 8960 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_3518
timestamp 1668089732
transform 1 0 8960 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_3519
timestamp 1668089732
transform 1 0 8960 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_3520
timestamp 1668089732
transform 1 0 8960 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_3521
timestamp 1668089732
transform 1 0 8960 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_3522
timestamp 1668089732
transform 1 0 8960 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_3523
timestamp 1668089732
transform 1 0 8960 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_3524
timestamp 1668089732
transform 1 0 8960 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_3525
timestamp 1668089732
transform 1 0 8960 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_3526
timestamp 1668089732
transform 1 0 8960 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_3527
timestamp 1668089732
transform 1 0 8960 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_3528
timestamp 1668089732
transform 1 0 8960 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_3529
timestamp 1668089732
transform 1 0 8960 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_3530
timestamp 1668089732
transform 1 0 8960 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_3531
timestamp 1668089732
transform 1 0 8960 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_3532
timestamp 1668089732
transform 1 0 8960 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_3533
timestamp 1668089732
transform 1 0 8960 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_3534
timestamp 1668089732
transform 1 0 9120 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_3535
timestamp 1668089732
transform 1 0 9120 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_3536
timestamp 1668089732
transform 1 0 9120 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_3537
timestamp 1668089732
transform 1 0 9120 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_3538
timestamp 1668089732
transform 1 0 9120 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_3539
timestamp 1668089732
transform 1 0 9120 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_3540
timestamp 1668089732
transform 1 0 9120 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_3541
timestamp 1668089732
transform 1 0 9120 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_3542
timestamp 1668089732
transform 1 0 9120 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_3543
timestamp 1668089732
transform 1 0 9120 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_3544
timestamp 1668089732
transform 1 0 9120 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_3545
timestamp 1668089732
transform 1 0 9120 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_3546
timestamp 1668089732
transform 1 0 9120 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_3547
timestamp 1668089732
transform 1 0 9120 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_3548
timestamp 1668089732
transform 1 0 9120 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_3549
timestamp 1668089732
transform 1 0 9120 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_3550
timestamp 1668089732
transform 1 0 9120 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_3551
timestamp 1668089732
transform 1 0 9120 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_3552
timestamp 1668089732
transform 1 0 9120 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_3553
timestamp 1668089732
transform 1 0 9120 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_3554
timestamp 1668089732
transform 1 0 9120 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_3555
timestamp 1668089732
transform 1 0 9120 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_3556
timestamp 1668089732
transform 1 0 9120 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_3557
timestamp 1668089732
transform 1 0 9120 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_3558
timestamp 1668089732
transform 1 0 9120 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_3559
timestamp 1668089732
transform 1 0 9120 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_3560
timestamp 1668089732
transform 1 0 9120 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_3561
timestamp 1668089732
transform 1 0 9120 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_3562
timestamp 1668089732
transform 1 0 9120 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_3563
timestamp 1668089732
transform 1 0 9120 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_3564
timestamp 1668089732
transform 1 0 9120 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_3565
timestamp 1668089732
transform 1 0 9120 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_3566
timestamp 1668089732
transform 1 0 9120 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_3567
timestamp 1668089732
transform 1 0 9120 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_3568
timestamp 1668089732
transform 1 0 9120 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_3569
timestamp 1668089732
transform 1 0 9120 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_3570
timestamp 1668089732
transform 1 0 9120 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_3571
timestamp 1668089732
transform 1 0 9120 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_3572
timestamp 1668089732
transform 1 0 9120 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_3573
timestamp 1668089732
transform 1 0 9120 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_3574
timestamp 1668089732
transform 1 0 9120 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_3575
timestamp 1668089732
transform 1 0 9120 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_3576
timestamp 1668089732
transform 1 0 9120 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_3577
timestamp 1668089732
transform 1 0 9120 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_3578
timestamp 1668089732
transform 1 0 9120 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_3579
timestamp 1668089732
transform 1 0 9120 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_3580
timestamp 1668089732
transform 1 0 9120 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_3581
timestamp 1668089732
transform 1 0 9120 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_3582
timestamp 1668089732
transform 1 0 9120 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_3583
timestamp 1668089732
transform 1 0 9120 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_3584
timestamp 1668089732
transform 1 0 9120 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_3585
timestamp 1668089732
transform 1 0 9120 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_3586
timestamp 1668089732
transform 1 0 9120 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_3587
timestamp 1668089732
transform 1 0 9120 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_3588
timestamp 1668089732
transform 1 0 9120 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_3589
timestamp 1668089732
transform 1 0 9120 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_3590
timestamp 1668089732
transform 1 0 9120 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_3591
timestamp 1668089732
transform 1 0 9120 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_3592
timestamp 1668089732
transform 1 0 9120 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_3593
timestamp 1668089732
transform 1 0 9120 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_3594
timestamp 1668089732
transform 1 0 9120 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_3595
timestamp 1668089732
transform 1 0 9120 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_3596
timestamp 1668089732
transform 1 0 9280 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_3597
timestamp 1668089732
transform 1 0 9280 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_3598
timestamp 1668089732
transform 1 0 9280 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_3599
timestamp 1668089732
transform 1 0 9280 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_3600
timestamp 1668089732
transform 1 0 9280 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_3601
timestamp 1668089732
transform 1 0 9280 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_3602
timestamp 1668089732
transform 1 0 9280 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_3603
timestamp 1668089732
transform 1 0 9280 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_3604
timestamp 1668089732
transform 1 0 9280 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_3605
timestamp 1668089732
transform 1 0 9280 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_3606
timestamp 1668089732
transform 1 0 9280 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_3607
timestamp 1668089732
transform 1 0 9280 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_3608
timestamp 1668089732
transform 1 0 9280 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_3609
timestamp 1668089732
transform 1 0 9280 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_3610
timestamp 1668089732
transform 1 0 9280 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_3611
timestamp 1668089732
transform 1 0 9280 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_3612
timestamp 1668089732
transform 1 0 9280 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_3613
timestamp 1668089732
transform 1 0 9280 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_3614
timestamp 1668089732
transform 1 0 9280 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_3615
timestamp 1668089732
transform 1 0 9280 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_3616
timestamp 1668089732
transform 1 0 9280 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_3617
timestamp 1668089732
transform 1 0 9280 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_3618
timestamp 1668089732
transform 1 0 9280 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_3619
timestamp 1668089732
transform 1 0 9280 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_3620
timestamp 1668089732
transform 1 0 9280 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_3621
timestamp 1668089732
transform 1 0 9280 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_3622
timestamp 1668089732
transform 1 0 9280 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_3623
timestamp 1668089732
transform 1 0 9280 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_3624
timestamp 1668089732
transform 1 0 9280 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_3625
timestamp 1668089732
transform 1 0 9280 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_3626
timestamp 1668089732
transform 1 0 9280 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_3627
timestamp 1668089732
transform 1 0 9280 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_3628
timestamp 1668089732
transform 1 0 9280 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_3629
timestamp 1668089732
transform 1 0 9280 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_3630
timestamp 1668089732
transform 1 0 9280 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_3631
timestamp 1668089732
transform 1 0 9280 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_3632
timestamp 1668089732
transform 1 0 9280 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_3633
timestamp 1668089732
transform 1 0 9280 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_3634
timestamp 1668089732
transform 1 0 9280 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_3635
timestamp 1668089732
transform 1 0 9280 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_3636
timestamp 1668089732
transform 1 0 9280 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_3637
timestamp 1668089732
transform 1 0 9280 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_3638
timestamp 1668089732
transform 1 0 9280 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_3639
timestamp 1668089732
transform 1 0 9280 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_3640
timestamp 1668089732
transform 1 0 9280 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_3641
timestamp 1668089732
transform 1 0 9280 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_3642
timestamp 1668089732
transform 1 0 9280 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_3643
timestamp 1668089732
transform 1 0 9280 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_3644
timestamp 1668089732
transform 1 0 9280 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_3645
timestamp 1668089732
transform 1 0 9280 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_3646
timestamp 1668089732
transform 1 0 9280 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_3647
timestamp 1668089732
transform 1 0 9280 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_3648
timestamp 1668089732
transform 1 0 9280 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_3649
timestamp 1668089732
transform 1 0 9280 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_3650
timestamp 1668089732
transform 1 0 9280 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_3651
timestamp 1668089732
transform 1 0 9280 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_3652
timestamp 1668089732
transform 1 0 9280 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_3653
timestamp 1668089732
transform 1 0 9280 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_3654
timestamp 1668089732
transform 1 0 9280 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_3655
timestamp 1668089732
transform 1 0 9280 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_3656
timestamp 1668089732
transform 1 0 9280 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_3657
timestamp 1668089732
transform 1 0 9280 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_3658
timestamp 1668089732
transform 1 0 9440 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_3659
timestamp 1668089732
transform 1 0 9440 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_3660
timestamp 1668089732
transform 1 0 9440 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_3661
timestamp 1668089732
transform 1 0 9440 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_3662
timestamp 1668089732
transform 1 0 9440 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_3663
timestamp 1668089732
transform 1 0 9440 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_3664
timestamp 1668089732
transform 1 0 9440 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_3665
timestamp 1668089732
transform 1 0 9440 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_3666
timestamp 1668089732
transform 1 0 9440 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_3667
timestamp 1668089732
transform 1 0 9440 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_3668
timestamp 1668089732
transform 1 0 9440 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_3669
timestamp 1668089732
transform 1 0 9440 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_3670
timestamp 1668089732
transform 1 0 9440 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_3671
timestamp 1668089732
transform 1 0 9440 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_3672
timestamp 1668089732
transform 1 0 9440 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_3673
timestamp 1668089732
transform 1 0 9440 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_3674
timestamp 1668089732
transform 1 0 9440 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_3675
timestamp 1668089732
transform 1 0 9440 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_3676
timestamp 1668089732
transform 1 0 9440 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_3677
timestamp 1668089732
transform 1 0 9440 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_3678
timestamp 1668089732
transform 1 0 9440 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_3679
timestamp 1668089732
transform 1 0 9440 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_3680
timestamp 1668089732
transform 1 0 9440 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_3681
timestamp 1668089732
transform 1 0 9440 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_3682
timestamp 1668089732
transform 1 0 9440 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_3683
timestamp 1668089732
transform 1 0 9440 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_3684
timestamp 1668089732
transform 1 0 9440 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_3685
timestamp 1668089732
transform 1 0 9440 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_3686
timestamp 1668089732
transform 1 0 9440 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_3687
timestamp 1668089732
transform 1 0 9440 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_3688
timestamp 1668089732
transform 1 0 9440 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_3689
timestamp 1668089732
transform 1 0 9440 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_3690
timestamp 1668089732
transform 1 0 9440 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_3691
timestamp 1668089732
transform 1 0 9440 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_3692
timestamp 1668089732
transform 1 0 9440 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_3693
timestamp 1668089732
transform 1 0 9440 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_3694
timestamp 1668089732
transform 1 0 9440 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_3695
timestamp 1668089732
transform 1 0 9440 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_3696
timestamp 1668089732
transform 1 0 9440 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_3697
timestamp 1668089732
transform 1 0 9440 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_3698
timestamp 1668089732
transform 1 0 9440 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_3699
timestamp 1668089732
transform 1 0 9440 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_3700
timestamp 1668089732
transform 1 0 9440 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_3701
timestamp 1668089732
transform 1 0 9440 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_3702
timestamp 1668089732
transform 1 0 9440 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_3703
timestamp 1668089732
transform 1 0 9440 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_3704
timestamp 1668089732
transform 1 0 9440 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_3705
timestamp 1668089732
transform 1 0 9440 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_3706
timestamp 1668089732
transform 1 0 9440 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_3707
timestamp 1668089732
transform 1 0 9440 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_3708
timestamp 1668089732
transform 1 0 9440 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_3709
timestamp 1668089732
transform 1 0 9440 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_3710
timestamp 1668089732
transform 1 0 9440 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_3711
timestamp 1668089732
transform 1 0 9440 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_3712
timestamp 1668089732
transform 1 0 9440 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_3713
timestamp 1668089732
transform 1 0 9440 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_3714
timestamp 1668089732
transform 1 0 9440 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_3715
timestamp 1668089732
transform 1 0 9440 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_3716
timestamp 1668089732
transform 1 0 9440 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_3717
timestamp 1668089732
transform 1 0 9440 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_3718
timestamp 1668089732
transform 1 0 9440 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_3719
timestamp 1668089732
transform 1 0 9440 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_3720
timestamp 1668089732
transform 1 0 9600 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_3721
timestamp 1668089732
transform 1 0 9600 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_3722
timestamp 1668089732
transform 1 0 9600 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_3723
timestamp 1668089732
transform 1 0 9600 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_3724
timestamp 1668089732
transform 1 0 9600 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_3725
timestamp 1668089732
transform 1 0 9600 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_3726
timestamp 1668089732
transform 1 0 9600 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_3727
timestamp 1668089732
transform 1 0 9600 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_3728
timestamp 1668089732
transform 1 0 9600 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_3729
timestamp 1668089732
transform 1 0 9600 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_3730
timestamp 1668089732
transform 1 0 9600 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_3731
timestamp 1668089732
transform 1 0 9600 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_3732
timestamp 1668089732
transform 1 0 9600 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_3733
timestamp 1668089732
transform 1 0 9600 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_3734
timestamp 1668089732
transform 1 0 9600 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_3735
timestamp 1668089732
transform 1 0 9600 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_3736
timestamp 1668089732
transform 1 0 9600 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_3737
timestamp 1668089732
transform 1 0 9600 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_3738
timestamp 1668089732
transform 1 0 9600 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_3739
timestamp 1668089732
transform 1 0 9600 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_3740
timestamp 1668089732
transform 1 0 9600 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_3741
timestamp 1668089732
transform 1 0 9600 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_3742
timestamp 1668089732
transform 1 0 9600 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_3743
timestamp 1668089732
transform 1 0 9600 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_3744
timestamp 1668089732
transform 1 0 9600 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_3745
timestamp 1668089732
transform 1 0 9600 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_3746
timestamp 1668089732
transform 1 0 9600 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_3747
timestamp 1668089732
transform 1 0 9600 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_3748
timestamp 1668089732
transform 1 0 9600 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_3749
timestamp 1668089732
transform 1 0 9600 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_3750
timestamp 1668089732
transform 1 0 9600 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_3751
timestamp 1668089732
transform 1 0 9600 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_3752
timestamp 1668089732
transform 1 0 9600 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_3753
timestamp 1668089732
transform 1 0 9600 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_3754
timestamp 1668089732
transform 1 0 9600 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_3755
timestamp 1668089732
transform 1 0 9600 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_3756
timestamp 1668089732
transform 1 0 9600 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_3757
timestamp 1668089732
transform 1 0 9600 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_3758
timestamp 1668089732
transform 1 0 9600 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_3759
timestamp 1668089732
transform 1 0 9600 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_3760
timestamp 1668089732
transform 1 0 9600 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_3761
timestamp 1668089732
transform 1 0 9600 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_3762
timestamp 1668089732
transform 1 0 9600 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_3763
timestamp 1668089732
transform 1 0 9600 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_3764
timestamp 1668089732
transform 1 0 9600 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_3765
timestamp 1668089732
transform 1 0 9600 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_3766
timestamp 1668089732
transform 1 0 9600 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_3767
timestamp 1668089732
transform 1 0 9600 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_3768
timestamp 1668089732
transform 1 0 9600 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_3769
timestamp 1668089732
transform 1 0 9600 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_3770
timestamp 1668089732
transform 1 0 9600 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_3771
timestamp 1668089732
transform 1 0 9600 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_3772
timestamp 1668089732
transform 1 0 9600 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_3773
timestamp 1668089732
transform 1 0 9600 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_3774
timestamp 1668089732
transform 1 0 9600 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_3775
timestamp 1668089732
transform 1 0 9600 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_3776
timestamp 1668089732
transform 1 0 9600 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_3777
timestamp 1668089732
transform 1 0 9600 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_3778
timestamp 1668089732
transform 1 0 9600 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_3779
timestamp 1668089732
transform 1 0 9600 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_3780
timestamp 1668089732
transform 1 0 9600 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_3781
timestamp 1668089732
transform 1 0 9600 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_3782
timestamp 1668089732
transform 1 0 9760 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_3783
timestamp 1668089732
transform 1 0 9760 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_3784
timestamp 1668089732
transform 1 0 9760 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_3785
timestamp 1668089732
transform 1 0 9760 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_3786
timestamp 1668089732
transform 1 0 9760 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_3787
timestamp 1668089732
transform 1 0 9760 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_3788
timestamp 1668089732
transform 1 0 9760 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_3789
timestamp 1668089732
transform 1 0 9760 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_3790
timestamp 1668089732
transform 1 0 9760 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_3791
timestamp 1668089732
transform 1 0 9760 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_3792
timestamp 1668089732
transform 1 0 9760 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_3793
timestamp 1668089732
transform 1 0 9760 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_3794
timestamp 1668089732
transform 1 0 9760 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_3795
timestamp 1668089732
transform 1 0 9760 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_3796
timestamp 1668089732
transform 1 0 9760 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_3797
timestamp 1668089732
transform 1 0 9760 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_3798
timestamp 1668089732
transform 1 0 9760 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_3799
timestamp 1668089732
transform 1 0 9760 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_3800
timestamp 1668089732
transform 1 0 9760 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_3801
timestamp 1668089732
transform 1 0 9760 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_3802
timestamp 1668089732
transform 1 0 9760 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_3803
timestamp 1668089732
transform 1 0 9760 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_3804
timestamp 1668089732
transform 1 0 9760 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_3805
timestamp 1668089732
transform 1 0 9760 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_3806
timestamp 1668089732
transform 1 0 9760 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_3807
timestamp 1668089732
transform 1 0 9760 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_3808
timestamp 1668089732
transform 1 0 9760 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_3809
timestamp 1668089732
transform 1 0 9760 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_3810
timestamp 1668089732
transform 1 0 9760 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_3811
timestamp 1668089732
transform 1 0 9760 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_3812
timestamp 1668089732
transform 1 0 9760 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_3813
timestamp 1668089732
transform 1 0 9760 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_3814
timestamp 1668089732
transform 1 0 9760 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_3815
timestamp 1668089732
transform 1 0 9760 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_3816
timestamp 1668089732
transform 1 0 9760 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_3817
timestamp 1668089732
transform 1 0 9760 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_3818
timestamp 1668089732
transform 1 0 9760 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_3819
timestamp 1668089732
transform 1 0 9760 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_3820
timestamp 1668089732
transform 1 0 9760 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_3821
timestamp 1668089732
transform 1 0 9760 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_3822
timestamp 1668089732
transform 1 0 9760 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_3823
timestamp 1668089732
transform 1 0 9760 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_3824
timestamp 1668089732
transform 1 0 9760 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_3825
timestamp 1668089732
transform 1 0 9760 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_3826
timestamp 1668089732
transform 1 0 9760 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_3827
timestamp 1668089732
transform 1 0 9760 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_3828
timestamp 1668089732
transform 1 0 9760 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_3829
timestamp 1668089732
transform 1 0 9760 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_3830
timestamp 1668089732
transform 1 0 9760 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_3831
timestamp 1668089732
transform 1 0 9760 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_3832
timestamp 1668089732
transform 1 0 9760 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_3833
timestamp 1668089732
transform 1 0 9760 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_3834
timestamp 1668089732
transform 1 0 9760 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_3835
timestamp 1668089732
transform 1 0 9760 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_3836
timestamp 1668089732
transform 1 0 9760 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_3837
timestamp 1668089732
transform 1 0 9760 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_3838
timestamp 1668089732
transform 1 0 9760 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_3839
timestamp 1668089732
transform 1 0 9760 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_3840
timestamp 1668089732
transform 1 0 9760 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_3841
timestamp 1668089732
transform 1 0 9760 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_3842
timestamp 1668089732
transform 1 0 9760 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_3843
timestamp 1668089732
transform 1 0 9760 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_3844
timestamp 1668089732
transform 1 0 9920 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_3845
timestamp 1668089732
transform 1 0 9920 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_3846
timestamp 1668089732
transform 1 0 9920 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_3847
timestamp 1668089732
transform 1 0 9920 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_3848
timestamp 1668089732
transform 1 0 9920 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_3849
timestamp 1668089732
transform 1 0 9920 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_3850
timestamp 1668089732
transform 1 0 9920 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_3851
timestamp 1668089732
transform 1 0 9920 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_3852
timestamp 1668089732
transform 1 0 9920 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_3853
timestamp 1668089732
transform 1 0 9920 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_3854
timestamp 1668089732
transform 1 0 9920 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_3855
timestamp 1668089732
transform 1 0 9920 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_3856
timestamp 1668089732
transform 1 0 9920 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_3857
timestamp 1668089732
transform 1 0 9920 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_3858
timestamp 1668089732
transform 1 0 9920 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_3859
timestamp 1668089732
transform 1 0 9920 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_3860
timestamp 1668089732
transform 1 0 9920 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_3861
timestamp 1668089732
transform 1 0 9920 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_3862
timestamp 1668089732
transform 1 0 9920 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_3863
timestamp 1668089732
transform 1 0 9920 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_3864
timestamp 1668089732
transform 1 0 9920 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_3865
timestamp 1668089732
transform 1 0 9920 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_3866
timestamp 1668089732
transform 1 0 9920 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_3867
timestamp 1668089732
transform 1 0 9920 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_3868
timestamp 1668089732
transform 1 0 9920 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_3869
timestamp 1668089732
transform 1 0 9920 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_3870
timestamp 1668089732
transform 1 0 9920 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_3871
timestamp 1668089732
transform 1 0 9920 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_3872
timestamp 1668089732
transform 1 0 9920 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_3873
timestamp 1668089732
transform 1 0 9920 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_3874
timestamp 1668089732
transform 1 0 9920 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_3875
timestamp 1668089732
transform 1 0 9920 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_3876
timestamp 1668089732
transform 1 0 9920 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_3877
timestamp 1668089732
transform 1 0 9920 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_3878
timestamp 1668089732
transform 1 0 9920 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_3879
timestamp 1668089732
transform 1 0 9920 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_3880
timestamp 1668089732
transform 1 0 9920 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_3881
timestamp 1668089732
transform 1 0 9920 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_3882
timestamp 1668089732
transform 1 0 9920 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_3883
timestamp 1668089732
transform 1 0 9920 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_3884
timestamp 1668089732
transform 1 0 9920 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_3885
timestamp 1668089732
transform 1 0 9920 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_3886
timestamp 1668089732
transform 1 0 9920 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_3887
timestamp 1668089732
transform 1 0 9920 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_3888
timestamp 1668089732
transform 1 0 9920 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_3889
timestamp 1668089732
transform 1 0 9920 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_3890
timestamp 1668089732
transform 1 0 9920 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_3891
timestamp 1668089732
transform 1 0 9920 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_3892
timestamp 1668089732
transform 1 0 9920 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_3893
timestamp 1668089732
transform 1 0 9920 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_3894
timestamp 1668089732
transform 1 0 9920 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_3895
timestamp 1668089732
transform 1 0 9920 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_3896
timestamp 1668089732
transform 1 0 9920 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_3897
timestamp 1668089732
transform 1 0 9920 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_3898
timestamp 1668089732
transform 1 0 9920 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_3899
timestamp 1668089732
transform 1 0 9920 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_3900
timestamp 1668089732
transform 1 0 9920 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_3901
timestamp 1668089732
transform 1 0 9920 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_3902
timestamp 1668089732
transform 1 0 9920 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_3903
timestamp 1668089732
transform 1 0 9920 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_3904
timestamp 1668089732
transform 1 0 9920 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_3905
timestamp 1668089732
transform 1 0 9920 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_3906
timestamp 1668089732
transform 1 0 10080 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_3907
timestamp 1668089732
transform 1 0 10080 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_3908
timestamp 1668089732
transform 1 0 10080 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_3909
timestamp 1668089732
transform 1 0 10080 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_3910
timestamp 1668089732
transform 1 0 10080 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_3911
timestamp 1668089732
transform 1 0 10080 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_3912
timestamp 1668089732
transform 1 0 10080 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_3913
timestamp 1668089732
transform 1 0 10080 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_3914
timestamp 1668089732
transform 1 0 10080 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_3915
timestamp 1668089732
transform 1 0 10080 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_3916
timestamp 1668089732
transform 1 0 10080 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_3917
timestamp 1668089732
transform 1 0 10080 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_3918
timestamp 1668089732
transform 1 0 10080 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_3919
timestamp 1668089732
transform 1 0 10080 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_3920
timestamp 1668089732
transform 1 0 10080 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_3921
timestamp 1668089732
transform 1 0 10080 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_3922
timestamp 1668089732
transform 1 0 10080 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_3923
timestamp 1668089732
transform 1 0 10080 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_3924
timestamp 1668089732
transform 1 0 10080 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_3925
timestamp 1668089732
transform 1 0 10080 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_3926
timestamp 1668089732
transform 1 0 10080 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_3927
timestamp 1668089732
transform 1 0 10080 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_3928
timestamp 1668089732
transform 1 0 10080 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_3929
timestamp 1668089732
transform 1 0 10080 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_3930
timestamp 1668089732
transform 1 0 10080 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_3931
timestamp 1668089732
transform 1 0 10080 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_3932
timestamp 1668089732
transform 1 0 10080 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_3933
timestamp 1668089732
transform 1 0 10080 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_3934
timestamp 1668089732
transform 1 0 10080 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_3935
timestamp 1668089732
transform 1 0 10080 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_3936
timestamp 1668089732
transform 1 0 10080 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_3937
timestamp 1668089732
transform 1 0 10080 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_3938
timestamp 1668089732
transform 1 0 10080 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_3939
timestamp 1668089732
transform 1 0 10080 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_3940
timestamp 1668089732
transform 1 0 10080 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_3941
timestamp 1668089732
transform 1 0 10080 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_3942
timestamp 1668089732
transform 1 0 10080 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_3943
timestamp 1668089732
transform 1 0 10080 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_3944
timestamp 1668089732
transform 1 0 10080 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_3945
timestamp 1668089732
transform 1 0 10080 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_3946
timestamp 1668089732
transform 1 0 10080 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_3947
timestamp 1668089732
transform 1 0 10080 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_3948
timestamp 1668089732
transform 1 0 10080 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_3949
timestamp 1668089732
transform 1 0 10080 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_3950
timestamp 1668089732
transform 1 0 10080 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_3951
timestamp 1668089732
transform 1 0 10080 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_3952
timestamp 1668089732
transform 1 0 10080 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_3953
timestamp 1668089732
transform 1 0 10080 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_3954
timestamp 1668089732
transform 1 0 10080 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_3955
timestamp 1668089732
transform 1 0 10080 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_3956
timestamp 1668089732
transform 1 0 10080 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_3957
timestamp 1668089732
transform 1 0 10080 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_3958
timestamp 1668089732
transform 1 0 10080 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_3959
timestamp 1668089732
transform 1 0 10080 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_3960
timestamp 1668089732
transform 1 0 10080 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_3961
timestamp 1668089732
transform 1 0 10080 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_3962
timestamp 1668089732
transform 1 0 10080 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_3963
timestamp 1668089732
transform 1 0 10080 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_3964
timestamp 1668089732
transform 1 0 10080 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_3965
timestamp 1668089732
transform 1 0 10080 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_3966
timestamp 1668089732
transform 1 0 10080 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_3967
timestamp 1668089732
transform 1 0 10080 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_3968
timestamp 1668089732
transform 1 0 10240 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_3969
timestamp 1668089732
transform 1 0 10240 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_3970
timestamp 1668089732
transform 1 0 10240 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_3971
timestamp 1668089732
transform 1 0 10240 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_3972
timestamp 1668089732
transform 1 0 10240 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_3973
timestamp 1668089732
transform 1 0 10240 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_3974
timestamp 1668089732
transform 1 0 10240 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_3975
timestamp 1668089732
transform 1 0 10240 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_3976
timestamp 1668089732
transform 1 0 10240 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_3977
timestamp 1668089732
transform 1 0 10240 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_3978
timestamp 1668089732
transform 1 0 10240 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_3979
timestamp 1668089732
transform 1 0 10240 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_3980
timestamp 1668089732
transform 1 0 10240 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_3981
timestamp 1668089732
transform 1 0 10240 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_3982
timestamp 1668089732
transform 1 0 10240 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_3983
timestamp 1668089732
transform 1 0 10240 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_3984
timestamp 1668089732
transform 1 0 10240 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_3985
timestamp 1668089732
transform 1 0 10240 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_3986
timestamp 1668089732
transform 1 0 10240 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_3987
timestamp 1668089732
transform 1 0 10240 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_3988
timestamp 1668089732
transform 1 0 10240 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_3989
timestamp 1668089732
transform 1 0 10240 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_3990
timestamp 1668089732
transform 1 0 10240 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_3991
timestamp 1668089732
transform 1 0 10240 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_3992
timestamp 1668089732
transform 1 0 10240 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_3993
timestamp 1668089732
transform 1 0 10240 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_3994
timestamp 1668089732
transform 1 0 10240 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_3995
timestamp 1668089732
transform 1 0 10240 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_3996
timestamp 1668089732
transform 1 0 10240 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_3997
timestamp 1668089732
transform 1 0 10240 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_3998
timestamp 1668089732
transform 1 0 10240 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_3999
timestamp 1668089732
transform 1 0 10240 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_4000
timestamp 1668089732
transform 1 0 10240 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_4001
timestamp 1668089732
transform 1 0 10240 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_4002
timestamp 1668089732
transform 1 0 10240 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_4003
timestamp 1668089732
transform 1 0 10240 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_4004
timestamp 1668089732
transform 1 0 10240 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_4005
timestamp 1668089732
transform 1 0 10240 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_4006
timestamp 1668089732
transform 1 0 10240 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_4007
timestamp 1668089732
transform 1 0 10240 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_4008
timestamp 1668089732
transform 1 0 10240 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_4009
timestamp 1668089732
transform 1 0 10240 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_4010
timestamp 1668089732
transform 1 0 10240 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_4011
timestamp 1668089732
transform 1 0 10240 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_4012
timestamp 1668089732
transform 1 0 10240 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_4013
timestamp 1668089732
transform 1 0 10240 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_4014
timestamp 1668089732
transform 1 0 10240 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_4015
timestamp 1668089732
transform 1 0 10240 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_4016
timestamp 1668089732
transform 1 0 10240 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_4017
timestamp 1668089732
transform 1 0 10240 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_4018
timestamp 1668089732
transform 1 0 10240 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_4019
timestamp 1668089732
transform 1 0 10240 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_4020
timestamp 1668089732
transform 1 0 10240 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_4021
timestamp 1668089732
transform 1 0 10240 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_4022
timestamp 1668089732
transform 1 0 10240 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_4023
timestamp 1668089732
transform 1 0 10240 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_4024
timestamp 1668089732
transform 1 0 10240 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_4025
timestamp 1668089732
transform 1 0 10240 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_4026
timestamp 1668089732
transform 1 0 10240 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_4027
timestamp 1668089732
transform 1 0 10240 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_4028
timestamp 1668089732
transform 1 0 10240 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_4029
timestamp 1668089732
transform 1 0 10240 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_4030
timestamp 1668089732
transform 1 0 10400 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_4031
timestamp 1668089732
transform 1 0 10400 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_4032
timestamp 1668089732
transform 1 0 10400 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_4033
timestamp 1668089732
transform 1 0 10400 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_4034
timestamp 1668089732
transform 1 0 10400 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_4035
timestamp 1668089732
transform 1 0 10400 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_4036
timestamp 1668089732
transform 1 0 10400 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_4037
timestamp 1668089732
transform 1 0 10400 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_4038
timestamp 1668089732
transform 1 0 10400 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_4039
timestamp 1668089732
transform 1 0 10400 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_4040
timestamp 1668089732
transform 1 0 10400 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_4041
timestamp 1668089732
transform 1 0 10400 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_4042
timestamp 1668089732
transform 1 0 10400 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_4043
timestamp 1668089732
transform 1 0 10400 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_4044
timestamp 1668089732
transform 1 0 10400 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_4045
timestamp 1668089732
transform 1 0 10400 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_4046
timestamp 1668089732
transform 1 0 10400 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_4047
timestamp 1668089732
transform 1 0 10400 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_4048
timestamp 1668089732
transform 1 0 10400 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_4049
timestamp 1668089732
transform 1 0 10400 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_4050
timestamp 1668089732
transform 1 0 10400 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_4051
timestamp 1668089732
transform 1 0 10400 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_4052
timestamp 1668089732
transform 1 0 10400 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_4053
timestamp 1668089732
transform 1 0 10400 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_4054
timestamp 1668089732
transform 1 0 10400 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_4055
timestamp 1668089732
transform 1 0 10400 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_4056
timestamp 1668089732
transform 1 0 10400 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_4057
timestamp 1668089732
transform 1 0 10400 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_4058
timestamp 1668089732
transform 1 0 10400 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_4059
timestamp 1668089732
transform 1 0 10400 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_4060
timestamp 1668089732
transform 1 0 10400 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_4061
timestamp 1668089732
transform 1 0 10400 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_4062
timestamp 1668089732
transform 1 0 10400 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_4063
timestamp 1668089732
transform 1 0 10400 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_4064
timestamp 1668089732
transform 1 0 10400 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_4065
timestamp 1668089732
transform 1 0 10400 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_4066
timestamp 1668089732
transform 1 0 10400 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_4067
timestamp 1668089732
transform 1 0 10400 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_4068
timestamp 1668089732
transform 1 0 10400 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_4069
timestamp 1668089732
transform 1 0 10400 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_4070
timestamp 1668089732
transform 1 0 10400 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_4071
timestamp 1668089732
transform 1 0 10400 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_4072
timestamp 1668089732
transform 1 0 10400 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_4073
timestamp 1668089732
transform 1 0 10400 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_4074
timestamp 1668089732
transform 1 0 10400 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_4075
timestamp 1668089732
transform 1 0 10400 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_4076
timestamp 1668089732
transform 1 0 10400 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_4077
timestamp 1668089732
transform 1 0 10400 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_4078
timestamp 1668089732
transform 1 0 10400 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_4079
timestamp 1668089732
transform 1 0 10400 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_4080
timestamp 1668089732
transform 1 0 10400 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_4081
timestamp 1668089732
transform 1 0 10400 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_4082
timestamp 1668089732
transform 1 0 10400 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_4083
timestamp 1668089732
transform 1 0 10400 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_4084
timestamp 1668089732
transform 1 0 10400 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_4085
timestamp 1668089732
transform 1 0 10400 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_4086
timestamp 1668089732
transform 1 0 10400 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_4087
timestamp 1668089732
transform 1 0 10400 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_4088
timestamp 1668089732
transform 1 0 10400 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_4089
timestamp 1668089732
transform 1 0 10400 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_4090
timestamp 1668089732
transform 1 0 10400 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_4091
timestamp 1668089732
transform 1 0 10400 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_4092
timestamp 1668089732
transform 1 0 10560 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_4093
timestamp 1668089732
transform 1 0 10560 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_4094
timestamp 1668089732
transform 1 0 10560 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_4095
timestamp 1668089732
transform 1 0 10560 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_4096
timestamp 1668089732
transform 1 0 10560 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_4097
timestamp 1668089732
transform 1 0 10560 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_4098
timestamp 1668089732
transform 1 0 10560 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_4099
timestamp 1668089732
transform 1 0 10560 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_4100
timestamp 1668089732
transform 1 0 10560 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_4101
timestamp 1668089732
transform 1 0 10560 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_4102
timestamp 1668089732
transform 1 0 10560 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_4103
timestamp 1668089732
transform 1 0 10560 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_4104
timestamp 1668089732
transform 1 0 10560 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_4105
timestamp 1668089732
transform 1 0 10560 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_4106
timestamp 1668089732
transform 1 0 10560 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_4107
timestamp 1668089732
transform 1 0 10560 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_4108
timestamp 1668089732
transform 1 0 10560 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_4109
timestamp 1668089732
transform 1 0 10560 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_4110
timestamp 1668089732
transform 1 0 10560 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_4111
timestamp 1668089732
transform 1 0 10560 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_4112
timestamp 1668089732
transform 1 0 10560 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_4113
timestamp 1668089732
transform 1 0 10560 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_4114
timestamp 1668089732
transform 1 0 10560 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_4115
timestamp 1668089732
transform 1 0 10560 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_4116
timestamp 1668089732
transform 1 0 10560 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_4117
timestamp 1668089732
transform 1 0 10560 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_4118
timestamp 1668089732
transform 1 0 10560 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_4119
timestamp 1668089732
transform 1 0 10560 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_4120
timestamp 1668089732
transform 1 0 10560 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_4121
timestamp 1668089732
transform 1 0 10560 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_4122
timestamp 1668089732
transform 1 0 10560 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_4123
timestamp 1668089732
transform 1 0 10560 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_4124
timestamp 1668089732
transform 1 0 10560 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_4125
timestamp 1668089732
transform 1 0 10560 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_4126
timestamp 1668089732
transform 1 0 10560 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_4127
timestamp 1668089732
transform 1 0 10560 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_4128
timestamp 1668089732
transform 1 0 10560 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_4129
timestamp 1668089732
transform 1 0 10560 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_4130
timestamp 1668089732
transform 1 0 10560 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_4131
timestamp 1668089732
transform 1 0 10560 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_4132
timestamp 1668089732
transform 1 0 10560 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_4133
timestamp 1668089732
transform 1 0 10560 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_4134
timestamp 1668089732
transform 1 0 10560 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_4135
timestamp 1668089732
transform 1 0 10560 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_4136
timestamp 1668089732
transform 1 0 10560 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_4137
timestamp 1668089732
transform 1 0 10560 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_4138
timestamp 1668089732
transform 1 0 10560 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_4139
timestamp 1668089732
transform 1 0 10560 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_4140
timestamp 1668089732
transform 1 0 10560 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_4141
timestamp 1668089732
transform 1 0 10560 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_4142
timestamp 1668089732
transform 1 0 10560 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_4143
timestamp 1668089732
transform 1 0 10560 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_4144
timestamp 1668089732
transform 1 0 10560 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_4145
timestamp 1668089732
transform 1 0 10560 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_4146
timestamp 1668089732
transform 1 0 10560 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_4147
timestamp 1668089732
transform 1 0 10560 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_4148
timestamp 1668089732
transform 1 0 10560 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_4149
timestamp 1668089732
transform 1 0 10560 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_4150
timestamp 1668089732
transform 1 0 10560 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_4151
timestamp 1668089732
transform 1 0 10560 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_4152
timestamp 1668089732
transform 1 0 10560 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_4153
timestamp 1668089732
transform 1 0 10560 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_4154
timestamp 1668089732
transform 1 0 10720 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_4155
timestamp 1668089732
transform 1 0 10720 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_4156
timestamp 1668089732
transform 1 0 10720 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_4157
timestamp 1668089732
transform 1 0 10720 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_4158
timestamp 1668089732
transform 1 0 10720 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_4159
timestamp 1668089732
transform 1 0 10720 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_4160
timestamp 1668089732
transform 1 0 10720 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_4161
timestamp 1668089732
transform 1 0 10720 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_4162
timestamp 1668089732
transform 1 0 10720 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_4163
timestamp 1668089732
transform 1 0 10720 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_4164
timestamp 1668089732
transform 1 0 10720 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_4165
timestamp 1668089732
transform 1 0 10720 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_4166
timestamp 1668089732
transform 1 0 10720 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_4167
timestamp 1668089732
transform 1 0 10720 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_4168
timestamp 1668089732
transform 1 0 10720 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_4169
timestamp 1668089732
transform 1 0 10720 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_4170
timestamp 1668089732
transform 1 0 10720 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_4171
timestamp 1668089732
transform 1 0 10720 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_4172
timestamp 1668089732
transform 1 0 10720 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_4173
timestamp 1668089732
transform 1 0 10720 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_4174
timestamp 1668089732
transform 1 0 10720 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_4175
timestamp 1668089732
transform 1 0 10720 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_4176
timestamp 1668089732
transform 1 0 10720 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_4177
timestamp 1668089732
transform 1 0 10720 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_4178
timestamp 1668089732
transform 1 0 10720 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_4179
timestamp 1668089732
transform 1 0 10720 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_4180
timestamp 1668089732
transform 1 0 10720 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_4181
timestamp 1668089732
transform 1 0 10720 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_4182
timestamp 1668089732
transform 1 0 10720 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_4183
timestamp 1668089732
transform 1 0 10720 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_4184
timestamp 1668089732
transform 1 0 10720 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_4185
timestamp 1668089732
transform 1 0 10720 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_4186
timestamp 1668089732
transform 1 0 10720 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_4187
timestamp 1668089732
transform 1 0 10720 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_4188
timestamp 1668089732
transform 1 0 10720 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_4189
timestamp 1668089732
transform 1 0 10720 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_4190
timestamp 1668089732
transform 1 0 10720 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_4191
timestamp 1668089732
transform 1 0 10720 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_4192
timestamp 1668089732
transform 1 0 10720 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_4193
timestamp 1668089732
transform 1 0 10720 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_4194
timestamp 1668089732
transform 1 0 10720 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_4195
timestamp 1668089732
transform 1 0 10720 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_4196
timestamp 1668089732
transform 1 0 10720 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_4197
timestamp 1668089732
transform 1 0 10720 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_4198
timestamp 1668089732
transform 1 0 10720 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_4199
timestamp 1668089732
transform 1 0 10720 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_4200
timestamp 1668089732
transform 1 0 10720 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_4201
timestamp 1668089732
transform 1 0 10720 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_4202
timestamp 1668089732
transform 1 0 10720 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_4203
timestamp 1668089732
transform 1 0 10720 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_4204
timestamp 1668089732
transform 1 0 10720 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_4205
timestamp 1668089732
transform 1 0 10720 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_4206
timestamp 1668089732
transform 1 0 10720 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_4207
timestamp 1668089732
transform 1 0 10720 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_4208
timestamp 1668089732
transform 1 0 10720 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_4209
timestamp 1668089732
transform 1 0 10720 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_4210
timestamp 1668089732
transform 1 0 10720 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_4211
timestamp 1668089732
transform 1 0 10720 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_4212
timestamp 1668089732
transform 1 0 10720 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_4213
timestamp 1668089732
transform 1 0 10720 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_4214
timestamp 1668089732
transform 1 0 10720 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_4215
timestamp 1668089732
transform 1 0 10720 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_4216
timestamp 1668089732
transform 1 0 10880 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_4217
timestamp 1668089732
transform 1 0 10880 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_4218
timestamp 1668089732
transform 1 0 10880 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_4219
timestamp 1668089732
transform 1 0 10880 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_4220
timestamp 1668089732
transform 1 0 10880 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_4221
timestamp 1668089732
transform 1 0 10880 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_4222
timestamp 1668089732
transform 1 0 10880 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_4223
timestamp 1668089732
transform 1 0 10880 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_4224
timestamp 1668089732
transform 1 0 10880 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_4225
timestamp 1668089732
transform 1 0 10880 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_4226
timestamp 1668089732
transform 1 0 10880 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_4227
timestamp 1668089732
transform 1 0 10880 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_4228
timestamp 1668089732
transform 1 0 10880 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_4229
timestamp 1668089732
transform 1 0 10880 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_4230
timestamp 1668089732
transform 1 0 10880 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_4231
timestamp 1668089732
transform 1 0 10880 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_4232
timestamp 1668089732
transform 1 0 10880 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_4233
timestamp 1668089732
transform 1 0 10880 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_4234
timestamp 1668089732
transform 1 0 10880 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_4235
timestamp 1668089732
transform 1 0 10880 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_4236
timestamp 1668089732
transform 1 0 10880 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_4237
timestamp 1668089732
transform 1 0 10880 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_4238
timestamp 1668089732
transform 1 0 10880 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_4239
timestamp 1668089732
transform 1 0 10880 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_4240
timestamp 1668089732
transform 1 0 10880 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_4241
timestamp 1668089732
transform 1 0 10880 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_4242
timestamp 1668089732
transform 1 0 10880 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_4243
timestamp 1668089732
transform 1 0 10880 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_4244
timestamp 1668089732
transform 1 0 10880 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_4245
timestamp 1668089732
transform 1 0 10880 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_4246
timestamp 1668089732
transform 1 0 10880 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_4247
timestamp 1668089732
transform 1 0 10880 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_4248
timestamp 1668089732
transform 1 0 10880 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_4249
timestamp 1668089732
transform 1 0 10880 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_4250
timestamp 1668089732
transform 1 0 10880 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_4251
timestamp 1668089732
transform 1 0 10880 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_4252
timestamp 1668089732
transform 1 0 10880 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_4253
timestamp 1668089732
transform 1 0 10880 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_4254
timestamp 1668089732
transform 1 0 10880 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_4255
timestamp 1668089732
transform 1 0 10880 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_4256
timestamp 1668089732
transform 1 0 10880 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_4257
timestamp 1668089732
transform 1 0 10880 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_4258
timestamp 1668089732
transform 1 0 10880 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_4259
timestamp 1668089732
transform 1 0 10880 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_4260
timestamp 1668089732
transform 1 0 10880 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_4261
timestamp 1668089732
transform 1 0 10880 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_4262
timestamp 1668089732
transform 1 0 10880 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_4263
timestamp 1668089732
transform 1 0 10880 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_4264
timestamp 1668089732
transform 1 0 10880 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_4265
timestamp 1668089732
transform 1 0 10880 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_4266
timestamp 1668089732
transform 1 0 10880 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_4267
timestamp 1668089732
transform 1 0 10880 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_4268
timestamp 1668089732
transform 1 0 10880 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_4269
timestamp 1668089732
transform 1 0 10880 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_4270
timestamp 1668089732
transform 1 0 10880 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_4271
timestamp 1668089732
transform 1 0 10880 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_4272
timestamp 1668089732
transform 1 0 10880 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_4273
timestamp 1668089732
transform 1 0 10880 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_4274
timestamp 1668089732
transform 1 0 10880 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_4275
timestamp 1668089732
transform 1 0 10880 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_4276
timestamp 1668089732
transform 1 0 10880 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_4277
timestamp 1668089732
transform 1 0 10880 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_4278
timestamp 1668089732
transform 1 0 11040 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_4279
timestamp 1668089732
transform 1 0 11040 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_4280
timestamp 1668089732
transform 1 0 11040 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_4281
timestamp 1668089732
transform 1 0 11040 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_4282
timestamp 1668089732
transform 1 0 11040 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_4283
timestamp 1668089732
transform 1 0 11040 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_4284
timestamp 1668089732
transform 1 0 11040 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_4285
timestamp 1668089732
transform 1 0 11040 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_4286
timestamp 1668089732
transform 1 0 11040 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_4287
timestamp 1668089732
transform 1 0 11040 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_4288
timestamp 1668089732
transform 1 0 11040 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_4289
timestamp 1668089732
transform 1 0 11040 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_4290
timestamp 1668089732
transform 1 0 11040 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_4291
timestamp 1668089732
transform 1 0 11040 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_4292
timestamp 1668089732
transform 1 0 11040 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_4293
timestamp 1668089732
transform 1 0 11040 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_4294
timestamp 1668089732
transform 1 0 11040 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_4295
timestamp 1668089732
transform 1 0 11040 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_4296
timestamp 1668089732
transform 1 0 11040 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_4297
timestamp 1668089732
transform 1 0 11040 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_4298
timestamp 1668089732
transform 1 0 11040 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_4299
timestamp 1668089732
transform 1 0 11040 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_4300
timestamp 1668089732
transform 1 0 11040 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_4301
timestamp 1668089732
transform 1 0 11040 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_4302
timestamp 1668089732
transform 1 0 11040 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_4303
timestamp 1668089732
transform 1 0 11040 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_4304
timestamp 1668089732
transform 1 0 11040 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_4305
timestamp 1668089732
transform 1 0 11040 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_4306
timestamp 1668089732
transform 1 0 11040 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_4307
timestamp 1668089732
transform 1 0 11040 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_4308
timestamp 1668089732
transform 1 0 11040 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_4309
timestamp 1668089732
transform 1 0 11040 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_4310
timestamp 1668089732
transform 1 0 11040 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_4311
timestamp 1668089732
transform 1 0 11040 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_4312
timestamp 1668089732
transform 1 0 11040 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_4313
timestamp 1668089732
transform 1 0 11040 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_4314
timestamp 1668089732
transform 1 0 11040 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_4315
timestamp 1668089732
transform 1 0 11040 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_4316
timestamp 1668089732
transform 1 0 11040 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_4317
timestamp 1668089732
transform 1 0 11040 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_4318
timestamp 1668089732
transform 1 0 11040 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_4319
timestamp 1668089732
transform 1 0 11040 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_4320
timestamp 1668089732
transform 1 0 11040 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_4321
timestamp 1668089732
transform 1 0 11040 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_4322
timestamp 1668089732
transform 1 0 11040 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_4323
timestamp 1668089732
transform 1 0 11040 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_4324
timestamp 1668089732
transform 1 0 11040 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_4325
timestamp 1668089732
transform 1 0 11040 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_4326
timestamp 1668089732
transform 1 0 11040 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_4327
timestamp 1668089732
transform 1 0 11040 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_4328
timestamp 1668089732
transform 1 0 11040 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_4329
timestamp 1668089732
transform 1 0 11040 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_4330
timestamp 1668089732
transform 1 0 11040 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_4331
timestamp 1668089732
transform 1 0 11040 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_4332
timestamp 1668089732
transform 1 0 11040 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_4333
timestamp 1668089732
transform 1 0 11040 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_4334
timestamp 1668089732
transform 1 0 11040 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_4335
timestamp 1668089732
transform 1 0 11040 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_4336
timestamp 1668089732
transform 1 0 11040 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_4337
timestamp 1668089732
transform 1 0 11040 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_4338
timestamp 1668089732
transform 1 0 11040 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_4339
timestamp 1668089732
transform 1 0 11040 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_4340
timestamp 1668089732
transform 1 0 11200 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_4341
timestamp 1668089732
transform 1 0 11200 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_4342
timestamp 1668089732
transform 1 0 11200 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_4343
timestamp 1668089732
transform 1 0 11200 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_4344
timestamp 1668089732
transform 1 0 11200 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_4345
timestamp 1668089732
transform 1 0 11200 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_4346
timestamp 1668089732
transform 1 0 11200 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_4347
timestamp 1668089732
transform 1 0 11200 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_4348
timestamp 1668089732
transform 1 0 11200 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_4349
timestamp 1668089732
transform 1 0 11200 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_4350
timestamp 1668089732
transform 1 0 11200 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_4351
timestamp 1668089732
transform 1 0 11200 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_4352
timestamp 1668089732
transform 1 0 11200 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_4353
timestamp 1668089732
transform 1 0 11200 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_4354
timestamp 1668089732
transform 1 0 11200 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_4355
timestamp 1668089732
transform 1 0 11200 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_4356
timestamp 1668089732
transform 1 0 11200 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_4357
timestamp 1668089732
transform 1 0 11200 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_4358
timestamp 1668089732
transform 1 0 11200 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_4359
timestamp 1668089732
transform 1 0 11200 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_4360
timestamp 1668089732
transform 1 0 11200 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_4361
timestamp 1668089732
transform 1 0 11200 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_4362
timestamp 1668089732
transform 1 0 11200 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_4363
timestamp 1668089732
transform 1 0 11200 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_4364
timestamp 1668089732
transform 1 0 11200 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_4365
timestamp 1668089732
transform 1 0 11200 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_4366
timestamp 1668089732
transform 1 0 11200 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_4367
timestamp 1668089732
transform 1 0 11200 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_4368
timestamp 1668089732
transform 1 0 11200 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_4369
timestamp 1668089732
transform 1 0 11200 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_4370
timestamp 1668089732
transform 1 0 11200 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_4371
timestamp 1668089732
transform 1 0 11200 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_4372
timestamp 1668089732
transform 1 0 11200 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_4373
timestamp 1668089732
transform 1 0 11200 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_4374
timestamp 1668089732
transform 1 0 11200 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_4375
timestamp 1668089732
transform 1 0 11200 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_4376
timestamp 1668089732
transform 1 0 11200 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_4377
timestamp 1668089732
transform 1 0 11200 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_4378
timestamp 1668089732
transform 1 0 11200 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_4379
timestamp 1668089732
transform 1 0 11200 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_4380
timestamp 1668089732
transform 1 0 11200 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_4381
timestamp 1668089732
transform 1 0 11200 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_4382
timestamp 1668089732
transform 1 0 11200 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_4383
timestamp 1668089732
transform 1 0 11200 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_4384
timestamp 1668089732
transform 1 0 11200 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_4385
timestamp 1668089732
transform 1 0 11200 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_4386
timestamp 1668089732
transform 1 0 11200 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_4387
timestamp 1668089732
transform 1 0 11200 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_4388
timestamp 1668089732
transform 1 0 11200 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_4389
timestamp 1668089732
transform 1 0 11200 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_4390
timestamp 1668089732
transform 1 0 11200 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_4391
timestamp 1668089732
transform 1 0 11200 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_4392
timestamp 1668089732
transform 1 0 11200 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_4393
timestamp 1668089732
transform 1 0 11200 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_4394
timestamp 1668089732
transform 1 0 11200 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_4395
timestamp 1668089732
transform 1 0 11200 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_4396
timestamp 1668089732
transform 1 0 11200 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_4397
timestamp 1668089732
transform 1 0 11200 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_4398
timestamp 1668089732
transform 1 0 11200 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_4399
timestamp 1668089732
transform 1 0 11200 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_4400
timestamp 1668089732
transform 1 0 11200 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_4401
timestamp 1668089732
transform 1 0 11200 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_4402
timestamp 1668089732
transform 1 0 11360 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_4403
timestamp 1668089732
transform 1 0 11360 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_4404
timestamp 1668089732
transform 1 0 11360 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_4405
timestamp 1668089732
transform 1 0 11360 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_4406
timestamp 1668089732
transform 1 0 11360 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_4407
timestamp 1668089732
transform 1 0 11360 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_4408
timestamp 1668089732
transform 1 0 11360 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_4409
timestamp 1668089732
transform 1 0 11360 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_4410
timestamp 1668089732
transform 1 0 11360 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_4411
timestamp 1668089732
transform 1 0 11360 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_4412
timestamp 1668089732
transform 1 0 11360 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_4413
timestamp 1668089732
transform 1 0 11360 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_4414
timestamp 1668089732
transform 1 0 11360 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_4415
timestamp 1668089732
transform 1 0 11360 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_4416
timestamp 1668089732
transform 1 0 11360 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_4417
timestamp 1668089732
transform 1 0 11360 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_4418
timestamp 1668089732
transform 1 0 11360 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_4419
timestamp 1668089732
transform 1 0 11360 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_4420
timestamp 1668089732
transform 1 0 11360 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_4421
timestamp 1668089732
transform 1 0 11360 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_4422
timestamp 1668089732
transform 1 0 11360 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_4423
timestamp 1668089732
transform 1 0 11360 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_4424
timestamp 1668089732
transform 1 0 11360 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_4425
timestamp 1668089732
transform 1 0 11360 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_4426
timestamp 1668089732
transform 1 0 11360 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_4427
timestamp 1668089732
transform 1 0 11360 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_4428
timestamp 1668089732
transform 1 0 11360 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_4429
timestamp 1668089732
transform 1 0 11360 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_4430
timestamp 1668089732
transform 1 0 11360 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_4431
timestamp 1668089732
transform 1 0 11360 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_4432
timestamp 1668089732
transform 1 0 11360 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_4433
timestamp 1668089732
transform 1 0 11360 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_4434
timestamp 1668089732
transform 1 0 11360 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_4435
timestamp 1668089732
transform 1 0 11360 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_4436
timestamp 1668089732
transform 1 0 11360 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_4437
timestamp 1668089732
transform 1 0 11360 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_4438
timestamp 1668089732
transform 1 0 11360 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_4439
timestamp 1668089732
transform 1 0 11360 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_4440
timestamp 1668089732
transform 1 0 11360 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_4441
timestamp 1668089732
transform 1 0 11360 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_4442
timestamp 1668089732
transform 1 0 11360 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_4443
timestamp 1668089732
transform 1 0 11360 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_4444
timestamp 1668089732
transform 1 0 11360 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_4445
timestamp 1668089732
transform 1 0 11360 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_4446
timestamp 1668089732
transform 1 0 11360 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_4447
timestamp 1668089732
transform 1 0 11360 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_4448
timestamp 1668089732
transform 1 0 11360 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_4449
timestamp 1668089732
transform 1 0 11360 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_4450
timestamp 1668089732
transform 1 0 11360 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_4451
timestamp 1668089732
transform 1 0 11360 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_4452
timestamp 1668089732
transform 1 0 11360 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_4453
timestamp 1668089732
transform 1 0 11360 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_4454
timestamp 1668089732
transform 1 0 11360 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_4455
timestamp 1668089732
transform 1 0 11360 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_4456
timestamp 1668089732
transform 1 0 11360 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_4457
timestamp 1668089732
transform 1 0 11360 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_4458
timestamp 1668089732
transform 1 0 11360 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_4459
timestamp 1668089732
transform 1 0 11360 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_4460
timestamp 1668089732
transform 1 0 11360 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_4461
timestamp 1668089732
transform 1 0 11360 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_4462
timestamp 1668089732
transform 1 0 11360 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_4463
timestamp 1668089732
transform 1 0 11360 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_4464
timestamp 1668089732
transform 1 0 11520 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_4465
timestamp 1668089732
transform 1 0 11520 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_4466
timestamp 1668089732
transform 1 0 11520 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_4467
timestamp 1668089732
transform 1 0 11520 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_4468
timestamp 1668089732
transform 1 0 11520 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_4469
timestamp 1668089732
transform 1 0 11520 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_4470
timestamp 1668089732
transform 1 0 11520 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_4471
timestamp 1668089732
transform 1 0 11520 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_4472
timestamp 1668089732
transform 1 0 11520 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_4473
timestamp 1668089732
transform 1 0 11520 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_4474
timestamp 1668089732
transform 1 0 11520 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_4475
timestamp 1668089732
transform 1 0 11520 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_4476
timestamp 1668089732
transform 1 0 11520 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_4477
timestamp 1668089732
transform 1 0 11520 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_4478
timestamp 1668089732
transform 1 0 11520 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_4479
timestamp 1668089732
transform 1 0 11520 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_4480
timestamp 1668089732
transform 1 0 11520 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_4481
timestamp 1668089732
transform 1 0 11520 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_4482
timestamp 1668089732
transform 1 0 11520 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_4483
timestamp 1668089732
transform 1 0 11520 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_4484
timestamp 1668089732
transform 1 0 11520 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_4485
timestamp 1668089732
transform 1 0 11520 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_4486
timestamp 1668089732
transform 1 0 11520 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_4487
timestamp 1668089732
transform 1 0 11520 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_4488
timestamp 1668089732
transform 1 0 11520 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_4489
timestamp 1668089732
transform 1 0 11520 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_4490
timestamp 1668089732
transform 1 0 11520 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_4491
timestamp 1668089732
transform 1 0 11520 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_4492
timestamp 1668089732
transform 1 0 11520 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_4493
timestamp 1668089732
transform 1 0 11520 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_4494
timestamp 1668089732
transform 1 0 11520 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_4495
timestamp 1668089732
transform 1 0 11520 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_4496
timestamp 1668089732
transform 1 0 11520 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_4497
timestamp 1668089732
transform 1 0 11520 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_4498
timestamp 1668089732
transform 1 0 11520 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_4499
timestamp 1668089732
transform 1 0 11520 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_4500
timestamp 1668089732
transform 1 0 11520 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_4501
timestamp 1668089732
transform 1 0 11520 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_4502
timestamp 1668089732
transform 1 0 11520 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_4503
timestamp 1668089732
transform 1 0 11520 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_4504
timestamp 1668089732
transform 1 0 11520 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_4505
timestamp 1668089732
transform 1 0 11520 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_4506
timestamp 1668089732
transform 1 0 11520 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_4507
timestamp 1668089732
transform 1 0 11520 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_4508
timestamp 1668089732
transform 1 0 11520 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_4509
timestamp 1668089732
transform 1 0 11520 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_4510
timestamp 1668089732
transform 1 0 11520 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_4511
timestamp 1668089732
transform 1 0 11520 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_4512
timestamp 1668089732
transform 1 0 11520 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_4513
timestamp 1668089732
transform 1 0 11520 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_4514
timestamp 1668089732
transform 1 0 11520 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_4515
timestamp 1668089732
transform 1 0 11520 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_4516
timestamp 1668089732
transform 1 0 11520 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_4517
timestamp 1668089732
transform 1 0 11520 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_4518
timestamp 1668089732
transform 1 0 11520 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_4519
timestamp 1668089732
transform 1 0 11520 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_4520
timestamp 1668089732
transform 1 0 11520 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_4521
timestamp 1668089732
transform 1 0 11520 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_4522
timestamp 1668089732
transform 1 0 11520 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_4523
timestamp 1668089732
transform 1 0 11520 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_4524
timestamp 1668089732
transform 1 0 11520 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_4525
timestamp 1668089732
transform 1 0 11520 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_4526
timestamp 1668089732
transform 1 0 11680 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_4527
timestamp 1668089732
transform 1 0 11680 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_4528
timestamp 1668089732
transform 1 0 11680 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_4529
timestamp 1668089732
transform 1 0 11680 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_4530
timestamp 1668089732
transform 1 0 11680 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_4531
timestamp 1668089732
transform 1 0 11680 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_4532
timestamp 1668089732
transform 1 0 11680 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_4533
timestamp 1668089732
transform 1 0 11680 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_4534
timestamp 1668089732
transform 1 0 11680 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_4535
timestamp 1668089732
transform 1 0 11680 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_4536
timestamp 1668089732
transform 1 0 11680 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_4537
timestamp 1668089732
transform 1 0 11680 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_4538
timestamp 1668089732
transform 1 0 11680 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_4539
timestamp 1668089732
transform 1 0 11680 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_4540
timestamp 1668089732
transform 1 0 11680 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_4541
timestamp 1668089732
transform 1 0 11680 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_4542
timestamp 1668089732
transform 1 0 11680 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_4543
timestamp 1668089732
transform 1 0 11680 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_4544
timestamp 1668089732
transform 1 0 11680 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_4545
timestamp 1668089732
transform 1 0 11680 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_4546
timestamp 1668089732
transform 1 0 11680 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_4547
timestamp 1668089732
transform 1 0 11680 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_4548
timestamp 1668089732
transform 1 0 11680 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_4549
timestamp 1668089732
transform 1 0 11680 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_4550
timestamp 1668089732
transform 1 0 11680 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_4551
timestamp 1668089732
transform 1 0 11680 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_4552
timestamp 1668089732
transform 1 0 11680 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_4553
timestamp 1668089732
transform 1 0 11680 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_4554
timestamp 1668089732
transform 1 0 11680 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_4555
timestamp 1668089732
transform 1 0 11680 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_4556
timestamp 1668089732
transform 1 0 11680 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_4557
timestamp 1668089732
transform 1 0 11680 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_4558
timestamp 1668089732
transform 1 0 11680 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_4559
timestamp 1668089732
transform 1 0 11680 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_4560
timestamp 1668089732
transform 1 0 11680 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_4561
timestamp 1668089732
transform 1 0 11680 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_4562
timestamp 1668089732
transform 1 0 11680 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_4563
timestamp 1668089732
transform 1 0 11680 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_4564
timestamp 1668089732
transform 1 0 11680 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_4565
timestamp 1668089732
transform 1 0 11680 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_4566
timestamp 1668089732
transform 1 0 11680 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_4567
timestamp 1668089732
transform 1 0 11680 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_4568
timestamp 1668089732
transform 1 0 11680 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_4569
timestamp 1668089732
transform 1 0 11680 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_4570
timestamp 1668089732
transform 1 0 11680 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_4571
timestamp 1668089732
transform 1 0 11680 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_4572
timestamp 1668089732
transform 1 0 11680 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_4573
timestamp 1668089732
transform 1 0 11680 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_4574
timestamp 1668089732
transform 1 0 11680 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_4575
timestamp 1668089732
transform 1 0 11680 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_4576
timestamp 1668089732
transform 1 0 11680 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_4577
timestamp 1668089732
transform 1 0 11680 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_4578
timestamp 1668089732
transform 1 0 11680 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_4579
timestamp 1668089732
transform 1 0 11680 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_4580
timestamp 1668089732
transform 1 0 11680 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_4581
timestamp 1668089732
transform 1 0 11680 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_4582
timestamp 1668089732
transform 1 0 11680 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_4583
timestamp 1668089732
transform 1 0 11680 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_4584
timestamp 1668089732
transform 1 0 11680 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_4585
timestamp 1668089732
transform 1 0 11680 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_4586
timestamp 1668089732
transform 1 0 11680 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_4587
timestamp 1668089732
transform 1 0 11680 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_4588
timestamp 1668089732
transform 1 0 11840 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_4589
timestamp 1668089732
transform 1 0 11840 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_4590
timestamp 1668089732
transform 1 0 11840 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_4591
timestamp 1668089732
transform 1 0 11840 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_4592
timestamp 1668089732
transform 1 0 11840 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_4593
timestamp 1668089732
transform 1 0 11840 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_4594
timestamp 1668089732
transform 1 0 11840 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_4595
timestamp 1668089732
transform 1 0 11840 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_4596
timestamp 1668089732
transform 1 0 11840 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_4597
timestamp 1668089732
transform 1 0 11840 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_4598
timestamp 1668089732
transform 1 0 11840 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_4599
timestamp 1668089732
transform 1 0 11840 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_4600
timestamp 1668089732
transform 1 0 11840 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_4601
timestamp 1668089732
transform 1 0 11840 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_4602
timestamp 1668089732
transform 1 0 11840 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_4603
timestamp 1668089732
transform 1 0 11840 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_4604
timestamp 1668089732
transform 1 0 11840 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_4605
timestamp 1668089732
transform 1 0 11840 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_4606
timestamp 1668089732
transform 1 0 11840 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_4607
timestamp 1668089732
transform 1 0 11840 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_4608
timestamp 1668089732
transform 1 0 11840 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_4609
timestamp 1668089732
transform 1 0 11840 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_4610
timestamp 1668089732
transform 1 0 11840 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_4611
timestamp 1668089732
transform 1 0 11840 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_4612
timestamp 1668089732
transform 1 0 11840 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_4613
timestamp 1668089732
transform 1 0 11840 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_4614
timestamp 1668089732
transform 1 0 11840 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_4615
timestamp 1668089732
transform 1 0 11840 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_4616
timestamp 1668089732
transform 1 0 11840 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_4617
timestamp 1668089732
transform 1 0 11840 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_4618
timestamp 1668089732
transform 1 0 11840 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_4619
timestamp 1668089732
transform 1 0 11840 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_4620
timestamp 1668089732
transform 1 0 11840 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_4621
timestamp 1668089732
transform 1 0 11840 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_4622
timestamp 1668089732
transform 1 0 11840 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_4623
timestamp 1668089732
transform 1 0 11840 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_4624
timestamp 1668089732
transform 1 0 11840 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_4625
timestamp 1668089732
transform 1 0 11840 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_4626
timestamp 1668089732
transform 1 0 11840 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_4627
timestamp 1668089732
transform 1 0 11840 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_4628
timestamp 1668089732
transform 1 0 11840 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_4629
timestamp 1668089732
transform 1 0 11840 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_4630
timestamp 1668089732
transform 1 0 11840 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_4631
timestamp 1668089732
transform 1 0 11840 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_4632
timestamp 1668089732
transform 1 0 11840 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_4633
timestamp 1668089732
transform 1 0 11840 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_4634
timestamp 1668089732
transform 1 0 11840 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_4635
timestamp 1668089732
transform 1 0 11840 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_4636
timestamp 1668089732
transform 1 0 11840 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_4637
timestamp 1668089732
transform 1 0 11840 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_4638
timestamp 1668089732
transform 1 0 11840 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_4639
timestamp 1668089732
transform 1 0 11840 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_4640
timestamp 1668089732
transform 1 0 11840 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_4641
timestamp 1668089732
transform 1 0 11840 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_4642
timestamp 1668089732
transform 1 0 11840 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_4643
timestamp 1668089732
transform 1 0 11840 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_4644
timestamp 1668089732
transform 1 0 11840 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_4645
timestamp 1668089732
transform 1 0 11840 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_4646
timestamp 1668089732
transform 1 0 11840 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_4647
timestamp 1668089732
transform 1 0 11840 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_4648
timestamp 1668089732
transform 1 0 11840 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_4649
timestamp 1668089732
transform 1 0 11840 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_4650
timestamp 1668089732
transform 1 0 12000 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_4651
timestamp 1668089732
transform 1 0 12000 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_4652
timestamp 1668089732
transform 1 0 12000 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_4653
timestamp 1668089732
transform 1 0 12000 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_4654
timestamp 1668089732
transform 1 0 12000 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_4655
timestamp 1668089732
transform 1 0 12000 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_4656
timestamp 1668089732
transform 1 0 12000 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_4657
timestamp 1668089732
transform 1 0 12000 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_4658
timestamp 1668089732
transform 1 0 12000 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_4659
timestamp 1668089732
transform 1 0 12000 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_4660
timestamp 1668089732
transform 1 0 12000 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_4661
timestamp 1668089732
transform 1 0 12000 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_4662
timestamp 1668089732
transform 1 0 12000 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_4663
timestamp 1668089732
transform 1 0 12000 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_4664
timestamp 1668089732
transform 1 0 12000 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_4665
timestamp 1668089732
transform 1 0 12000 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_4666
timestamp 1668089732
transform 1 0 12000 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_4667
timestamp 1668089732
transform 1 0 12000 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_4668
timestamp 1668089732
transform 1 0 12000 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_4669
timestamp 1668089732
transform 1 0 12000 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_4670
timestamp 1668089732
transform 1 0 12000 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_4671
timestamp 1668089732
transform 1 0 12000 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_4672
timestamp 1668089732
transform 1 0 12000 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_4673
timestamp 1668089732
transform 1 0 12000 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_4674
timestamp 1668089732
transform 1 0 12000 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_4675
timestamp 1668089732
transform 1 0 12000 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_4676
timestamp 1668089732
transform 1 0 12000 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_4677
timestamp 1668089732
transform 1 0 12000 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_4678
timestamp 1668089732
transform 1 0 12000 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_4679
timestamp 1668089732
transform 1 0 12000 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_4680
timestamp 1668089732
transform 1 0 12000 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_4681
timestamp 1668089732
transform 1 0 12000 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_4682
timestamp 1668089732
transform 1 0 12000 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_4683
timestamp 1668089732
transform 1 0 12000 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_4684
timestamp 1668089732
transform 1 0 12000 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_4685
timestamp 1668089732
transform 1 0 12000 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_4686
timestamp 1668089732
transform 1 0 12000 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_4687
timestamp 1668089732
transform 1 0 12000 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_4688
timestamp 1668089732
transform 1 0 12000 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_4689
timestamp 1668089732
transform 1 0 12000 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_4690
timestamp 1668089732
transform 1 0 12000 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_4691
timestamp 1668089732
transform 1 0 12000 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_4692
timestamp 1668089732
transform 1 0 12000 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_4693
timestamp 1668089732
transform 1 0 12000 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_4694
timestamp 1668089732
transform 1 0 12000 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_4695
timestamp 1668089732
transform 1 0 12000 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_4696
timestamp 1668089732
transform 1 0 12000 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_4697
timestamp 1668089732
transform 1 0 12000 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_4698
timestamp 1668089732
transform 1 0 12000 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_4699
timestamp 1668089732
transform 1 0 12000 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_4700
timestamp 1668089732
transform 1 0 12000 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_4701
timestamp 1668089732
transform 1 0 12000 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_4702
timestamp 1668089732
transform 1 0 12000 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_4703
timestamp 1668089732
transform 1 0 12000 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_4704
timestamp 1668089732
transform 1 0 12000 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_4705
timestamp 1668089732
transform 1 0 12000 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_4706
timestamp 1668089732
transform 1 0 12000 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_4707
timestamp 1668089732
transform 1 0 12000 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_4708
timestamp 1668089732
transform 1 0 12000 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_4709
timestamp 1668089732
transform 1 0 12000 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_4710
timestamp 1668089732
transform 1 0 12000 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_4711
timestamp 1668089732
transform 1 0 12000 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_4712
timestamp 1668089732
transform 1 0 12160 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_4713
timestamp 1668089732
transform 1 0 12160 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_4714
timestamp 1668089732
transform 1 0 12160 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_4715
timestamp 1668089732
transform 1 0 12160 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_4716
timestamp 1668089732
transform 1 0 12160 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_4717
timestamp 1668089732
transform 1 0 12160 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_4718
timestamp 1668089732
transform 1 0 12160 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_4719
timestamp 1668089732
transform 1 0 12160 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_4720
timestamp 1668089732
transform 1 0 12160 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_4721
timestamp 1668089732
transform 1 0 12160 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_4722
timestamp 1668089732
transform 1 0 12160 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_4723
timestamp 1668089732
transform 1 0 12160 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_4724
timestamp 1668089732
transform 1 0 12160 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_4725
timestamp 1668089732
transform 1 0 12160 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_4726
timestamp 1668089732
transform 1 0 12160 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_4727
timestamp 1668089732
transform 1 0 12160 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_4728
timestamp 1668089732
transform 1 0 12160 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_4729
timestamp 1668089732
transform 1 0 12160 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_4730
timestamp 1668089732
transform 1 0 12160 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_4731
timestamp 1668089732
transform 1 0 12160 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_4732
timestamp 1668089732
transform 1 0 12160 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_4733
timestamp 1668089732
transform 1 0 12160 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_4734
timestamp 1668089732
transform 1 0 12160 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_4735
timestamp 1668089732
transform 1 0 12160 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_4736
timestamp 1668089732
transform 1 0 12160 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_4737
timestamp 1668089732
transform 1 0 12160 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_4738
timestamp 1668089732
transform 1 0 12160 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_4739
timestamp 1668089732
transform 1 0 12160 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_4740
timestamp 1668089732
transform 1 0 12160 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_4741
timestamp 1668089732
transform 1 0 12160 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_4742
timestamp 1668089732
transform 1 0 12160 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_4743
timestamp 1668089732
transform 1 0 12160 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_4744
timestamp 1668089732
transform 1 0 12160 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_4745
timestamp 1668089732
transform 1 0 12160 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_4746
timestamp 1668089732
transform 1 0 12160 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_4747
timestamp 1668089732
transform 1 0 12160 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_4748
timestamp 1668089732
transform 1 0 12160 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_4749
timestamp 1668089732
transform 1 0 12160 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_4750
timestamp 1668089732
transform 1 0 12160 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_4751
timestamp 1668089732
transform 1 0 12160 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_4752
timestamp 1668089732
transform 1 0 12160 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_4753
timestamp 1668089732
transform 1 0 12160 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_4754
timestamp 1668089732
transform 1 0 12160 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_4755
timestamp 1668089732
transform 1 0 12160 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_4756
timestamp 1668089732
transform 1 0 12160 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_4757
timestamp 1668089732
transform 1 0 12160 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_4758
timestamp 1668089732
transform 1 0 12160 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_4759
timestamp 1668089732
transform 1 0 12160 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_4760
timestamp 1668089732
transform 1 0 12160 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_4761
timestamp 1668089732
transform 1 0 12160 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_4762
timestamp 1668089732
transform 1 0 12160 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_4763
timestamp 1668089732
transform 1 0 12160 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_4764
timestamp 1668089732
transform 1 0 12160 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_4765
timestamp 1668089732
transform 1 0 12160 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_4766
timestamp 1668089732
transform 1 0 12160 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_4767
timestamp 1668089732
transform 1 0 12160 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_4768
timestamp 1668089732
transform 1 0 12160 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_4769
timestamp 1668089732
transform 1 0 12160 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_4770
timestamp 1668089732
transform 1 0 12160 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_4771
timestamp 1668089732
transform 1 0 12160 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_4772
timestamp 1668089732
transform 1 0 12160 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_4773
timestamp 1668089732
transform 1 0 12160 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_4774
timestamp 1668089732
transform 1 0 12320 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_4775
timestamp 1668089732
transform 1 0 12320 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_4776
timestamp 1668089732
transform 1 0 12320 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_4777
timestamp 1668089732
transform 1 0 12320 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_4778
timestamp 1668089732
transform 1 0 12320 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_4779
timestamp 1668089732
transform 1 0 12320 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_4780
timestamp 1668089732
transform 1 0 12320 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_4781
timestamp 1668089732
transform 1 0 12320 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_4782
timestamp 1668089732
transform 1 0 12320 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_4783
timestamp 1668089732
transform 1 0 12320 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_4784
timestamp 1668089732
transform 1 0 12320 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_4785
timestamp 1668089732
transform 1 0 12320 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_4786
timestamp 1668089732
transform 1 0 12320 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_4787
timestamp 1668089732
transform 1 0 12320 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_4788
timestamp 1668089732
transform 1 0 12320 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_4789
timestamp 1668089732
transform 1 0 12320 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_4790
timestamp 1668089732
transform 1 0 12320 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_4791
timestamp 1668089732
transform 1 0 12320 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_4792
timestamp 1668089732
transform 1 0 12320 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_4793
timestamp 1668089732
transform 1 0 12320 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_4794
timestamp 1668089732
transform 1 0 12320 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_4795
timestamp 1668089732
transform 1 0 12320 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_4796
timestamp 1668089732
transform 1 0 12320 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_4797
timestamp 1668089732
transform 1 0 12320 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_4798
timestamp 1668089732
transform 1 0 12320 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_4799
timestamp 1668089732
transform 1 0 12320 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_4800
timestamp 1668089732
transform 1 0 12320 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_4801
timestamp 1668089732
transform 1 0 12320 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_4802
timestamp 1668089732
transform 1 0 12320 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_4803
timestamp 1668089732
transform 1 0 12320 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_4804
timestamp 1668089732
transform 1 0 12320 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_4805
timestamp 1668089732
transform 1 0 12320 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_4806
timestamp 1668089732
transform 1 0 12320 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_4807
timestamp 1668089732
transform 1 0 12320 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_4808
timestamp 1668089732
transform 1 0 12320 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_4809
timestamp 1668089732
transform 1 0 12320 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_4810
timestamp 1668089732
transform 1 0 12320 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_4811
timestamp 1668089732
transform 1 0 12320 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_4812
timestamp 1668089732
transform 1 0 12320 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_4813
timestamp 1668089732
transform 1 0 12320 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_4814
timestamp 1668089732
transform 1 0 12320 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_4815
timestamp 1668089732
transform 1 0 12320 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_4816
timestamp 1668089732
transform 1 0 12320 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_4817
timestamp 1668089732
transform 1 0 12320 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_4818
timestamp 1668089732
transform 1 0 12320 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_4819
timestamp 1668089732
transform 1 0 12320 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_4820
timestamp 1668089732
transform 1 0 12320 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_4821
timestamp 1668089732
transform 1 0 12320 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_4822
timestamp 1668089732
transform 1 0 12320 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_4823
timestamp 1668089732
transform 1 0 12320 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_4824
timestamp 1668089732
transform 1 0 12320 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_4825
timestamp 1668089732
transform 1 0 12320 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_4826
timestamp 1668089732
transform 1 0 12320 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_4827
timestamp 1668089732
transform 1 0 12320 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_4828
timestamp 1668089732
transform 1 0 12320 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_4829
timestamp 1668089732
transform 1 0 12320 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_4830
timestamp 1668089732
transform 1 0 12320 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_4831
timestamp 1668089732
transform 1 0 12320 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_4832
timestamp 1668089732
transform 1 0 12320 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_4833
timestamp 1668089732
transform 1 0 12320 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_4834
timestamp 1668089732
transform 1 0 12320 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_4835
timestamp 1668089732
transform 1 0 12320 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_4836
timestamp 1668089732
transform 1 0 12480 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_4837
timestamp 1668089732
transform 1 0 12480 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_4838
timestamp 1668089732
transform 1 0 12480 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_4839
timestamp 1668089732
transform 1 0 12480 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_4840
timestamp 1668089732
transform 1 0 12480 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_4841
timestamp 1668089732
transform 1 0 12480 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_4842
timestamp 1668089732
transform 1 0 12480 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_4843
timestamp 1668089732
transform 1 0 12480 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_4844
timestamp 1668089732
transform 1 0 12480 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_4845
timestamp 1668089732
transform 1 0 12480 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_4846
timestamp 1668089732
transform 1 0 12480 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_4847
timestamp 1668089732
transform 1 0 12480 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_4848
timestamp 1668089732
transform 1 0 12480 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_4849
timestamp 1668089732
transform 1 0 12480 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_4850
timestamp 1668089732
transform 1 0 12480 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_4851
timestamp 1668089732
transform 1 0 12480 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_4852
timestamp 1668089732
transform 1 0 12480 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_4853
timestamp 1668089732
transform 1 0 12480 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_4854
timestamp 1668089732
transform 1 0 12480 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_4855
timestamp 1668089732
transform 1 0 12480 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_4856
timestamp 1668089732
transform 1 0 12480 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_4857
timestamp 1668089732
transform 1 0 12480 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_4858
timestamp 1668089732
transform 1 0 12480 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_4859
timestamp 1668089732
transform 1 0 12480 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_4860
timestamp 1668089732
transform 1 0 12480 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_4861
timestamp 1668089732
transform 1 0 12480 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_4862
timestamp 1668089732
transform 1 0 12480 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_4863
timestamp 1668089732
transform 1 0 12480 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_4864
timestamp 1668089732
transform 1 0 12480 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_4865
timestamp 1668089732
transform 1 0 12480 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_4866
timestamp 1668089732
transform 1 0 12480 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_4867
timestamp 1668089732
transform 1 0 12480 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_4868
timestamp 1668089732
transform 1 0 12480 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_4869
timestamp 1668089732
transform 1 0 12480 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_4870
timestamp 1668089732
transform 1 0 12480 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_4871
timestamp 1668089732
transform 1 0 12480 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_4872
timestamp 1668089732
transform 1 0 12480 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_4873
timestamp 1668089732
transform 1 0 12480 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_4874
timestamp 1668089732
transform 1 0 12480 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_4875
timestamp 1668089732
transform 1 0 12480 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_4876
timestamp 1668089732
transform 1 0 12480 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_4877
timestamp 1668089732
transform 1 0 12480 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_4878
timestamp 1668089732
transform 1 0 12480 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_4879
timestamp 1668089732
transform 1 0 12480 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_4880
timestamp 1668089732
transform 1 0 12480 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_4881
timestamp 1668089732
transform 1 0 12480 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_4882
timestamp 1668089732
transform 1 0 12480 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_4883
timestamp 1668089732
transform 1 0 12480 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_4884
timestamp 1668089732
transform 1 0 12480 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_4885
timestamp 1668089732
transform 1 0 12480 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_4886
timestamp 1668089732
transform 1 0 12480 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_4887
timestamp 1668089732
transform 1 0 12480 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_4888
timestamp 1668089732
transform 1 0 12480 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_4889
timestamp 1668089732
transform 1 0 12480 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_4890
timestamp 1668089732
transform 1 0 12480 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_4891
timestamp 1668089732
transform 1 0 12480 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_4892
timestamp 1668089732
transform 1 0 12480 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_4893
timestamp 1668089732
transform 1 0 12480 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_4894
timestamp 1668089732
transform 1 0 12480 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_4895
timestamp 1668089732
transform 1 0 12480 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_4896
timestamp 1668089732
transform 1 0 12480 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_4897
timestamp 1668089732
transform 1 0 12480 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_4898
timestamp 1668089732
transform 1 0 12640 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_4899
timestamp 1668089732
transform 1 0 12640 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_4900
timestamp 1668089732
transform 1 0 12640 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_4901
timestamp 1668089732
transform 1 0 12640 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_4902
timestamp 1668089732
transform 1 0 12640 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_4903
timestamp 1668089732
transform 1 0 12640 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_4904
timestamp 1668089732
transform 1 0 12640 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_4905
timestamp 1668089732
transform 1 0 12640 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_4906
timestamp 1668089732
transform 1 0 12640 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_4907
timestamp 1668089732
transform 1 0 12640 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_4908
timestamp 1668089732
transform 1 0 12640 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_4909
timestamp 1668089732
transform 1 0 12640 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_4910
timestamp 1668089732
transform 1 0 12640 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_4911
timestamp 1668089732
transform 1 0 12640 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_4912
timestamp 1668089732
transform 1 0 12640 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_4913
timestamp 1668089732
transform 1 0 12640 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_4914
timestamp 1668089732
transform 1 0 12640 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_4915
timestamp 1668089732
transform 1 0 12640 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_4916
timestamp 1668089732
transform 1 0 12640 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_4917
timestamp 1668089732
transform 1 0 12640 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_4918
timestamp 1668089732
transform 1 0 12640 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_4919
timestamp 1668089732
transform 1 0 12640 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_4920
timestamp 1668089732
transform 1 0 12640 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_4921
timestamp 1668089732
transform 1 0 12640 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_4922
timestamp 1668089732
transform 1 0 12640 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_4923
timestamp 1668089732
transform 1 0 12640 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_4924
timestamp 1668089732
transform 1 0 12640 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_4925
timestamp 1668089732
transform 1 0 12640 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_4926
timestamp 1668089732
transform 1 0 12640 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_4927
timestamp 1668089732
transform 1 0 12640 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_4928
timestamp 1668089732
transform 1 0 12640 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_4929
timestamp 1668089732
transform 1 0 12640 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_4930
timestamp 1668089732
transform 1 0 12640 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_4931
timestamp 1668089732
transform 1 0 12640 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_4932
timestamp 1668089732
transform 1 0 12640 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_4933
timestamp 1668089732
transform 1 0 12640 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_4934
timestamp 1668089732
transform 1 0 12640 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_4935
timestamp 1668089732
transform 1 0 12640 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_4936
timestamp 1668089732
transform 1 0 12640 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_4937
timestamp 1668089732
transform 1 0 12640 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_4938
timestamp 1668089732
transform 1 0 12640 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_4939
timestamp 1668089732
transform 1 0 12640 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_4940
timestamp 1668089732
transform 1 0 12640 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_4941
timestamp 1668089732
transform 1 0 12640 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_4942
timestamp 1668089732
transform 1 0 12640 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_4943
timestamp 1668089732
transform 1 0 12640 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_4944
timestamp 1668089732
transform 1 0 12640 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_4945
timestamp 1668089732
transform 1 0 12640 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_4946
timestamp 1668089732
transform 1 0 12640 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_4947
timestamp 1668089732
transform 1 0 12640 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_4948
timestamp 1668089732
transform 1 0 12640 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_4949
timestamp 1668089732
transform 1 0 12640 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_4950
timestamp 1668089732
transform 1 0 12640 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_4951
timestamp 1668089732
transform 1 0 12640 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_4952
timestamp 1668089732
transform 1 0 12640 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_4953
timestamp 1668089732
transform 1 0 12640 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_4954
timestamp 1668089732
transform 1 0 12640 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_4955
timestamp 1668089732
transform 1 0 12640 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_4956
timestamp 1668089732
transform 1 0 12640 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_4957
timestamp 1668089732
transform 1 0 12640 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_4958
timestamp 1668089732
transform 1 0 12640 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_4959
timestamp 1668089732
transform 1 0 12640 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_4960
timestamp 1668089732
transform 1 0 12800 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_4961
timestamp 1668089732
transform 1 0 12800 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_4962
timestamp 1668089732
transform 1 0 12800 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_4963
timestamp 1668089732
transform 1 0 12800 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_4964
timestamp 1668089732
transform 1 0 12800 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_4965
timestamp 1668089732
transform 1 0 12800 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_4966
timestamp 1668089732
transform 1 0 12800 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_4967
timestamp 1668089732
transform 1 0 12800 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_4968
timestamp 1668089732
transform 1 0 12800 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_4969
timestamp 1668089732
transform 1 0 12800 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_4970
timestamp 1668089732
transform 1 0 12800 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_4971
timestamp 1668089732
transform 1 0 12800 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_4972
timestamp 1668089732
transform 1 0 12800 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_4973
timestamp 1668089732
transform 1 0 12800 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_4974
timestamp 1668089732
transform 1 0 12800 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_4975
timestamp 1668089732
transform 1 0 12800 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_4976
timestamp 1668089732
transform 1 0 12800 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_4977
timestamp 1668089732
transform 1 0 12800 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_4978
timestamp 1668089732
transform 1 0 12800 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_4979
timestamp 1668089732
transform 1 0 12800 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_4980
timestamp 1668089732
transform 1 0 12800 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_4981
timestamp 1668089732
transform 1 0 12800 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_4982
timestamp 1668089732
transform 1 0 12800 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_4983
timestamp 1668089732
transform 1 0 12800 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_4984
timestamp 1668089732
transform 1 0 12800 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_4985
timestamp 1668089732
transform 1 0 12800 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_4986
timestamp 1668089732
transform 1 0 12800 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_4987
timestamp 1668089732
transform 1 0 12800 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_4988
timestamp 1668089732
transform 1 0 12800 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_4989
timestamp 1668089732
transform 1 0 12800 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_4990
timestamp 1668089732
transform 1 0 12800 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_4991
timestamp 1668089732
transform 1 0 12800 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_4992
timestamp 1668089732
transform 1 0 12800 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_4993
timestamp 1668089732
transform 1 0 12800 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_4994
timestamp 1668089732
transform 1 0 12800 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_4995
timestamp 1668089732
transform 1 0 12800 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_4996
timestamp 1668089732
transform 1 0 12800 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_4997
timestamp 1668089732
transform 1 0 12800 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_4998
timestamp 1668089732
transform 1 0 12800 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_4999
timestamp 1668089732
transform 1 0 12800 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_5000
timestamp 1668089732
transform 1 0 12800 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_5001
timestamp 1668089732
transform 1 0 12800 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_5002
timestamp 1668089732
transform 1 0 12800 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_5003
timestamp 1668089732
transform 1 0 12800 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_5004
timestamp 1668089732
transform 1 0 12800 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_5005
timestamp 1668089732
transform 1 0 12800 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_5006
timestamp 1668089732
transform 1 0 12800 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_5007
timestamp 1668089732
transform 1 0 12800 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_5008
timestamp 1668089732
transform 1 0 12800 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_5009
timestamp 1668089732
transform 1 0 12800 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_5010
timestamp 1668089732
transform 1 0 12800 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_5011
timestamp 1668089732
transform 1 0 12800 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_5012
timestamp 1668089732
transform 1 0 12800 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_5013
timestamp 1668089732
transform 1 0 12800 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_5014
timestamp 1668089732
transform 1 0 12800 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_5015
timestamp 1668089732
transform 1 0 12800 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_5016
timestamp 1668089732
transform 1 0 12800 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_5017
timestamp 1668089732
transform 1 0 12800 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_5018
timestamp 1668089732
transform 1 0 12800 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_5019
timestamp 1668089732
transform 1 0 12800 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_5020
timestamp 1668089732
transform 1 0 12800 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_5021
timestamp 1668089732
transform 1 0 12800 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_5022
timestamp 1668089732
transform 1 0 12960 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_5023
timestamp 1668089732
transform 1 0 12960 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_5024
timestamp 1668089732
transform 1 0 12960 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_5025
timestamp 1668089732
transform 1 0 12960 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_5026
timestamp 1668089732
transform 1 0 12960 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_5027
timestamp 1668089732
transform 1 0 12960 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_5028
timestamp 1668089732
transform 1 0 12960 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_5029
timestamp 1668089732
transform 1 0 12960 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_5030
timestamp 1668089732
transform 1 0 12960 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_5031
timestamp 1668089732
transform 1 0 12960 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_5032
timestamp 1668089732
transform 1 0 12960 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_5033
timestamp 1668089732
transform 1 0 12960 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_5034
timestamp 1668089732
transform 1 0 12960 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_5035
timestamp 1668089732
transform 1 0 12960 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_5036
timestamp 1668089732
transform 1 0 12960 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_5037
timestamp 1668089732
transform 1 0 12960 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_5038
timestamp 1668089732
transform 1 0 12960 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_5039
timestamp 1668089732
transform 1 0 12960 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_5040
timestamp 1668089732
transform 1 0 12960 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_5041
timestamp 1668089732
transform 1 0 12960 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_5042
timestamp 1668089732
transform 1 0 12960 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_5043
timestamp 1668089732
transform 1 0 12960 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_5044
timestamp 1668089732
transform 1 0 12960 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_5045
timestamp 1668089732
transform 1 0 12960 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_5046
timestamp 1668089732
transform 1 0 12960 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_5047
timestamp 1668089732
transform 1 0 12960 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_5048
timestamp 1668089732
transform 1 0 12960 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_5049
timestamp 1668089732
transform 1 0 12960 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_5050
timestamp 1668089732
transform 1 0 12960 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_5051
timestamp 1668089732
transform 1 0 12960 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_5052
timestamp 1668089732
transform 1 0 12960 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_5053
timestamp 1668089732
transform 1 0 12960 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_5054
timestamp 1668089732
transform 1 0 12960 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_5055
timestamp 1668089732
transform 1 0 12960 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_5056
timestamp 1668089732
transform 1 0 12960 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_5057
timestamp 1668089732
transform 1 0 12960 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_5058
timestamp 1668089732
transform 1 0 12960 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_5059
timestamp 1668089732
transform 1 0 12960 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_5060
timestamp 1668089732
transform 1 0 12960 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_5061
timestamp 1668089732
transform 1 0 12960 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_5062
timestamp 1668089732
transform 1 0 12960 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_5063
timestamp 1668089732
transform 1 0 12960 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_5064
timestamp 1668089732
transform 1 0 12960 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_5065
timestamp 1668089732
transform 1 0 12960 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_5066
timestamp 1668089732
transform 1 0 12960 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_5067
timestamp 1668089732
transform 1 0 12960 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_5068
timestamp 1668089732
transform 1 0 12960 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_5069
timestamp 1668089732
transform 1 0 12960 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_5070
timestamp 1668089732
transform 1 0 12960 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_5071
timestamp 1668089732
transform 1 0 12960 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_5072
timestamp 1668089732
transform 1 0 12960 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_5073
timestamp 1668089732
transform 1 0 12960 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_5074
timestamp 1668089732
transform 1 0 12960 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_5075
timestamp 1668089732
transform 1 0 12960 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_5076
timestamp 1668089732
transform 1 0 12960 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_5077
timestamp 1668089732
transform 1 0 12960 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_5078
timestamp 1668089732
transform 1 0 12960 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_5079
timestamp 1668089732
transform 1 0 12960 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_5080
timestamp 1668089732
transform 1 0 12960 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_5081
timestamp 1668089732
transform 1 0 12960 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_5082
timestamp 1668089732
transform 1 0 12960 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_5083
timestamp 1668089732
transform 1 0 12960 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_5084
timestamp 1668089732
transform 1 0 13120 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_5085
timestamp 1668089732
transform 1 0 13120 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_5086
timestamp 1668089732
transform 1 0 13120 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_5087
timestamp 1668089732
transform 1 0 13120 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_5088
timestamp 1668089732
transform 1 0 13120 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_5089
timestamp 1668089732
transform 1 0 13120 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_5090
timestamp 1668089732
transform 1 0 13120 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_5091
timestamp 1668089732
transform 1 0 13120 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_5092
timestamp 1668089732
transform 1 0 13120 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_5093
timestamp 1668089732
transform 1 0 13120 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_5094
timestamp 1668089732
transform 1 0 13120 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_5095
timestamp 1668089732
transform 1 0 13120 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_5096
timestamp 1668089732
transform 1 0 13120 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_5097
timestamp 1668089732
transform 1 0 13120 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_5098
timestamp 1668089732
transform 1 0 13120 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_5099
timestamp 1668089732
transform 1 0 13120 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_5100
timestamp 1668089732
transform 1 0 13120 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_5101
timestamp 1668089732
transform 1 0 13120 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_5102
timestamp 1668089732
transform 1 0 13120 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_5103
timestamp 1668089732
transform 1 0 13120 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_5104
timestamp 1668089732
transform 1 0 13120 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_5105
timestamp 1668089732
transform 1 0 13120 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_5106
timestamp 1668089732
transform 1 0 13120 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_5107
timestamp 1668089732
transform 1 0 13120 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_5108
timestamp 1668089732
transform 1 0 13120 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_5109
timestamp 1668089732
transform 1 0 13120 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_5110
timestamp 1668089732
transform 1 0 13120 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_5111
timestamp 1668089732
transform 1 0 13120 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_5112
timestamp 1668089732
transform 1 0 13120 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_5113
timestamp 1668089732
transform 1 0 13120 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_5114
timestamp 1668089732
transform 1 0 13120 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_5115
timestamp 1668089732
transform 1 0 13120 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_5116
timestamp 1668089732
transform 1 0 13120 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_5117
timestamp 1668089732
transform 1 0 13120 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_5118
timestamp 1668089732
transform 1 0 13120 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_5119
timestamp 1668089732
transform 1 0 13120 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_5120
timestamp 1668089732
transform 1 0 13120 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_5121
timestamp 1668089732
transform 1 0 13120 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_5122
timestamp 1668089732
transform 1 0 13120 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_5123
timestamp 1668089732
transform 1 0 13120 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_5124
timestamp 1668089732
transform 1 0 13120 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_5125
timestamp 1668089732
transform 1 0 13120 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_5126
timestamp 1668089732
transform 1 0 13120 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_5127
timestamp 1668089732
transform 1 0 13120 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_5128
timestamp 1668089732
transform 1 0 13120 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_5129
timestamp 1668089732
transform 1 0 13120 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_5130
timestamp 1668089732
transform 1 0 13120 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_5131
timestamp 1668089732
transform 1 0 13120 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_5132
timestamp 1668089732
transform 1 0 13120 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_5133
timestamp 1668089732
transform 1 0 13120 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_5134
timestamp 1668089732
transform 1 0 13120 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_5135
timestamp 1668089732
transform 1 0 13120 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_5136
timestamp 1668089732
transform 1 0 13120 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_5137
timestamp 1668089732
transform 1 0 13120 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_5138
timestamp 1668089732
transform 1 0 13120 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_5139
timestamp 1668089732
transform 1 0 13120 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_5140
timestamp 1668089732
transform 1 0 13120 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_5141
timestamp 1668089732
transform 1 0 13120 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_5142
timestamp 1668089732
transform 1 0 13120 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_5143
timestamp 1668089732
transform 1 0 13120 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_5144
timestamp 1668089732
transform 1 0 13120 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_5145
timestamp 1668089732
transform 1 0 13120 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_5146
timestamp 1668089732
transform 1 0 13280 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_5147
timestamp 1668089732
transform 1 0 13280 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_5148
timestamp 1668089732
transform 1 0 13280 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_5149
timestamp 1668089732
transform 1 0 13280 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_5150
timestamp 1668089732
transform 1 0 13280 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_5151
timestamp 1668089732
transform 1 0 13280 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_5152
timestamp 1668089732
transform 1 0 13280 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_5153
timestamp 1668089732
transform 1 0 13280 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_5154
timestamp 1668089732
transform 1 0 13280 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_5155
timestamp 1668089732
transform 1 0 13280 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_5156
timestamp 1668089732
transform 1 0 13280 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_5157
timestamp 1668089732
transform 1 0 13280 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_5158
timestamp 1668089732
transform 1 0 13280 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_5159
timestamp 1668089732
transform 1 0 13280 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_5160
timestamp 1668089732
transform 1 0 13280 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_5161
timestamp 1668089732
transform 1 0 13280 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_5162
timestamp 1668089732
transform 1 0 13280 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_5163
timestamp 1668089732
transform 1 0 13280 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_5164
timestamp 1668089732
transform 1 0 13280 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_5165
timestamp 1668089732
transform 1 0 13280 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_5166
timestamp 1668089732
transform 1 0 13280 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_5167
timestamp 1668089732
transform 1 0 13280 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_5168
timestamp 1668089732
transform 1 0 13280 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_5169
timestamp 1668089732
transform 1 0 13280 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_5170
timestamp 1668089732
transform 1 0 13280 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_5171
timestamp 1668089732
transform 1 0 13280 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_5172
timestamp 1668089732
transform 1 0 13280 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_5173
timestamp 1668089732
transform 1 0 13280 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_5174
timestamp 1668089732
transform 1 0 13280 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_5175
timestamp 1668089732
transform 1 0 13280 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_5176
timestamp 1668089732
transform 1 0 13280 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_5177
timestamp 1668089732
transform 1 0 13280 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_5178
timestamp 1668089732
transform 1 0 13280 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_5179
timestamp 1668089732
transform 1 0 13280 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_5180
timestamp 1668089732
transform 1 0 13280 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_5181
timestamp 1668089732
transform 1 0 13280 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_5182
timestamp 1668089732
transform 1 0 13280 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_5183
timestamp 1668089732
transform 1 0 13280 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_5184
timestamp 1668089732
transform 1 0 13280 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_5185
timestamp 1668089732
transform 1 0 13280 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_5186
timestamp 1668089732
transform 1 0 13280 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_5187
timestamp 1668089732
transform 1 0 13280 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_5188
timestamp 1668089732
transform 1 0 13280 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_5189
timestamp 1668089732
transform 1 0 13280 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_5190
timestamp 1668089732
transform 1 0 13280 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_5191
timestamp 1668089732
transform 1 0 13280 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_5192
timestamp 1668089732
transform 1 0 13280 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_5193
timestamp 1668089732
transform 1 0 13280 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_5194
timestamp 1668089732
transform 1 0 13280 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_5195
timestamp 1668089732
transform 1 0 13280 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_5196
timestamp 1668089732
transform 1 0 13280 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_5197
timestamp 1668089732
transform 1 0 13280 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_5198
timestamp 1668089732
transform 1 0 13280 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_5199
timestamp 1668089732
transform 1 0 13280 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_5200
timestamp 1668089732
transform 1 0 13280 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_5201
timestamp 1668089732
transform 1 0 13280 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_5202
timestamp 1668089732
transform 1 0 13280 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_5203
timestamp 1668089732
transform 1 0 13280 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_5204
timestamp 1668089732
transform 1 0 13280 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_5205
timestamp 1668089732
transform 1 0 13280 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_5206
timestamp 1668089732
transform 1 0 13280 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_5207
timestamp 1668089732
transform 1 0 13280 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_5208
timestamp 1668089732
transform 1 0 13440 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_5209
timestamp 1668089732
transform 1 0 13440 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_5210
timestamp 1668089732
transform 1 0 13440 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_5211
timestamp 1668089732
transform 1 0 13440 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_5212
timestamp 1668089732
transform 1 0 13440 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_5213
timestamp 1668089732
transform 1 0 13440 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_5214
timestamp 1668089732
transform 1 0 13440 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_5215
timestamp 1668089732
transform 1 0 13440 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_5216
timestamp 1668089732
transform 1 0 13440 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_5217
timestamp 1668089732
transform 1 0 13440 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_5218
timestamp 1668089732
transform 1 0 13440 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_5219
timestamp 1668089732
transform 1 0 13440 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_5220
timestamp 1668089732
transform 1 0 13440 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_5221
timestamp 1668089732
transform 1 0 13440 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_5222
timestamp 1668089732
transform 1 0 13440 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_5223
timestamp 1668089732
transform 1 0 13440 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_5224
timestamp 1668089732
transform 1 0 13440 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_5225
timestamp 1668089732
transform 1 0 13440 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_5226
timestamp 1668089732
transform 1 0 13440 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_5227
timestamp 1668089732
transform 1 0 13440 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_5228
timestamp 1668089732
transform 1 0 13440 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_5229
timestamp 1668089732
transform 1 0 13440 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_5230
timestamp 1668089732
transform 1 0 13440 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_5231
timestamp 1668089732
transform 1 0 13440 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_5232
timestamp 1668089732
transform 1 0 13440 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_5233
timestamp 1668089732
transform 1 0 13440 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_5234
timestamp 1668089732
transform 1 0 13440 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_5235
timestamp 1668089732
transform 1 0 13440 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_5236
timestamp 1668089732
transform 1 0 13440 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_5237
timestamp 1668089732
transform 1 0 13440 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_5238
timestamp 1668089732
transform 1 0 13440 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_5239
timestamp 1668089732
transform 1 0 13440 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_5240
timestamp 1668089732
transform 1 0 13440 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_5241
timestamp 1668089732
transform 1 0 13440 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_5242
timestamp 1668089732
transform 1 0 13440 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_5243
timestamp 1668089732
transform 1 0 13440 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_5244
timestamp 1668089732
transform 1 0 13440 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_5245
timestamp 1668089732
transform 1 0 13440 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_5246
timestamp 1668089732
transform 1 0 13440 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_5247
timestamp 1668089732
transform 1 0 13440 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_5248
timestamp 1668089732
transform 1 0 13440 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_5249
timestamp 1668089732
transform 1 0 13440 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_5250
timestamp 1668089732
transform 1 0 13440 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_5251
timestamp 1668089732
transform 1 0 13440 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_5252
timestamp 1668089732
transform 1 0 13440 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_5253
timestamp 1668089732
transform 1 0 13440 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_5254
timestamp 1668089732
transform 1 0 13440 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_5255
timestamp 1668089732
transform 1 0 13440 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_5256
timestamp 1668089732
transform 1 0 13440 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_5257
timestamp 1668089732
transform 1 0 13440 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_5258
timestamp 1668089732
transform 1 0 13440 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_5259
timestamp 1668089732
transform 1 0 13440 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_5260
timestamp 1668089732
transform 1 0 13440 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_5261
timestamp 1668089732
transform 1 0 13440 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_5262
timestamp 1668089732
transform 1 0 13440 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_5263
timestamp 1668089732
transform 1 0 13440 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_5264
timestamp 1668089732
transform 1 0 13440 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_5265
timestamp 1668089732
transform 1 0 13440 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_5266
timestamp 1668089732
transform 1 0 13440 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_5267
timestamp 1668089732
transform 1 0 13440 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_5268
timestamp 1668089732
transform 1 0 13440 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_5269
timestamp 1668089732
transform 1 0 13440 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_5270
timestamp 1668089732
transform 1 0 13600 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_5271
timestamp 1668089732
transform 1 0 13600 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_5272
timestamp 1668089732
transform 1 0 13600 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_5273
timestamp 1668089732
transform 1 0 13600 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_5274
timestamp 1668089732
transform 1 0 13600 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_5275
timestamp 1668089732
transform 1 0 13600 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_5276
timestamp 1668089732
transform 1 0 13600 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_5277
timestamp 1668089732
transform 1 0 13600 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_5278
timestamp 1668089732
transform 1 0 13600 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_5279
timestamp 1668089732
transform 1 0 13600 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_5280
timestamp 1668089732
transform 1 0 13600 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_5281
timestamp 1668089732
transform 1 0 13600 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_5282
timestamp 1668089732
transform 1 0 13600 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_5283
timestamp 1668089732
transform 1 0 13600 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_5284
timestamp 1668089732
transform 1 0 13600 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_5285
timestamp 1668089732
transform 1 0 13600 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_5286
timestamp 1668089732
transform 1 0 13600 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_5287
timestamp 1668089732
transform 1 0 13600 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_5288
timestamp 1668089732
transform 1 0 13600 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_5289
timestamp 1668089732
transform 1 0 13600 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_5290
timestamp 1668089732
transform 1 0 13600 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_5291
timestamp 1668089732
transform 1 0 13600 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_5292
timestamp 1668089732
transform 1 0 13600 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_5293
timestamp 1668089732
transform 1 0 13600 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_5294
timestamp 1668089732
transform 1 0 13600 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_5295
timestamp 1668089732
transform 1 0 13600 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_5296
timestamp 1668089732
transform 1 0 13600 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_5297
timestamp 1668089732
transform 1 0 13600 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_5298
timestamp 1668089732
transform 1 0 13600 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_5299
timestamp 1668089732
transform 1 0 13600 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_5300
timestamp 1668089732
transform 1 0 13600 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_5301
timestamp 1668089732
transform 1 0 13600 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_5302
timestamp 1668089732
transform 1 0 13600 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_5303
timestamp 1668089732
transform 1 0 13600 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_5304
timestamp 1668089732
transform 1 0 13600 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_5305
timestamp 1668089732
transform 1 0 13600 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_5306
timestamp 1668089732
transform 1 0 13600 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_5307
timestamp 1668089732
transform 1 0 13600 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_5308
timestamp 1668089732
transform 1 0 13600 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_5309
timestamp 1668089732
transform 1 0 13600 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_5310
timestamp 1668089732
transform 1 0 13600 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_5311
timestamp 1668089732
transform 1 0 13600 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_5312
timestamp 1668089732
transform 1 0 13600 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_5313
timestamp 1668089732
transform 1 0 13600 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_5314
timestamp 1668089732
transform 1 0 13600 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_5315
timestamp 1668089732
transform 1 0 13600 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_5316
timestamp 1668089732
transform 1 0 13600 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_5317
timestamp 1668089732
transform 1 0 13600 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_5318
timestamp 1668089732
transform 1 0 13600 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_5319
timestamp 1668089732
transform 1 0 13600 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_5320
timestamp 1668089732
transform 1 0 13600 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_5321
timestamp 1668089732
transform 1 0 13600 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_5322
timestamp 1668089732
transform 1 0 13600 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_5323
timestamp 1668089732
transform 1 0 13600 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_5324
timestamp 1668089732
transform 1 0 13600 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_5325
timestamp 1668089732
transform 1 0 13600 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_5326
timestamp 1668089732
transform 1 0 13600 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_5327
timestamp 1668089732
transform 1 0 13600 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_5328
timestamp 1668089732
transform 1 0 13600 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_5329
timestamp 1668089732
transform 1 0 13600 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_5330
timestamp 1668089732
transform 1 0 13600 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_5331
timestamp 1668089732
transform 1 0 13600 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_5332
timestamp 1668089732
transform 1 0 13760 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_5333
timestamp 1668089732
transform 1 0 13760 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_5334
timestamp 1668089732
transform 1 0 13760 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_5335
timestamp 1668089732
transform 1 0 13760 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_5336
timestamp 1668089732
transform 1 0 13760 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_5337
timestamp 1668089732
transform 1 0 13760 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_5338
timestamp 1668089732
transform 1 0 13760 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_5339
timestamp 1668089732
transform 1 0 13760 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_5340
timestamp 1668089732
transform 1 0 13760 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_5341
timestamp 1668089732
transform 1 0 13760 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_5342
timestamp 1668089732
transform 1 0 13760 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_5343
timestamp 1668089732
transform 1 0 13760 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_5344
timestamp 1668089732
transform 1 0 13760 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_5345
timestamp 1668089732
transform 1 0 13760 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_5346
timestamp 1668089732
transform 1 0 13760 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_5347
timestamp 1668089732
transform 1 0 13760 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_5348
timestamp 1668089732
transform 1 0 13760 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_5349
timestamp 1668089732
transform 1 0 13760 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_5350
timestamp 1668089732
transform 1 0 13760 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_5351
timestamp 1668089732
transform 1 0 13760 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_5352
timestamp 1668089732
transform 1 0 13760 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_5353
timestamp 1668089732
transform 1 0 13760 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_5354
timestamp 1668089732
transform 1 0 13760 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_5355
timestamp 1668089732
transform 1 0 13760 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_5356
timestamp 1668089732
transform 1 0 13760 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_5357
timestamp 1668089732
transform 1 0 13760 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_5358
timestamp 1668089732
transform 1 0 13760 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_5359
timestamp 1668089732
transform 1 0 13760 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_5360
timestamp 1668089732
transform 1 0 13760 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_5361
timestamp 1668089732
transform 1 0 13760 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_5362
timestamp 1668089732
transform 1 0 13760 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_5363
timestamp 1668089732
transform 1 0 13760 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_5364
timestamp 1668089732
transform 1 0 13760 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_5365
timestamp 1668089732
transform 1 0 13760 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_5366
timestamp 1668089732
transform 1 0 13760 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_5367
timestamp 1668089732
transform 1 0 13760 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_5368
timestamp 1668089732
transform 1 0 13760 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_5369
timestamp 1668089732
transform 1 0 13760 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_5370
timestamp 1668089732
transform 1 0 13760 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_5371
timestamp 1668089732
transform 1 0 13760 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_5372
timestamp 1668089732
transform 1 0 13760 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_5373
timestamp 1668089732
transform 1 0 13760 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_5374
timestamp 1668089732
transform 1 0 13760 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_5375
timestamp 1668089732
transform 1 0 13760 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_5376
timestamp 1668089732
transform 1 0 13760 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_5377
timestamp 1668089732
transform 1 0 13760 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_5378
timestamp 1668089732
transform 1 0 13760 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_5379
timestamp 1668089732
transform 1 0 13760 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_5380
timestamp 1668089732
transform 1 0 13760 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_5381
timestamp 1668089732
transform 1 0 13760 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_5382
timestamp 1668089732
transform 1 0 13760 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_5383
timestamp 1668089732
transform 1 0 13760 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_5384
timestamp 1668089732
transform 1 0 13760 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_5385
timestamp 1668089732
transform 1 0 13760 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_5386
timestamp 1668089732
transform 1 0 13760 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_5387
timestamp 1668089732
transform 1 0 13760 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_5388
timestamp 1668089732
transform 1 0 13760 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_5389
timestamp 1668089732
transform 1 0 13760 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_5390
timestamp 1668089732
transform 1 0 13760 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_5391
timestamp 1668089732
transform 1 0 13760 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_5392
timestamp 1668089732
transform 1 0 13760 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_5393
timestamp 1668089732
transform 1 0 13760 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_5394
timestamp 1668089732
transform 1 0 13920 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_5395
timestamp 1668089732
transform 1 0 13920 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_5396
timestamp 1668089732
transform 1 0 13920 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_5397
timestamp 1668089732
transform 1 0 13920 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_5398
timestamp 1668089732
transform 1 0 13920 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_5399
timestamp 1668089732
transform 1 0 13920 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_5400
timestamp 1668089732
transform 1 0 13920 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_5401
timestamp 1668089732
transform 1 0 13920 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_5402
timestamp 1668089732
transform 1 0 13920 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_5403
timestamp 1668089732
transform 1 0 13920 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_5404
timestamp 1668089732
transform 1 0 13920 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_5405
timestamp 1668089732
transform 1 0 13920 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_5406
timestamp 1668089732
transform 1 0 13920 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_5407
timestamp 1668089732
transform 1 0 13920 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_5408
timestamp 1668089732
transform 1 0 13920 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_5409
timestamp 1668089732
transform 1 0 13920 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_5410
timestamp 1668089732
transform 1 0 13920 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_5411
timestamp 1668089732
transform 1 0 13920 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_5412
timestamp 1668089732
transform 1 0 13920 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_5413
timestamp 1668089732
transform 1 0 13920 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_5414
timestamp 1668089732
transform 1 0 13920 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_5415
timestamp 1668089732
transform 1 0 13920 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_5416
timestamp 1668089732
transform 1 0 13920 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_5417
timestamp 1668089732
transform 1 0 13920 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_5418
timestamp 1668089732
transform 1 0 13920 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_5419
timestamp 1668089732
transform 1 0 13920 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_5420
timestamp 1668089732
transform 1 0 13920 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_5421
timestamp 1668089732
transform 1 0 13920 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_5422
timestamp 1668089732
transform 1 0 13920 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_5423
timestamp 1668089732
transform 1 0 13920 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_5424
timestamp 1668089732
transform 1 0 13920 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_5425
timestamp 1668089732
transform 1 0 13920 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_5426
timestamp 1668089732
transform 1 0 13920 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_5427
timestamp 1668089732
transform 1 0 13920 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_5428
timestamp 1668089732
transform 1 0 13920 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_5429
timestamp 1668089732
transform 1 0 13920 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_5430
timestamp 1668089732
transform 1 0 13920 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_5431
timestamp 1668089732
transform 1 0 13920 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_5432
timestamp 1668089732
transform 1 0 13920 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_5433
timestamp 1668089732
transform 1 0 13920 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_5434
timestamp 1668089732
transform 1 0 13920 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_5435
timestamp 1668089732
transform 1 0 13920 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_5436
timestamp 1668089732
transform 1 0 13920 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_5437
timestamp 1668089732
transform 1 0 13920 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_5438
timestamp 1668089732
transform 1 0 13920 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_5439
timestamp 1668089732
transform 1 0 13920 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_5440
timestamp 1668089732
transform 1 0 13920 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_5441
timestamp 1668089732
transform 1 0 13920 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_5442
timestamp 1668089732
transform 1 0 13920 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_5443
timestamp 1668089732
transform 1 0 13920 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_5444
timestamp 1668089732
transform 1 0 13920 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_5445
timestamp 1668089732
transform 1 0 13920 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_5446
timestamp 1668089732
transform 1 0 13920 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_5447
timestamp 1668089732
transform 1 0 13920 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_5448
timestamp 1668089732
transform 1 0 13920 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_5449
timestamp 1668089732
transform 1 0 13920 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_5450
timestamp 1668089732
transform 1 0 13920 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_5451
timestamp 1668089732
transform 1 0 13920 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_5452
timestamp 1668089732
transform 1 0 13920 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_5453
timestamp 1668089732
transform 1 0 13920 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_5454
timestamp 1668089732
transform 1 0 13920 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_5455
timestamp 1668089732
transform 1 0 13920 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_5456
timestamp 1668089732
transform 1 0 14080 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_5457
timestamp 1668089732
transform 1 0 14080 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_5458
timestamp 1668089732
transform 1 0 14080 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_5459
timestamp 1668089732
transform 1 0 14080 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_5460
timestamp 1668089732
transform 1 0 14080 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_5461
timestamp 1668089732
transform 1 0 14080 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_5462
timestamp 1668089732
transform 1 0 14080 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_5463
timestamp 1668089732
transform 1 0 14080 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_5464
timestamp 1668089732
transform 1 0 14080 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_5465
timestamp 1668089732
transform 1 0 14080 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_5466
timestamp 1668089732
transform 1 0 14080 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_5467
timestamp 1668089732
transform 1 0 14080 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_5468
timestamp 1668089732
transform 1 0 14080 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_5469
timestamp 1668089732
transform 1 0 14080 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_5470
timestamp 1668089732
transform 1 0 14080 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_5471
timestamp 1668089732
transform 1 0 14080 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_5472
timestamp 1668089732
transform 1 0 14080 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_5473
timestamp 1668089732
transform 1 0 14080 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_5474
timestamp 1668089732
transform 1 0 14080 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_5475
timestamp 1668089732
transform 1 0 14080 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_5476
timestamp 1668089732
transform 1 0 14080 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_5477
timestamp 1668089732
transform 1 0 14080 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_5478
timestamp 1668089732
transform 1 0 14080 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_5479
timestamp 1668089732
transform 1 0 14080 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_5480
timestamp 1668089732
transform 1 0 14080 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_5481
timestamp 1668089732
transform 1 0 14080 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_5482
timestamp 1668089732
transform 1 0 14080 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_5483
timestamp 1668089732
transform 1 0 14080 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_5484
timestamp 1668089732
transform 1 0 14080 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_5485
timestamp 1668089732
transform 1 0 14080 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_5486
timestamp 1668089732
transform 1 0 14080 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_5487
timestamp 1668089732
transform 1 0 14080 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_5488
timestamp 1668089732
transform 1 0 14080 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_5489
timestamp 1668089732
transform 1 0 14080 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_5490
timestamp 1668089732
transform 1 0 14080 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_5491
timestamp 1668089732
transform 1 0 14080 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_5492
timestamp 1668089732
transform 1 0 14080 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_5493
timestamp 1668089732
transform 1 0 14080 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_5494
timestamp 1668089732
transform 1 0 14080 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_5495
timestamp 1668089732
transform 1 0 14080 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_5496
timestamp 1668089732
transform 1 0 14080 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_5497
timestamp 1668089732
transform 1 0 14080 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_5498
timestamp 1668089732
transform 1 0 14080 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_5499
timestamp 1668089732
transform 1 0 14080 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_5500
timestamp 1668089732
transform 1 0 14080 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_5501
timestamp 1668089732
transform 1 0 14080 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_5502
timestamp 1668089732
transform 1 0 14080 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_5503
timestamp 1668089732
transform 1 0 14080 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_5504
timestamp 1668089732
transform 1 0 14080 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_5505
timestamp 1668089732
transform 1 0 14080 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_5506
timestamp 1668089732
transform 1 0 14080 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_5507
timestamp 1668089732
transform 1 0 14080 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_5508
timestamp 1668089732
transform 1 0 14080 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_5509
timestamp 1668089732
transform 1 0 14080 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_5510
timestamp 1668089732
transform 1 0 14080 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_5511
timestamp 1668089732
transform 1 0 14080 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_5512
timestamp 1668089732
transform 1 0 14080 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_5513
timestamp 1668089732
transform 1 0 14080 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_5514
timestamp 1668089732
transform 1 0 14080 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_5515
timestamp 1668089732
transform 1 0 14080 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_5516
timestamp 1668089732
transform 1 0 14080 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_5517
timestamp 1668089732
transform 1 0 14080 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_5518
timestamp 1668089732
transform 1 0 14240 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_5519
timestamp 1668089732
transform 1 0 14240 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_5520
timestamp 1668089732
transform 1 0 14240 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_5521
timestamp 1668089732
transform 1 0 14240 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_5522
timestamp 1668089732
transform 1 0 14240 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_5523
timestamp 1668089732
transform 1 0 14240 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_5524
timestamp 1668089732
transform 1 0 14240 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_5525
timestamp 1668089732
transform 1 0 14240 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_5526
timestamp 1668089732
transform 1 0 14240 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_5527
timestamp 1668089732
transform 1 0 14240 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_5528
timestamp 1668089732
transform 1 0 14240 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_5529
timestamp 1668089732
transform 1 0 14240 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_5530
timestamp 1668089732
transform 1 0 14240 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_5531
timestamp 1668089732
transform 1 0 14240 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_5532
timestamp 1668089732
transform 1 0 14240 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_5533
timestamp 1668089732
transform 1 0 14240 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_5534
timestamp 1668089732
transform 1 0 14240 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_5535
timestamp 1668089732
transform 1 0 14240 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_5536
timestamp 1668089732
transform 1 0 14240 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_5537
timestamp 1668089732
transform 1 0 14240 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_5538
timestamp 1668089732
transform 1 0 14240 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_5539
timestamp 1668089732
transform 1 0 14240 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_5540
timestamp 1668089732
transform 1 0 14240 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_5541
timestamp 1668089732
transform 1 0 14240 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_5542
timestamp 1668089732
transform 1 0 14240 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_5543
timestamp 1668089732
transform 1 0 14240 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_5544
timestamp 1668089732
transform 1 0 14240 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_5545
timestamp 1668089732
transform 1 0 14240 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_5546
timestamp 1668089732
transform 1 0 14240 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_5547
timestamp 1668089732
transform 1 0 14240 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_5548
timestamp 1668089732
transform 1 0 14240 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_5549
timestamp 1668089732
transform 1 0 14240 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_5550
timestamp 1668089732
transform 1 0 14240 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_5551
timestamp 1668089732
transform 1 0 14240 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_5552
timestamp 1668089732
transform 1 0 14240 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_5553
timestamp 1668089732
transform 1 0 14240 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_5554
timestamp 1668089732
transform 1 0 14240 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_5555
timestamp 1668089732
transform 1 0 14240 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_5556
timestamp 1668089732
transform 1 0 14240 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_5557
timestamp 1668089732
transform 1 0 14240 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_5558
timestamp 1668089732
transform 1 0 14240 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_5559
timestamp 1668089732
transform 1 0 14240 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_5560
timestamp 1668089732
transform 1 0 14240 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_5561
timestamp 1668089732
transform 1 0 14240 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_5562
timestamp 1668089732
transform 1 0 14240 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_5563
timestamp 1668089732
transform 1 0 14240 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_5564
timestamp 1668089732
transform 1 0 14240 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_5565
timestamp 1668089732
transform 1 0 14240 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_5566
timestamp 1668089732
transform 1 0 14240 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_5567
timestamp 1668089732
transform 1 0 14240 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_5568
timestamp 1668089732
transform 1 0 14240 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_5569
timestamp 1668089732
transform 1 0 14240 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_5570
timestamp 1668089732
transform 1 0 14240 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_5571
timestamp 1668089732
transform 1 0 14240 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_5572
timestamp 1668089732
transform 1 0 14240 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_5573
timestamp 1668089732
transform 1 0 14240 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_5574
timestamp 1668089732
transform 1 0 14240 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_5575
timestamp 1668089732
transform 1 0 14240 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_5576
timestamp 1668089732
transform 1 0 14240 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_5577
timestamp 1668089732
transform 1 0 14240 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_5578
timestamp 1668089732
transform 1 0 14240 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_5579
timestamp 1668089732
transform 1 0 14240 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_5580
timestamp 1668089732
transform 1 0 14400 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_5581
timestamp 1668089732
transform 1 0 14400 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_5582
timestamp 1668089732
transform 1 0 14400 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_5583
timestamp 1668089732
transform 1 0 14400 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_5584
timestamp 1668089732
transform 1 0 14400 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_5585
timestamp 1668089732
transform 1 0 14400 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_5586
timestamp 1668089732
transform 1 0 14400 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_5587
timestamp 1668089732
transform 1 0 14400 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_5588
timestamp 1668089732
transform 1 0 14400 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_5589
timestamp 1668089732
transform 1 0 14400 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_5590
timestamp 1668089732
transform 1 0 14400 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_5591
timestamp 1668089732
transform 1 0 14400 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_5592
timestamp 1668089732
transform 1 0 14400 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_5593
timestamp 1668089732
transform 1 0 14400 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_5594
timestamp 1668089732
transform 1 0 14400 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_5595
timestamp 1668089732
transform 1 0 14400 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_5596
timestamp 1668089732
transform 1 0 14400 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_5597
timestamp 1668089732
transform 1 0 14400 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_5598
timestamp 1668089732
transform 1 0 14400 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_5599
timestamp 1668089732
transform 1 0 14400 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_5600
timestamp 1668089732
transform 1 0 14400 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_5601
timestamp 1668089732
transform 1 0 14400 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_5602
timestamp 1668089732
transform 1 0 14400 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_5603
timestamp 1668089732
transform 1 0 14400 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_5604
timestamp 1668089732
transform 1 0 14400 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_5605
timestamp 1668089732
transform 1 0 14400 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_5606
timestamp 1668089732
transform 1 0 14400 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_5607
timestamp 1668089732
transform 1 0 14400 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_5608
timestamp 1668089732
transform 1 0 14400 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_5609
timestamp 1668089732
transform 1 0 14400 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_5610
timestamp 1668089732
transform 1 0 14400 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_5611
timestamp 1668089732
transform 1 0 14400 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_5612
timestamp 1668089732
transform 1 0 14400 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_5613
timestamp 1668089732
transform 1 0 14400 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_5614
timestamp 1668089732
transform 1 0 14400 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_5615
timestamp 1668089732
transform 1 0 14400 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_5616
timestamp 1668089732
transform 1 0 14400 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_5617
timestamp 1668089732
transform 1 0 14400 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_5618
timestamp 1668089732
transform 1 0 14400 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_5619
timestamp 1668089732
transform 1 0 14400 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_5620
timestamp 1668089732
transform 1 0 14400 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_5621
timestamp 1668089732
transform 1 0 14400 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_5622
timestamp 1668089732
transform 1 0 14400 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_5623
timestamp 1668089732
transform 1 0 14400 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_5624
timestamp 1668089732
transform 1 0 14400 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_5625
timestamp 1668089732
transform 1 0 14400 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_5626
timestamp 1668089732
transform 1 0 14400 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_5627
timestamp 1668089732
transform 1 0 14400 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_5628
timestamp 1668089732
transform 1 0 14400 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_5629
timestamp 1668089732
transform 1 0 14400 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_5630
timestamp 1668089732
transform 1 0 14400 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_5631
timestamp 1668089732
transform 1 0 14400 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_5632
timestamp 1668089732
transform 1 0 14400 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_5633
timestamp 1668089732
transform 1 0 14400 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_5634
timestamp 1668089732
transform 1 0 14400 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_5635
timestamp 1668089732
transform 1 0 14400 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_5636
timestamp 1668089732
transform 1 0 14400 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_5637
timestamp 1668089732
transform 1 0 14400 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_5638
timestamp 1668089732
transform 1 0 14400 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_5639
timestamp 1668089732
transform 1 0 14400 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_5640
timestamp 1668089732
transform 1 0 14400 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_5641
timestamp 1668089732
transform 1 0 14400 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_5642
timestamp 1668089732
transform 1 0 14560 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_5643
timestamp 1668089732
transform 1 0 14560 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_5644
timestamp 1668089732
transform 1 0 14560 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_5645
timestamp 1668089732
transform 1 0 14560 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_5646
timestamp 1668089732
transform 1 0 14560 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_5647
timestamp 1668089732
transform 1 0 14560 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_5648
timestamp 1668089732
transform 1 0 14560 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_5649
timestamp 1668089732
transform 1 0 14560 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_5650
timestamp 1668089732
transform 1 0 14560 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_5651
timestamp 1668089732
transform 1 0 14560 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_5652
timestamp 1668089732
transform 1 0 14560 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_5653
timestamp 1668089732
transform 1 0 14560 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_5654
timestamp 1668089732
transform 1 0 14560 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_5655
timestamp 1668089732
transform 1 0 14560 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_5656
timestamp 1668089732
transform 1 0 14560 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_5657
timestamp 1668089732
transform 1 0 14560 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_5658
timestamp 1668089732
transform 1 0 14560 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_5659
timestamp 1668089732
transform 1 0 14560 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_5660
timestamp 1668089732
transform 1 0 14560 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_5661
timestamp 1668089732
transform 1 0 14560 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_5662
timestamp 1668089732
transform 1 0 14560 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_5663
timestamp 1668089732
transform 1 0 14560 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_5664
timestamp 1668089732
transform 1 0 14560 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_5665
timestamp 1668089732
transform 1 0 14560 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_5666
timestamp 1668089732
transform 1 0 14560 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_5667
timestamp 1668089732
transform 1 0 14560 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_5668
timestamp 1668089732
transform 1 0 14560 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_5669
timestamp 1668089732
transform 1 0 14560 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_5670
timestamp 1668089732
transform 1 0 14560 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_5671
timestamp 1668089732
transform 1 0 14560 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_5672
timestamp 1668089732
transform 1 0 14560 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_5673
timestamp 1668089732
transform 1 0 14560 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_5674
timestamp 1668089732
transform 1 0 14560 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_5675
timestamp 1668089732
transform 1 0 14560 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_5676
timestamp 1668089732
transform 1 0 14560 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_5677
timestamp 1668089732
transform 1 0 14560 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_5678
timestamp 1668089732
transform 1 0 14560 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_5679
timestamp 1668089732
transform 1 0 14560 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_5680
timestamp 1668089732
transform 1 0 14560 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_5681
timestamp 1668089732
transform 1 0 14560 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_5682
timestamp 1668089732
transform 1 0 14560 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_5683
timestamp 1668089732
transform 1 0 14560 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_5684
timestamp 1668089732
transform 1 0 14560 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_5685
timestamp 1668089732
transform 1 0 14560 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_5686
timestamp 1668089732
transform 1 0 14560 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_5687
timestamp 1668089732
transform 1 0 14560 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_5688
timestamp 1668089732
transform 1 0 14560 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_5689
timestamp 1668089732
transform 1 0 14560 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_5690
timestamp 1668089732
transform 1 0 14560 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_5691
timestamp 1668089732
transform 1 0 14560 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_5692
timestamp 1668089732
transform 1 0 14560 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_5693
timestamp 1668089732
transform 1 0 14560 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_5694
timestamp 1668089732
transform 1 0 14560 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_5695
timestamp 1668089732
transform 1 0 14560 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_5696
timestamp 1668089732
transform 1 0 14560 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_5697
timestamp 1668089732
transform 1 0 14560 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_5698
timestamp 1668089732
transform 1 0 14560 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_5699
timestamp 1668089732
transform 1 0 14560 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_5700
timestamp 1668089732
transform 1 0 14560 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_5701
timestamp 1668089732
transform 1 0 14560 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_5702
timestamp 1668089732
transform 1 0 14560 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_5703
timestamp 1668089732
transform 1 0 14560 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_5704
timestamp 1668089732
transform 1 0 14720 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_5705
timestamp 1668089732
transform 1 0 14720 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_5706
timestamp 1668089732
transform 1 0 14720 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_5707
timestamp 1668089732
transform 1 0 14720 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_5708
timestamp 1668089732
transform 1 0 14720 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_5709
timestamp 1668089732
transform 1 0 14720 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_5710
timestamp 1668089732
transform 1 0 14720 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_5711
timestamp 1668089732
transform 1 0 14720 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_5712
timestamp 1668089732
transform 1 0 14720 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_5713
timestamp 1668089732
transform 1 0 14720 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_5714
timestamp 1668089732
transform 1 0 14720 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_5715
timestamp 1668089732
transform 1 0 14720 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_5716
timestamp 1668089732
transform 1 0 14720 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_5717
timestamp 1668089732
transform 1 0 14720 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_5718
timestamp 1668089732
transform 1 0 14720 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_5719
timestamp 1668089732
transform 1 0 14720 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_5720
timestamp 1668089732
transform 1 0 14720 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_5721
timestamp 1668089732
transform 1 0 14720 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_5722
timestamp 1668089732
transform 1 0 14720 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_5723
timestamp 1668089732
transform 1 0 14720 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_5724
timestamp 1668089732
transform 1 0 14720 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_5725
timestamp 1668089732
transform 1 0 14720 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_5726
timestamp 1668089732
transform 1 0 14720 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_5727
timestamp 1668089732
transform 1 0 14720 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_5728
timestamp 1668089732
transform 1 0 14720 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_5729
timestamp 1668089732
transform 1 0 14720 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_5730
timestamp 1668089732
transform 1 0 14720 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_5731
timestamp 1668089732
transform 1 0 14720 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_5732
timestamp 1668089732
transform 1 0 14720 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_5733
timestamp 1668089732
transform 1 0 14720 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_5734
timestamp 1668089732
transform 1 0 14720 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_5735
timestamp 1668089732
transform 1 0 14720 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_5736
timestamp 1668089732
transform 1 0 14720 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_5737
timestamp 1668089732
transform 1 0 14720 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_5738
timestamp 1668089732
transform 1 0 14720 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_5739
timestamp 1668089732
transform 1 0 14720 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_5740
timestamp 1668089732
transform 1 0 14720 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_5741
timestamp 1668089732
transform 1 0 14720 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_5742
timestamp 1668089732
transform 1 0 14720 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_5743
timestamp 1668089732
transform 1 0 14720 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_5744
timestamp 1668089732
transform 1 0 14720 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_5745
timestamp 1668089732
transform 1 0 14720 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_5746
timestamp 1668089732
transform 1 0 14720 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_5747
timestamp 1668089732
transform 1 0 14720 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_5748
timestamp 1668089732
transform 1 0 14720 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_5749
timestamp 1668089732
transform 1 0 14720 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_5750
timestamp 1668089732
transform 1 0 14720 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_5751
timestamp 1668089732
transform 1 0 14720 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_5752
timestamp 1668089732
transform 1 0 14720 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_5753
timestamp 1668089732
transform 1 0 14720 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_5754
timestamp 1668089732
transform 1 0 14720 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_5755
timestamp 1668089732
transform 1 0 14720 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_5756
timestamp 1668089732
transform 1 0 14720 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_5757
timestamp 1668089732
transform 1 0 14720 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_5758
timestamp 1668089732
transform 1 0 14720 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_5759
timestamp 1668089732
transform 1 0 14720 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_5760
timestamp 1668089732
transform 1 0 14720 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_5761
timestamp 1668089732
transform 1 0 14720 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_5762
timestamp 1668089732
transform 1 0 14720 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_5763
timestamp 1668089732
transform 1 0 14720 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_5764
timestamp 1668089732
transform 1 0 14720 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_5765
timestamp 1668089732
transform 1 0 14720 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_5766
timestamp 1668089732
transform 1 0 14880 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_5767
timestamp 1668089732
transform 1 0 14880 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_5768
timestamp 1668089732
transform 1 0 14880 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_5769
timestamp 1668089732
transform 1 0 14880 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_5770
timestamp 1668089732
transform 1 0 14880 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_5771
timestamp 1668089732
transform 1 0 14880 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_5772
timestamp 1668089732
transform 1 0 14880 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_5773
timestamp 1668089732
transform 1 0 14880 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_5774
timestamp 1668089732
transform 1 0 14880 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_5775
timestamp 1668089732
transform 1 0 14880 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_5776
timestamp 1668089732
transform 1 0 14880 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_5777
timestamp 1668089732
transform 1 0 14880 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_5778
timestamp 1668089732
transform 1 0 14880 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_5779
timestamp 1668089732
transform 1 0 14880 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_5780
timestamp 1668089732
transform 1 0 14880 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_5781
timestamp 1668089732
transform 1 0 14880 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_5782
timestamp 1668089732
transform 1 0 14880 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_5783
timestamp 1668089732
transform 1 0 14880 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_5784
timestamp 1668089732
transform 1 0 14880 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_5785
timestamp 1668089732
transform 1 0 14880 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_5786
timestamp 1668089732
transform 1 0 14880 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_5787
timestamp 1668089732
transform 1 0 14880 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_5788
timestamp 1668089732
transform 1 0 14880 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_5789
timestamp 1668089732
transform 1 0 14880 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_5790
timestamp 1668089732
transform 1 0 14880 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_5791
timestamp 1668089732
transform 1 0 14880 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_5792
timestamp 1668089732
transform 1 0 14880 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_5793
timestamp 1668089732
transform 1 0 14880 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_5794
timestamp 1668089732
transform 1 0 14880 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_5795
timestamp 1668089732
transform 1 0 14880 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_5796
timestamp 1668089732
transform 1 0 14880 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_5797
timestamp 1668089732
transform 1 0 14880 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_5798
timestamp 1668089732
transform 1 0 14880 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_5799
timestamp 1668089732
transform 1 0 14880 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_5800
timestamp 1668089732
transform 1 0 14880 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_5801
timestamp 1668089732
transform 1 0 14880 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_5802
timestamp 1668089732
transform 1 0 14880 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_5803
timestamp 1668089732
transform 1 0 14880 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_5804
timestamp 1668089732
transform 1 0 14880 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_5805
timestamp 1668089732
transform 1 0 14880 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_5806
timestamp 1668089732
transform 1 0 14880 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_5807
timestamp 1668089732
transform 1 0 14880 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_5808
timestamp 1668089732
transform 1 0 14880 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_5809
timestamp 1668089732
transform 1 0 14880 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_5810
timestamp 1668089732
transform 1 0 14880 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_5811
timestamp 1668089732
transform 1 0 14880 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_5812
timestamp 1668089732
transform 1 0 14880 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_5813
timestamp 1668089732
transform 1 0 14880 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_5814
timestamp 1668089732
transform 1 0 14880 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_5815
timestamp 1668089732
transform 1 0 14880 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_5816
timestamp 1668089732
transform 1 0 14880 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_5817
timestamp 1668089732
transform 1 0 14880 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_5818
timestamp 1668089732
transform 1 0 14880 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_5819
timestamp 1668089732
transform 1 0 14880 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_5820
timestamp 1668089732
transform 1 0 14880 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_5821
timestamp 1668089732
transform 1 0 14880 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_5822
timestamp 1668089732
transform 1 0 14880 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_5823
timestamp 1668089732
transform 1 0 14880 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_5824
timestamp 1668089732
transform 1 0 14880 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_5825
timestamp 1668089732
transform 1 0 14880 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_5826
timestamp 1668089732
transform 1 0 14880 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_5827
timestamp 1668089732
transform 1 0 14880 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_5828
timestamp 1668089732
transform 1 0 15040 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_5829
timestamp 1668089732
transform 1 0 15040 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_5830
timestamp 1668089732
transform 1 0 15040 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_5831
timestamp 1668089732
transform 1 0 15040 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_5832
timestamp 1668089732
transform 1 0 15040 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_5833
timestamp 1668089732
transform 1 0 15040 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_5834
timestamp 1668089732
transform 1 0 15040 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_5835
timestamp 1668089732
transform 1 0 15040 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_5836
timestamp 1668089732
transform 1 0 15040 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_5837
timestamp 1668089732
transform 1 0 15040 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_5838
timestamp 1668089732
transform 1 0 15040 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_5839
timestamp 1668089732
transform 1 0 15040 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_5840
timestamp 1668089732
transform 1 0 15040 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_5841
timestamp 1668089732
transform 1 0 15040 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_5842
timestamp 1668089732
transform 1 0 15040 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_5843
timestamp 1668089732
transform 1 0 15040 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_5844
timestamp 1668089732
transform 1 0 15040 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_5845
timestamp 1668089732
transform 1 0 15040 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_5846
timestamp 1668089732
transform 1 0 15040 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_5847
timestamp 1668089732
transform 1 0 15040 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_5848
timestamp 1668089732
transform 1 0 15040 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_5849
timestamp 1668089732
transform 1 0 15040 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_5850
timestamp 1668089732
transform 1 0 15040 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_5851
timestamp 1668089732
transform 1 0 15040 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_5852
timestamp 1668089732
transform 1 0 15040 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_5853
timestamp 1668089732
transform 1 0 15040 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_5854
timestamp 1668089732
transform 1 0 15040 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_5855
timestamp 1668089732
transform 1 0 15040 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_5856
timestamp 1668089732
transform 1 0 15040 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_5857
timestamp 1668089732
transform 1 0 15040 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_5858
timestamp 1668089732
transform 1 0 15040 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_5859
timestamp 1668089732
transform 1 0 15040 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_5860
timestamp 1668089732
transform 1 0 15040 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_5861
timestamp 1668089732
transform 1 0 15040 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_5862
timestamp 1668089732
transform 1 0 15040 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_5863
timestamp 1668089732
transform 1 0 15040 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_5864
timestamp 1668089732
transform 1 0 15040 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_5865
timestamp 1668089732
transform 1 0 15040 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_5866
timestamp 1668089732
transform 1 0 15040 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_5867
timestamp 1668089732
transform 1 0 15040 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_5868
timestamp 1668089732
transform 1 0 15040 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_5869
timestamp 1668089732
transform 1 0 15040 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_5870
timestamp 1668089732
transform 1 0 15040 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_5871
timestamp 1668089732
transform 1 0 15040 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_5872
timestamp 1668089732
transform 1 0 15040 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_5873
timestamp 1668089732
transform 1 0 15040 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_5874
timestamp 1668089732
transform 1 0 15040 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_5875
timestamp 1668089732
transform 1 0 15040 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_5876
timestamp 1668089732
transform 1 0 15040 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_5877
timestamp 1668089732
transform 1 0 15040 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_5878
timestamp 1668089732
transform 1 0 15040 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_5879
timestamp 1668089732
transform 1 0 15040 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_5880
timestamp 1668089732
transform 1 0 15040 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_5881
timestamp 1668089732
transform 1 0 15040 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_5882
timestamp 1668089732
transform 1 0 15040 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_5883
timestamp 1668089732
transform 1 0 15040 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_5884
timestamp 1668089732
transform 1 0 15040 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_5885
timestamp 1668089732
transform 1 0 15040 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_5886
timestamp 1668089732
transform 1 0 15040 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_5887
timestamp 1668089732
transform 1 0 15040 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_5888
timestamp 1668089732
transform 1 0 15040 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_5889
timestamp 1668089732
transform 1 0 15040 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_5890
timestamp 1668089732
transform 1 0 15200 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_5891
timestamp 1668089732
transform 1 0 15200 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_5892
timestamp 1668089732
transform 1 0 15200 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_5893
timestamp 1668089732
transform 1 0 15200 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_5894
timestamp 1668089732
transform 1 0 15200 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_5895
timestamp 1668089732
transform 1 0 15200 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_5896
timestamp 1668089732
transform 1 0 15200 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_5897
timestamp 1668089732
transform 1 0 15200 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_5898
timestamp 1668089732
transform 1 0 15200 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_5899
timestamp 1668089732
transform 1 0 15200 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_5900
timestamp 1668089732
transform 1 0 15200 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_5901
timestamp 1668089732
transform 1 0 15200 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_5902
timestamp 1668089732
transform 1 0 15200 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_5903
timestamp 1668089732
transform 1 0 15200 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_5904
timestamp 1668089732
transform 1 0 15200 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_5905
timestamp 1668089732
transform 1 0 15200 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_5906
timestamp 1668089732
transform 1 0 15200 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_5907
timestamp 1668089732
transform 1 0 15200 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_5908
timestamp 1668089732
transform 1 0 15200 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_5909
timestamp 1668089732
transform 1 0 15200 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_5910
timestamp 1668089732
transform 1 0 15200 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_5911
timestamp 1668089732
transform 1 0 15200 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_5912
timestamp 1668089732
transform 1 0 15200 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_5913
timestamp 1668089732
transform 1 0 15200 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_5914
timestamp 1668089732
transform 1 0 15200 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_5915
timestamp 1668089732
transform 1 0 15200 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_5916
timestamp 1668089732
transform 1 0 15200 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_5917
timestamp 1668089732
transform 1 0 15200 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_5918
timestamp 1668089732
transform 1 0 15200 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_5919
timestamp 1668089732
transform 1 0 15200 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_5920
timestamp 1668089732
transform 1 0 15200 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_5921
timestamp 1668089732
transform 1 0 15200 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_5922
timestamp 1668089732
transform 1 0 15200 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_5923
timestamp 1668089732
transform 1 0 15200 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_5924
timestamp 1668089732
transform 1 0 15200 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_5925
timestamp 1668089732
transform 1 0 15200 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_5926
timestamp 1668089732
transform 1 0 15200 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_5927
timestamp 1668089732
transform 1 0 15200 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_5928
timestamp 1668089732
transform 1 0 15200 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_5929
timestamp 1668089732
transform 1 0 15200 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_5930
timestamp 1668089732
transform 1 0 15200 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_5931
timestamp 1668089732
transform 1 0 15200 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_5932
timestamp 1668089732
transform 1 0 15200 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_5933
timestamp 1668089732
transform 1 0 15200 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_5934
timestamp 1668089732
transform 1 0 15200 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_5935
timestamp 1668089732
transform 1 0 15200 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_5936
timestamp 1668089732
transform 1 0 15200 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_5937
timestamp 1668089732
transform 1 0 15200 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_5938
timestamp 1668089732
transform 1 0 15200 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_5939
timestamp 1668089732
transform 1 0 15200 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_5940
timestamp 1668089732
transform 1 0 15200 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_5941
timestamp 1668089732
transform 1 0 15200 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_5942
timestamp 1668089732
transform 1 0 15200 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_5943
timestamp 1668089732
transform 1 0 15200 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_5944
timestamp 1668089732
transform 1 0 15200 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_5945
timestamp 1668089732
transform 1 0 15200 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_5946
timestamp 1668089732
transform 1 0 15200 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_5947
timestamp 1668089732
transform 1 0 15200 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_5948
timestamp 1668089732
transform 1 0 15200 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_5949
timestamp 1668089732
transform 1 0 15200 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_5950
timestamp 1668089732
transform 1 0 15200 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_5951
timestamp 1668089732
transform 1 0 15200 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_5952
timestamp 1668089732
transform 1 0 15360 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_5953
timestamp 1668089732
transform 1 0 15360 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_5954
timestamp 1668089732
transform 1 0 15360 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_5955
timestamp 1668089732
transform 1 0 15360 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_5956
timestamp 1668089732
transform 1 0 15360 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_5957
timestamp 1668089732
transform 1 0 15360 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_5958
timestamp 1668089732
transform 1 0 15360 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_5959
timestamp 1668089732
transform 1 0 15360 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_5960
timestamp 1668089732
transform 1 0 15360 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_5961
timestamp 1668089732
transform 1 0 15360 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_5962
timestamp 1668089732
transform 1 0 15360 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_5963
timestamp 1668089732
transform 1 0 15360 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_5964
timestamp 1668089732
transform 1 0 15360 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_5965
timestamp 1668089732
transform 1 0 15360 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_5966
timestamp 1668089732
transform 1 0 15360 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_5967
timestamp 1668089732
transform 1 0 15360 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_5968
timestamp 1668089732
transform 1 0 15360 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_5969
timestamp 1668089732
transform 1 0 15360 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_5970
timestamp 1668089732
transform 1 0 15360 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_5971
timestamp 1668089732
transform 1 0 15360 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_5972
timestamp 1668089732
transform 1 0 15360 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_5973
timestamp 1668089732
transform 1 0 15360 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_5974
timestamp 1668089732
transform 1 0 15360 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_5975
timestamp 1668089732
transform 1 0 15360 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_5976
timestamp 1668089732
transform 1 0 15360 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_5977
timestamp 1668089732
transform 1 0 15360 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_5978
timestamp 1668089732
transform 1 0 15360 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_5979
timestamp 1668089732
transform 1 0 15360 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_5980
timestamp 1668089732
transform 1 0 15360 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_5981
timestamp 1668089732
transform 1 0 15360 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_5982
timestamp 1668089732
transform 1 0 15360 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_5983
timestamp 1668089732
transform 1 0 15360 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_5984
timestamp 1668089732
transform 1 0 15360 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_5985
timestamp 1668089732
transform 1 0 15360 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_5986
timestamp 1668089732
transform 1 0 15360 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_5987
timestamp 1668089732
transform 1 0 15360 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_5988
timestamp 1668089732
transform 1 0 15360 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_5989
timestamp 1668089732
transform 1 0 15360 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_5990
timestamp 1668089732
transform 1 0 15360 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_5991
timestamp 1668089732
transform 1 0 15360 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_5992
timestamp 1668089732
transform 1 0 15360 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_5993
timestamp 1668089732
transform 1 0 15360 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_5994
timestamp 1668089732
transform 1 0 15360 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_5995
timestamp 1668089732
transform 1 0 15360 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_5996
timestamp 1668089732
transform 1 0 15360 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_5997
timestamp 1668089732
transform 1 0 15360 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_5998
timestamp 1668089732
transform 1 0 15360 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_5999
timestamp 1668089732
transform 1 0 15360 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_6000
timestamp 1668089732
transform 1 0 15360 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_6001
timestamp 1668089732
transform 1 0 15360 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_6002
timestamp 1668089732
transform 1 0 15360 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_6003
timestamp 1668089732
transform 1 0 15360 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_6004
timestamp 1668089732
transform 1 0 15360 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_6005
timestamp 1668089732
transform 1 0 15360 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_6006
timestamp 1668089732
transform 1 0 15360 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_6007
timestamp 1668089732
transform 1 0 15360 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_6008
timestamp 1668089732
transform 1 0 15360 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_6009
timestamp 1668089732
transform 1 0 15360 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_6010
timestamp 1668089732
transform 1 0 15360 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_6011
timestamp 1668089732
transform 1 0 15360 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_6012
timestamp 1668089732
transform 1 0 15360 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_6013
timestamp 1668089732
transform 1 0 15360 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_6014
timestamp 1668089732
transform 1 0 15520 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_6015
timestamp 1668089732
transform 1 0 15520 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_6016
timestamp 1668089732
transform 1 0 15520 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_6017
timestamp 1668089732
transform 1 0 15520 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_6018
timestamp 1668089732
transform 1 0 15520 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_6019
timestamp 1668089732
transform 1 0 15520 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_6020
timestamp 1668089732
transform 1 0 15520 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_6021
timestamp 1668089732
transform 1 0 15520 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_6022
timestamp 1668089732
transform 1 0 15520 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_6023
timestamp 1668089732
transform 1 0 15520 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_6024
timestamp 1668089732
transform 1 0 15520 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_6025
timestamp 1668089732
transform 1 0 15520 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_6026
timestamp 1668089732
transform 1 0 15520 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_6027
timestamp 1668089732
transform 1 0 15520 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_6028
timestamp 1668089732
transform 1 0 15520 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_6029
timestamp 1668089732
transform 1 0 15520 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_6030
timestamp 1668089732
transform 1 0 15520 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_6031
timestamp 1668089732
transform 1 0 15520 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_6032
timestamp 1668089732
transform 1 0 15520 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_6033
timestamp 1668089732
transform 1 0 15520 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_6034
timestamp 1668089732
transform 1 0 15520 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_6035
timestamp 1668089732
transform 1 0 15520 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_6036
timestamp 1668089732
transform 1 0 15520 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_6037
timestamp 1668089732
transform 1 0 15520 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_6038
timestamp 1668089732
transform 1 0 15520 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_6039
timestamp 1668089732
transform 1 0 15520 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_6040
timestamp 1668089732
transform 1 0 15520 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_6041
timestamp 1668089732
transform 1 0 15520 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_6042
timestamp 1668089732
transform 1 0 15520 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_6043
timestamp 1668089732
transform 1 0 15520 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_6044
timestamp 1668089732
transform 1 0 15520 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_6045
timestamp 1668089732
transform 1 0 15520 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_6046
timestamp 1668089732
transform 1 0 15520 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_6047
timestamp 1668089732
transform 1 0 15520 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_6048
timestamp 1668089732
transform 1 0 15520 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_6049
timestamp 1668089732
transform 1 0 15520 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_6050
timestamp 1668089732
transform 1 0 15520 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_6051
timestamp 1668089732
transform 1 0 15520 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_6052
timestamp 1668089732
transform 1 0 15520 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_6053
timestamp 1668089732
transform 1 0 15520 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_6054
timestamp 1668089732
transform 1 0 15520 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_6055
timestamp 1668089732
transform 1 0 15520 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_6056
timestamp 1668089732
transform 1 0 15520 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_6057
timestamp 1668089732
transform 1 0 15520 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_6058
timestamp 1668089732
transform 1 0 15520 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_6059
timestamp 1668089732
transform 1 0 15520 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_6060
timestamp 1668089732
transform 1 0 15520 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_6061
timestamp 1668089732
transform 1 0 15520 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_6062
timestamp 1668089732
transform 1 0 15520 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_6063
timestamp 1668089732
transform 1 0 15520 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_6064
timestamp 1668089732
transform 1 0 15520 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_6065
timestamp 1668089732
transform 1 0 15520 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_6066
timestamp 1668089732
transform 1 0 15520 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_6067
timestamp 1668089732
transform 1 0 15520 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_6068
timestamp 1668089732
transform 1 0 15520 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_6069
timestamp 1668089732
transform 1 0 15520 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_6070
timestamp 1668089732
transform 1 0 15520 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_6071
timestamp 1668089732
transform 1 0 15520 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_6072
timestamp 1668089732
transform 1 0 15520 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_6073
timestamp 1668089732
transform 1 0 15520 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_6074
timestamp 1668089732
transform 1 0 15520 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_6075
timestamp 1668089732
transform 1 0 15520 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_6076
timestamp 1668089732
transform 1 0 15680 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_6077
timestamp 1668089732
transform 1 0 15680 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_6078
timestamp 1668089732
transform 1 0 15680 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_6079
timestamp 1668089732
transform 1 0 15680 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_6080
timestamp 1668089732
transform 1 0 15680 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_6081
timestamp 1668089732
transform 1 0 15680 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_6082
timestamp 1668089732
transform 1 0 15680 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_6083
timestamp 1668089732
transform 1 0 15680 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_6084
timestamp 1668089732
transform 1 0 15680 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_6085
timestamp 1668089732
transform 1 0 15680 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_6086
timestamp 1668089732
transform 1 0 15680 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_6087
timestamp 1668089732
transform 1 0 15680 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_6088
timestamp 1668089732
transform 1 0 15680 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_6089
timestamp 1668089732
transform 1 0 15680 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_6090
timestamp 1668089732
transform 1 0 15680 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_6091
timestamp 1668089732
transform 1 0 15680 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_6092
timestamp 1668089732
transform 1 0 15680 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_6093
timestamp 1668089732
transform 1 0 15680 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_6094
timestamp 1668089732
transform 1 0 15680 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_6095
timestamp 1668089732
transform 1 0 15680 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_6096
timestamp 1668089732
transform 1 0 15680 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_6097
timestamp 1668089732
transform 1 0 15680 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_6098
timestamp 1668089732
transform 1 0 15680 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_6099
timestamp 1668089732
transform 1 0 15680 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_6100
timestamp 1668089732
transform 1 0 15680 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_6101
timestamp 1668089732
transform 1 0 15680 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_6102
timestamp 1668089732
transform 1 0 15680 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_6103
timestamp 1668089732
transform 1 0 15680 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_6104
timestamp 1668089732
transform 1 0 15680 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_6105
timestamp 1668089732
transform 1 0 15680 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_6106
timestamp 1668089732
transform 1 0 15680 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_6107
timestamp 1668089732
transform 1 0 15680 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_6108
timestamp 1668089732
transform 1 0 15680 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_6109
timestamp 1668089732
transform 1 0 15680 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_6110
timestamp 1668089732
transform 1 0 15680 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_6111
timestamp 1668089732
transform 1 0 15680 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_6112
timestamp 1668089732
transform 1 0 15680 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_6113
timestamp 1668089732
transform 1 0 15680 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_6114
timestamp 1668089732
transform 1 0 15680 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_6115
timestamp 1668089732
transform 1 0 15680 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_6116
timestamp 1668089732
transform 1 0 15680 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_6117
timestamp 1668089732
transform 1 0 15680 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_6118
timestamp 1668089732
transform 1 0 15680 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_6119
timestamp 1668089732
transform 1 0 15680 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_6120
timestamp 1668089732
transform 1 0 15680 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_6121
timestamp 1668089732
transform 1 0 15680 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_6122
timestamp 1668089732
transform 1 0 15680 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_6123
timestamp 1668089732
transform 1 0 15680 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_6124
timestamp 1668089732
transform 1 0 15680 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_6125
timestamp 1668089732
transform 1 0 15680 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_6126
timestamp 1668089732
transform 1 0 15680 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_6127
timestamp 1668089732
transform 1 0 15680 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_6128
timestamp 1668089732
transform 1 0 15680 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_6129
timestamp 1668089732
transform 1 0 15680 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_6130
timestamp 1668089732
transform 1 0 15680 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_6131
timestamp 1668089732
transform 1 0 15680 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_6132
timestamp 1668089732
transform 1 0 15680 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_6133
timestamp 1668089732
transform 1 0 15680 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_6134
timestamp 1668089732
transform 1 0 15680 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_6135
timestamp 1668089732
transform 1 0 15680 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_6136
timestamp 1668089732
transform 1 0 15680 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_6137
timestamp 1668089732
transform 1 0 15680 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_6138
timestamp 1668089732
transform 1 0 15840 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_6139
timestamp 1668089732
transform 1 0 15840 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_6140
timestamp 1668089732
transform 1 0 15840 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_6141
timestamp 1668089732
transform 1 0 15840 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_6142
timestamp 1668089732
transform 1 0 15840 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_6143
timestamp 1668089732
transform 1 0 15840 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_6144
timestamp 1668089732
transform 1 0 15840 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_6145
timestamp 1668089732
transform 1 0 15840 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_6146
timestamp 1668089732
transform 1 0 15840 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_6147
timestamp 1668089732
transform 1 0 15840 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_6148
timestamp 1668089732
transform 1 0 15840 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_6149
timestamp 1668089732
transform 1 0 15840 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_6150
timestamp 1668089732
transform 1 0 15840 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_6151
timestamp 1668089732
transform 1 0 15840 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_6152
timestamp 1668089732
transform 1 0 15840 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_6153
timestamp 1668089732
transform 1 0 15840 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_6154
timestamp 1668089732
transform 1 0 15840 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_6155
timestamp 1668089732
transform 1 0 15840 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_6156
timestamp 1668089732
transform 1 0 15840 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_6157
timestamp 1668089732
transform 1 0 15840 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_6158
timestamp 1668089732
transform 1 0 15840 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_6159
timestamp 1668089732
transform 1 0 15840 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_6160
timestamp 1668089732
transform 1 0 15840 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_6161
timestamp 1668089732
transform 1 0 15840 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_6162
timestamp 1668089732
transform 1 0 15840 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_6163
timestamp 1668089732
transform 1 0 15840 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_6164
timestamp 1668089732
transform 1 0 15840 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_6165
timestamp 1668089732
transform 1 0 15840 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_6166
timestamp 1668089732
transform 1 0 15840 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_6167
timestamp 1668089732
transform 1 0 15840 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_6168
timestamp 1668089732
transform 1 0 15840 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_6169
timestamp 1668089732
transform 1 0 15840 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_6170
timestamp 1668089732
transform 1 0 15840 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_6171
timestamp 1668089732
transform 1 0 15840 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_6172
timestamp 1668089732
transform 1 0 15840 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_6173
timestamp 1668089732
transform 1 0 15840 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_6174
timestamp 1668089732
transform 1 0 15840 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_6175
timestamp 1668089732
transform 1 0 15840 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_6176
timestamp 1668089732
transform 1 0 15840 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_6177
timestamp 1668089732
transform 1 0 15840 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_6178
timestamp 1668089732
transform 1 0 15840 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_6179
timestamp 1668089732
transform 1 0 15840 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_6180
timestamp 1668089732
transform 1 0 15840 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_6181
timestamp 1668089732
transform 1 0 15840 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_6182
timestamp 1668089732
transform 1 0 15840 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_6183
timestamp 1668089732
transform 1 0 15840 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_6184
timestamp 1668089732
transform 1 0 15840 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_6185
timestamp 1668089732
transform 1 0 15840 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_6186
timestamp 1668089732
transform 1 0 15840 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_6187
timestamp 1668089732
transform 1 0 15840 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_6188
timestamp 1668089732
transform 1 0 15840 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_6189
timestamp 1668089732
transform 1 0 15840 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_6190
timestamp 1668089732
transform 1 0 15840 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_6191
timestamp 1668089732
transform 1 0 15840 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_6192
timestamp 1668089732
transform 1 0 15840 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_6193
timestamp 1668089732
transform 1 0 15840 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_6194
timestamp 1668089732
transform 1 0 15840 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_6195
timestamp 1668089732
transform 1 0 15840 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_6196
timestamp 1668089732
transform 1 0 15840 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_6197
timestamp 1668089732
transform 1 0 15840 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_6198
timestamp 1668089732
transform 1 0 15840 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_6199
timestamp 1668089732
transform 1 0 15840 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_6200
timestamp 1668089732
transform 1 0 16000 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_6201
timestamp 1668089732
transform 1 0 16000 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_6202
timestamp 1668089732
transform 1 0 16000 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_6203
timestamp 1668089732
transform 1 0 16000 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_6204
timestamp 1668089732
transform 1 0 16000 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_6205
timestamp 1668089732
transform 1 0 16000 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_6206
timestamp 1668089732
transform 1 0 16000 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_6207
timestamp 1668089732
transform 1 0 16000 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_6208
timestamp 1668089732
transform 1 0 16000 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_6209
timestamp 1668089732
transform 1 0 16000 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_6210
timestamp 1668089732
transform 1 0 16000 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_6211
timestamp 1668089732
transform 1 0 16000 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_6212
timestamp 1668089732
transform 1 0 16000 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_6213
timestamp 1668089732
transform 1 0 16000 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_6214
timestamp 1668089732
transform 1 0 16000 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_6215
timestamp 1668089732
transform 1 0 16000 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_6216
timestamp 1668089732
transform 1 0 16000 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_6217
timestamp 1668089732
transform 1 0 16000 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_6218
timestamp 1668089732
transform 1 0 16000 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_6219
timestamp 1668089732
transform 1 0 16000 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_6220
timestamp 1668089732
transform 1 0 16000 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_6221
timestamp 1668089732
transform 1 0 16000 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_6222
timestamp 1668089732
transform 1 0 16000 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_6223
timestamp 1668089732
transform 1 0 16000 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_6224
timestamp 1668089732
transform 1 0 16000 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_6225
timestamp 1668089732
transform 1 0 16000 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_6226
timestamp 1668089732
transform 1 0 16000 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_6227
timestamp 1668089732
transform 1 0 16000 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_6228
timestamp 1668089732
transform 1 0 16000 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_6229
timestamp 1668089732
transform 1 0 16000 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_6230
timestamp 1668089732
transform 1 0 16000 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_6231
timestamp 1668089732
transform 1 0 16000 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_6232
timestamp 1668089732
transform 1 0 16000 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_6233
timestamp 1668089732
transform 1 0 16000 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_6234
timestamp 1668089732
transform 1 0 16000 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_6235
timestamp 1668089732
transform 1 0 16000 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_6236
timestamp 1668089732
transform 1 0 16000 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_6237
timestamp 1668089732
transform 1 0 16000 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_6238
timestamp 1668089732
transform 1 0 16000 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_6239
timestamp 1668089732
transform 1 0 16000 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_6240
timestamp 1668089732
transform 1 0 16000 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_6241
timestamp 1668089732
transform 1 0 16000 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_6242
timestamp 1668089732
transform 1 0 16000 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_6243
timestamp 1668089732
transform 1 0 16000 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_6244
timestamp 1668089732
transform 1 0 16000 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_6245
timestamp 1668089732
transform 1 0 16000 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_6246
timestamp 1668089732
transform 1 0 16000 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_6247
timestamp 1668089732
transform 1 0 16000 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_6248
timestamp 1668089732
transform 1 0 16000 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_6249
timestamp 1668089732
transform 1 0 16000 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_6250
timestamp 1668089732
transform 1 0 16000 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_6251
timestamp 1668089732
transform 1 0 16000 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_6252
timestamp 1668089732
transform 1 0 16000 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_6253
timestamp 1668089732
transform 1 0 16000 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_6254
timestamp 1668089732
transform 1 0 16000 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_6255
timestamp 1668089732
transform 1 0 16000 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_6256
timestamp 1668089732
transform 1 0 16000 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_6257
timestamp 1668089732
transform 1 0 16000 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_6258
timestamp 1668089732
transform 1 0 16000 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_6259
timestamp 1668089732
transform 1 0 16000 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_6260
timestamp 1668089732
transform 1 0 16000 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_6261
timestamp 1668089732
transform 1 0 16000 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_6262
timestamp 1668089732
transform 1 0 16160 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_6263
timestamp 1668089732
transform 1 0 16160 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_6264
timestamp 1668089732
transform 1 0 16160 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_6265
timestamp 1668089732
transform 1 0 16160 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_6266
timestamp 1668089732
transform 1 0 16160 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_6267
timestamp 1668089732
transform 1 0 16160 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_6268
timestamp 1668089732
transform 1 0 16160 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_6269
timestamp 1668089732
transform 1 0 16160 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_6270
timestamp 1668089732
transform 1 0 16160 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_6271
timestamp 1668089732
transform 1 0 16160 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_6272
timestamp 1668089732
transform 1 0 16160 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_6273
timestamp 1668089732
transform 1 0 16160 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_6274
timestamp 1668089732
transform 1 0 16160 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_6275
timestamp 1668089732
transform 1 0 16160 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_6276
timestamp 1668089732
transform 1 0 16160 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_6277
timestamp 1668089732
transform 1 0 16160 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_6278
timestamp 1668089732
transform 1 0 16160 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_6279
timestamp 1668089732
transform 1 0 16160 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_6280
timestamp 1668089732
transform 1 0 16160 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_6281
timestamp 1668089732
transform 1 0 16160 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_6282
timestamp 1668089732
transform 1 0 16160 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_6283
timestamp 1668089732
transform 1 0 16160 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_6284
timestamp 1668089732
transform 1 0 16160 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_6285
timestamp 1668089732
transform 1 0 16160 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_6286
timestamp 1668089732
transform 1 0 16160 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_6287
timestamp 1668089732
transform 1 0 16160 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_6288
timestamp 1668089732
transform 1 0 16160 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_6289
timestamp 1668089732
transform 1 0 16160 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_6290
timestamp 1668089732
transform 1 0 16160 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_6291
timestamp 1668089732
transform 1 0 16160 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_6292
timestamp 1668089732
transform 1 0 16160 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_6293
timestamp 1668089732
transform 1 0 16160 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_6294
timestamp 1668089732
transform 1 0 16160 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_6295
timestamp 1668089732
transform 1 0 16160 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_6296
timestamp 1668089732
transform 1 0 16160 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_6297
timestamp 1668089732
transform 1 0 16160 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_6298
timestamp 1668089732
transform 1 0 16160 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_6299
timestamp 1668089732
transform 1 0 16160 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_6300
timestamp 1668089732
transform 1 0 16160 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_6301
timestamp 1668089732
transform 1 0 16160 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_6302
timestamp 1668089732
transform 1 0 16160 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_6303
timestamp 1668089732
transform 1 0 16160 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_6304
timestamp 1668089732
transform 1 0 16160 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_6305
timestamp 1668089732
transform 1 0 16160 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_6306
timestamp 1668089732
transform 1 0 16160 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_6307
timestamp 1668089732
transform 1 0 16160 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_6308
timestamp 1668089732
transform 1 0 16160 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_6309
timestamp 1668089732
transform 1 0 16160 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_6310
timestamp 1668089732
transform 1 0 16160 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_6311
timestamp 1668089732
transform 1 0 16160 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_6312
timestamp 1668089732
transform 1 0 16160 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_6313
timestamp 1668089732
transform 1 0 16160 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_6314
timestamp 1668089732
transform 1 0 16160 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_6315
timestamp 1668089732
transform 1 0 16160 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_6316
timestamp 1668089732
transform 1 0 16160 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_6317
timestamp 1668089732
transform 1 0 16160 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_6318
timestamp 1668089732
transform 1 0 16160 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_6319
timestamp 1668089732
transform 1 0 16160 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_6320
timestamp 1668089732
transform 1 0 16160 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_6321
timestamp 1668089732
transform 1 0 16160 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_6322
timestamp 1668089732
transform 1 0 16160 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_6323
timestamp 1668089732
transform 1 0 16160 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_6324
timestamp 1668089732
transform 1 0 16320 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_6325
timestamp 1668089732
transform 1 0 16320 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_6326
timestamp 1668089732
transform 1 0 16320 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_6327
timestamp 1668089732
transform 1 0 16320 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_6328
timestamp 1668089732
transform 1 0 16320 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_6329
timestamp 1668089732
transform 1 0 16320 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_6330
timestamp 1668089732
transform 1 0 16320 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_6331
timestamp 1668089732
transform 1 0 16320 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_6332
timestamp 1668089732
transform 1 0 16320 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_6333
timestamp 1668089732
transform 1 0 16320 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_6334
timestamp 1668089732
transform 1 0 16320 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_6335
timestamp 1668089732
transform 1 0 16320 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_6336
timestamp 1668089732
transform 1 0 16320 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_6337
timestamp 1668089732
transform 1 0 16320 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_6338
timestamp 1668089732
transform 1 0 16320 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_6339
timestamp 1668089732
transform 1 0 16320 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_6340
timestamp 1668089732
transform 1 0 16320 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_6341
timestamp 1668089732
transform 1 0 16320 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_6342
timestamp 1668089732
transform 1 0 16320 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_6343
timestamp 1668089732
transform 1 0 16320 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_6344
timestamp 1668089732
transform 1 0 16320 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_6345
timestamp 1668089732
transform 1 0 16320 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_6346
timestamp 1668089732
transform 1 0 16320 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_6347
timestamp 1668089732
transform 1 0 16320 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_6348
timestamp 1668089732
transform 1 0 16320 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_6349
timestamp 1668089732
transform 1 0 16320 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_6350
timestamp 1668089732
transform 1 0 16320 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_6351
timestamp 1668089732
transform 1 0 16320 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_6352
timestamp 1668089732
transform 1 0 16320 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_6353
timestamp 1668089732
transform 1 0 16320 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_6354
timestamp 1668089732
transform 1 0 16320 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_6355
timestamp 1668089732
transform 1 0 16320 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_6356
timestamp 1668089732
transform 1 0 16320 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_6357
timestamp 1668089732
transform 1 0 16320 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_6358
timestamp 1668089732
transform 1 0 16320 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_6359
timestamp 1668089732
transform 1 0 16320 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_6360
timestamp 1668089732
transform 1 0 16320 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_6361
timestamp 1668089732
transform 1 0 16320 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_6362
timestamp 1668089732
transform 1 0 16320 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_6363
timestamp 1668089732
transform 1 0 16320 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_6364
timestamp 1668089732
transform 1 0 16320 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_6365
timestamp 1668089732
transform 1 0 16320 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_6366
timestamp 1668089732
transform 1 0 16320 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_6367
timestamp 1668089732
transform 1 0 16320 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_6368
timestamp 1668089732
transform 1 0 16320 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_6369
timestamp 1668089732
transform 1 0 16320 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_6370
timestamp 1668089732
transform 1 0 16320 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_6371
timestamp 1668089732
transform 1 0 16320 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_6372
timestamp 1668089732
transform 1 0 16320 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_6373
timestamp 1668089732
transform 1 0 16320 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_6374
timestamp 1668089732
transform 1 0 16320 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_6375
timestamp 1668089732
transform 1 0 16320 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_6376
timestamp 1668089732
transform 1 0 16320 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_6377
timestamp 1668089732
transform 1 0 16320 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_6378
timestamp 1668089732
transform 1 0 16320 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_6379
timestamp 1668089732
transform 1 0 16320 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_6380
timestamp 1668089732
transform 1 0 16320 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_6381
timestamp 1668089732
transform 1 0 16320 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_6382
timestamp 1668089732
transform 1 0 16320 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_6383
timestamp 1668089732
transform 1 0 16320 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_6384
timestamp 1668089732
transform 1 0 16320 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_6385
timestamp 1668089732
transform 1 0 16320 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_6386
timestamp 1668089732
transform 1 0 16480 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_6387
timestamp 1668089732
transform 1 0 16480 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_6388
timestamp 1668089732
transform 1 0 16480 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_6389
timestamp 1668089732
transform 1 0 16480 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_6390
timestamp 1668089732
transform 1 0 16480 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_6391
timestamp 1668089732
transform 1 0 16480 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_6392
timestamp 1668089732
transform 1 0 16480 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_6393
timestamp 1668089732
transform 1 0 16480 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_6394
timestamp 1668089732
transform 1 0 16480 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_6395
timestamp 1668089732
transform 1 0 16480 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_6396
timestamp 1668089732
transform 1 0 16480 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_6397
timestamp 1668089732
transform 1 0 16480 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_6398
timestamp 1668089732
transform 1 0 16480 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_6399
timestamp 1668089732
transform 1 0 16480 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_6400
timestamp 1668089732
transform 1 0 16480 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_6401
timestamp 1668089732
transform 1 0 16480 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_6402
timestamp 1668089732
transform 1 0 16480 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_6403
timestamp 1668089732
transform 1 0 16480 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_6404
timestamp 1668089732
transform 1 0 16480 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_6405
timestamp 1668089732
transform 1 0 16480 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_6406
timestamp 1668089732
transform 1 0 16480 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_6407
timestamp 1668089732
transform 1 0 16480 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_6408
timestamp 1668089732
transform 1 0 16480 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_6409
timestamp 1668089732
transform 1 0 16480 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_6410
timestamp 1668089732
transform 1 0 16480 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_6411
timestamp 1668089732
transform 1 0 16480 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_6412
timestamp 1668089732
transform 1 0 16480 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_6413
timestamp 1668089732
transform 1 0 16480 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_6414
timestamp 1668089732
transform 1 0 16480 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_6415
timestamp 1668089732
transform 1 0 16480 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_6416
timestamp 1668089732
transform 1 0 16480 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_6417
timestamp 1668089732
transform 1 0 16480 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_6418
timestamp 1668089732
transform 1 0 16480 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_6419
timestamp 1668089732
transform 1 0 16480 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_6420
timestamp 1668089732
transform 1 0 16480 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_6421
timestamp 1668089732
transform 1 0 16480 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_6422
timestamp 1668089732
transform 1 0 16480 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_6423
timestamp 1668089732
transform 1 0 16480 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_6424
timestamp 1668089732
transform 1 0 16480 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_6425
timestamp 1668089732
transform 1 0 16480 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_6426
timestamp 1668089732
transform 1 0 16480 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_6427
timestamp 1668089732
transform 1 0 16480 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_6428
timestamp 1668089732
transform 1 0 16480 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_6429
timestamp 1668089732
transform 1 0 16480 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_6430
timestamp 1668089732
transform 1 0 16480 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_6431
timestamp 1668089732
transform 1 0 16480 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_6432
timestamp 1668089732
transform 1 0 16480 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_6433
timestamp 1668089732
transform 1 0 16480 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_6434
timestamp 1668089732
transform 1 0 16480 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_6435
timestamp 1668089732
transform 1 0 16480 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_6436
timestamp 1668089732
transform 1 0 16480 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_6437
timestamp 1668089732
transform 1 0 16480 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_6438
timestamp 1668089732
transform 1 0 16480 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_6439
timestamp 1668089732
transform 1 0 16480 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_6440
timestamp 1668089732
transform 1 0 16480 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_6441
timestamp 1668089732
transform 1 0 16480 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_6442
timestamp 1668089732
transform 1 0 16480 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_6443
timestamp 1668089732
transform 1 0 16480 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_6444
timestamp 1668089732
transform 1 0 16480 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_6445
timestamp 1668089732
transform 1 0 16480 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_6446
timestamp 1668089732
transform 1 0 16480 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_6447
timestamp 1668089732
transform 1 0 16480 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_6448
timestamp 1668089732
transform 1 0 16640 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_6449
timestamp 1668089732
transform 1 0 16640 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_6450
timestamp 1668089732
transform 1 0 16640 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_6451
timestamp 1668089732
transform 1 0 16640 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_6452
timestamp 1668089732
transform 1 0 16640 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_6453
timestamp 1668089732
transform 1 0 16640 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_6454
timestamp 1668089732
transform 1 0 16640 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_6455
timestamp 1668089732
transform 1 0 16640 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_6456
timestamp 1668089732
transform 1 0 16640 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_6457
timestamp 1668089732
transform 1 0 16640 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_6458
timestamp 1668089732
transform 1 0 16640 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_6459
timestamp 1668089732
transform 1 0 16640 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_6460
timestamp 1668089732
transform 1 0 16640 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_6461
timestamp 1668089732
transform 1 0 16640 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_6462
timestamp 1668089732
transform 1 0 16640 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_6463
timestamp 1668089732
transform 1 0 16640 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_6464
timestamp 1668089732
transform 1 0 16640 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_6465
timestamp 1668089732
transform 1 0 16640 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_6466
timestamp 1668089732
transform 1 0 16640 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_6467
timestamp 1668089732
transform 1 0 16640 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_6468
timestamp 1668089732
transform 1 0 16640 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_6469
timestamp 1668089732
transform 1 0 16640 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_6470
timestamp 1668089732
transform 1 0 16640 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_6471
timestamp 1668089732
transform 1 0 16640 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_6472
timestamp 1668089732
transform 1 0 16640 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_6473
timestamp 1668089732
transform 1 0 16640 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_6474
timestamp 1668089732
transform 1 0 16640 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_6475
timestamp 1668089732
transform 1 0 16640 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_6476
timestamp 1668089732
transform 1 0 16640 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_6477
timestamp 1668089732
transform 1 0 16640 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_6478
timestamp 1668089732
transform 1 0 16640 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_6479
timestamp 1668089732
transform 1 0 16640 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_6480
timestamp 1668089732
transform 1 0 16640 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_6481
timestamp 1668089732
transform 1 0 16640 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_6482
timestamp 1668089732
transform 1 0 16640 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_6483
timestamp 1668089732
transform 1 0 16640 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_6484
timestamp 1668089732
transform 1 0 16640 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_6485
timestamp 1668089732
transform 1 0 16640 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_6486
timestamp 1668089732
transform 1 0 16640 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_6487
timestamp 1668089732
transform 1 0 16640 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_6488
timestamp 1668089732
transform 1 0 16640 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_6489
timestamp 1668089732
transform 1 0 16640 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_6490
timestamp 1668089732
transform 1 0 16640 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_6491
timestamp 1668089732
transform 1 0 16640 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_6492
timestamp 1668089732
transform 1 0 16640 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_6493
timestamp 1668089732
transform 1 0 16640 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_6494
timestamp 1668089732
transform 1 0 16640 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_6495
timestamp 1668089732
transform 1 0 16640 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_6496
timestamp 1668089732
transform 1 0 16640 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_6497
timestamp 1668089732
transform 1 0 16640 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_6498
timestamp 1668089732
transform 1 0 16640 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_6499
timestamp 1668089732
transform 1 0 16640 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_6500
timestamp 1668089732
transform 1 0 16640 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_6501
timestamp 1668089732
transform 1 0 16640 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_6502
timestamp 1668089732
transform 1 0 16640 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_6503
timestamp 1668089732
transform 1 0 16640 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_6504
timestamp 1668089732
transform 1 0 16640 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_6505
timestamp 1668089732
transform 1 0 16640 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_6506
timestamp 1668089732
transform 1 0 16640 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_6507
timestamp 1668089732
transform 1 0 16640 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_6508
timestamp 1668089732
transform 1 0 16640 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_6509
timestamp 1668089732
transform 1 0 16640 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_6510
timestamp 1668089732
transform 1 0 16800 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_6511
timestamp 1668089732
transform 1 0 16800 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_6512
timestamp 1668089732
transform 1 0 16800 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_6513
timestamp 1668089732
transform 1 0 16800 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_6514
timestamp 1668089732
transform 1 0 16800 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_6515
timestamp 1668089732
transform 1 0 16800 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_6516
timestamp 1668089732
transform 1 0 16800 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_6517
timestamp 1668089732
transform 1 0 16800 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_6518
timestamp 1668089732
transform 1 0 16800 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_6519
timestamp 1668089732
transform 1 0 16800 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_6520
timestamp 1668089732
transform 1 0 16800 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_6521
timestamp 1668089732
transform 1 0 16800 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_6522
timestamp 1668089732
transform 1 0 16800 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_6523
timestamp 1668089732
transform 1 0 16800 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_6524
timestamp 1668089732
transform 1 0 16800 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_6525
timestamp 1668089732
transform 1 0 16800 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_6526
timestamp 1668089732
transform 1 0 16800 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_6527
timestamp 1668089732
transform 1 0 16800 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_6528
timestamp 1668089732
transform 1 0 16800 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_6529
timestamp 1668089732
transform 1 0 16800 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_6530
timestamp 1668089732
transform 1 0 16800 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_6531
timestamp 1668089732
transform 1 0 16800 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_6532
timestamp 1668089732
transform 1 0 16800 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_6533
timestamp 1668089732
transform 1 0 16800 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_6534
timestamp 1668089732
transform 1 0 16800 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_6535
timestamp 1668089732
transform 1 0 16800 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_6536
timestamp 1668089732
transform 1 0 16800 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_6537
timestamp 1668089732
transform 1 0 16800 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_6538
timestamp 1668089732
transform 1 0 16800 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_6539
timestamp 1668089732
transform 1 0 16800 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_6540
timestamp 1668089732
transform 1 0 16800 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_6541
timestamp 1668089732
transform 1 0 16800 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_6542
timestamp 1668089732
transform 1 0 16800 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_6543
timestamp 1668089732
transform 1 0 16800 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_6544
timestamp 1668089732
transform 1 0 16800 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_6545
timestamp 1668089732
transform 1 0 16800 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_6546
timestamp 1668089732
transform 1 0 16800 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_6547
timestamp 1668089732
transform 1 0 16800 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_6548
timestamp 1668089732
transform 1 0 16800 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_6549
timestamp 1668089732
transform 1 0 16800 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_6550
timestamp 1668089732
transform 1 0 16800 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_6551
timestamp 1668089732
transform 1 0 16800 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_6552
timestamp 1668089732
transform 1 0 16800 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_6553
timestamp 1668089732
transform 1 0 16800 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_6554
timestamp 1668089732
transform 1 0 16800 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_6555
timestamp 1668089732
transform 1 0 16800 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_6556
timestamp 1668089732
transform 1 0 16800 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_6557
timestamp 1668089732
transform 1 0 16800 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_6558
timestamp 1668089732
transform 1 0 16800 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_6559
timestamp 1668089732
transform 1 0 16800 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_6560
timestamp 1668089732
transform 1 0 16800 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_6561
timestamp 1668089732
transform 1 0 16800 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_6562
timestamp 1668089732
transform 1 0 16800 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_6563
timestamp 1668089732
transform 1 0 16800 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_6564
timestamp 1668089732
transform 1 0 16800 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_6565
timestamp 1668089732
transform 1 0 16800 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_6566
timestamp 1668089732
transform 1 0 16800 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_6567
timestamp 1668089732
transform 1 0 16800 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_6568
timestamp 1668089732
transform 1 0 16800 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_6569
timestamp 1668089732
transform 1 0 16800 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_6570
timestamp 1668089732
transform 1 0 16800 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_6571
timestamp 1668089732
transform 1 0 16800 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_6572
timestamp 1668089732
transform 1 0 16960 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_6573
timestamp 1668089732
transform 1 0 16960 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_6574
timestamp 1668089732
transform 1 0 16960 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_6575
timestamp 1668089732
transform 1 0 16960 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_6576
timestamp 1668089732
transform 1 0 16960 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_6577
timestamp 1668089732
transform 1 0 16960 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_6578
timestamp 1668089732
transform 1 0 16960 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_6579
timestamp 1668089732
transform 1 0 16960 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_6580
timestamp 1668089732
transform 1 0 16960 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_6581
timestamp 1668089732
transform 1 0 16960 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_6582
timestamp 1668089732
transform 1 0 16960 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_6583
timestamp 1668089732
transform 1 0 16960 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_6584
timestamp 1668089732
transform 1 0 16960 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_6585
timestamp 1668089732
transform 1 0 16960 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_6586
timestamp 1668089732
transform 1 0 16960 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_6587
timestamp 1668089732
transform 1 0 16960 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_6588
timestamp 1668089732
transform 1 0 16960 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_6589
timestamp 1668089732
transform 1 0 16960 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_6590
timestamp 1668089732
transform 1 0 16960 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_6591
timestamp 1668089732
transform 1 0 16960 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_6592
timestamp 1668089732
transform 1 0 16960 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_6593
timestamp 1668089732
transform 1 0 16960 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_6594
timestamp 1668089732
transform 1 0 16960 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_6595
timestamp 1668089732
transform 1 0 16960 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_6596
timestamp 1668089732
transform 1 0 16960 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_6597
timestamp 1668089732
transform 1 0 16960 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_6598
timestamp 1668089732
transform 1 0 16960 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_6599
timestamp 1668089732
transform 1 0 16960 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_6600
timestamp 1668089732
transform 1 0 16960 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_6601
timestamp 1668089732
transform 1 0 16960 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_6602
timestamp 1668089732
transform 1 0 16960 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_6603
timestamp 1668089732
transform 1 0 16960 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_6604
timestamp 1668089732
transform 1 0 16960 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_6605
timestamp 1668089732
transform 1 0 16960 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_6606
timestamp 1668089732
transform 1 0 16960 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_6607
timestamp 1668089732
transform 1 0 16960 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_6608
timestamp 1668089732
transform 1 0 16960 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_6609
timestamp 1668089732
transform 1 0 16960 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_6610
timestamp 1668089732
transform 1 0 16960 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_6611
timestamp 1668089732
transform 1 0 16960 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_6612
timestamp 1668089732
transform 1 0 16960 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_6613
timestamp 1668089732
transform 1 0 16960 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_6614
timestamp 1668089732
transform 1 0 16960 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_6615
timestamp 1668089732
transform 1 0 16960 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_6616
timestamp 1668089732
transform 1 0 16960 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_6617
timestamp 1668089732
transform 1 0 16960 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_6618
timestamp 1668089732
transform 1 0 16960 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_6619
timestamp 1668089732
transform 1 0 16960 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_6620
timestamp 1668089732
transform 1 0 16960 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_6621
timestamp 1668089732
transform 1 0 16960 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_6622
timestamp 1668089732
transform 1 0 16960 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_6623
timestamp 1668089732
transform 1 0 16960 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_6624
timestamp 1668089732
transform 1 0 16960 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_6625
timestamp 1668089732
transform 1 0 16960 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_6626
timestamp 1668089732
transform 1 0 16960 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_6627
timestamp 1668089732
transform 1 0 16960 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_6628
timestamp 1668089732
transform 1 0 16960 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_6629
timestamp 1668089732
transform 1 0 16960 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_6630
timestamp 1668089732
transform 1 0 16960 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_6631
timestamp 1668089732
transform 1 0 16960 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_6632
timestamp 1668089732
transform 1 0 16960 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_6633
timestamp 1668089732
transform 1 0 16960 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_6634
timestamp 1668089732
transform 1 0 17120 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_6635
timestamp 1668089732
transform 1 0 17120 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_6636
timestamp 1668089732
transform 1 0 17120 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_6637
timestamp 1668089732
transform 1 0 17120 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_6638
timestamp 1668089732
transform 1 0 17120 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_6639
timestamp 1668089732
transform 1 0 17120 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_6640
timestamp 1668089732
transform 1 0 17120 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_6641
timestamp 1668089732
transform 1 0 17120 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_6642
timestamp 1668089732
transform 1 0 17120 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_6643
timestamp 1668089732
transform 1 0 17120 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_6644
timestamp 1668089732
transform 1 0 17120 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_6645
timestamp 1668089732
transform 1 0 17120 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_6646
timestamp 1668089732
transform 1 0 17120 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_6647
timestamp 1668089732
transform 1 0 17120 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_6648
timestamp 1668089732
transform 1 0 17120 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_6649
timestamp 1668089732
transform 1 0 17120 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_6650
timestamp 1668089732
transform 1 0 17120 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_6651
timestamp 1668089732
transform 1 0 17120 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_6652
timestamp 1668089732
transform 1 0 17120 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_6653
timestamp 1668089732
transform 1 0 17120 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_6654
timestamp 1668089732
transform 1 0 17120 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_6655
timestamp 1668089732
transform 1 0 17120 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_6656
timestamp 1668089732
transform 1 0 17120 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_6657
timestamp 1668089732
transform 1 0 17120 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_6658
timestamp 1668089732
transform 1 0 17120 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_6659
timestamp 1668089732
transform 1 0 17120 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_6660
timestamp 1668089732
transform 1 0 17120 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_6661
timestamp 1668089732
transform 1 0 17120 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_6662
timestamp 1668089732
transform 1 0 17120 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_6663
timestamp 1668089732
transform 1 0 17120 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_6664
timestamp 1668089732
transform 1 0 17120 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_6665
timestamp 1668089732
transform 1 0 17120 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_6666
timestamp 1668089732
transform 1 0 17120 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_6667
timestamp 1668089732
transform 1 0 17120 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_6668
timestamp 1668089732
transform 1 0 17120 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_6669
timestamp 1668089732
transform 1 0 17120 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_6670
timestamp 1668089732
transform 1 0 17120 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_6671
timestamp 1668089732
transform 1 0 17120 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_6672
timestamp 1668089732
transform 1 0 17120 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_6673
timestamp 1668089732
transform 1 0 17120 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_6674
timestamp 1668089732
transform 1 0 17120 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_6675
timestamp 1668089732
transform 1 0 17120 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_6676
timestamp 1668089732
transform 1 0 17120 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_6677
timestamp 1668089732
transform 1 0 17120 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_6678
timestamp 1668089732
transform 1 0 17120 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_6679
timestamp 1668089732
transform 1 0 17120 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_6680
timestamp 1668089732
transform 1 0 17120 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_6681
timestamp 1668089732
transform 1 0 17120 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_6682
timestamp 1668089732
transform 1 0 17120 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_6683
timestamp 1668089732
transform 1 0 17120 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_6684
timestamp 1668089732
transform 1 0 17120 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_6685
timestamp 1668089732
transform 1 0 17120 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_6686
timestamp 1668089732
transform 1 0 17120 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_6687
timestamp 1668089732
transform 1 0 17120 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_6688
timestamp 1668089732
transform 1 0 17120 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_6689
timestamp 1668089732
transform 1 0 17120 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_6690
timestamp 1668089732
transform 1 0 17120 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_6691
timestamp 1668089732
transform 1 0 17120 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_6692
timestamp 1668089732
transform 1 0 17120 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_6693
timestamp 1668089732
transform 1 0 17120 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_6694
timestamp 1668089732
transform 1 0 17120 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_6695
timestamp 1668089732
transform 1 0 17120 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_6696
timestamp 1668089732
transform 1 0 17280 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_6697
timestamp 1668089732
transform 1 0 17280 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_6698
timestamp 1668089732
transform 1 0 17280 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_6699
timestamp 1668089732
transform 1 0 17280 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_6700
timestamp 1668089732
transform 1 0 17280 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_6701
timestamp 1668089732
transform 1 0 17280 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_6702
timestamp 1668089732
transform 1 0 17280 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_6703
timestamp 1668089732
transform 1 0 17280 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_6704
timestamp 1668089732
transform 1 0 17280 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_6705
timestamp 1668089732
transform 1 0 17280 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_6706
timestamp 1668089732
transform 1 0 17280 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_6707
timestamp 1668089732
transform 1 0 17280 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_6708
timestamp 1668089732
transform 1 0 17280 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_6709
timestamp 1668089732
transform 1 0 17280 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_6710
timestamp 1668089732
transform 1 0 17280 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_6711
timestamp 1668089732
transform 1 0 17280 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_6712
timestamp 1668089732
transform 1 0 17280 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_6713
timestamp 1668089732
transform 1 0 17280 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_6714
timestamp 1668089732
transform 1 0 17280 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_6715
timestamp 1668089732
transform 1 0 17280 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_6716
timestamp 1668089732
transform 1 0 17280 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_6717
timestamp 1668089732
transform 1 0 17280 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_6718
timestamp 1668089732
transform 1 0 17280 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_6719
timestamp 1668089732
transform 1 0 17280 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_6720
timestamp 1668089732
transform 1 0 17280 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_6721
timestamp 1668089732
transform 1 0 17280 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_6722
timestamp 1668089732
transform 1 0 17280 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_6723
timestamp 1668089732
transform 1 0 17280 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_6724
timestamp 1668089732
transform 1 0 17280 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_6725
timestamp 1668089732
transform 1 0 17280 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_6726
timestamp 1668089732
transform 1 0 17280 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_6727
timestamp 1668089732
transform 1 0 17280 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_6728
timestamp 1668089732
transform 1 0 17280 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_6729
timestamp 1668089732
transform 1 0 17280 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_6730
timestamp 1668089732
transform 1 0 17280 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_6731
timestamp 1668089732
transform 1 0 17280 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_6732
timestamp 1668089732
transform 1 0 17280 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_6733
timestamp 1668089732
transform 1 0 17280 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_6734
timestamp 1668089732
transform 1 0 17280 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_6735
timestamp 1668089732
transform 1 0 17280 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_6736
timestamp 1668089732
transform 1 0 17280 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_6737
timestamp 1668089732
transform 1 0 17280 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_6738
timestamp 1668089732
transform 1 0 17280 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_6739
timestamp 1668089732
transform 1 0 17280 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_6740
timestamp 1668089732
transform 1 0 17280 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_6741
timestamp 1668089732
transform 1 0 17280 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_6742
timestamp 1668089732
transform 1 0 17280 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_6743
timestamp 1668089732
transform 1 0 17280 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_6744
timestamp 1668089732
transform 1 0 17280 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_6745
timestamp 1668089732
transform 1 0 17280 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_6746
timestamp 1668089732
transform 1 0 17280 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_6747
timestamp 1668089732
transform 1 0 17280 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_6748
timestamp 1668089732
transform 1 0 17280 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_6749
timestamp 1668089732
transform 1 0 17280 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_6750
timestamp 1668089732
transform 1 0 17280 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_6751
timestamp 1668089732
transform 1 0 17280 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_6752
timestamp 1668089732
transform 1 0 17280 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_6753
timestamp 1668089732
transform 1 0 17280 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_6754
timestamp 1668089732
transform 1 0 17280 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_6755
timestamp 1668089732
transform 1 0 17280 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_6756
timestamp 1668089732
transform 1 0 17280 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_6757
timestamp 1668089732
transform 1 0 17280 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_6758
timestamp 1668089732
transform 1 0 17440 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_6759
timestamp 1668089732
transform 1 0 17440 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_6760
timestamp 1668089732
transform 1 0 17440 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_6761
timestamp 1668089732
transform 1 0 17440 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_6762
timestamp 1668089732
transform 1 0 17440 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_6763
timestamp 1668089732
transform 1 0 17440 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_6764
timestamp 1668089732
transform 1 0 17440 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_6765
timestamp 1668089732
transform 1 0 17440 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_6766
timestamp 1668089732
transform 1 0 17440 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_6767
timestamp 1668089732
transform 1 0 17440 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_6768
timestamp 1668089732
transform 1 0 17440 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_6769
timestamp 1668089732
transform 1 0 17440 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_6770
timestamp 1668089732
transform 1 0 17440 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_6771
timestamp 1668089732
transform 1 0 17440 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_6772
timestamp 1668089732
transform 1 0 17440 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_6773
timestamp 1668089732
transform 1 0 17440 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_6774
timestamp 1668089732
transform 1 0 17440 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_6775
timestamp 1668089732
transform 1 0 17440 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_6776
timestamp 1668089732
transform 1 0 17440 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_6777
timestamp 1668089732
transform 1 0 17440 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_6778
timestamp 1668089732
transform 1 0 17440 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_6779
timestamp 1668089732
transform 1 0 17440 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_6780
timestamp 1668089732
transform 1 0 17440 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_6781
timestamp 1668089732
transform 1 0 17440 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_6782
timestamp 1668089732
transform 1 0 17440 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_6783
timestamp 1668089732
transform 1 0 17440 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_6784
timestamp 1668089732
transform 1 0 17440 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_6785
timestamp 1668089732
transform 1 0 17440 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_6786
timestamp 1668089732
transform 1 0 17440 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_6787
timestamp 1668089732
transform 1 0 17440 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_6788
timestamp 1668089732
transform 1 0 17440 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_6789
timestamp 1668089732
transform 1 0 17440 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_6790
timestamp 1668089732
transform 1 0 17440 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_6791
timestamp 1668089732
transform 1 0 17440 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_6792
timestamp 1668089732
transform 1 0 17440 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_6793
timestamp 1668089732
transform 1 0 17440 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_6794
timestamp 1668089732
transform 1 0 17440 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_6795
timestamp 1668089732
transform 1 0 17440 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_6796
timestamp 1668089732
transform 1 0 17440 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_6797
timestamp 1668089732
transform 1 0 17440 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_6798
timestamp 1668089732
transform 1 0 17440 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_6799
timestamp 1668089732
transform 1 0 17440 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_6800
timestamp 1668089732
transform 1 0 17440 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_6801
timestamp 1668089732
transform 1 0 17440 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_6802
timestamp 1668089732
transform 1 0 17440 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_6803
timestamp 1668089732
transform 1 0 17440 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_6804
timestamp 1668089732
transform 1 0 17440 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_6805
timestamp 1668089732
transform 1 0 17440 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_6806
timestamp 1668089732
transform 1 0 17440 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_6807
timestamp 1668089732
transform 1 0 17440 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_6808
timestamp 1668089732
transform 1 0 17440 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_6809
timestamp 1668089732
transform 1 0 17440 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_6810
timestamp 1668089732
transform 1 0 17440 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_6811
timestamp 1668089732
transform 1 0 17440 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_6812
timestamp 1668089732
transform 1 0 17440 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_6813
timestamp 1668089732
transform 1 0 17440 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_6814
timestamp 1668089732
transform 1 0 17440 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_6815
timestamp 1668089732
transform 1 0 17440 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_6816
timestamp 1668089732
transform 1 0 17440 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_6817
timestamp 1668089732
transform 1 0 17440 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_6818
timestamp 1668089732
transform 1 0 17440 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_6819
timestamp 1668089732
transform 1 0 17440 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_6820
timestamp 1668089732
transform 1 0 17600 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_6821
timestamp 1668089732
transform 1 0 17600 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_6822
timestamp 1668089732
transform 1 0 17600 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_6823
timestamp 1668089732
transform 1 0 17600 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_6824
timestamp 1668089732
transform 1 0 17600 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_6825
timestamp 1668089732
transform 1 0 17600 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_6826
timestamp 1668089732
transform 1 0 17600 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_6827
timestamp 1668089732
transform 1 0 17600 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_6828
timestamp 1668089732
transform 1 0 17600 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_6829
timestamp 1668089732
transform 1 0 17600 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_6830
timestamp 1668089732
transform 1 0 17600 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_6831
timestamp 1668089732
transform 1 0 17600 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_6832
timestamp 1668089732
transform 1 0 17600 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_6833
timestamp 1668089732
transform 1 0 17600 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_6834
timestamp 1668089732
transform 1 0 17600 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_6835
timestamp 1668089732
transform 1 0 17600 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_6836
timestamp 1668089732
transform 1 0 17600 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_6837
timestamp 1668089732
transform 1 0 17600 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_6838
timestamp 1668089732
transform 1 0 17600 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_6839
timestamp 1668089732
transform 1 0 17600 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_6840
timestamp 1668089732
transform 1 0 17600 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_6841
timestamp 1668089732
transform 1 0 17600 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_6842
timestamp 1668089732
transform 1 0 17600 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_6843
timestamp 1668089732
transform 1 0 17600 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_6844
timestamp 1668089732
transform 1 0 17600 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_6845
timestamp 1668089732
transform 1 0 17600 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_6846
timestamp 1668089732
transform 1 0 17600 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_6847
timestamp 1668089732
transform 1 0 17600 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_6848
timestamp 1668089732
transform 1 0 17600 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_6849
timestamp 1668089732
transform 1 0 17600 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_6850
timestamp 1668089732
transform 1 0 17600 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_6851
timestamp 1668089732
transform 1 0 17600 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_6852
timestamp 1668089732
transform 1 0 17600 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_6853
timestamp 1668089732
transform 1 0 17600 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_6854
timestamp 1668089732
transform 1 0 17600 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_6855
timestamp 1668089732
transform 1 0 17600 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_6856
timestamp 1668089732
transform 1 0 17600 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_6857
timestamp 1668089732
transform 1 0 17600 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_6858
timestamp 1668089732
transform 1 0 17600 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_6859
timestamp 1668089732
transform 1 0 17600 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_6860
timestamp 1668089732
transform 1 0 17600 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_6861
timestamp 1668089732
transform 1 0 17600 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_6862
timestamp 1668089732
transform 1 0 17600 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_6863
timestamp 1668089732
transform 1 0 17600 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_6864
timestamp 1668089732
transform 1 0 17600 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_6865
timestamp 1668089732
transform 1 0 17600 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_6866
timestamp 1668089732
transform 1 0 17600 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_6867
timestamp 1668089732
transform 1 0 17600 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_6868
timestamp 1668089732
transform 1 0 17600 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_6869
timestamp 1668089732
transform 1 0 17600 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_6870
timestamp 1668089732
transform 1 0 17600 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_6871
timestamp 1668089732
transform 1 0 17600 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_6872
timestamp 1668089732
transform 1 0 17600 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_6873
timestamp 1668089732
transform 1 0 17600 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_6874
timestamp 1668089732
transform 1 0 17600 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_6875
timestamp 1668089732
transform 1 0 17600 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_6876
timestamp 1668089732
transform 1 0 17600 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_6877
timestamp 1668089732
transform 1 0 17600 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_6878
timestamp 1668089732
transform 1 0 17600 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_6879
timestamp 1668089732
transform 1 0 17600 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_6880
timestamp 1668089732
transform 1 0 17600 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_6881
timestamp 1668089732
transform 1 0 17600 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_6882
timestamp 1668089732
transform 1 0 17760 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_6883
timestamp 1668089732
transform 1 0 17760 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_6884
timestamp 1668089732
transform 1 0 17760 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_6885
timestamp 1668089732
transform 1 0 17760 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_6886
timestamp 1668089732
transform 1 0 17760 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_6887
timestamp 1668089732
transform 1 0 17760 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_6888
timestamp 1668089732
transform 1 0 17760 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_6889
timestamp 1668089732
transform 1 0 17760 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_6890
timestamp 1668089732
transform 1 0 17760 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_6891
timestamp 1668089732
transform 1 0 17760 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_6892
timestamp 1668089732
transform 1 0 17760 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_6893
timestamp 1668089732
transform 1 0 17760 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_6894
timestamp 1668089732
transform 1 0 17760 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_6895
timestamp 1668089732
transform 1 0 17760 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_6896
timestamp 1668089732
transform 1 0 17760 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_6897
timestamp 1668089732
transform 1 0 17760 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_6898
timestamp 1668089732
transform 1 0 17760 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_6899
timestamp 1668089732
transform 1 0 17760 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_6900
timestamp 1668089732
transform 1 0 17760 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_6901
timestamp 1668089732
transform 1 0 17760 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_6902
timestamp 1668089732
transform 1 0 17760 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_6903
timestamp 1668089732
transform 1 0 17760 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_6904
timestamp 1668089732
transform 1 0 17760 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_6905
timestamp 1668089732
transform 1 0 17760 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_6906
timestamp 1668089732
transform 1 0 17760 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_6907
timestamp 1668089732
transform 1 0 17760 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_6908
timestamp 1668089732
transform 1 0 17760 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_6909
timestamp 1668089732
transform 1 0 17760 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_6910
timestamp 1668089732
transform 1 0 17760 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_6911
timestamp 1668089732
transform 1 0 17760 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_6912
timestamp 1668089732
transform 1 0 17760 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_6913
timestamp 1668089732
transform 1 0 17760 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_6914
timestamp 1668089732
transform 1 0 17760 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_6915
timestamp 1668089732
transform 1 0 17760 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_6916
timestamp 1668089732
transform 1 0 17760 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_6917
timestamp 1668089732
transform 1 0 17760 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_6918
timestamp 1668089732
transform 1 0 17760 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_6919
timestamp 1668089732
transform 1 0 17760 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_6920
timestamp 1668089732
transform 1 0 17760 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_6921
timestamp 1668089732
transform 1 0 17760 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_6922
timestamp 1668089732
transform 1 0 17760 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_6923
timestamp 1668089732
transform 1 0 17760 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_6924
timestamp 1668089732
transform 1 0 17760 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_6925
timestamp 1668089732
transform 1 0 17760 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_6926
timestamp 1668089732
transform 1 0 17760 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_6927
timestamp 1668089732
transform 1 0 17760 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_6928
timestamp 1668089732
transform 1 0 17760 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_6929
timestamp 1668089732
transform 1 0 17760 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_6930
timestamp 1668089732
transform 1 0 17760 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_6931
timestamp 1668089732
transform 1 0 17760 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_6932
timestamp 1668089732
transform 1 0 17760 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_6933
timestamp 1668089732
transform 1 0 17760 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_6934
timestamp 1668089732
transform 1 0 17760 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_6935
timestamp 1668089732
transform 1 0 17760 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_6936
timestamp 1668089732
transform 1 0 17760 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_6937
timestamp 1668089732
transform 1 0 17760 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_6938
timestamp 1668089732
transform 1 0 17760 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_6939
timestamp 1668089732
transform 1 0 17760 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_6940
timestamp 1668089732
transform 1 0 17760 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_6941
timestamp 1668089732
transform 1 0 17760 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_6942
timestamp 1668089732
transform 1 0 17760 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_6943
timestamp 1668089732
transform 1 0 17760 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_6944
timestamp 1668089732
transform 1 0 17920 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_6945
timestamp 1668089732
transform 1 0 17920 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_6946
timestamp 1668089732
transform 1 0 17920 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_6947
timestamp 1668089732
transform 1 0 17920 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_6948
timestamp 1668089732
transform 1 0 17920 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_6949
timestamp 1668089732
transform 1 0 17920 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_6950
timestamp 1668089732
transform 1 0 17920 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_6951
timestamp 1668089732
transform 1 0 17920 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_6952
timestamp 1668089732
transform 1 0 17920 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_6953
timestamp 1668089732
transform 1 0 17920 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_6954
timestamp 1668089732
transform 1 0 17920 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_6955
timestamp 1668089732
transform 1 0 17920 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_6956
timestamp 1668089732
transform 1 0 17920 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_6957
timestamp 1668089732
transform 1 0 17920 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_6958
timestamp 1668089732
transform 1 0 17920 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_6959
timestamp 1668089732
transform 1 0 17920 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_6960
timestamp 1668089732
transform 1 0 17920 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_6961
timestamp 1668089732
transform 1 0 17920 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_6962
timestamp 1668089732
transform 1 0 17920 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_6963
timestamp 1668089732
transform 1 0 17920 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_6964
timestamp 1668089732
transform 1 0 17920 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_6965
timestamp 1668089732
transform 1 0 17920 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_6966
timestamp 1668089732
transform 1 0 17920 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_6967
timestamp 1668089732
transform 1 0 17920 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_6968
timestamp 1668089732
transform 1 0 17920 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_6969
timestamp 1668089732
transform 1 0 17920 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_6970
timestamp 1668089732
transform 1 0 17920 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_6971
timestamp 1668089732
transform 1 0 17920 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_6972
timestamp 1668089732
transform 1 0 17920 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_6973
timestamp 1668089732
transform 1 0 17920 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_6974
timestamp 1668089732
transform 1 0 17920 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_6975
timestamp 1668089732
transform 1 0 17920 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_6976
timestamp 1668089732
transform 1 0 17920 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_6977
timestamp 1668089732
transform 1 0 17920 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_6978
timestamp 1668089732
transform 1 0 17920 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_6979
timestamp 1668089732
transform 1 0 17920 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_6980
timestamp 1668089732
transform 1 0 17920 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_6981
timestamp 1668089732
transform 1 0 17920 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_6982
timestamp 1668089732
transform 1 0 17920 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_6983
timestamp 1668089732
transform 1 0 17920 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_6984
timestamp 1668089732
transform 1 0 17920 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_6985
timestamp 1668089732
transform 1 0 17920 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_6986
timestamp 1668089732
transform 1 0 17920 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_6987
timestamp 1668089732
transform 1 0 17920 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_6988
timestamp 1668089732
transform 1 0 17920 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_6989
timestamp 1668089732
transform 1 0 17920 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_6990
timestamp 1668089732
transform 1 0 17920 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_6991
timestamp 1668089732
transform 1 0 17920 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_6992
timestamp 1668089732
transform 1 0 17920 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_6993
timestamp 1668089732
transform 1 0 17920 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_6994
timestamp 1668089732
transform 1 0 17920 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_6995
timestamp 1668089732
transform 1 0 17920 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_6996
timestamp 1668089732
transform 1 0 17920 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_6997
timestamp 1668089732
transform 1 0 17920 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_6998
timestamp 1668089732
transform 1 0 17920 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_6999
timestamp 1668089732
transform 1 0 17920 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_7000
timestamp 1668089732
transform 1 0 17920 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_7001
timestamp 1668089732
transform 1 0 17920 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_7002
timestamp 1668089732
transform 1 0 17920 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_7003
timestamp 1668089732
transform 1 0 17920 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_7004
timestamp 1668089732
transform 1 0 17920 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_7005
timestamp 1668089732
transform 1 0 17920 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_7006
timestamp 1668089732
transform 1 0 18080 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_7007
timestamp 1668089732
transform 1 0 18080 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_7008
timestamp 1668089732
transform 1 0 18080 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_7009
timestamp 1668089732
transform 1 0 18080 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_7010
timestamp 1668089732
transform 1 0 18080 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_7011
timestamp 1668089732
transform 1 0 18080 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_7012
timestamp 1668089732
transform 1 0 18080 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_7013
timestamp 1668089732
transform 1 0 18080 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_7014
timestamp 1668089732
transform 1 0 18080 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_7015
timestamp 1668089732
transform 1 0 18080 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_7016
timestamp 1668089732
transform 1 0 18080 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_7017
timestamp 1668089732
transform 1 0 18080 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_7018
timestamp 1668089732
transform 1 0 18080 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_7019
timestamp 1668089732
transform 1 0 18080 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_7020
timestamp 1668089732
transform 1 0 18080 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_7021
timestamp 1668089732
transform 1 0 18080 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_7022
timestamp 1668089732
transform 1 0 18080 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_7023
timestamp 1668089732
transform 1 0 18080 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_7024
timestamp 1668089732
transform 1 0 18080 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_7025
timestamp 1668089732
transform 1 0 18080 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_7026
timestamp 1668089732
transform 1 0 18080 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_7027
timestamp 1668089732
transform 1 0 18080 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_7028
timestamp 1668089732
transform 1 0 18080 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_7029
timestamp 1668089732
transform 1 0 18080 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_7030
timestamp 1668089732
transform 1 0 18080 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_7031
timestamp 1668089732
transform 1 0 18080 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_7032
timestamp 1668089732
transform 1 0 18080 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_7033
timestamp 1668089732
transform 1 0 18080 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_7034
timestamp 1668089732
transform 1 0 18080 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_7035
timestamp 1668089732
transform 1 0 18080 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_7036
timestamp 1668089732
transform 1 0 18080 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_7037
timestamp 1668089732
transform 1 0 18080 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_7038
timestamp 1668089732
transform 1 0 18080 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_7039
timestamp 1668089732
transform 1 0 18080 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_7040
timestamp 1668089732
transform 1 0 18080 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_7041
timestamp 1668089732
transform 1 0 18080 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_7042
timestamp 1668089732
transform 1 0 18080 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_7043
timestamp 1668089732
transform 1 0 18080 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_7044
timestamp 1668089732
transform 1 0 18080 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_7045
timestamp 1668089732
transform 1 0 18080 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_7046
timestamp 1668089732
transform 1 0 18080 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_7047
timestamp 1668089732
transform 1 0 18080 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_7048
timestamp 1668089732
transform 1 0 18080 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_7049
timestamp 1668089732
transform 1 0 18080 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_7050
timestamp 1668089732
transform 1 0 18080 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_7051
timestamp 1668089732
transform 1 0 18080 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_7052
timestamp 1668089732
transform 1 0 18080 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_7053
timestamp 1668089732
transform 1 0 18080 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_7054
timestamp 1668089732
transform 1 0 18080 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_7055
timestamp 1668089732
transform 1 0 18080 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_7056
timestamp 1668089732
transform 1 0 18080 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_7057
timestamp 1668089732
transform 1 0 18080 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_7058
timestamp 1668089732
transform 1 0 18080 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_7059
timestamp 1668089732
transform 1 0 18080 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_7060
timestamp 1668089732
transform 1 0 18080 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_7061
timestamp 1668089732
transform 1 0 18080 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_7062
timestamp 1668089732
transform 1 0 18080 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_7063
timestamp 1668089732
transform 1 0 18080 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_7064
timestamp 1668089732
transform 1 0 18080 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_7065
timestamp 1668089732
transform 1 0 18080 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_7066
timestamp 1668089732
transform 1 0 18080 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_7067
timestamp 1668089732
transform 1 0 18080 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_7068
timestamp 1668089732
transform 1 0 18240 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_7069
timestamp 1668089732
transform 1 0 18240 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_7070
timestamp 1668089732
transform 1 0 18240 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_7071
timestamp 1668089732
transform 1 0 18240 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_7072
timestamp 1668089732
transform 1 0 18240 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_7073
timestamp 1668089732
transform 1 0 18240 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_7074
timestamp 1668089732
transform 1 0 18240 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_7075
timestamp 1668089732
transform 1 0 18240 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_7076
timestamp 1668089732
transform 1 0 18240 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_7077
timestamp 1668089732
transform 1 0 18240 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_7078
timestamp 1668089732
transform 1 0 18240 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_7079
timestamp 1668089732
transform 1 0 18240 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_7080
timestamp 1668089732
transform 1 0 18240 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_7081
timestamp 1668089732
transform 1 0 18240 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_7082
timestamp 1668089732
transform 1 0 18240 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_7083
timestamp 1668089732
transform 1 0 18240 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_7084
timestamp 1668089732
transform 1 0 18240 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_7085
timestamp 1668089732
transform 1 0 18240 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_7086
timestamp 1668089732
transform 1 0 18240 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_7087
timestamp 1668089732
transform 1 0 18240 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_7088
timestamp 1668089732
transform 1 0 18240 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_7089
timestamp 1668089732
transform 1 0 18240 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_7090
timestamp 1668089732
transform 1 0 18240 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_7091
timestamp 1668089732
transform 1 0 18240 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_7092
timestamp 1668089732
transform 1 0 18240 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_7093
timestamp 1668089732
transform 1 0 18240 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_7094
timestamp 1668089732
transform 1 0 18240 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_7095
timestamp 1668089732
transform 1 0 18240 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_7096
timestamp 1668089732
transform 1 0 18240 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_7097
timestamp 1668089732
transform 1 0 18240 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_7098
timestamp 1668089732
transform 1 0 18240 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_7099
timestamp 1668089732
transform 1 0 18240 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_7100
timestamp 1668089732
transform 1 0 18240 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_7101
timestamp 1668089732
transform 1 0 18240 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_7102
timestamp 1668089732
transform 1 0 18240 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_7103
timestamp 1668089732
transform 1 0 18240 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_7104
timestamp 1668089732
transform 1 0 18240 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_7105
timestamp 1668089732
transform 1 0 18240 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_7106
timestamp 1668089732
transform 1 0 18240 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_7107
timestamp 1668089732
transform 1 0 18240 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_7108
timestamp 1668089732
transform 1 0 18240 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_7109
timestamp 1668089732
transform 1 0 18240 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_7110
timestamp 1668089732
transform 1 0 18240 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_7111
timestamp 1668089732
transform 1 0 18240 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_7112
timestamp 1668089732
transform 1 0 18240 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_7113
timestamp 1668089732
transform 1 0 18240 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_7114
timestamp 1668089732
transform 1 0 18240 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_7115
timestamp 1668089732
transform 1 0 18240 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_7116
timestamp 1668089732
transform 1 0 18240 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_7117
timestamp 1668089732
transform 1 0 18240 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_7118
timestamp 1668089732
transform 1 0 18240 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_7119
timestamp 1668089732
transform 1 0 18240 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_7120
timestamp 1668089732
transform 1 0 18240 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_7121
timestamp 1668089732
transform 1 0 18240 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_7122
timestamp 1668089732
transform 1 0 18240 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_7123
timestamp 1668089732
transform 1 0 18240 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_7124
timestamp 1668089732
transform 1 0 18240 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_7125
timestamp 1668089732
transform 1 0 18240 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_7126
timestamp 1668089732
transform 1 0 18240 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_7127
timestamp 1668089732
transform 1 0 18240 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_7128
timestamp 1668089732
transform 1 0 18240 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_7129
timestamp 1668089732
transform 1 0 18240 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_7130
timestamp 1668089732
transform 1 0 18400 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_7131
timestamp 1668089732
transform 1 0 18400 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_7132
timestamp 1668089732
transform 1 0 18400 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_7133
timestamp 1668089732
transform 1 0 18400 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_7134
timestamp 1668089732
transform 1 0 18400 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_7135
timestamp 1668089732
transform 1 0 18400 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_7136
timestamp 1668089732
transform 1 0 18400 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_7137
timestamp 1668089732
transform 1 0 18400 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_7138
timestamp 1668089732
transform 1 0 18400 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_7139
timestamp 1668089732
transform 1 0 18400 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_7140
timestamp 1668089732
transform 1 0 18400 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_7141
timestamp 1668089732
transform 1 0 18400 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_7142
timestamp 1668089732
transform 1 0 18400 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_7143
timestamp 1668089732
transform 1 0 18400 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_7144
timestamp 1668089732
transform 1 0 18400 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_7145
timestamp 1668089732
transform 1 0 18400 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_7146
timestamp 1668089732
transform 1 0 18400 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_7147
timestamp 1668089732
transform 1 0 18400 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_7148
timestamp 1668089732
transform 1 0 18400 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_7149
timestamp 1668089732
transform 1 0 18400 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_7150
timestamp 1668089732
transform 1 0 18400 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_7151
timestamp 1668089732
transform 1 0 18400 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_7152
timestamp 1668089732
transform 1 0 18400 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_7153
timestamp 1668089732
transform 1 0 18400 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_7154
timestamp 1668089732
transform 1 0 18400 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_7155
timestamp 1668089732
transform 1 0 18400 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_7156
timestamp 1668089732
transform 1 0 18400 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_7157
timestamp 1668089732
transform 1 0 18400 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_7158
timestamp 1668089732
transform 1 0 18400 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_7159
timestamp 1668089732
transform 1 0 18400 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_7160
timestamp 1668089732
transform 1 0 18400 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_7161
timestamp 1668089732
transform 1 0 18400 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_7162
timestamp 1668089732
transform 1 0 18400 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_7163
timestamp 1668089732
transform 1 0 18400 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_7164
timestamp 1668089732
transform 1 0 18400 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_7165
timestamp 1668089732
transform 1 0 18400 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_7166
timestamp 1668089732
transform 1 0 18400 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_7167
timestamp 1668089732
transform 1 0 18400 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_7168
timestamp 1668089732
transform 1 0 18400 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_7169
timestamp 1668089732
transform 1 0 18400 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_7170
timestamp 1668089732
transform 1 0 18400 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_7171
timestamp 1668089732
transform 1 0 18400 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_7172
timestamp 1668089732
transform 1 0 18400 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_7173
timestamp 1668089732
transform 1 0 18400 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_7174
timestamp 1668089732
transform 1 0 18400 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_7175
timestamp 1668089732
transform 1 0 18400 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_7176
timestamp 1668089732
transform 1 0 18400 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_7177
timestamp 1668089732
transform 1 0 18400 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_7178
timestamp 1668089732
transform 1 0 18400 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_7179
timestamp 1668089732
transform 1 0 18400 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_7180
timestamp 1668089732
transform 1 0 18400 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_7181
timestamp 1668089732
transform 1 0 18400 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_7182
timestamp 1668089732
transform 1 0 18400 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_7183
timestamp 1668089732
transform 1 0 18400 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_7184
timestamp 1668089732
transform 1 0 18400 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_7185
timestamp 1668089732
transform 1 0 18400 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_7186
timestamp 1668089732
transform 1 0 18400 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_7187
timestamp 1668089732
transform 1 0 18400 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_7188
timestamp 1668089732
transform 1 0 18400 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_7189
timestamp 1668089732
transform 1 0 18400 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_7190
timestamp 1668089732
transform 1 0 18400 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_7191
timestamp 1668089732
transform 1 0 18400 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_7192
timestamp 1668089732
transform 1 0 18560 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_7193
timestamp 1668089732
transform 1 0 18560 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_7194
timestamp 1668089732
transform 1 0 18560 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_7195
timestamp 1668089732
transform 1 0 18560 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_7196
timestamp 1668089732
transform 1 0 18560 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_7197
timestamp 1668089732
transform 1 0 18560 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_7198
timestamp 1668089732
transform 1 0 18560 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_7199
timestamp 1668089732
transform 1 0 18560 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_7200
timestamp 1668089732
transform 1 0 18560 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_7201
timestamp 1668089732
transform 1 0 18560 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_7202
timestamp 1668089732
transform 1 0 18560 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_7203
timestamp 1668089732
transform 1 0 18560 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_7204
timestamp 1668089732
transform 1 0 18560 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_7205
timestamp 1668089732
transform 1 0 18560 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_7206
timestamp 1668089732
transform 1 0 18560 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_7207
timestamp 1668089732
transform 1 0 18560 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_7208
timestamp 1668089732
transform 1 0 18560 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_7209
timestamp 1668089732
transform 1 0 18560 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_7210
timestamp 1668089732
transform 1 0 18560 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_7211
timestamp 1668089732
transform 1 0 18560 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_7212
timestamp 1668089732
transform 1 0 18560 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_7213
timestamp 1668089732
transform 1 0 18560 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_7214
timestamp 1668089732
transform 1 0 18560 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_7215
timestamp 1668089732
transform 1 0 18560 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_7216
timestamp 1668089732
transform 1 0 18560 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_7217
timestamp 1668089732
transform 1 0 18560 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_7218
timestamp 1668089732
transform 1 0 18560 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_7219
timestamp 1668089732
transform 1 0 18560 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_7220
timestamp 1668089732
transform 1 0 18560 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_7221
timestamp 1668089732
transform 1 0 18560 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_7222
timestamp 1668089732
transform 1 0 18560 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_7223
timestamp 1668089732
transform 1 0 18560 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_7224
timestamp 1668089732
transform 1 0 18560 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_7225
timestamp 1668089732
transform 1 0 18560 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_7226
timestamp 1668089732
transform 1 0 18560 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_7227
timestamp 1668089732
transform 1 0 18560 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_7228
timestamp 1668089732
transform 1 0 18560 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_7229
timestamp 1668089732
transform 1 0 18560 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_7230
timestamp 1668089732
transform 1 0 18560 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_7231
timestamp 1668089732
transform 1 0 18560 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_7232
timestamp 1668089732
transform 1 0 18560 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_7233
timestamp 1668089732
transform 1 0 18560 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_7234
timestamp 1668089732
transform 1 0 18560 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_7235
timestamp 1668089732
transform 1 0 18560 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_7236
timestamp 1668089732
transform 1 0 18560 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_7237
timestamp 1668089732
transform 1 0 18560 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_7238
timestamp 1668089732
transform 1 0 18560 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_7239
timestamp 1668089732
transform 1 0 18560 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_7240
timestamp 1668089732
transform 1 0 18560 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_7241
timestamp 1668089732
transform 1 0 18560 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_7242
timestamp 1668089732
transform 1 0 18560 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_7243
timestamp 1668089732
transform 1 0 18560 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_7244
timestamp 1668089732
transform 1 0 18560 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_7245
timestamp 1668089732
transform 1 0 18560 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_7246
timestamp 1668089732
transform 1 0 18560 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_7247
timestamp 1668089732
transform 1 0 18560 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_7248
timestamp 1668089732
transform 1 0 18560 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_7249
timestamp 1668089732
transform 1 0 18560 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_7250
timestamp 1668089732
transform 1 0 18560 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_7251
timestamp 1668089732
transform 1 0 18560 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_7252
timestamp 1668089732
transform 1 0 18560 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_7253
timestamp 1668089732
transform 1 0 18560 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_7254
timestamp 1668089732
transform 1 0 18720 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_7255
timestamp 1668089732
transform 1 0 18720 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_7256
timestamp 1668089732
transform 1 0 18720 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_7257
timestamp 1668089732
transform 1 0 18720 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_7258
timestamp 1668089732
transform 1 0 18720 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_7259
timestamp 1668089732
transform 1 0 18720 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_7260
timestamp 1668089732
transform 1 0 18720 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_7261
timestamp 1668089732
transform 1 0 18720 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_7262
timestamp 1668089732
transform 1 0 18720 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_7263
timestamp 1668089732
transform 1 0 18720 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_7264
timestamp 1668089732
transform 1 0 18720 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_7265
timestamp 1668089732
transform 1 0 18720 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_7266
timestamp 1668089732
transform 1 0 18720 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_7267
timestamp 1668089732
transform 1 0 18720 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_7268
timestamp 1668089732
transform 1 0 18720 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_7269
timestamp 1668089732
transform 1 0 18720 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_7270
timestamp 1668089732
transform 1 0 18720 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_7271
timestamp 1668089732
transform 1 0 18720 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_7272
timestamp 1668089732
transform 1 0 18720 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_7273
timestamp 1668089732
transform 1 0 18720 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_7274
timestamp 1668089732
transform 1 0 18720 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_7275
timestamp 1668089732
transform 1 0 18720 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_7276
timestamp 1668089732
transform 1 0 18720 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_7277
timestamp 1668089732
transform 1 0 18720 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_7278
timestamp 1668089732
transform 1 0 18720 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_7279
timestamp 1668089732
transform 1 0 18720 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_7280
timestamp 1668089732
transform 1 0 18720 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_7281
timestamp 1668089732
transform 1 0 18720 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_7282
timestamp 1668089732
transform 1 0 18720 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_7283
timestamp 1668089732
transform 1 0 18720 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_7284
timestamp 1668089732
transform 1 0 18720 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_7285
timestamp 1668089732
transform 1 0 18720 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_7286
timestamp 1668089732
transform 1 0 18720 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_7287
timestamp 1668089732
transform 1 0 18720 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_7288
timestamp 1668089732
transform 1 0 18720 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_7289
timestamp 1668089732
transform 1 0 18720 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_7290
timestamp 1668089732
transform 1 0 18720 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_7291
timestamp 1668089732
transform 1 0 18720 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_7292
timestamp 1668089732
transform 1 0 18720 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_7293
timestamp 1668089732
transform 1 0 18720 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_7294
timestamp 1668089732
transform 1 0 18720 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_7295
timestamp 1668089732
transform 1 0 18720 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_7296
timestamp 1668089732
transform 1 0 18720 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_7297
timestamp 1668089732
transform 1 0 18720 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_7298
timestamp 1668089732
transform 1 0 18720 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_7299
timestamp 1668089732
transform 1 0 18720 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_7300
timestamp 1668089732
transform 1 0 18720 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_7301
timestamp 1668089732
transform 1 0 18720 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_7302
timestamp 1668089732
transform 1 0 18720 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_7303
timestamp 1668089732
transform 1 0 18720 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_7304
timestamp 1668089732
transform 1 0 18720 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_7305
timestamp 1668089732
transform 1 0 18720 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_7306
timestamp 1668089732
transform 1 0 18720 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_7307
timestamp 1668089732
transform 1 0 18720 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_7308
timestamp 1668089732
transform 1 0 18720 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_7309
timestamp 1668089732
transform 1 0 18720 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_7310
timestamp 1668089732
transform 1 0 18720 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_7311
timestamp 1668089732
transform 1 0 18720 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_7312
timestamp 1668089732
transform 1 0 18720 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_7313
timestamp 1668089732
transform 1 0 18720 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_7314
timestamp 1668089732
transform 1 0 18720 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_7315
timestamp 1668089732
transform 1 0 18720 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_7316
timestamp 1668089732
transform 1 0 18880 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_7317
timestamp 1668089732
transform 1 0 18880 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_7318
timestamp 1668089732
transform 1 0 18880 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_7319
timestamp 1668089732
transform 1 0 18880 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_7320
timestamp 1668089732
transform 1 0 18880 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_7321
timestamp 1668089732
transform 1 0 18880 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_7322
timestamp 1668089732
transform 1 0 18880 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_7323
timestamp 1668089732
transform 1 0 18880 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_7324
timestamp 1668089732
transform 1 0 18880 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_7325
timestamp 1668089732
transform 1 0 18880 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_7326
timestamp 1668089732
transform 1 0 18880 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_7327
timestamp 1668089732
transform 1 0 18880 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_7328
timestamp 1668089732
transform 1 0 18880 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_7329
timestamp 1668089732
transform 1 0 18880 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_7330
timestamp 1668089732
transform 1 0 18880 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_7331
timestamp 1668089732
transform 1 0 18880 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_7332
timestamp 1668089732
transform 1 0 18880 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_7333
timestamp 1668089732
transform 1 0 18880 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_7334
timestamp 1668089732
transform 1 0 18880 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_7335
timestamp 1668089732
transform 1 0 18880 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_7336
timestamp 1668089732
transform 1 0 18880 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_7337
timestamp 1668089732
transform 1 0 18880 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_7338
timestamp 1668089732
transform 1 0 18880 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_7339
timestamp 1668089732
transform 1 0 18880 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_7340
timestamp 1668089732
transform 1 0 18880 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_7341
timestamp 1668089732
transform 1 0 18880 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_7342
timestamp 1668089732
transform 1 0 18880 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_7343
timestamp 1668089732
transform 1 0 18880 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_7344
timestamp 1668089732
transform 1 0 18880 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_7345
timestamp 1668089732
transform 1 0 18880 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_7346
timestamp 1668089732
transform 1 0 18880 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_7347
timestamp 1668089732
transform 1 0 18880 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_7348
timestamp 1668089732
transform 1 0 18880 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_7349
timestamp 1668089732
transform 1 0 18880 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_7350
timestamp 1668089732
transform 1 0 18880 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_7351
timestamp 1668089732
transform 1 0 18880 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_7352
timestamp 1668089732
transform 1 0 18880 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_7353
timestamp 1668089732
transform 1 0 18880 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_7354
timestamp 1668089732
transform 1 0 18880 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_7355
timestamp 1668089732
transform 1 0 18880 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_7356
timestamp 1668089732
transform 1 0 18880 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_7357
timestamp 1668089732
transform 1 0 18880 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_7358
timestamp 1668089732
transform 1 0 18880 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_7359
timestamp 1668089732
transform 1 0 18880 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_7360
timestamp 1668089732
transform 1 0 18880 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_7361
timestamp 1668089732
transform 1 0 18880 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_7362
timestamp 1668089732
transform 1 0 18880 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_7363
timestamp 1668089732
transform 1 0 18880 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_7364
timestamp 1668089732
transform 1 0 18880 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_7365
timestamp 1668089732
transform 1 0 18880 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_7366
timestamp 1668089732
transform 1 0 18880 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_7367
timestamp 1668089732
transform 1 0 18880 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_7368
timestamp 1668089732
transform 1 0 18880 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_7369
timestamp 1668089732
transform 1 0 18880 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_7370
timestamp 1668089732
transform 1 0 18880 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_7371
timestamp 1668089732
transform 1 0 18880 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_7372
timestamp 1668089732
transform 1 0 18880 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_7373
timestamp 1668089732
transform 1 0 18880 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_7374
timestamp 1668089732
transform 1 0 18880 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_7375
timestamp 1668089732
transform 1 0 18880 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_7376
timestamp 1668089732
transform 1 0 18880 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_7377
timestamp 1668089732
transform 1 0 18880 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_7378
timestamp 1668089732
transform 1 0 19040 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_7379
timestamp 1668089732
transform 1 0 19040 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_7380
timestamp 1668089732
transform 1 0 19040 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_7381
timestamp 1668089732
transform 1 0 19040 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_7382
timestamp 1668089732
transform 1 0 19040 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_7383
timestamp 1668089732
transform 1 0 19040 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_7384
timestamp 1668089732
transform 1 0 19040 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_7385
timestamp 1668089732
transform 1 0 19040 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_7386
timestamp 1668089732
transform 1 0 19040 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_7387
timestamp 1668089732
transform 1 0 19040 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_7388
timestamp 1668089732
transform 1 0 19040 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_7389
timestamp 1668089732
transform 1 0 19040 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_7390
timestamp 1668089732
transform 1 0 19040 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_7391
timestamp 1668089732
transform 1 0 19040 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_7392
timestamp 1668089732
transform 1 0 19040 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_7393
timestamp 1668089732
transform 1 0 19040 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_7394
timestamp 1668089732
transform 1 0 19040 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_7395
timestamp 1668089732
transform 1 0 19040 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_7396
timestamp 1668089732
transform 1 0 19040 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_7397
timestamp 1668089732
transform 1 0 19040 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_7398
timestamp 1668089732
transform 1 0 19040 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_7399
timestamp 1668089732
transform 1 0 19040 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_7400
timestamp 1668089732
transform 1 0 19040 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_7401
timestamp 1668089732
transform 1 0 19040 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_7402
timestamp 1668089732
transform 1 0 19040 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_7403
timestamp 1668089732
transform 1 0 19040 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_7404
timestamp 1668089732
transform 1 0 19040 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_7405
timestamp 1668089732
transform 1 0 19040 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_7406
timestamp 1668089732
transform 1 0 19040 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_7407
timestamp 1668089732
transform 1 0 19040 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_7408
timestamp 1668089732
transform 1 0 19040 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_7409
timestamp 1668089732
transform 1 0 19040 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_7410
timestamp 1668089732
transform 1 0 19040 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_7411
timestamp 1668089732
transform 1 0 19040 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_7412
timestamp 1668089732
transform 1 0 19040 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_7413
timestamp 1668089732
transform 1 0 19040 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_7414
timestamp 1668089732
transform 1 0 19040 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_7415
timestamp 1668089732
transform 1 0 19040 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_7416
timestamp 1668089732
transform 1 0 19040 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_7417
timestamp 1668089732
transform 1 0 19040 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_7418
timestamp 1668089732
transform 1 0 19040 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_7419
timestamp 1668089732
transform 1 0 19040 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_7420
timestamp 1668089732
transform 1 0 19040 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_7421
timestamp 1668089732
transform 1 0 19040 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_7422
timestamp 1668089732
transform 1 0 19040 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_7423
timestamp 1668089732
transform 1 0 19040 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_7424
timestamp 1668089732
transform 1 0 19040 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_7425
timestamp 1668089732
transform 1 0 19040 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_7426
timestamp 1668089732
transform 1 0 19040 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_7427
timestamp 1668089732
transform 1 0 19040 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_7428
timestamp 1668089732
transform 1 0 19040 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_7429
timestamp 1668089732
transform 1 0 19040 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_7430
timestamp 1668089732
transform 1 0 19040 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_7431
timestamp 1668089732
transform 1 0 19040 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_7432
timestamp 1668089732
transform 1 0 19040 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_7433
timestamp 1668089732
transform 1 0 19040 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_7434
timestamp 1668089732
transform 1 0 19040 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_7435
timestamp 1668089732
transform 1 0 19040 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_7436
timestamp 1668089732
transform 1 0 19040 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_7437
timestamp 1668089732
transform 1 0 19040 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_7438
timestamp 1668089732
transform 1 0 19040 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_7439
timestamp 1668089732
transform 1 0 19040 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_7440
timestamp 1668089732
transform 1 0 19200 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_7441
timestamp 1668089732
transform 1 0 19200 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_7442
timestamp 1668089732
transform 1 0 19200 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_7443
timestamp 1668089732
transform 1 0 19200 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_7444
timestamp 1668089732
transform 1 0 19200 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_7445
timestamp 1668089732
transform 1 0 19200 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_7446
timestamp 1668089732
transform 1 0 19200 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_7447
timestamp 1668089732
transform 1 0 19200 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_7448
timestamp 1668089732
transform 1 0 19200 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_7449
timestamp 1668089732
transform 1 0 19200 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_7450
timestamp 1668089732
transform 1 0 19200 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_7451
timestamp 1668089732
transform 1 0 19200 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_7452
timestamp 1668089732
transform 1 0 19200 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_7453
timestamp 1668089732
transform 1 0 19200 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_7454
timestamp 1668089732
transform 1 0 19200 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_7455
timestamp 1668089732
transform 1 0 19200 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_7456
timestamp 1668089732
transform 1 0 19200 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_7457
timestamp 1668089732
transform 1 0 19200 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_7458
timestamp 1668089732
transform 1 0 19200 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_7459
timestamp 1668089732
transform 1 0 19200 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_7460
timestamp 1668089732
transform 1 0 19200 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_7461
timestamp 1668089732
transform 1 0 19200 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_7462
timestamp 1668089732
transform 1 0 19200 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_7463
timestamp 1668089732
transform 1 0 19200 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_7464
timestamp 1668089732
transform 1 0 19200 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_7465
timestamp 1668089732
transform 1 0 19200 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_7466
timestamp 1668089732
transform 1 0 19200 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_7467
timestamp 1668089732
transform 1 0 19200 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_7468
timestamp 1668089732
transform 1 0 19200 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_7469
timestamp 1668089732
transform 1 0 19200 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_7470
timestamp 1668089732
transform 1 0 19200 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_7471
timestamp 1668089732
transform 1 0 19200 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_7472
timestamp 1668089732
transform 1 0 19200 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_7473
timestamp 1668089732
transform 1 0 19200 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_7474
timestamp 1668089732
transform 1 0 19200 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_7475
timestamp 1668089732
transform 1 0 19200 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_7476
timestamp 1668089732
transform 1 0 19200 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_7477
timestamp 1668089732
transform 1 0 19200 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_7478
timestamp 1668089732
transform 1 0 19200 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_7479
timestamp 1668089732
transform 1 0 19200 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_7480
timestamp 1668089732
transform 1 0 19200 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_7481
timestamp 1668089732
transform 1 0 19200 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_7482
timestamp 1668089732
transform 1 0 19200 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_7483
timestamp 1668089732
transform 1 0 19200 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_7484
timestamp 1668089732
transform 1 0 19200 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_7485
timestamp 1668089732
transform 1 0 19200 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_7486
timestamp 1668089732
transform 1 0 19200 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_7487
timestamp 1668089732
transform 1 0 19200 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_7488
timestamp 1668089732
transform 1 0 19200 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_7489
timestamp 1668089732
transform 1 0 19200 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_7490
timestamp 1668089732
transform 1 0 19200 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_7491
timestamp 1668089732
transform 1 0 19200 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_7492
timestamp 1668089732
transform 1 0 19200 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_7493
timestamp 1668089732
transform 1 0 19200 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_7494
timestamp 1668089732
transform 1 0 19200 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_7495
timestamp 1668089732
transform 1 0 19200 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_7496
timestamp 1668089732
transform 1 0 19200 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_7497
timestamp 1668089732
transform 1 0 19200 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_7498
timestamp 1668089732
transform 1 0 19200 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_7499
timestamp 1668089732
transform 1 0 19200 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_7500
timestamp 1668089732
transform 1 0 19200 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_7501
timestamp 1668089732
transform 1 0 19200 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_7502
timestamp 1668089732
transform 1 0 19360 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_7503
timestamp 1668089732
transform 1 0 19360 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_7504
timestamp 1668089732
transform 1 0 19360 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_7505
timestamp 1668089732
transform 1 0 19360 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_7506
timestamp 1668089732
transform 1 0 19360 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_7507
timestamp 1668089732
transform 1 0 19360 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_7508
timestamp 1668089732
transform 1 0 19360 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_7509
timestamp 1668089732
transform 1 0 19360 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_7510
timestamp 1668089732
transform 1 0 19360 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_7511
timestamp 1668089732
transform 1 0 19360 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_7512
timestamp 1668089732
transform 1 0 19360 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_7513
timestamp 1668089732
transform 1 0 19360 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_7514
timestamp 1668089732
transform 1 0 19360 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_7515
timestamp 1668089732
transform 1 0 19360 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_7516
timestamp 1668089732
transform 1 0 19360 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_7517
timestamp 1668089732
transform 1 0 19360 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_7518
timestamp 1668089732
transform 1 0 19360 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_7519
timestamp 1668089732
transform 1 0 19360 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_7520
timestamp 1668089732
transform 1 0 19360 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_7521
timestamp 1668089732
transform 1 0 19360 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_7522
timestamp 1668089732
transform 1 0 19360 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_7523
timestamp 1668089732
transform 1 0 19360 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_7524
timestamp 1668089732
transform 1 0 19360 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_7525
timestamp 1668089732
transform 1 0 19360 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_7526
timestamp 1668089732
transform 1 0 19360 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_7527
timestamp 1668089732
transform 1 0 19360 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_7528
timestamp 1668089732
transform 1 0 19360 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_7529
timestamp 1668089732
transform 1 0 19360 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_7530
timestamp 1668089732
transform 1 0 19360 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_7531
timestamp 1668089732
transform 1 0 19360 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_7532
timestamp 1668089732
transform 1 0 19360 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_7533
timestamp 1668089732
transform 1 0 19360 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_7534
timestamp 1668089732
transform 1 0 19360 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_7535
timestamp 1668089732
transform 1 0 19360 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_7536
timestamp 1668089732
transform 1 0 19360 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_7537
timestamp 1668089732
transform 1 0 19360 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_7538
timestamp 1668089732
transform 1 0 19360 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_7539
timestamp 1668089732
transform 1 0 19360 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_7540
timestamp 1668089732
transform 1 0 19360 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_7541
timestamp 1668089732
transform 1 0 19360 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_7542
timestamp 1668089732
transform 1 0 19360 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_7543
timestamp 1668089732
transform 1 0 19360 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_7544
timestamp 1668089732
transform 1 0 19360 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_7545
timestamp 1668089732
transform 1 0 19360 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_7546
timestamp 1668089732
transform 1 0 19360 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_7547
timestamp 1668089732
transform 1 0 19360 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_7548
timestamp 1668089732
transform 1 0 19360 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_7549
timestamp 1668089732
transform 1 0 19360 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_7550
timestamp 1668089732
transform 1 0 19360 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_7551
timestamp 1668089732
transform 1 0 19360 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_7552
timestamp 1668089732
transform 1 0 19360 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_7553
timestamp 1668089732
transform 1 0 19360 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_7554
timestamp 1668089732
transform 1 0 19360 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_7555
timestamp 1668089732
transform 1 0 19360 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_7556
timestamp 1668089732
transform 1 0 19360 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_7557
timestamp 1668089732
transform 1 0 19360 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_7558
timestamp 1668089732
transform 1 0 19360 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_7559
timestamp 1668089732
transform 1 0 19360 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_7560
timestamp 1668089732
transform 1 0 19360 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_7561
timestamp 1668089732
transform 1 0 19360 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_7562
timestamp 1668089732
transform 1 0 19360 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_7563
timestamp 1668089732
transform 1 0 19360 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_7564
timestamp 1668089732
transform 1 0 19520 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_7565
timestamp 1668089732
transform 1 0 19520 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_7566
timestamp 1668089732
transform 1 0 19520 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_7567
timestamp 1668089732
transform 1 0 19520 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_7568
timestamp 1668089732
transform 1 0 19520 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_7569
timestamp 1668089732
transform 1 0 19520 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_7570
timestamp 1668089732
transform 1 0 19520 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_7571
timestamp 1668089732
transform 1 0 19520 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_7572
timestamp 1668089732
transform 1 0 19520 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_7573
timestamp 1668089732
transform 1 0 19520 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_7574
timestamp 1668089732
transform 1 0 19520 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_7575
timestamp 1668089732
transform 1 0 19520 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_7576
timestamp 1668089732
transform 1 0 19520 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_7577
timestamp 1668089732
transform 1 0 19520 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_7578
timestamp 1668089732
transform 1 0 19520 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_7579
timestamp 1668089732
transform 1 0 19520 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_7580
timestamp 1668089732
transform 1 0 19520 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_7581
timestamp 1668089732
transform 1 0 19520 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_7582
timestamp 1668089732
transform 1 0 19520 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_7583
timestamp 1668089732
transform 1 0 19520 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_7584
timestamp 1668089732
transform 1 0 19520 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_7585
timestamp 1668089732
transform 1 0 19520 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_7586
timestamp 1668089732
transform 1 0 19520 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_7587
timestamp 1668089732
transform 1 0 19520 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_7588
timestamp 1668089732
transform 1 0 19520 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_7589
timestamp 1668089732
transform 1 0 19520 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_7590
timestamp 1668089732
transform 1 0 19520 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_7591
timestamp 1668089732
transform 1 0 19520 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_7592
timestamp 1668089732
transform 1 0 19520 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_7593
timestamp 1668089732
transform 1 0 19520 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_7594
timestamp 1668089732
transform 1 0 19520 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_7595
timestamp 1668089732
transform 1 0 19520 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_7596
timestamp 1668089732
transform 1 0 19520 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_7597
timestamp 1668089732
transform 1 0 19520 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_7598
timestamp 1668089732
transform 1 0 19520 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_7599
timestamp 1668089732
transform 1 0 19520 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_7600
timestamp 1668089732
transform 1 0 19520 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_7601
timestamp 1668089732
transform 1 0 19520 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_7602
timestamp 1668089732
transform 1 0 19520 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_7603
timestamp 1668089732
transform 1 0 19520 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_7604
timestamp 1668089732
transform 1 0 19520 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_7605
timestamp 1668089732
transform 1 0 19520 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_7606
timestamp 1668089732
transform 1 0 19520 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_7607
timestamp 1668089732
transform 1 0 19520 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_7608
timestamp 1668089732
transform 1 0 19520 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_7609
timestamp 1668089732
transform 1 0 19520 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_7610
timestamp 1668089732
transform 1 0 19520 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_7611
timestamp 1668089732
transform 1 0 19520 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_7612
timestamp 1668089732
transform 1 0 19520 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_7613
timestamp 1668089732
transform 1 0 19520 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_7614
timestamp 1668089732
transform 1 0 19520 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_7615
timestamp 1668089732
transform 1 0 19520 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_7616
timestamp 1668089732
transform 1 0 19520 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_7617
timestamp 1668089732
transform 1 0 19520 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_7618
timestamp 1668089732
transform 1 0 19520 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_7619
timestamp 1668089732
transform 1 0 19520 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_7620
timestamp 1668089732
transform 1 0 19520 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_7621
timestamp 1668089732
transform 1 0 19520 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_7622
timestamp 1668089732
transform 1 0 19520 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_7623
timestamp 1668089732
transform 1 0 19520 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_7624
timestamp 1668089732
transform 1 0 19520 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_7625
timestamp 1668089732
transform 1 0 19520 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_7626
timestamp 1668089732
transform 1 0 19680 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_7627
timestamp 1668089732
transform 1 0 19680 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_7628
timestamp 1668089732
transform 1 0 19680 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_7629
timestamp 1668089732
transform 1 0 19680 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_7630
timestamp 1668089732
transform 1 0 19680 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_7631
timestamp 1668089732
transform 1 0 19680 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_7632
timestamp 1668089732
transform 1 0 19680 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_7633
timestamp 1668089732
transform 1 0 19680 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_7634
timestamp 1668089732
transform 1 0 19680 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_7635
timestamp 1668089732
transform 1 0 19680 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_7636
timestamp 1668089732
transform 1 0 19680 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_7637
timestamp 1668089732
transform 1 0 19680 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_7638
timestamp 1668089732
transform 1 0 19680 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_7639
timestamp 1668089732
transform 1 0 19680 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_7640
timestamp 1668089732
transform 1 0 19680 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_7641
timestamp 1668089732
transform 1 0 19680 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_7642
timestamp 1668089732
transform 1 0 19680 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_7643
timestamp 1668089732
transform 1 0 19680 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_7644
timestamp 1668089732
transform 1 0 19680 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_7645
timestamp 1668089732
transform 1 0 19680 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_7646
timestamp 1668089732
transform 1 0 19680 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_7647
timestamp 1668089732
transform 1 0 19680 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_7648
timestamp 1668089732
transform 1 0 19680 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_7649
timestamp 1668089732
transform 1 0 19680 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_7650
timestamp 1668089732
transform 1 0 19680 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_7651
timestamp 1668089732
transform 1 0 19680 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_7652
timestamp 1668089732
transform 1 0 19680 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_7653
timestamp 1668089732
transform 1 0 19680 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_7654
timestamp 1668089732
transform 1 0 19680 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_7655
timestamp 1668089732
transform 1 0 19680 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_7656
timestamp 1668089732
transform 1 0 19680 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_7657
timestamp 1668089732
transform 1 0 19680 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_7658
timestamp 1668089732
transform 1 0 19680 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_7659
timestamp 1668089732
transform 1 0 19680 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_7660
timestamp 1668089732
transform 1 0 19680 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_7661
timestamp 1668089732
transform 1 0 19680 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_7662
timestamp 1668089732
transform 1 0 19680 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_7663
timestamp 1668089732
transform 1 0 19680 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_7664
timestamp 1668089732
transform 1 0 19680 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_7665
timestamp 1668089732
transform 1 0 19680 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_7666
timestamp 1668089732
transform 1 0 19680 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_7667
timestamp 1668089732
transform 1 0 19680 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_7668
timestamp 1668089732
transform 1 0 19680 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_7669
timestamp 1668089732
transform 1 0 19680 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_7670
timestamp 1668089732
transform 1 0 19680 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_7671
timestamp 1668089732
transform 1 0 19680 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_7672
timestamp 1668089732
transform 1 0 19680 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_7673
timestamp 1668089732
transform 1 0 19680 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_7674
timestamp 1668089732
transform 1 0 19680 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_7675
timestamp 1668089732
transform 1 0 19680 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_7676
timestamp 1668089732
transform 1 0 19680 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_7677
timestamp 1668089732
transform 1 0 19680 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_7678
timestamp 1668089732
transform 1 0 19680 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_7679
timestamp 1668089732
transform 1 0 19680 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_7680
timestamp 1668089732
transform 1 0 19680 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_7681
timestamp 1668089732
transform 1 0 19680 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_7682
timestamp 1668089732
transform 1 0 19680 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_7683
timestamp 1668089732
transform 1 0 19680 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_7684
timestamp 1668089732
transform 1 0 19680 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_7685
timestamp 1668089732
transform 1 0 19680 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_7686
timestamp 1668089732
transform 1 0 19680 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_7687
timestamp 1668089732
transform 1 0 19680 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_7688
timestamp 1668089732
transform 1 0 19840 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_7689
timestamp 1668089732
transform 1 0 19840 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_7690
timestamp 1668089732
transform 1 0 19840 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_7691
timestamp 1668089732
transform 1 0 19840 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_7692
timestamp 1668089732
transform 1 0 19840 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_7693
timestamp 1668089732
transform 1 0 19840 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_7694
timestamp 1668089732
transform 1 0 19840 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_7695
timestamp 1668089732
transform 1 0 19840 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_7696
timestamp 1668089732
transform 1 0 19840 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_7697
timestamp 1668089732
transform 1 0 19840 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_7698
timestamp 1668089732
transform 1 0 19840 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_7699
timestamp 1668089732
transform 1 0 19840 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_7700
timestamp 1668089732
transform 1 0 19840 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_7701
timestamp 1668089732
transform 1 0 19840 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_7702
timestamp 1668089732
transform 1 0 19840 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_7703
timestamp 1668089732
transform 1 0 19840 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_7704
timestamp 1668089732
transform 1 0 19840 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_7705
timestamp 1668089732
transform 1 0 19840 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_7706
timestamp 1668089732
transform 1 0 19840 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_7707
timestamp 1668089732
transform 1 0 19840 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_7708
timestamp 1668089732
transform 1 0 19840 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_7709
timestamp 1668089732
transform 1 0 19840 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_7710
timestamp 1668089732
transform 1 0 19840 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_7711
timestamp 1668089732
transform 1 0 19840 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_7712
timestamp 1668089732
transform 1 0 19840 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_7713
timestamp 1668089732
transform 1 0 19840 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_7714
timestamp 1668089732
transform 1 0 19840 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_7715
timestamp 1668089732
transform 1 0 19840 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_7716
timestamp 1668089732
transform 1 0 19840 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_7717
timestamp 1668089732
transform 1 0 19840 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_7718
timestamp 1668089732
transform 1 0 19840 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_7719
timestamp 1668089732
transform 1 0 19840 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_7720
timestamp 1668089732
transform 1 0 19840 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_7721
timestamp 1668089732
transform 1 0 19840 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_7722
timestamp 1668089732
transform 1 0 19840 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_7723
timestamp 1668089732
transform 1 0 19840 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_7724
timestamp 1668089732
transform 1 0 19840 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_7725
timestamp 1668089732
transform 1 0 19840 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_7726
timestamp 1668089732
transform 1 0 19840 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_7727
timestamp 1668089732
transform 1 0 19840 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_7728
timestamp 1668089732
transform 1 0 19840 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_7729
timestamp 1668089732
transform 1 0 19840 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_7730
timestamp 1668089732
transform 1 0 19840 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_7731
timestamp 1668089732
transform 1 0 19840 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_7732
timestamp 1668089732
transform 1 0 19840 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_7733
timestamp 1668089732
transform 1 0 19840 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_7734
timestamp 1668089732
transform 1 0 19840 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_7735
timestamp 1668089732
transform 1 0 19840 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_7736
timestamp 1668089732
transform 1 0 19840 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_7737
timestamp 1668089732
transform 1 0 19840 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_7738
timestamp 1668089732
transform 1 0 19840 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_7739
timestamp 1668089732
transform 1 0 19840 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_7740
timestamp 1668089732
transform 1 0 19840 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_7741
timestamp 1668089732
transform 1 0 19840 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_7742
timestamp 1668089732
transform 1 0 19840 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_7743
timestamp 1668089732
transform 1 0 19840 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_7744
timestamp 1668089732
transform 1 0 19840 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_7745
timestamp 1668089732
transform 1 0 19840 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_7746
timestamp 1668089732
transform 1 0 19840 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_7747
timestamp 1668089732
transform 1 0 19840 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_7748
timestamp 1668089732
transform 1 0 19840 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_7749
timestamp 1668089732
transform 1 0 19840 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_7750
timestamp 1668089732
transform 1 0 20000 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_7751
timestamp 1668089732
transform 1 0 20000 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_7752
timestamp 1668089732
transform 1 0 20000 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_7753
timestamp 1668089732
transform 1 0 20000 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_7754
timestamp 1668089732
transform 1 0 20000 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_7755
timestamp 1668089732
transform 1 0 20000 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_7756
timestamp 1668089732
transform 1 0 20000 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_7757
timestamp 1668089732
transform 1 0 20000 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_7758
timestamp 1668089732
transform 1 0 20000 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_7759
timestamp 1668089732
transform 1 0 20000 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_7760
timestamp 1668089732
transform 1 0 20000 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_7761
timestamp 1668089732
transform 1 0 20000 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_7762
timestamp 1668089732
transform 1 0 20000 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_7763
timestamp 1668089732
transform 1 0 20000 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_7764
timestamp 1668089732
transform 1 0 20000 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_7765
timestamp 1668089732
transform 1 0 20000 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_7766
timestamp 1668089732
transform 1 0 20000 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_7767
timestamp 1668089732
transform 1 0 20000 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_7768
timestamp 1668089732
transform 1 0 20000 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_7769
timestamp 1668089732
transform 1 0 20000 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_7770
timestamp 1668089732
transform 1 0 20000 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_7771
timestamp 1668089732
transform 1 0 20000 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_7772
timestamp 1668089732
transform 1 0 20000 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_7773
timestamp 1668089732
transform 1 0 20000 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_7774
timestamp 1668089732
transform 1 0 20000 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_7775
timestamp 1668089732
transform 1 0 20000 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_7776
timestamp 1668089732
transform 1 0 20000 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_7777
timestamp 1668089732
transform 1 0 20000 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_7778
timestamp 1668089732
transform 1 0 20000 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_7779
timestamp 1668089732
transform 1 0 20000 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_7780
timestamp 1668089732
transform 1 0 20000 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_7781
timestamp 1668089732
transform 1 0 20000 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_7782
timestamp 1668089732
transform 1 0 20000 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_7783
timestamp 1668089732
transform 1 0 20000 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_7784
timestamp 1668089732
transform 1 0 20000 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_7785
timestamp 1668089732
transform 1 0 20000 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_7786
timestamp 1668089732
transform 1 0 20000 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_7787
timestamp 1668089732
transform 1 0 20000 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_7788
timestamp 1668089732
transform 1 0 20000 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_7789
timestamp 1668089732
transform 1 0 20000 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_7790
timestamp 1668089732
transform 1 0 20000 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_7791
timestamp 1668089732
transform 1 0 20000 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_7792
timestamp 1668089732
transform 1 0 20000 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_7793
timestamp 1668089732
transform 1 0 20000 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_7794
timestamp 1668089732
transform 1 0 20000 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_7795
timestamp 1668089732
transform 1 0 20000 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_7796
timestamp 1668089732
transform 1 0 20000 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_7797
timestamp 1668089732
transform 1 0 20000 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_7798
timestamp 1668089732
transform 1 0 20000 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_7799
timestamp 1668089732
transform 1 0 20000 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_7800
timestamp 1668089732
transform 1 0 20000 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_7801
timestamp 1668089732
transform 1 0 20000 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_7802
timestamp 1668089732
transform 1 0 20000 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_7803
timestamp 1668089732
transform 1 0 20000 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_7804
timestamp 1668089732
transform 1 0 20000 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_7805
timestamp 1668089732
transform 1 0 20000 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_7806
timestamp 1668089732
transform 1 0 20000 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_7807
timestamp 1668089732
transform 1 0 20000 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_7808
timestamp 1668089732
transform 1 0 20000 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_7809
timestamp 1668089732
transform 1 0 20000 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_7810
timestamp 1668089732
transform 1 0 20000 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_7811
timestamp 1668089732
transform 1 0 20000 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_7812
timestamp 1668089732
transform 1 0 20160 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_7813
timestamp 1668089732
transform 1 0 20160 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_7814
timestamp 1668089732
transform 1 0 20160 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_7815
timestamp 1668089732
transform 1 0 20160 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_7816
timestamp 1668089732
transform 1 0 20160 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_7817
timestamp 1668089732
transform 1 0 20160 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_7818
timestamp 1668089732
transform 1 0 20160 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_7819
timestamp 1668089732
transform 1 0 20160 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_7820
timestamp 1668089732
transform 1 0 20160 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_7821
timestamp 1668089732
transform 1 0 20160 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_7822
timestamp 1668089732
transform 1 0 20160 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_7823
timestamp 1668089732
transform 1 0 20160 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_7824
timestamp 1668089732
transform 1 0 20160 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_7825
timestamp 1668089732
transform 1 0 20160 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_7826
timestamp 1668089732
transform 1 0 20160 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_7827
timestamp 1668089732
transform 1 0 20160 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_7828
timestamp 1668089732
transform 1 0 20160 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_7829
timestamp 1668089732
transform 1 0 20160 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_7830
timestamp 1668089732
transform 1 0 20160 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_7831
timestamp 1668089732
transform 1 0 20160 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_7832
timestamp 1668089732
transform 1 0 20160 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_7833
timestamp 1668089732
transform 1 0 20160 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_7834
timestamp 1668089732
transform 1 0 20160 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_7835
timestamp 1668089732
transform 1 0 20160 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_7836
timestamp 1668089732
transform 1 0 20160 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_7837
timestamp 1668089732
transform 1 0 20160 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_7838
timestamp 1668089732
transform 1 0 20160 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_7839
timestamp 1668089732
transform 1 0 20160 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_7840
timestamp 1668089732
transform 1 0 20160 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_7841
timestamp 1668089732
transform 1 0 20160 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_7842
timestamp 1668089732
transform 1 0 20160 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_7843
timestamp 1668089732
transform 1 0 20160 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_7844
timestamp 1668089732
transform 1 0 20160 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_7845
timestamp 1668089732
transform 1 0 20160 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_7846
timestamp 1668089732
transform 1 0 20160 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_7847
timestamp 1668089732
transform 1 0 20160 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_7848
timestamp 1668089732
transform 1 0 20160 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_7849
timestamp 1668089732
transform 1 0 20160 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_7850
timestamp 1668089732
transform 1 0 20160 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_7851
timestamp 1668089732
transform 1 0 20160 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_7852
timestamp 1668089732
transform 1 0 20160 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_7853
timestamp 1668089732
transform 1 0 20160 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_7854
timestamp 1668089732
transform 1 0 20160 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_7855
timestamp 1668089732
transform 1 0 20160 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_7856
timestamp 1668089732
transform 1 0 20160 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_7857
timestamp 1668089732
transform 1 0 20160 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_7858
timestamp 1668089732
transform 1 0 20160 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_7859
timestamp 1668089732
transform 1 0 20160 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_7860
timestamp 1668089732
transform 1 0 20160 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_7861
timestamp 1668089732
transform 1 0 20160 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_7862
timestamp 1668089732
transform 1 0 20160 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_7863
timestamp 1668089732
transform 1 0 20160 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_7864
timestamp 1668089732
transform 1 0 20160 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_7865
timestamp 1668089732
transform 1 0 20160 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_7866
timestamp 1668089732
transform 1 0 20160 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_7867
timestamp 1668089732
transform 1 0 20160 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_7868
timestamp 1668089732
transform 1 0 20160 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_7869
timestamp 1668089732
transform 1 0 20160 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_7870
timestamp 1668089732
transform 1 0 20160 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_7871
timestamp 1668089732
transform 1 0 20160 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_7872
timestamp 1668089732
transform 1 0 20160 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_7873
timestamp 1668089732
transform 1 0 20160 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_7874
timestamp 1668089732
transform 1 0 20320 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_7875
timestamp 1668089732
transform 1 0 20320 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_7876
timestamp 1668089732
transform 1 0 20320 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_7877
timestamp 1668089732
transform 1 0 20320 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_7878
timestamp 1668089732
transform 1 0 20320 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_7879
timestamp 1668089732
transform 1 0 20320 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_7880
timestamp 1668089732
transform 1 0 20320 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_7881
timestamp 1668089732
transform 1 0 20320 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_7882
timestamp 1668089732
transform 1 0 20320 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_7883
timestamp 1668089732
transform 1 0 20320 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_7884
timestamp 1668089732
transform 1 0 20320 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_7885
timestamp 1668089732
transform 1 0 20320 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_7886
timestamp 1668089732
transform 1 0 20320 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_7887
timestamp 1668089732
transform 1 0 20320 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_7888
timestamp 1668089732
transform 1 0 20320 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_7889
timestamp 1668089732
transform 1 0 20320 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_7890
timestamp 1668089732
transform 1 0 20320 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_7891
timestamp 1668089732
transform 1 0 20320 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_7892
timestamp 1668089732
transform 1 0 20320 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_7893
timestamp 1668089732
transform 1 0 20320 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_7894
timestamp 1668089732
transform 1 0 20320 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_7895
timestamp 1668089732
transform 1 0 20320 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_7896
timestamp 1668089732
transform 1 0 20320 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_7897
timestamp 1668089732
transform 1 0 20320 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_7898
timestamp 1668089732
transform 1 0 20320 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_7899
timestamp 1668089732
transform 1 0 20320 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_7900
timestamp 1668089732
transform 1 0 20320 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_7901
timestamp 1668089732
transform 1 0 20320 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_7902
timestamp 1668089732
transform 1 0 20320 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_7903
timestamp 1668089732
transform 1 0 20320 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_7904
timestamp 1668089732
transform 1 0 20320 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_7905
timestamp 1668089732
transform 1 0 20320 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_7906
timestamp 1668089732
transform 1 0 20320 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_7907
timestamp 1668089732
transform 1 0 20320 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_7908
timestamp 1668089732
transform 1 0 20320 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_7909
timestamp 1668089732
transform 1 0 20320 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_7910
timestamp 1668089732
transform 1 0 20320 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_7911
timestamp 1668089732
transform 1 0 20320 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_7912
timestamp 1668089732
transform 1 0 20320 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_7913
timestamp 1668089732
transform 1 0 20320 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_7914
timestamp 1668089732
transform 1 0 20320 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_7915
timestamp 1668089732
transform 1 0 20320 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_7916
timestamp 1668089732
transform 1 0 20320 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_7917
timestamp 1668089732
transform 1 0 20320 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_7918
timestamp 1668089732
transform 1 0 20320 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_7919
timestamp 1668089732
transform 1 0 20320 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_7920
timestamp 1668089732
transform 1 0 20320 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_7921
timestamp 1668089732
transform 1 0 20320 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_7922
timestamp 1668089732
transform 1 0 20320 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_7923
timestamp 1668089732
transform 1 0 20320 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_7924
timestamp 1668089732
transform 1 0 20320 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_7925
timestamp 1668089732
transform 1 0 20320 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_7926
timestamp 1668089732
transform 1 0 20320 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_7927
timestamp 1668089732
transform 1 0 20320 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_7928
timestamp 1668089732
transform 1 0 20320 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_7929
timestamp 1668089732
transform 1 0 20320 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_7930
timestamp 1668089732
transform 1 0 20320 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_7931
timestamp 1668089732
transform 1 0 20320 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_7932
timestamp 1668089732
transform 1 0 20320 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_7933
timestamp 1668089732
transform 1 0 20320 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_7934
timestamp 1668089732
transform 1 0 20320 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_7935
timestamp 1668089732
transform 1 0 20320 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_7936
timestamp 1668089732
transform 1 0 20480 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_7937
timestamp 1668089732
transform 1 0 20480 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_7938
timestamp 1668089732
transform 1 0 20480 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_7939
timestamp 1668089732
transform 1 0 20480 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_7940
timestamp 1668089732
transform 1 0 20480 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_7941
timestamp 1668089732
transform 1 0 20480 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_7942
timestamp 1668089732
transform 1 0 20480 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_7943
timestamp 1668089732
transform 1 0 20480 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_7944
timestamp 1668089732
transform 1 0 20480 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_7945
timestamp 1668089732
transform 1 0 20480 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_7946
timestamp 1668089732
transform 1 0 20480 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_7947
timestamp 1668089732
transform 1 0 20480 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_7948
timestamp 1668089732
transform 1 0 20480 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_7949
timestamp 1668089732
transform 1 0 20480 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_7950
timestamp 1668089732
transform 1 0 20480 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_7951
timestamp 1668089732
transform 1 0 20480 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_7952
timestamp 1668089732
transform 1 0 20480 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_7953
timestamp 1668089732
transform 1 0 20480 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_7954
timestamp 1668089732
transform 1 0 20480 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_7955
timestamp 1668089732
transform 1 0 20480 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_7956
timestamp 1668089732
transform 1 0 20480 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_7957
timestamp 1668089732
transform 1 0 20480 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_7958
timestamp 1668089732
transform 1 0 20480 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_7959
timestamp 1668089732
transform 1 0 20480 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_7960
timestamp 1668089732
transform 1 0 20480 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_7961
timestamp 1668089732
transform 1 0 20480 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_7962
timestamp 1668089732
transform 1 0 20480 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_7963
timestamp 1668089732
transform 1 0 20480 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_7964
timestamp 1668089732
transform 1 0 20480 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_7965
timestamp 1668089732
transform 1 0 20480 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_7966
timestamp 1668089732
transform 1 0 20480 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_7967
timestamp 1668089732
transform 1 0 20480 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_7968
timestamp 1668089732
transform 1 0 20480 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_7969
timestamp 1668089732
transform 1 0 20480 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_7970
timestamp 1668089732
transform 1 0 20480 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_7971
timestamp 1668089732
transform 1 0 20480 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_7972
timestamp 1668089732
transform 1 0 20480 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_7973
timestamp 1668089732
transform 1 0 20480 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_7974
timestamp 1668089732
transform 1 0 20480 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_7975
timestamp 1668089732
transform 1 0 20480 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_7976
timestamp 1668089732
transform 1 0 20480 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_7977
timestamp 1668089732
transform 1 0 20480 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_7978
timestamp 1668089732
transform 1 0 20480 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_7979
timestamp 1668089732
transform 1 0 20480 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_7980
timestamp 1668089732
transform 1 0 20480 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_7981
timestamp 1668089732
transform 1 0 20480 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_7982
timestamp 1668089732
transform 1 0 20480 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_7983
timestamp 1668089732
transform 1 0 20480 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_7984
timestamp 1668089732
transform 1 0 20480 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_7985
timestamp 1668089732
transform 1 0 20480 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_7986
timestamp 1668089732
transform 1 0 20480 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_7987
timestamp 1668089732
transform 1 0 20480 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_7988
timestamp 1668089732
transform 1 0 20480 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_7989
timestamp 1668089732
transform 1 0 20480 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_7990
timestamp 1668089732
transform 1 0 20480 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_7991
timestamp 1668089732
transform 1 0 20480 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_7992
timestamp 1668089732
transform 1 0 20480 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_7993
timestamp 1668089732
transform 1 0 20480 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_7994
timestamp 1668089732
transform 1 0 20480 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_7995
timestamp 1668089732
transform 1 0 20480 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_7996
timestamp 1668089732
transform 1 0 20480 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_7997
timestamp 1668089732
transform 1 0 20480 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_7998
timestamp 1668089732
transform 1 0 20640 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_7999
timestamp 1668089732
transform 1 0 20640 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_8000
timestamp 1668089732
transform 1 0 20640 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_8001
timestamp 1668089732
transform 1 0 20640 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_8002
timestamp 1668089732
transform 1 0 20640 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_8003
timestamp 1668089732
transform 1 0 20640 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_8004
timestamp 1668089732
transform 1 0 20640 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_8005
timestamp 1668089732
transform 1 0 20640 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_8006
timestamp 1668089732
transform 1 0 20640 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_8007
timestamp 1668089732
transform 1 0 20640 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_8008
timestamp 1668089732
transform 1 0 20640 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_8009
timestamp 1668089732
transform 1 0 20640 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_8010
timestamp 1668089732
transform 1 0 20640 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_8011
timestamp 1668089732
transform 1 0 20640 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_8012
timestamp 1668089732
transform 1 0 20640 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_8013
timestamp 1668089732
transform 1 0 20640 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_8014
timestamp 1668089732
transform 1 0 20640 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_8015
timestamp 1668089732
transform 1 0 20640 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_8016
timestamp 1668089732
transform 1 0 20640 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_8017
timestamp 1668089732
transform 1 0 20640 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_8018
timestamp 1668089732
transform 1 0 20640 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_8019
timestamp 1668089732
transform 1 0 20640 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_8020
timestamp 1668089732
transform 1 0 20640 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_8021
timestamp 1668089732
transform 1 0 20640 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_8022
timestamp 1668089732
transform 1 0 20640 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_8023
timestamp 1668089732
transform 1 0 20640 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_8024
timestamp 1668089732
transform 1 0 20640 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_8025
timestamp 1668089732
transform 1 0 20640 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_8026
timestamp 1668089732
transform 1 0 20640 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_8027
timestamp 1668089732
transform 1 0 20640 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_8028
timestamp 1668089732
transform 1 0 20640 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_8029
timestamp 1668089732
transform 1 0 20640 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_8030
timestamp 1668089732
transform 1 0 20640 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_8031
timestamp 1668089732
transform 1 0 20640 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_8032
timestamp 1668089732
transform 1 0 20640 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_8033
timestamp 1668089732
transform 1 0 20640 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_8034
timestamp 1668089732
transform 1 0 20640 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_8035
timestamp 1668089732
transform 1 0 20640 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_8036
timestamp 1668089732
transform 1 0 20640 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_8037
timestamp 1668089732
transform 1 0 20640 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_8038
timestamp 1668089732
transform 1 0 20640 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_8039
timestamp 1668089732
transform 1 0 20640 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_8040
timestamp 1668089732
transform 1 0 20640 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_8041
timestamp 1668089732
transform 1 0 20640 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_8042
timestamp 1668089732
transform 1 0 20640 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_8043
timestamp 1668089732
transform 1 0 20640 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_8044
timestamp 1668089732
transform 1 0 20640 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_8045
timestamp 1668089732
transform 1 0 20640 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_8046
timestamp 1668089732
transform 1 0 20640 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_8047
timestamp 1668089732
transform 1 0 20640 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_8048
timestamp 1668089732
transform 1 0 20640 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_8049
timestamp 1668089732
transform 1 0 20640 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_8050
timestamp 1668089732
transform 1 0 20640 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_8051
timestamp 1668089732
transform 1 0 20640 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_8052
timestamp 1668089732
transform 1 0 20640 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_8053
timestamp 1668089732
transform 1 0 20640 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_8054
timestamp 1668089732
transform 1 0 20640 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_8055
timestamp 1668089732
transform 1 0 20640 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_8056
timestamp 1668089732
transform 1 0 20640 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_8057
timestamp 1668089732
transform 1 0 20640 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_8058
timestamp 1668089732
transform 1 0 20640 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_8059
timestamp 1668089732
transform 1 0 20640 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_8060
timestamp 1668089732
transform 1 0 20800 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_8061
timestamp 1668089732
transform 1 0 20800 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_8062
timestamp 1668089732
transform 1 0 20800 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_8063
timestamp 1668089732
transform 1 0 20800 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_8064
timestamp 1668089732
transform 1 0 20800 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_8065
timestamp 1668089732
transform 1 0 20800 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_8066
timestamp 1668089732
transform 1 0 20800 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_8067
timestamp 1668089732
transform 1 0 20800 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_8068
timestamp 1668089732
transform 1 0 20800 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_8069
timestamp 1668089732
transform 1 0 20800 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_8070
timestamp 1668089732
transform 1 0 20800 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_8071
timestamp 1668089732
transform 1 0 20800 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_8072
timestamp 1668089732
transform 1 0 20800 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_8073
timestamp 1668089732
transform 1 0 20800 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_8074
timestamp 1668089732
transform 1 0 20800 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_8075
timestamp 1668089732
transform 1 0 20800 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_8076
timestamp 1668089732
transform 1 0 20800 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_8077
timestamp 1668089732
transform 1 0 20800 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_8078
timestamp 1668089732
transform 1 0 20800 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_8079
timestamp 1668089732
transform 1 0 20800 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_8080
timestamp 1668089732
transform 1 0 20800 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_8081
timestamp 1668089732
transform 1 0 20800 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_8082
timestamp 1668089732
transform 1 0 20800 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_8083
timestamp 1668089732
transform 1 0 20800 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_8084
timestamp 1668089732
transform 1 0 20800 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_8085
timestamp 1668089732
transform 1 0 20800 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_8086
timestamp 1668089732
transform 1 0 20800 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_8087
timestamp 1668089732
transform 1 0 20800 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_8088
timestamp 1668089732
transform 1 0 20800 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_8089
timestamp 1668089732
transform 1 0 20800 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_8090
timestamp 1668089732
transform 1 0 20800 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_8091
timestamp 1668089732
transform 1 0 20800 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_8092
timestamp 1668089732
transform 1 0 20800 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_8093
timestamp 1668089732
transform 1 0 20800 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_8094
timestamp 1668089732
transform 1 0 20800 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_8095
timestamp 1668089732
transform 1 0 20800 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_8096
timestamp 1668089732
transform 1 0 20800 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_8097
timestamp 1668089732
transform 1 0 20800 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_8098
timestamp 1668089732
transform 1 0 20800 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_8099
timestamp 1668089732
transform 1 0 20800 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_8100
timestamp 1668089732
transform 1 0 20800 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_8101
timestamp 1668089732
transform 1 0 20800 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_8102
timestamp 1668089732
transform 1 0 20800 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_8103
timestamp 1668089732
transform 1 0 20800 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_8104
timestamp 1668089732
transform 1 0 20800 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_8105
timestamp 1668089732
transform 1 0 20800 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_8106
timestamp 1668089732
transform 1 0 20800 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_8107
timestamp 1668089732
transform 1 0 20800 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_8108
timestamp 1668089732
transform 1 0 20800 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_8109
timestamp 1668089732
transform 1 0 20800 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_8110
timestamp 1668089732
transform 1 0 20800 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_8111
timestamp 1668089732
transform 1 0 20800 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_8112
timestamp 1668089732
transform 1 0 20800 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_8113
timestamp 1668089732
transform 1 0 20800 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_8114
timestamp 1668089732
transform 1 0 20800 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_8115
timestamp 1668089732
transform 1 0 20800 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_8116
timestamp 1668089732
transform 1 0 20800 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_8117
timestamp 1668089732
transform 1 0 20800 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_8118
timestamp 1668089732
transform 1 0 20800 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_8119
timestamp 1668089732
transform 1 0 20800 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_8120
timestamp 1668089732
transform 1 0 20800 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_8121
timestamp 1668089732
transform 1 0 20800 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_8122
timestamp 1668089732
transform 1 0 20960 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_8123
timestamp 1668089732
transform 1 0 20960 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_8124
timestamp 1668089732
transform 1 0 20960 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_8125
timestamp 1668089732
transform 1 0 20960 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_8126
timestamp 1668089732
transform 1 0 20960 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_8127
timestamp 1668089732
transform 1 0 20960 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_8128
timestamp 1668089732
transform 1 0 20960 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_8129
timestamp 1668089732
transform 1 0 20960 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_8130
timestamp 1668089732
transform 1 0 20960 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_8131
timestamp 1668089732
transform 1 0 20960 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_8132
timestamp 1668089732
transform 1 0 20960 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_8133
timestamp 1668089732
transform 1 0 20960 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_8134
timestamp 1668089732
transform 1 0 20960 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_8135
timestamp 1668089732
transform 1 0 20960 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_8136
timestamp 1668089732
transform 1 0 20960 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_8137
timestamp 1668089732
transform 1 0 20960 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_8138
timestamp 1668089732
transform 1 0 20960 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_8139
timestamp 1668089732
transform 1 0 20960 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_8140
timestamp 1668089732
transform 1 0 20960 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_8141
timestamp 1668089732
transform 1 0 20960 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_8142
timestamp 1668089732
transform 1 0 20960 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_8143
timestamp 1668089732
transform 1 0 20960 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_8144
timestamp 1668089732
transform 1 0 20960 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_8145
timestamp 1668089732
transform 1 0 20960 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_8146
timestamp 1668089732
transform 1 0 20960 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_8147
timestamp 1668089732
transform 1 0 20960 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_8148
timestamp 1668089732
transform 1 0 20960 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_8149
timestamp 1668089732
transform 1 0 20960 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_8150
timestamp 1668089732
transform 1 0 20960 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_8151
timestamp 1668089732
transform 1 0 20960 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_8152
timestamp 1668089732
transform 1 0 20960 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_8153
timestamp 1668089732
transform 1 0 20960 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_8154
timestamp 1668089732
transform 1 0 20960 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_8155
timestamp 1668089732
transform 1 0 20960 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_8156
timestamp 1668089732
transform 1 0 20960 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_8157
timestamp 1668089732
transform 1 0 20960 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_8158
timestamp 1668089732
transform 1 0 20960 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_8159
timestamp 1668089732
transform 1 0 20960 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_8160
timestamp 1668089732
transform 1 0 20960 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_8161
timestamp 1668089732
transform 1 0 20960 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_8162
timestamp 1668089732
transform 1 0 20960 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_8163
timestamp 1668089732
transform 1 0 20960 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_8164
timestamp 1668089732
transform 1 0 20960 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_8165
timestamp 1668089732
transform 1 0 20960 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_8166
timestamp 1668089732
transform 1 0 20960 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_8167
timestamp 1668089732
transform 1 0 20960 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_8168
timestamp 1668089732
transform 1 0 20960 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_8169
timestamp 1668089732
transform 1 0 20960 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_8170
timestamp 1668089732
transform 1 0 20960 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_8171
timestamp 1668089732
transform 1 0 20960 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_8172
timestamp 1668089732
transform 1 0 20960 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_8173
timestamp 1668089732
transform 1 0 20960 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_8174
timestamp 1668089732
transform 1 0 20960 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_8175
timestamp 1668089732
transform 1 0 20960 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_8176
timestamp 1668089732
transform 1 0 20960 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_8177
timestamp 1668089732
transform 1 0 20960 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_8178
timestamp 1668089732
transform 1 0 20960 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_8179
timestamp 1668089732
transform 1 0 20960 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_8180
timestamp 1668089732
transform 1 0 20960 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_8181
timestamp 1668089732
transform 1 0 20960 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_8182
timestamp 1668089732
transform 1 0 20960 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_8183
timestamp 1668089732
transform 1 0 20960 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_8184
timestamp 1668089732
transform 1 0 21120 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_8185
timestamp 1668089732
transform 1 0 21120 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_8186
timestamp 1668089732
transform 1 0 21120 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_8187
timestamp 1668089732
transform 1 0 21120 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_8188
timestamp 1668089732
transform 1 0 21120 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_8189
timestamp 1668089732
transform 1 0 21120 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_8190
timestamp 1668089732
transform 1 0 21120 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_8191
timestamp 1668089732
transform 1 0 21120 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_8192
timestamp 1668089732
transform 1 0 21120 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_8193
timestamp 1668089732
transform 1 0 21120 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_8194
timestamp 1668089732
transform 1 0 21120 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_8195
timestamp 1668089732
transform 1 0 21120 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_8196
timestamp 1668089732
transform 1 0 21120 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_8197
timestamp 1668089732
transform 1 0 21120 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_8198
timestamp 1668089732
transform 1 0 21120 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_8199
timestamp 1668089732
transform 1 0 21120 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_8200
timestamp 1668089732
transform 1 0 21120 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_8201
timestamp 1668089732
transform 1 0 21120 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_8202
timestamp 1668089732
transform 1 0 21120 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_8203
timestamp 1668089732
transform 1 0 21120 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_8204
timestamp 1668089732
transform 1 0 21120 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_8205
timestamp 1668089732
transform 1 0 21120 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_8206
timestamp 1668089732
transform 1 0 21120 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_8207
timestamp 1668089732
transform 1 0 21120 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_8208
timestamp 1668089732
transform 1 0 21120 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_8209
timestamp 1668089732
transform 1 0 21120 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_8210
timestamp 1668089732
transform 1 0 21120 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_8211
timestamp 1668089732
transform 1 0 21120 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_8212
timestamp 1668089732
transform 1 0 21120 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_8213
timestamp 1668089732
transform 1 0 21120 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_8214
timestamp 1668089732
transform 1 0 21120 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_8215
timestamp 1668089732
transform 1 0 21120 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_8216
timestamp 1668089732
transform 1 0 21120 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_8217
timestamp 1668089732
transform 1 0 21120 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_8218
timestamp 1668089732
transform 1 0 21120 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_8219
timestamp 1668089732
transform 1 0 21120 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_8220
timestamp 1668089732
transform 1 0 21120 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_8221
timestamp 1668089732
transform 1 0 21120 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_8222
timestamp 1668089732
transform 1 0 21120 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_8223
timestamp 1668089732
transform 1 0 21120 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_8224
timestamp 1668089732
transform 1 0 21120 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_8225
timestamp 1668089732
transform 1 0 21120 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_8226
timestamp 1668089732
transform 1 0 21120 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_8227
timestamp 1668089732
transform 1 0 21120 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_8228
timestamp 1668089732
transform 1 0 21120 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_8229
timestamp 1668089732
transform 1 0 21120 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_8230
timestamp 1668089732
transform 1 0 21120 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_8231
timestamp 1668089732
transform 1 0 21120 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_8232
timestamp 1668089732
transform 1 0 21120 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_8233
timestamp 1668089732
transform 1 0 21120 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_8234
timestamp 1668089732
transform 1 0 21120 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_8235
timestamp 1668089732
transform 1 0 21120 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_8236
timestamp 1668089732
transform 1 0 21120 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_8237
timestamp 1668089732
transform 1 0 21120 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_8238
timestamp 1668089732
transform 1 0 21120 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_8239
timestamp 1668089732
transform 1 0 21120 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_8240
timestamp 1668089732
transform 1 0 21120 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_8241
timestamp 1668089732
transform 1 0 21120 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_8242
timestamp 1668089732
transform 1 0 21120 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_8243
timestamp 1668089732
transform 1 0 21120 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_8244
timestamp 1668089732
transform 1 0 21120 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_8245
timestamp 1668089732
transform 1 0 21120 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_8246
timestamp 1668089732
transform 1 0 21280 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_8247
timestamp 1668089732
transform 1 0 21280 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_8248
timestamp 1668089732
transform 1 0 21280 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_8249
timestamp 1668089732
transform 1 0 21280 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_8250
timestamp 1668089732
transform 1 0 21280 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_8251
timestamp 1668089732
transform 1 0 21280 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_8252
timestamp 1668089732
transform 1 0 21280 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_8253
timestamp 1668089732
transform 1 0 21280 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_8254
timestamp 1668089732
transform 1 0 21280 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_8255
timestamp 1668089732
transform 1 0 21280 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_8256
timestamp 1668089732
transform 1 0 21280 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_8257
timestamp 1668089732
transform 1 0 21280 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_8258
timestamp 1668089732
transform 1 0 21280 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_8259
timestamp 1668089732
transform 1 0 21280 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_8260
timestamp 1668089732
transform 1 0 21280 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_8261
timestamp 1668089732
transform 1 0 21280 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_8262
timestamp 1668089732
transform 1 0 21280 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_8263
timestamp 1668089732
transform 1 0 21280 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_8264
timestamp 1668089732
transform 1 0 21280 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_8265
timestamp 1668089732
transform 1 0 21280 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_8266
timestamp 1668089732
transform 1 0 21280 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_8267
timestamp 1668089732
transform 1 0 21280 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_8268
timestamp 1668089732
transform 1 0 21280 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_8269
timestamp 1668089732
transform 1 0 21280 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_8270
timestamp 1668089732
transform 1 0 21280 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_8271
timestamp 1668089732
transform 1 0 21280 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_8272
timestamp 1668089732
transform 1 0 21280 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_8273
timestamp 1668089732
transform 1 0 21280 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_8274
timestamp 1668089732
transform 1 0 21280 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_8275
timestamp 1668089732
transform 1 0 21280 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_8276
timestamp 1668089732
transform 1 0 21280 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_8277
timestamp 1668089732
transform 1 0 21280 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_8278
timestamp 1668089732
transform 1 0 21280 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_8279
timestamp 1668089732
transform 1 0 21280 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_8280
timestamp 1668089732
transform 1 0 21280 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_8281
timestamp 1668089732
transform 1 0 21280 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_8282
timestamp 1668089732
transform 1 0 21280 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_8283
timestamp 1668089732
transform 1 0 21280 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_8284
timestamp 1668089732
transform 1 0 21280 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_8285
timestamp 1668089732
transform 1 0 21280 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_8286
timestamp 1668089732
transform 1 0 21280 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_8287
timestamp 1668089732
transform 1 0 21280 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_8288
timestamp 1668089732
transform 1 0 21280 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_8289
timestamp 1668089732
transform 1 0 21280 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_8290
timestamp 1668089732
transform 1 0 21280 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_8291
timestamp 1668089732
transform 1 0 21280 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_8292
timestamp 1668089732
transform 1 0 21280 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_8293
timestamp 1668089732
transform 1 0 21280 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_8294
timestamp 1668089732
transform 1 0 21280 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_8295
timestamp 1668089732
transform 1 0 21280 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_8296
timestamp 1668089732
transform 1 0 21280 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_8297
timestamp 1668089732
transform 1 0 21280 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_8298
timestamp 1668089732
transform 1 0 21280 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_8299
timestamp 1668089732
transform 1 0 21280 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_8300
timestamp 1668089732
transform 1 0 21280 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_8301
timestamp 1668089732
transform 1 0 21280 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_8302
timestamp 1668089732
transform 1 0 21280 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_8303
timestamp 1668089732
transform 1 0 21280 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_8304
timestamp 1668089732
transform 1 0 21280 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_8305
timestamp 1668089732
transform 1 0 21280 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_8306
timestamp 1668089732
transform 1 0 21280 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_8307
timestamp 1668089732
transform 1 0 21280 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_8308
timestamp 1668089732
transform 1 0 21440 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_8309
timestamp 1668089732
transform 1 0 21440 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_8310
timestamp 1668089732
transform 1 0 21440 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_8311
timestamp 1668089732
transform 1 0 21440 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_8312
timestamp 1668089732
transform 1 0 21440 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_8313
timestamp 1668089732
transform 1 0 21440 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_8314
timestamp 1668089732
transform 1 0 21440 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_8315
timestamp 1668089732
transform 1 0 21440 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_8316
timestamp 1668089732
transform 1 0 21440 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_8317
timestamp 1668089732
transform 1 0 21440 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_8318
timestamp 1668089732
transform 1 0 21440 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_8319
timestamp 1668089732
transform 1 0 21440 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_8320
timestamp 1668089732
transform 1 0 21440 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_8321
timestamp 1668089732
transform 1 0 21440 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_8322
timestamp 1668089732
transform 1 0 21440 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_8323
timestamp 1668089732
transform 1 0 21440 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_8324
timestamp 1668089732
transform 1 0 21440 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_8325
timestamp 1668089732
transform 1 0 21440 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_8326
timestamp 1668089732
transform 1 0 21440 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_8327
timestamp 1668089732
transform 1 0 21440 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_8328
timestamp 1668089732
transform 1 0 21440 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_8329
timestamp 1668089732
transform 1 0 21440 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_8330
timestamp 1668089732
transform 1 0 21440 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_8331
timestamp 1668089732
transform 1 0 21440 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_8332
timestamp 1668089732
transform 1 0 21440 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_8333
timestamp 1668089732
transform 1 0 21440 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_8334
timestamp 1668089732
transform 1 0 21440 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_8335
timestamp 1668089732
transform 1 0 21440 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_8336
timestamp 1668089732
transform 1 0 21440 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_8337
timestamp 1668089732
transform 1 0 21440 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_8338
timestamp 1668089732
transform 1 0 21440 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_8339
timestamp 1668089732
transform 1 0 21440 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_8340
timestamp 1668089732
transform 1 0 21440 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_8341
timestamp 1668089732
transform 1 0 21440 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_8342
timestamp 1668089732
transform 1 0 21440 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_8343
timestamp 1668089732
transform 1 0 21440 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_8344
timestamp 1668089732
transform 1 0 21440 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_8345
timestamp 1668089732
transform 1 0 21440 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_8346
timestamp 1668089732
transform 1 0 21440 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_8347
timestamp 1668089732
transform 1 0 21440 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_8348
timestamp 1668089732
transform 1 0 21440 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_8349
timestamp 1668089732
transform 1 0 21440 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_8350
timestamp 1668089732
transform 1 0 21440 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_8351
timestamp 1668089732
transform 1 0 21440 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_8352
timestamp 1668089732
transform 1 0 21440 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_8353
timestamp 1668089732
transform 1 0 21440 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_8354
timestamp 1668089732
transform 1 0 21440 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_8355
timestamp 1668089732
transform 1 0 21440 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_8356
timestamp 1668089732
transform 1 0 21440 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_8357
timestamp 1668089732
transform 1 0 21440 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_8358
timestamp 1668089732
transform 1 0 21440 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_8359
timestamp 1668089732
transform 1 0 21440 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_8360
timestamp 1668089732
transform 1 0 21440 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_8361
timestamp 1668089732
transform 1 0 21440 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_8362
timestamp 1668089732
transform 1 0 21440 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_8363
timestamp 1668089732
transform 1 0 21440 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_8364
timestamp 1668089732
transform 1 0 21440 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_8365
timestamp 1668089732
transform 1 0 21440 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_8366
timestamp 1668089732
transform 1 0 21440 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_8367
timestamp 1668089732
transform 1 0 21440 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_8368
timestamp 1668089732
transform 1 0 21440 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_8369
timestamp 1668089732
transform 1 0 21440 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_8370
timestamp 1668089732
transform 1 0 21600 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_8371
timestamp 1668089732
transform 1 0 21600 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_8372
timestamp 1668089732
transform 1 0 21600 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_8373
timestamp 1668089732
transform 1 0 21600 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_8374
timestamp 1668089732
transform 1 0 21600 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_8375
timestamp 1668089732
transform 1 0 21600 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_8376
timestamp 1668089732
transform 1 0 21600 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_8377
timestamp 1668089732
transform 1 0 21600 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_8378
timestamp 1668089732
transform 1 0 21600 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_8379
timestamp 1668089732
transform 1 0 21600 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_8380
timestamp 1668089732
transform 1 0 21600 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_8381
timestamp 1668089732
transform 1 0 21600 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_8382
timestamp 1668089732
transform 1 0 21600 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_8383
timestamp 1668089732
transform 1 0 21600 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_8384
timestamp 1668089732
transform 1 0 21600 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_8385
timestamp 1668089732
transform 1 0 21600 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_8386
timestamp 1668089732
transform 1 0 21600 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_8387
timestamp 1668089732
transform 1 0 21600 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_8388
timestamp 1668089732
transform 1 0 21600 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_8389
timestamp 1668089732
transform 1 0 21600 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_8390
timestamp 1668089732
transform 1 0 21600 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_8391
timestamp 1668089732
transform 1 0 21600 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_8392
timestamp 1668089732
transform 1 0 21600 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_8393
timestamp 1668089732
transform 1 0 21600 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_8394
timestamp 1668089732
transform 1 0 21600 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_8395
timestamp 1668089732
transform 1 0 21600 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_8396
timestamp 1668089732
transform 1 0 21600 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_8397
timestamp 1668089732
transform 1 0 21600 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_8398
timestamp 1668089732
transform 1 0 21600 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_8399
timestamp 1668089732
transform 1 0 21600 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_8400
timestamp 1668089732
transform 1 0 21600 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_8401
timestamp 1668089732
transform 1 0 21600 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_8402
timestamp 1668089732
transform 1 0 21600 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_8403
timestamp 1668089732
transform 1 0 21600 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_8404
timestamp 1668089732
transform 1 0 21600 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_8405
timestamp 1668089732
transform 1 0 21600 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_8406
timestamp 1668089732
transform 1 0 21600 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_8407
timestamp 1668089732
transform 1 0 21600 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_8408
timestamp 1668089732
transform 1 0 21600 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_8409
timestamp 1668089732
transform 1 0 21600 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_8410
timestamp 1668089732
transform 1 0 21600 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_8411
timestamp 1668089732
transform 1 0 21600 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_8412
timestamp 1668089732
transform 1 0 21600 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_8413
timestamp 1668089732
transform 1 0 21600 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_8414
timestamp 1668089732
transform 1 0 21600 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_8415
timestamp 1668089732
transform 1 0 21600 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_8416
timestamp 1668089732
transform 1 0 21600 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_8417
timestamp 1668089732
transform 1 0 21600 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_8418
timestamp 1668089732
transform 1 0 21600 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_8419
timestamp 1668089732
transform 1 0 21600 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_8420
timestamp 1668089732
transform 1 0 21600 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_8421
timestamp 1668089732
transform 1 0 21600 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_8422
timestamp 1668089732
transform 1 0 21600 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_8423
timestamp 1668089732
transform 1 0 21600 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_8424
timestamp 1668089732
transform 1 0 21600 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_8425
timestamp 1668089732
transform 1 0 21600 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_8426
timestamp 1668089732
transform 1 0 21600 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_8427
timestamp 1668089732
transform 1 0 21600 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_8428
timestamp 1668089732
transform 1 0 21600 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_8429
timestamp 1668089732
transform 1 0 21600 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_8430
timestamp 1668089732
transform 1 0 21600 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_8431
timestamp 1668089732
transform 1 0 21600 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_8432
timestamp 1668089732
transform 1 0 21760 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_8433
timestamp 1668089732
transform 1 0 21760 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_8434
timestamp 1668089732
transform 1 0 21760 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_8435
timestamp 1668089732
transform 1 0 21760 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_8436
timestamp 1668089732
transform 1 0 21760 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_8437
timestamp 1668089732
transform 1 0 21760 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_8438
timestamp 1668089732
transform 1 0 21760 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_8439
timestamp 1668089732
transform 1 0 21760 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_8440
timestamp 1668089732
transform 1 0 21760 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_8441
timestamp 1668089732
transform 1 0 21760 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_8442
timestamp 1668089732
transform 1 0 21760 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_8443
timestamp 1668089732
transform 1 0 21760 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_8444
timestamp 1668089732
transform 1 0 21760 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_8445
timestamp 1668089732
transform 1 0 21760 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_8446
timestamp 1668089732
transform 1 0 21760 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_8447
timestamp 1668089732
transform 1 0 21760 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_8448
timestamp 1668089732
transform 1 0 21760 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_8449
timestamp 1668089732
transform 1 0 21760 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_8450
timestamp 1668089732
transform 1 0 21760 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_8451
timestamp 1668089732
transform 1 0 21760 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_8452
timestamp 1668089732
transform 1 0 21760 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_8453
timestamp 1668089732
transform 1 0 21760 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_8454
timestamp 1668089732
transform 1 0 21760 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_8455
timestamp 1668089732
transform 1 0 21760 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_8456
timestamp 1668089732
transform 1 0 21760 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_8457
timestamp 1668089732
transform 1 0 21760 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_8458
timestamp 1668089732
transform 1 0 21760 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_8459
timestamp 1668089732
transform 1 0 21760 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_8460
timestamp 1668089732
transform 1 0 21760 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_8461
timestamp 1668089732
transform 1 0 21760 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_8462
timestamp 1668089732
transform 1 0 21760 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_8463
timestamp 1668089732
transform 1 0 21760 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_8464
timestamp 1668089732
transform 1 0 21760 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_8465
timestamp 1668089732
transform 1 0 21760 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_8466
timestamp 1668089732
transform 1 0 21760 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_8467
timestamp 1668089732
transform 1 0 21760 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_8468
timestamp 1668089732
transform 1 0 21760 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_8469
timestamp 1668089732
transform 1 0 21760 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_8470
timestamp 1668089732
transform 1 0 21760 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_8471
timestamp 1668089732
transform 1 0 21760 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_8472
timestamp 1668089732
transform 1 0 21760 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_8473
timestamp 1668089732
transform 1 0 21760 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_8474
timestamp 1668089732
transform 1 0 21760 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_8475
timestamp 1668089732
transform 1 0 21760 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_8476
timestamp 1668089732
transform 1 0 21760 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_8477
timestamp 1668089732
transform 1 0 21760 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_8478
timestamp 1668089732
transform 1 0 21760 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_8479
timestamp 1668089732
transform 1 0 21760 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_8480
timestamp 1668089732
transform 1 0 21760 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_8481
timestamp 1668089732
transform 1 0 21760 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_8482
timestamp 1668089732
transform 1 0 21760 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_8483
timestamp 1668089732
transform 1 0 21760 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_8484
timestamp 1668089732
transform 1 0 21760 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_8485
timestamp 1668089732
transform 1 0 21760 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_8486
timestamp 1668089732
transform 1 0 21760 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_8487
timestamp 1668089732
transform 1 0 21760 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_8488
timestamp 1668089732
transform 1 0 21760 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_8489
timestamp 1668089732
transform 1 0 21760 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_8490
timestamp 1668089732
transform 1 0 21760 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_8491
timestamp 1668089732
transform 1 0 21760 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_8492
timestamp 1668089732
transform 1 0 21760 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_8493
timestamp 1668089732
transform 1 0 21760 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_8494
timestamp 1668089732
transform 1 0 21920 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_8495
timestamp 1668089732
transform 1 0 21920 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_8496
timestamp 1668089732
transform 1 0 21920 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_8497
timestamp 1668089732
transform 1 0 21920 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_8498
timestamp 1668089732
transform 1 0 21920 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_8499
timestamp 1668089732
transform 1 0 21920 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_8500
timestamp 1668089732
transform 1 0 21920 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_8501
timestamp 1668089732
transform 1 0 21920 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_8502
timestamp 1668089732
transform 1 0 21920 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_8503
timestamp 1668089732
transform 1 0 21920 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_8504
timestamp 1668089732
transform 1 0 21920 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_8505
timestamp 1668089732
transform 1 0 21920 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_8506
timestamp 1668089732
transform 1 0 21920 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_8507
timestamp 1668089732
transform 1 0 21920 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_8508
timestamp 1668089732
transform 1 0 21920 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_8509
timestamp 1668089732
transform 1 0 21920 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_8510
timestamp 1668089732
transform 1 0 21920 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_8511
timestamp 1668089732
transform 1 0 21920 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_8512
timestamp 1668089732
transform 1 0 21920 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_8513
timestamp 1668089732
transform 1 0 21920 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_8514
timestamp 1668089732
transform 1 0 21920 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_8515
timestamp 1668089732
transform 1 0 21920 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_8516
timestamp 1668089732
transform 1 0 21920 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_8517
timestamp 1668089732
transform 1 0 21920 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_8518
timestamp 1668089732
transform 1 0 21920 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_8519
timestamp 1668089732
transform 1 0 21920 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_8520
timestamp 1668089732
transform 1 0 21920 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_8521
timestamp 1668089732
transform 1 0 21920 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_8522
timestamp 1668089732
transform 1 0 21920 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_8523
timestamp 1668089732
transform 1 0 21920 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_8524
timestamp 1668089732
transform 1 0 21920 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_8525
timestamp 1668089732
transform 1 0 21920 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_8526
timestamp 1668089732
transform 1 0 21920 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_8527
timestamp 1668089732
transform 1 0 21920 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_8528
timestamp 1668089732
transform 1 0 21920 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_8529
timestamp 1668089732
transform 1 0 21920 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_8530
timestamp 1668089732
transform 1 0 21920 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_8531
timestamp 1668089732
transform 1 0 21920 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_8532
timestamp 1668089732
transform 1 0 21920 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_8533
timestamp 1668089732
transform 1 0 21920 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_8534
timestamp 1668089732
transform 1 0 21920 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_8535
timestamp 1668089732
transform 1 0 21920 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_8536
timestamp 1668089732
transform 1 0 21920 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_8537
timestamp 1668089732
transform 1 0 21920 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_8538
timestamp 1668089732
transform 1 0 21920 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_8539
timestamp 1668089732
transform 1 0 21920 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_8540
timestamp 1668089732
transform 1 0 21920 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_8541
timestamp 1668089732
transform 1 0 21920 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_8542
timestamp 1668089732
transform 1 0 21920 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_8543
timestamp 1668089732
transform 1 0 21920 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_8544
timestamp 1668089732
transform 1 0 21920 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_8545
timestamp 1668089732
transform 1 0 21920 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_8546
timestamp 1668089732
transform 1 0 21920 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_8547
timestamp 1668089732
transform 1 0 21920 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_8548
timestamp 1668089732
transform 1 0 21920 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_8549
timestamp 1668089732
transform 1 0 21920 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_8550
timestamp 1668089732
transform 1 0 21920 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_8551
timestamp 1668089732
transform 1 0 21920 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_8552
timestamp 1668089732
transform 1 0 21920 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_8553
timestamp 1668089732
transform 1 0 21920 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_8554
timestamp 1668089732
transform 1 0 21920 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_8555
timestamp 1668089732
transform 1 0 21920 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_8556
timestamp 1668089732
transform 1 0 22080 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_8557
timestamp 1668089732
transform 1 0 22080 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_8558
timestamp 1668089732
transform 1 0 22080 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_8559
timestamp 1668089732
transform 1 0 22080 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_8560
timestamp 1668089732
transform 1 0 22080 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_8561
timestamp 1668089732
transform 1 0 22080 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_8562
timestamp 1668089732
transform 1 0 22080 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_8563
timestamp 1668089732
transform 1 0 22080 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_8564
timestamp 1668089732
transform 1 0 22080 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_8565
timestamp 1668089732
transform 1 0 22080 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_8566
timestamp 1668089732
transform 1 0 22080 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_8567
timestamp 1668089732
transform 1 0 22080 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_8568
timestamp 1668089732
transform 1 0 22080 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_8569
timestamp 1668089732
transform 1 0 22080 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_8570
timestamp 1668089732
transform 1 0 22080 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_8571
timestamp 1668089732
transform 1 0 22080 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_8572
timestamp 1668089732
transform 1 0 22080 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_8573
timestamp 1668089732
transform 1 0 22080 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_8574
timestamp 1668089732
transform 1 0 22080 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_8575
timestamp 1668089732
transform 1 0 22080 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_8576
timestamp 1668089732
transform 1 0 22080 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_8577
timestamp 1668089732
transform 1 0 22080 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_8578
timestamp 1668089732
transform 1 0 22080 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_8579
timestamp 1668089732
transform 1 0 22080 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_8580
timestamp 1668089732
transform 1 0 22080 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_8581
timestamp 1668089732
transform 1 0 22080 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_8582
timestamp 1668089732
transform 1 0 22080 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_8583
timestamp 1668089732
transform 1 0 22080 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_8584
timestamp 1668089732
transform 1 0 22080 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_8585
timestamp 1668089732
transform 1 0 22080 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_8586
timestamp 1668089732
transform 1 0 22080 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_8587
timestamp 1668089732
transform 1 0 22080 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_8588
timestamp 1668089732
transform 1 0 22080 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_8589
timestamp 1668089732
transform 1 0 22080 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_8590
timestamp 1668089732
transform 1 0 22080 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_8591
timestamp 1668089732
transform 1 0 22080 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_8592
timestamp 1668089732
transform 1 0 22080 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_8593
timestamp 1668089732
transform 1 0 22080 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_8594
timestamp 1668089732
transform 1 0 22080 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_8595
timestamp 1668089732
transform 1 0 22080 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_8596
timestamp 1668089732
transform 1 0 22080 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_8597
timestamp 1668089732
transform 1 0 22080 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_8598
timestamp 1668089732
transform 1 0 22080 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_8599
timestamp 1668089732
transform 1 0 22080 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_8600
timestamp 1668089732
transform 1 0 22080 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_8601
timestamp 1668089732
transform 1 0 22080 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_8602
timestamp 1668089732
transform 1 0 22080 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_8603
timestamp 1668089732
transform 1 0 22080 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_8604
timestamp 1668089732
transform 1 0 22080 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_8605
timestamp 1668089732
transform 1 0 22080 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_8606
timestamp 1668089732
transform 1 0 22080 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_8607
timestamp 1668089732
transform 1 0 22080 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_8608
timestamp 1668089732
transform 1 0 22080 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_8609
timestamp 1668089732
transform 1 0 22080 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_8610
timestamp 1668089732
transform 1 0 22080 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_8611
timestamp 1668089732
transform 1 0 22080 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_8612
timestamp 1668089732
transform 1 0 22080 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_8613
timestamp 1668089732
transform 1 0 22080 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_8614
timestamp 1668089732
transform 1 0 22080 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_8615
timestamp 1668089732
transform 1 0 22080 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_8616
timestamp 1668089732
transform 1 0 22080 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_8617
timestamp 1668089732
transform 1 0 22080 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_8618
timestamp 1668089732
transform 1 0 22240 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_8619
timestamp 1668089732
transform 1 0 22240 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_8620
timestamp 1668089732
transform 1 0 22240 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_8621
timestamp 1668089732
transform 1 0 22240 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_8622
timestamp 1668089732
transform 1 0 22240 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_8623
timestamp 1668089732
transform 1 0 22240 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_8624
timestamp 1668089732
transform 1 0 22240 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_8625
timestamp 1668089732
transform 1 0 22240 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_8626
timestamp 1668089732
transform 1 0 22240 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_8627
timestamp 1668089732
transform 1 0 22240 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_8628
timestamp 1668089732
transform 1 0 22240 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_8629
timestamp 1668089732
transform 1 0 22240 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_8630
timestamp 1668089732
transform 1 0 22240 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_8631
timestamp 1668089732
transform 1 0 22240 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_8632
timestamp 1668089732
transform 1 0 22240 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_8633
timestamp 1668089732
transform 1 0 22240 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_8634
timestamp 1668089732
transform 1 0 22240 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_8635
timestamp 1668089732
transform 1 0 22240 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_8636
timestamp 1668089732
transform 1 0 22240 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_8637
timestamp 1668089732
transform 1 0 22240 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_8638
timestamp 1668089732
transform 1 0 22240 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_8639
timestamp 1668089732
transform 1 0 22240 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_8640
timestamp 1668089732
transform 1 0 22240 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_8641
timestamp 1668089732
transform 1 0 22240 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_8642
timestamp 1668089732
transform 1 0 22240 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_8643
timestamp 1668089732
transform 1 0 22240 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_8644
timestamp 1668089732
transform 1 0 22240 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_8645
timestamp 1668089732
transform 1 0 22240 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_8646
timestamp 1668089732
transform 1 0 22240 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_8647
timestamp 1668089732
transform 1 0 22240 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_8648
timestamp 1668089732
transform 1 0 22240 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_8649
timestamp 1668089732
transform 1 0 22240 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_8650
timestamp 1668089732
transform 1 0 22240 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_8651
timestamp 1668089732
transform 1 0 22240 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_8652
timestamp 1668089732
transform 1 0 22240 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_8653
timestamp 1668089732
transform 1 0 22240 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_8654
timestamp 1668089732
transform 1 0 22240 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_8655
timestamp 1668089732
transform 1 0 22240 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_8656
timestamp 1668089732
transform 1 0 22240 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_8657
timestamp 1668089732
transform 1 0 22240 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_8658
timestamp 1668089732
transform 1 0 22240 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_8659
timestamp 1668089732
transform 1 0 22240 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_8660
timestamp 1668089732
transform 1 0 22240 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_8661
timestamp 1668089732
transform 1 0 22240 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_8662
timestamp 1668089732
transform 1 0 22240 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_8663
timestamp 1668089732
transform 1 0 22240 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_8664
timestamp 1668089732
transform 1 0 22240 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_8665
timestamp 1668089732
transform 1 0 22240 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_8666
timestamp 1668089732
transform 1 0 22240 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_8667
timestamp 1668089732
transform 1 0 22240 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_8668
timestamp 1668089732
transform 1 0 22240 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_8669
timestamp 1668089732
transform 1 0 22240 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_8670
timestamp 1668089732
transform 1 0 22240 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_8671
timestamp 1668089732
transform 1 0 22240 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_8672
timestamp 1668089732
transform 1 0 22240 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_8673
timestamp 1668089732
transform 1 0 22240 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_8674
timestamp 1668089732
transform 1 0 22240 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_8675
timestamp 1668089732
transform 1 0 22240 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_8676
timestamp 1668089732
transform 1 0 22240 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_8677
timestamp 1668089732
transform 1 0 22240 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_8678
timestamp 1668089732
transform 1 0 22240 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_8679
timestamp 1668089732
transform 1 0 22240 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_8680
timestamp 1668089732
transform 1 0 22400 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_8681
timestamp 1668089732
transform 1 0 22400 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_8682
timestamp 1668089732
transform 1 0 22400 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_8683
timestamp 1668089732
transform 1 0 22400 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_8684
timestamp 1668089732
transform 1 0 22400 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_8685
timestamp 1668089732
transform 1 0 22400 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_8686
timestamp 1668089732
transform 1 0 22400 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_8687
timestamp 1668089732
transform 1 0 22400 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_8688
timestamp 1668089732
transform 1 0 22400 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_8689
timestamp 1668089732
transform 1 0 22400 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_8690
timestamp 1668089732
transform 1 0 22400 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_8691
timestamp 1668089732
transform 1 0 22400 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_8692
timestamp 1668089732
transform 1 0 22400 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_8693
timestamp 1668089732
transform 1 0 22400 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_8694
timestamp 1668089732
transform 1 0 22400 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_8695
timestamp 1668089732
transform 1 0 22400 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_8696
timestamp 1668089732
transform 1 0 22400 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_8697
timestamp 1668089732
transform 1 0 22400 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_8698
timestamp 1668089732
transform 1 0 22400 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_8699
timestamp 1668089732
transform 1 0 22400 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_8700
timestamp 1668089732
transform 1 0 22400 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_8701
timestamp 1668089732
transform 1 0 22400 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_8702
timestamp 1668089732
transform 1 0 22400 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_8703
timestamp 1668089732
transform 1 0 22400 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_8704
timestamp 1668089732
transform 1 0 22400 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_8705
timestamp 1668089732
transform 1 0 22400 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_8706
timestamp 1668089732
transform 1 0 22400 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_8707
timestamp 1668089732
transform 1 0 22400 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_8708
timestamp 1668089732
transform 1 0 22400 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_8709
timestamp 1668089732
transform 1 0 22400 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_8710
timestamp 1668089732
transform 1 0 22400 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_8711
timestamp 1668089732
transform 1 0 22400 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_8712
timestamp 1668089732
transform 1 0 22400 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_8713
timestamp 1668089732
transform 1 0 22400 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_8714
timestamp 1668089732
transform 1 0 22400 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_8715
timestamp 1668089732
transform 1 0 22400 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_8716
timestamp 1668089732
transform 1 0 22400 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_8717
timestamp 1668089732
transform 1 0 22400 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_8718
timestamp 1668089732
transform 1 0 22400 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_8719
timestamp 1668089732
transform 1 0 22400 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_8720
timestamp 1668089732
transform 1 0 22400 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_8721
timestamp 1668089732
transform 1 0 22400 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_8722
timestamp 1668089732
transform 1 0 22400 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_8723
timestamp 1668089732
transform 1 0 22400 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_8724
timestamp 1668089732
transform 1 0 22400 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_8725
timestamp 1668089732
transform 1 0 22400 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_8726
timestamp 1668089732
transform 1 0 22400 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_8727
timestamp 1668089732
transform 1 0 22400 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_8728
timestamp 1668089732
transform 1 0 22400 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_8729
timestamp 1668089732
transform 1 0 22400 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_8730
timestamp 1668089732
transform 1 0 22400 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_8731
timestamp 1668089732
transform 1 0 22400 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_8732
timestamp 1668089732
transform 1 0 22400 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_8733
timestamp 1668089732
transform 1 0 22400 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_8734
timestamp 1668089732
transform 1 0 22400 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_8735
timestamp 1668089732
transform 1 0 22400 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_8736
timestamp 1668089732
transform 1 0 22400 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_8737
timestamp 1668089732
transform 1 0 22400 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_8738
timestamp 1668089732
transform 1 0 22400 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_8739
timestamp 1668089732
transform 1 0 22400 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_8740
timestamp 1668089732
transform 1 0 22400 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_8741
timestamp 1668089732
transform 1 0 22400 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_8742
timestamp 1668089732
transform 1 0 22560 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_8743
timestamp 1668089732
transform 1 0 22560 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_8744
timestamp 1668089732
transform 1 0 22560 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_8745
timestamp 1668089732
transform 1 0 22560 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_8746
timestamp 1668089732
transform 1 0 22560 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_8747
timestamp 1668089732
transform 1 0 22560 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_8748
timestamp 1668089732
transform 1 0 22560 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_8749
timestamp 1668089732
transform 1 0 22560 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_8750
timestamp 1668089732
transform 1 0 22560 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_8751
timestamp 1668089732
transform 1 0 22560 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_8752
timestamp 1668089732
transform 1 0 22560 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_8753
timestamp 1668089732
transform 1 0 22560 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_8754
timestamp 1668089732
transform 1 0 22560 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_8755
timestamp 1668089732
transform 1 0 22560 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_8756
timestamp 1668089732
transform 1 0 22560 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_8757
timestamp 1668089732
transform 1 0 22560 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_8758
timestamp 1668089732
transform 1 0 22560 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_8759
timestamp 1668089732
transform 1 0 22560 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_8760
timestamp 1668089732
transform 1 0 22560 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_8761
timestamp 1668089732
transform 1 0 22560 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_8762
timestamp 1668089732
transform 1 0 22560 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_8763
timestamp 1668089732
transform 1 0 22560 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_8764
timestamp 1668089732
transform 1 0 22560 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_8765
timestamp 1668089732
transform 1 0 22560 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_8766
timestamp 1668089732
transform 1 0 22560 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_8767
timestamp 1668089732
transform 1 0 22560 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_8768
timestamp 1668089732
transform 1 0 22560 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_8769
timestamp 1668089732
transform 1 0 22560 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_8770
timestamp 1668089732
transform 1 0 22560 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_8771
timestamp 1668089732
transform 1 0 22560 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_8772
timestamp 1668089732
transform 1 0 22560 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_8773
timestamp 1668089732
transform 1 0 22560 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_8774
timestamp 1668089732
transform 1 0 22560 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_8775
timestamp 1668089732
transform 1 0 22560 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_8776
timestamp 1668089732
transform 1 0 22560 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_8777
timestamp 1668089732
transform 1 0 22560 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_8778
timestamp 1668089732
transform 1 0 22560 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_8779
timestamp 1668089732
transform 1 0 22560 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_8780
timestamp 1668089732
transform 1 0 22560 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_8781
timestamp 1668089732
transform 1 0 22560 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_8782
timestamp 1668089732
transform 1 0 22560 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_8783
timestamp 1668089732
transform 1 0 22560 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_8784
timestamp 1668089732
transform 1 0 22560 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_8785
timestamp 1668089732
transform 1 0 22560 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_8786
timestamp 1668089732
transform 1 0 22560 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_8787
timestamp 1668089732
transform 1 0 22560 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_8788
timestamp 1668089732
transform 1 0 22560 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_8789
timestamp 1668089732
transform 1 0 22560 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_8790
timestamp 1668089732
transform 1 0 22560 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_8791
timestamp 1668089732
transform 1 0 22560 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_8792
timestamp 1668089732
transform 1 0 22560 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_8793
timestamp 1668089732
transform 1 0 22560 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_8794
timestamp 1668089732
transform 1 0 22560 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_8795
timestamp 1668089732
transform 1 0 22560 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_8796
timestamp 1668089732
transform 1 0 22560 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_8797
timestamp 1668089732
transform 1 0 22560 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_8798
timestamp 1668089732
transform 1 0 22560 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_8799
timestamp 1668089732
transform 1 0 22560 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_8800
timestamp 1668089732
transform 1 0 22560 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_8801
timestamp 1668089732
transform 1 0 22560 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_8802
timestamp 1668089732
transform 1 0 22560 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_8803
timestamp 1668089732
transform 1 0 22560 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_8804
timestamp 1668089732
transform 1 0 22720 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_8805
timestamp 1668089732
transform 1 0 22720 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_8806
timestamp 1668089732
transform 1 0 22720 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_8807
timestamp 1668089732
transform 1 0 22720 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_8808
timestamp 1668089732
transform 1 0 22720 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_8809
timestamp 1668089732
transform 1 0 22720 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_8810
timestamp 1668089732
transform 1 0 22720 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_8811
timestamp 1668089732
transform 1 0 22720 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_8812
timestamp 1668089732
transform 1 0 22720 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_8813
timestamp 1668089732
transform 1 0 22720 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_8814
timestamp 1668089732
transform 1 0 22720 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_8815
timestamp 1668089732
transform 1 0 22720 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_8816
timestamp 1668089732
transform 1 0 22720 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_8817
timestamp 1668089732
transform 1 0 22720 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_8818
timestamp 1668089732
transform 1 0 22720 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_8819
timestamp 1668089732
transform 1 0 22720 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_8820
timestamp 1668089732
transform 1 0 22720 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_8821
timestamp 1668089732
transform 1 0 22720 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_8822
timestamp 1668089732
transform 1 0 22720 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_8823
timestamp 1668089732
transform 1 0 22720 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_8824
timestamp 1668089732
transform 1 0 22720 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_8825
timestamp 1668089732
transform 1 0 22720 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_8826
timestamp 1668089732
transform 1 0 22720 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_8827
timestamp 1668089732
transform 1 0 22720 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_8828
timestamp 1668089732
transform 1 0 22720 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_8829
timestamp 1668089732
transform 1 0 22720 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_8830
timestamp 1668089732
transform 1 0 22720 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_8831
timestamp 1668089732
transform 1 0 22720 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_8832
timestamp 1668089732
transform 1 0 22720 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_8833
timestamp 1668089732
transform 1 0 22720 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_8834
timestamp 1668089732
transform 1 0 22720 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_8835
timestamp 1668089732
transform 1 0 22720 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_8836
timestamp 1668089732
transform 1 0 22720 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_8837
timestamp 1668089732
transform 1 0 22720 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_8838
timestamp 1668089732
transform 1 0 22720 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_8839
timestamp 1668089732
transform 1 0 22720 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_8840
timestamp 1668089732
transform 1 0 22720 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_8841
timestamp 1668089732
transform 1 0 22720 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_8842
timestamp 1668089732
transform 1 0 22720 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_8843
timestamp 1668089732
transform 1 0 22720 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_8844
timestamp 1668089732
transform 1 0 22720 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_8845
timestamp 1668089732
transform 1 0 22720 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_8846
timestamp 1668089732
transform 1 0 22720 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_8847
timestamp 1668089732
transform 1 0 22720 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_8848
timestamp 1668089732
transform 1 0 22720 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_8849
timestamp 1668089732
transform 1 0 22720 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_8850
timestamp 1668089732
transform 1 0 22720 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_8851
timestamp 1668089732
transform 1 0 22720 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_8852
timestamp 1668089732
transform 1 0 22720 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_8853
timestamp 1668089732
transform 1 0 22720 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_8854
timestamp 1668089732
transform 1 0 22720 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_8855
timestamp 1668089732
transform 1 0 22720 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_8856
timestamp 1668089732
transform 1 0 22720 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_8857
timestamp 1668089732
transform 1 0 22720 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_8858
timestamp 1668089732
transform 1 0 22720 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_8859
timestamp 1668089732
transform 1 0 22720 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_8860
timestamp 1668089732
transform 1 0 22720 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_8861
timestamp 1668089732
transform 1 0 22720 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_8862
timestamp 1668089732
transform 1 0 22720 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_8863
timestamp 1668089732
transform 1 0 22720 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_8864
timestamp 1668089732
transform 1 0 22720 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_8865
timestamp 1668089732
transform 1 0 22720 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_8866
timestamp 1668089732
transform 1 0 22880 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_8867
timestamp 1668089732
transform 1 0 22880 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_8868
timestamp 1668089732
transform 1 0 22880 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_8869
timestamp 1668089732
transform 1 0 22880 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_8870
timestamp 1668089732
transform 1 0 22880 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_8871
timestamp 1668089732
transform 1 0 22880 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_8872
timestamp 1668089732
transform 1 0 22880 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_8873
timestamp 1668089732
transform 1 0 22880 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_8874
timestamp 1668089732
transform 1 0 22880 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_8875
timestamp 1668089732
transform 1 0 22880 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_8876
timestamp 1668089732
transform 1 0 22880 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_8877
timestamp 1668089732
transform 1 0 22880 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_8878
timestamp 1668089732
transform 1 0 22880 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_8879
timestamp 1668089732
transform 1 0 22880 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_8880
timestamp 1668089732
transform 1 0 22880 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_8881
timestamp 1668089732
transform 1 0 22880 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_8882
timestamp 1668089732
transform 1 0 22880 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_8883
timestamp 1668089732
transform 1 0 22880 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_8884
timestamp 1668089732
transform 1 0 22880 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_8885
timestamp 1668089732
transform 1 0 22880 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_8886
timestamp 1668089732
transform 1 0 22880 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_8887
timestamp 1668089732
transform 1 0 22880 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_8888
timestamp 1668089732
transform 1 0 22880 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_8889
timestamp 1668089732
transform 1 0 22880 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_8890
timestamp 1668089732
transform 1 0 22880 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_8891
timestamp 1668089732
transform 1 0 22880 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_8892
timestamp 1668089732
transform 1 0 22880 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_8893
timestamp 1668089732
transform 1 0 22880 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_8894
timestamp 1668089732
transform 1 0 22880 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_8895
timestamp 1668089732
transform 1 0 22880 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_8896
timestamp 1668089732
transform 1 0 22880 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_8897
timestamp 1668089732
transform 1 0 22880 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_8898
timestamp 1668089732
transform 1 0 22880 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_8899
timestamp 1668089732
transform 1 0 22880 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_8900
timestamp 1668089732
transform 1 0 22880 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_8901
timestamp 1668089732
transform 1 0 22880 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_8902
timestamp 1668089732
transform 1 0 22880 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_8903
timestamp 1668089732
transform 1 0 22880 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_8904
timestamp 1668089732
transform 1 0 22880 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_8905
timestamp 1668089732
transform 1 0 22880 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_8906
timestamp 1668089732
transform 1 0 22880 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_8907
timestamp 1668089732
transform 1 0 22880 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_8908
timestamp 1668089732
transform 1 0 22880 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_8909
timestamp 1668089732
transform 1 0 22880 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_8910
timestamp 1668089732
transform 1 0 22880 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_8911
timestamp 1668089732
transform 1 0 22880 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_8912
timestamp 1668089732
transform 1 0 22880 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_8913
timestamp 1668089732
transform 1 0 22880 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_8914
timestamp 1668089732
transform 1 0 22880 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_8915
timestamp 1668089732
transform 1 0 22880 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_8916
timestamp 1668089732
transform 1 0 22880 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_8917
timestamp 1668089732
transform 1 0 22880 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_8918
timestamp 1668089732
transform 1 0 22880 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_8919
timestamp 1668089732
transform 1 0 22880 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_8920
timestamp 1668089732
transform 1 0 22880 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_8921
timestamp 1668089732
transform 1 0 22880 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_8922
timestamp 1668089732
transform 1 0 22880 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_8923
timestamp 1668089732
transform 1 0 22880 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_8924
timestamp 1668089732
transform 1 0 22880 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_8925
timestamp 1668089732
transform 1 0 22880 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_8926
timestamp 1668089732
transform 1 0 22880 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_8927
timestamp 1668089732
transform 1 0 22880 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_8928
timestamp 1668089732
transform 1 0 23040 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_8929
timestamp 1668089732
transform 1 0 23040 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_8930
timestamp 1668089732
transform 1 0 23040 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_8931
timestamp 1668089732
transform 1 0 23040 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_8932
timestamp 1668089732
transform 1 0 23040 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_8933
timestamp 1668089732
transform 1 0 23040 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_8934
timestamp 1668089732
transform 1 0 23040 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_8935
timestamp 1668089732
transform 1 0 23040 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_8936
timestamp 1668089732
transform 1 0 23040 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_8937
timestamp 1668089732
transform 1 0 23040 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_8938
timestamp 1668089732
transform 1 0 23040 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_8939
timestamp 1668089732
transform 1 0 23040 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_8940
timestamp 1668089732
transform 1 0 23040 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_8941
timestamp 1668089732
transform 1 0 23040 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_8942
timestamp 1668089732
transform 1 0 23040 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_8943
timestamp 1668089732
transform 1 0 23040 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_8944
timestamp 1668089732
transform 1 0 23040 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_8945
timestamp 1668089732
transform 1 0 23040 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_8946
timestamp 1668089732
transform 1 0 23040 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_8947
timestamp 1668089732
transform 1 0 23040 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_8948
timestamp 1668089732
transform 1 0 23040 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_8949
timestamp 1668089732
transform 1 0 23040 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_8950
timestamp 1668089732
transform 1 0 23040 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_8951
timestamp 1668089732
transform 1 0 23040 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_8952
timestamp 1668089732
transform 1 0 23040 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_8953
timestamp 1668089732
transform 1 0 23040 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_8954
timestamp 1668089732
transform 1 0 23040 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_8955
timestamp 1668089732
transform 1 0 23040 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_8956
timestamp 1668089732
transform 1 0 23040 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_8957
timestamp 1668089732
transform 1 0 23040 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_8958
timestamp 1668089732
transform 1 0 23040 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_8959
timestamp 1668089732
transform 1 0 23040 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_8960
timestamp 1668089732
transform 1 0 23040 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_8961
timestamp 1668089732
transform 1 0 23040 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_8962
timestamp 1668089732
transform 1 0 23040 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_8963
timestamp 1668089732
transform 1 0 23040 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_8964
timestamp 1668089732
transform 1 0 23040 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_8965
timestamp 1668089732
transform 1 0 23040 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_8966
timestamp 1668089732
transform 1 0 23040 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_8967
timestamp 1668089732
transform 1 0 23040 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_8968
timestamp 1668089732
transform 1 0 23040 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_8969
timestamp 1668089732
transform 1 0 23040 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_8970
timestamp 1668089732
transform 1 0 23040 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_8971
timestamp 1668089732
transform 1 0 23040 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_8972
timestamp 1668089732
transform 1 0 23040 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_8973
timestamp 1668089732
transform 1 0 23040 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_8974
timestamp 1668089732
transform 1 0 23040 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_8975
timestamp 1668089732
transform 1 0 23040 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_8976
timestamp 1668089732
transform 1 0 23040 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_8977
timestamp 1668089732
transform 1 0 23040 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_8978
timestamp 1668089732
transform 1 0 23040 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_8979
timestamp 1668089732
transform 1 0 23040 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_8980
timestamp 1668089732
transform 1 0 23040 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_8981
timestamp 1668089732
transform 1 0 23040 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_8982
timestamp 1668089732
transform 1 0 23040 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_8983
timestamp 1668089732
transform 1 0 23040 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_8984
timestamp 1668089732
transform 1 0 23040 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_8985
timestamp 1668089732
transform 1 0 23040 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_8986
timestamp 1668089732
transform 1 0 23040 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_8987
timestamp 1668089732
transform 1 0 23040 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_8988
timestamp 1668089732
transform 1 0 23040 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_8989
timestamp 1668089732
transform 1 0 23040 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_8990
timestamp 1668089732
transform 1 0 23200 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_8991
timestamp 1668089732
transform 1 0 23200 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_8992
timestamp 1668089732
transform 1 0 23200 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_8993
timestamp 1668089732
transform 1 0 23200 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_8994
timestamp 1668089732
transform 1 0 23200 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_8995
timestamp 1668089732
transform 1 0 23200 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_8996
timestamp 1668089732
transform 1 0 23200 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_8997
timestamp 1668089732
transform 1 0 23200 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_8998
timestamp 1668089732
transform 1 0 23200 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_8999
timestamp 1668089732
transform 1 0 23200 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_9000
timestamp 1668089732
transform 1 0 23200 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_9001
timestamp 1668089732
transform 1 0 23200 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_9002
timestamp 1668089732
transform 1 0 23200 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_9003
timestamp 1668089732
transform 1 0 23200 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_9004
timestamp 1668089732
transform 1 0 23200 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_9005
timestamp 1668089732
transform 1 0 23200 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_9006
timestamp 1668089732
transform 1 0 23200 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_9007
timestamp 1668089732
transform 1 0 23200 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_9008
timestamp 1668089732
transform 1 0 23200 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_9009
timestamp 1668089732
transform 1 0 23200 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_9010
timestamp 1668089732
transform 1 0 23200 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_9011
timestamp 1668089732
transform 1 0 23200 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_9012
timestamp 1668089732
transform 1 0 23200 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_9013
timestamp 1668089732
transform 1 0 23200 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_9014
timestamp 1668089732
transform 1 0 23200 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_9015
timestamp 1668089732
transform 1 0 23200 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_9016
timestamp 1668089732
transform 1 0 23200 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_9017
timestamp 1668089732
transform 1 0 23200 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_9018
timestamp 1668089732
transform 1 0 23200 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_9019
timestamp 1668089732
transform 1 0 23200 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_9020
timestamp 1668089732
transform 1 0 23200 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_9021
timestamp 1668089732
transform 1 0 23200 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_9022
timestamp 1668089732
transform 1 0 23200 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_9023
timestamp 1668089732
transform 1 0 23200 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_9024
timestamp 1668089732
transform 1 0 23200 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_9025
timestamp 1668089732
transform 1 0 23200 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_9026
timestamp 1668089732
transform 1 0 23200 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_9027
timestamp 1668089732
transform 1 0 23200 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_9028
timestamp 1668089732
transform 1 0 23200 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_9029
timestamp 1668089732
transform 1 0 23200 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_9030
timestamp 1668089732
transform 1 0 23200 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_9031
timestamp 1668089732
transform 1 0 23200 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_9032
timestamp 1668089732
transform 1 0 23200 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_9033
timestamp 1668089732
transform 1 0 23200 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_9034
timestamp 1668089732
transform 1 0 23200 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_9035
timestamp 1668089732
transform 1 0 23200 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_9036
timestamp 1668089732
transform 1 0 23200 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_9037
timestamp 1668089732
transform 1 0 23200 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_9038
timestamp 1668089732
transform 1 0 23200 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_9039
timestamp 1668089732
transform 1 0 23200 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_9040
timestamp 1668089732
transform 1 0 23200 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_9041
timestamp 1668089732
transform 1 0 23200 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_9042
timestamp 1668089732
transform 1 0 23200 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_9043
timestamp 1668089732
transform 1 0 23200 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_9044
timestamp 1668089732
transform 1 0 23200 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_9045
timestamp 1668089732
transform 1 0 23200 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_9046
timestamp 1668089732
transform 1 0 23200 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_9047
timestamp 1668089732
transform 1 0 23200 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_9048
timestamp 1668089732
transform 1 0 23200 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_9049
timestamp 1668089732
transform 1 0 23200 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_9050
timestamp 1668089732
transform 1 0 23200 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_9051
timestamp 1668089732
transform 1 0 23200 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_9052
timestamp 1668089732
transform 1 0 23360 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_9053
timestamp 1668089732
transform 1 0 23360 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_9054
timestamp 1668089732
transform 1 0 23360 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_9055
timestamp 1668089732
transform 1 0 23360 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_9056
timestamp 1668089732
transform 1 0 23360 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_9057
timestamp 1668089732
transform 1 0 23360 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_9058
timestamp 1668089732
transform 1 0 23360 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_9059
timestamp 1668089732
transform 1 0 23360 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_9060
timestamp 1668089732
transform 1 0 23360 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_9061
timestamp 1668089732
transform 1 0 23360 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_9062
timestamp 1668089732
transform 1 0 23360 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_9063
timestamp 1668089732
transform 1 0 23360 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_9064
timestamp 1668089732
transform 1 0 23360 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_9065
timestamp 1668089732
transform 1 0 23360 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_9066
timestamp 1668089732
transform 1 0 23360 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_9067
timestamp 1668089732
transform 1 0 23360 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_9068
timestamp 1668089732
transform 1 0 23360 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_9069
timestamp 1668089732
transform 1 0 23360 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_9070
timestamp 1668089732
transform 1 0 23360 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_9071
timestamp 1668089732
transform 1 0 23360 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_9072
timestamp 1668089732
transform 1 0 23360 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_9073
timestamp 1668089732
transform 1 0 23360 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_9074
timestamp 1668089732
transform 1 0 23360 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_9075
timestamp 1668089732
transform 1 0 23360 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_9076
timestamp 1668089732
transform 1 0 23360 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_9077
timestamp 1668089732
transform 1 0 23360 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_9078
timestamp 1668089732
transform 1 0 23360 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_9079
timestamp 1668089732
transform 1 0 23360 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_9080
timestamp 1668089732
transform 1 0 23360 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_9081
timestamp 1668089732
transform 1 0 23360 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_9082
timestamp 1668089732
transform 1 0 23360 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_9083
timestamp 1668089732
transform 1 0 23360 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_9084
timestamp 1668089732
transform 1 0 23360 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_9085
timestamp 1668089732
transform 1 0 23360 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_9086
timestamp 1668089732
transform 1 0 23360 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_9087
timestamp 1668089732
transform 1 0 23360 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_9088
timestamp 1668089732
transform 1 0 23360 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_9089
timestamp 1668089732
transform 1 0 23360 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_9090
timestamp 1668089732
transform 1 0 23360 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_9091
timestamp 1668089732
transform 1 0 23360 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_9092
timestamp 1668089732
transform 1 0 23360 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_9093
timestamp 1668089732
transform 1 0 23360 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_9094
timestamp 1668089732
transform 1 0 23360 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_9095
timestamp 1668089732
transform 1 0 23360 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_9096
timestamp 1668089732
transform 1 0 23360 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_9097
timestamp 1668089732
transform 1 0 23360 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_9098
timestamp 1668089732
transform 1 0 23360 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_9099
timestamp 1668089732
transform 1 0 23360 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_9100
timestamp 1668089732
transform 1 0 23360 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_9101
timestamp 1668089732
transform 1 0 23360 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_9102
timestamp 1668089732
transform 1 0 23360 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_9103
timestamp 1668089732
transform 1 0 23360 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_9104
timestamp 1668089732
transform 1 0 23360 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_9105
timestamp 1668089732
transform 1 0 23360 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_9106
timestamp 1668089732
transform 1 0 23360 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_9107
timestamp 1668089732
transform 1 0 23360 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_9108
timestamp 1668089732
transform 1 0 23360 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_9109
timestamp 1668089732
transform 1 0 23360 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_9110
timestamp 1668089732
transform 1 0 23360 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_9111
timestamp 1668089732
transform 1 0 23360 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_9112
timestamp 1668089732
transform 1 0 23360 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_9113
timestamp 1668089732
transform 1 0 23360 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_9114
timestamp 1668089732
transform 1 0 23520 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_9115
timestamp 1668089732
transform 1 0 23520 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_9116
timestamp 1668089732
transform 1 0 23520 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_9117
timestamp 1668089732
transform 1 0 23520 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_9118
timestamp 1668089732
transform 1 0 23520 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_9119
timestamp 1668089732
transform 1 0 23520 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_9120
timestamp 1668089732
transform 1 0 23520 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_9121
timestamp 1668089732
transform 1 0 23520 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_9122
timestamp 1668089732
transform 1 0 23520 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_9123
timestamp 1668089732
transform 1 0 23520 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_9124
timestamp 1668089732
transform 1 0 23520 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_9125
timestamp 1668089732
transform 1 0 23520 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_9126
timestamp 1668089732
transform 1 0 23520 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_9127
timestamp 1668089732
transform 1 0 23520 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_9128
timestamp 1668089732
transform 1 0 23520 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_9129
timestamp 1668089732
transform 1 0 23520 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_9130
timestamp 1668089732
transform 1 0 23520 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_9131
timestamp 1668089732
transform 1 0 23520 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_9132
timestamp 1668089732
transform 1 0 23520 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_9133
timestamp 1668089732
transform 1 0 23520 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_9134
timestamp 1668089732
transform 1 0 23520 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_9135
timestamp 1668089732
transform 1 0 23520 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_9136
timestamp 1668089732
transform 1 0 23520 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_9137
timestamp 1668089732
transform 1 0 23520 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_9138
timestamp 1668089732
transform 1 0 23520 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_9139
timestamp 1668089732
transform 1 0 23520 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_9140
timestamp 1668089732
transform 1 0 23520 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_9141
timestamp 1668089732
transform 1 0 23520 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_9142
timestamp 1668089732
transform 1 0 23520 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_9143
timestamp 1668089732
transform 1 0 23520 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_9144
timestamp 1668089732
transform 1 0 23520 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_9145
timestamp 1668089732
transform 1 0 23520 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_9146
timestamp 1668089732
transform 1 0 23520 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_9147
timestamp 1668089732
transform 1 0 23520 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_9148
timestamp 1668089732
transform 1 0 23520 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_9149
timestamp 1668089732
transform 1 0 23520 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_9150
timestamp 1668089732
transform 1 0 23520 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_9151
timestamp 1668089732
transform 1 0 23520 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_9152
timestamp 1668089732
transform 1 0 23520 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_9153
timestamp 1668089732
transform 1 0 23520 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_9154
timestamp 1668089732
transform 1 0 23520 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_9155
timestamp 1668089732
transform 1 0 23520 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_9156
timestamp 1668089732
transform 1 0 23520 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_9157
timestamp 1668089732
transform 1 0 23520 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_9158
timestamp 1668089732
transform 1 0 23520 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_9159
timestamp 1668089732
transform 1 0 23520 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_9160
timestamp 1668089732
transform 1 0 23520 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_9161
timestamp 1668089732
transform 1 0 23520 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_9162
timestamp 1668089732
transform 1 0 23520 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_9163
timestamp 1668089732
transform 1 0 23520 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_9164
timestamp 1668089732
transform 1 0 23520 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_9165
timestamp 1668089732
transform 1 0 23520 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_9166
timestamp 1668089732
transform 1 0 23520 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_9167
timestamp 1668089732
transform 1 0 23520 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_9168
timestamp 1668089732
transform 1 0 23520 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_9169
timestamp 1668089732
transform 1 0 23520 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_9170
timestamp 1668089732
transform 1 0 23520 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_9171
timestamp 1668089732
transform 1 0 23520 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_9172
timestamp 1668089732
transform 1 0 23520 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_9173
timestamp 1668089732
transform 1 0 23520 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_9174
timestamp 1668089732
transform 1 0 23520 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_9175
timestamp 1668089732
transform 1 0 23520 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_9176
timestamp 1668089732
transform 1 0 23680 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_9177
timestamp 1668089732
transform 1 0 23680 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_9178
timestamp 1668089732
transform 1 0 23680 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_9179
timestamp 1668089732
transform 1 0 23680 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_9180
timestamp 1668089732
transform 1 0 23680 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_9181
timestamp 1668089732
transform 1 0 23680 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_9182
timestamp 1668089732
transform 1 0 23680 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_9183
timestamp 1668089732
transform 1 0 23680 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_9184
timestamp 1668089732
transform 1 0 23680 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_9185
timestamp 1668089732
transform 1 0 23680 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_9186
timestamp 1668089732
transform 1 0 23680 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_9187
timestamp 1668089732
transform 1 0 23680 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_9188
timestamp 1668089732
transform 1 0 23680 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_9189
timestamp 1668089732
transform 1 0 23680 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_9190
timestamp 1668089732
transform 1 0 23680 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_9191
timestamp 1668089732
transform 1 0 23680 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_9192
timestamp 1668089732
transform 1 0 23680 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_9193
timestamp 1668089732
transform 1 0 23680 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_9194
timestamp 1668089732
transform 1 0 23680 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_9195
timestamp 1668089732
transform 1 0 23680 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_9196
timestamp 1668089732
transform 1 0 23680 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_9197
timestamp 1668089732
transform 1 0 23680 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_9198
timestamp 1668089732
transform 1 0 23680 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_9199
timestamp 1668089732
transform 1 0 23680 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_9200
timestamp 1668089732
transform 1 0 23680 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_9201
timestamp 1668089732
transform 1 0 23680 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_9202
timestamp 1668089732
transform 1 0 23680 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_9203
timestamp 1668089732
transform 1 0 23680 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_9204
timestamp 1668089732
transform 1 0 23680 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_9205
timestamp 1668089732
transform 1 0 23680 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_9206
timestamp 1668089732
transform 1 0 23680 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_9207
timestamp 1668089732
transform 1 0 23680 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_9208
timestamp 1668089732
transform 1 0 23680 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_9209
timestamp 1668089732
transform 1 0 23680 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_9210
timestamp 1668089732
transform 1 0 23680 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_9211
timestamp 1668089732
transform 1 0 23680 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_9212
timestamp 1668089732
transform 1 0 23680 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_9213
timestamp 1668089732
transform 1 0 23680 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_9214
timestamp 1668089732
transform 1 0 23680 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_9215
timestamp 1668089732
transform 1 0 23680 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_9216
timestamp 1668089732
transform 1 0 23680 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_9217
timestamp 1668089732
transform 1 0 23680 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_9218
timestamp 1668089732
transform 1 0 23680 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_9219
timestamp 1668089732
transform 1 0 23680 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_9220
timestamp 1668089732
transform 1 0 23680 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_9221
timestamp 1668089732
transform 1 0 23680 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_9222
timestamp 1668089732
transform 1 0 23680 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_9223
timestamp 1668089732
transform 1 0 23680 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_9224
timestamp 1668089732
transform 1 0 23680 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_9225
timestamp 1668089732
transform 1 0 23680 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_9226
timestamp 1668089732
transform 1 0 23680 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_9227
timestamp 1668089732
transform 1 0 23680 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_9228
timestamp 1668089732
transform 1 0 23680 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_9229
timestamp 1668089732
transform 1 0 23680 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_9230
timestamp 1668089732
transform 1 0 23680 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_9231
timestamp 1668089732
transform 1 0 23680 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_9232
timestamp 1668089732
transform 1 0 23680 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_9233
timestamp 1668089732
transform 1 0 23680 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_9234
timestamp 1668089732
transform 1 0 23680 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_9235
timestamp 1668089732
transform 1 0 23680 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_9236
timestamp 1668089732
transform 1 0 23680 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_9237
timestamp 1668089732
transform 1 0 23680 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_9238
timestamp 1668089732
transform 1 0 23840 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_9239
timestamp 1668089732
transform 1 0 23840 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_9240
timestamp 1668089732
transform 1 0 23840 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_9241
timestamp 1668089732
transform 1 0 23840 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_9242
timestamp 1668089732
transform 1 0 23840 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_9243
timestamp 1668089732
transform 1 0 23840 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_9244
timestamp 1668089732
transform 1 0 23840 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_9245
timestamp 1668089732
transform 1 0 23840 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_9246
timestamp 1668089732
transform 1 0 23840 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_9247
timestamp 1668089732
transform 1 0 23840 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_9248
timestamp 1668089732
transform 1 0 23840 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_9249
timestamp 1668089732
transform 1 0 23840 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_9250
timestamp 1668089732
transform 1 0 23840 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_9251
timestamp 1668089732
transform 1 0 23840 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_9252
timestamp 1668089732
transform 1 0 23840 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_9253
timestamp 1668089732
transform 1 0 23840 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_9254
timestamp 1668089732
transform 1 0 23840 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_9255
timestamp 1668089732
transform 1 0 23840 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_9256
timestamp 1668089732
transform 1 0 23840 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_9257
timestamp 1668089732
transform 1 0 23840 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_9258
timestamp 1668089732
transform 1 0 23840 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_9259
timestamp 1668089732
transform 1 0 23840 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_9260
timestamp 1668089732
transform 1 0 23840 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_9261
timestamp 1668089732
transform 1 0 23840 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_9262
timestamp 1668089732
transform 1 0 23840 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_9263
timestamp 1668089732
transform 1 0 23840 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_9264
timestamp 1668089732
transform 1 0 23840 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_9265
timestamp 1668089732
transform 1 0 23840 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_9266
timestamp 1668089732
transform 1 0 23840 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_9267
timestamp 1668089732
transform 1 0 23840 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_9268
timestamp 1668089732
transform 1 0 23840 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_9269
timestamp 1668089732
transform 1 0 23840 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_9270
timestamp 1668089732
transform 1 0 23840 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_9271
timestamp 1668089732
transform 1 0 23840 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_9272
timestamp 1668089732
transform 1 0 23840 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_9273
timestamp 1668089732
transform 1 0 23840 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_9274
timestamp 1668089732
transform 1 0 23840 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_9275
timestamp 1668089732
transform 1 0 23840 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_9276
timestamp 1668089732
transform 1 0 23840 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_9277
timestamp 1668089732
transform 1 0 23840 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_9278
timestamp 1668089732
transform 1 0 23840 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_9279
timestamp 1668089732
transform 1 0 23840 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_9280
timestamp 1668089732
transform 1 0 23840 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_9281
timestamp 1668089732
transform 1 0 23840 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_9282
timestamp 1668089732
transform 1 0 23840 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_9283
timestamp 1668089732
transform 1 0 23840 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_9284
timestamp 1668089732
transform 1 0 23840 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_9285
timestamp 1668089732
transform 1 0 23840 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_9286
timestamp 1668089732
transform 1 0 23840 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_9287
timestamp 1668089732
transform 1 0 23840 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_9288
timestamp 1668089732
transform 1 0 23840 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_9289
timestamp 1668089732
transform 1 0 23840 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_9290
timestamp 1668089732
transform 1 0 23840 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_9291
timestamp 1668089732
transform 1 0 23840 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_9292
timestamp 1668089732
transform 1 0 23840 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_9293
timestamp 1668089732
transform 1 0 23840 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_9294
timestamp 1668089732
transform 1 0 23840 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_9295
timestamp 1668089732
transform 1 0 23840 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_9296
timestamp 1668089732
transform 1 0 23840 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_9297
timestamp 1668089732
transform 1 0 23840 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_9298
timestamp 1668089732
transform 1 0 23840 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_9299
timestamp 1668089732
transform 1 0 23840 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_9300
timestamp 1668089732
transform 1 0 24000 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_9301
timestamp 1668089732
transform 1 0 24000 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_9302
timestamp 1668089732
transform 1 0 24000 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_9303
timestamp 1668089732
transform 1 0 24000 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_9304
timestamp 1668089732
transform 1 0 24000 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_9305
timestamp 1668089732
transform 1 0 24000 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_9306
timestamp 1668089732
transform 1 0 24000 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_9307
timestamp 1668089732
transform 1 0 24000 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_9308
timestamp 1668089732
transform 1 0 24000 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_9309
timestamp 1668089732
transform 1 0 24000 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_9310
timestamp 1668089732
transform 1 0 24000 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_9311
timestamp 1668089732
transform 1 0 24000 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_9312
timestamp 1668089732
transform 1 0 24000 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_9313
timestamp 1668089732
transform 1 0 24000 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_9314
timestamp 1668089732
transform 1 0 24000 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_9315
timestamp 1668089732
transform 1 0 24000 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_9316
timestamp 1668089732
transform 1 0 24000 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_9317
timestamp 1668089732
transform 1 0 24000 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_9318
timestamp 1668089732
transform 1 0 24000 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_9319
timestamp 1668089732
transform 1 0 24000 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_9320
timestamp 1668089732
transform 1 0 24000 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_9321
timestamp 1668089732
transform 1 0 24000 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_9322
timestamp 1668089732
transform 1 0 24000 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_9323
timestamp 1668089732
transform 1 0 24000 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_9324
timestamp 1668089732
transform 1 0 24000 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_9325
timestamp 1668089732
transform 1 0 24000 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_9326
timestamp 1668089732
transform 1 0 24000 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_9327
timestamp 1668089732
transform 1 0 24000 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_9328
timestamp 1668089732
transform 1 0 24000 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_9329
timestamp 1668089732
transform 1 0 24000 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_9330
timestamp 1668089732
transform 1 0 24000 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_9331
timestamp 1668089732
transform 1 0 24000 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_9332
timestamp 1668089732
transform 1 0 24000 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_9333
timestamp 1668089732
transform 1 0 24000 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_9334
timestamp 1668089732
transform 1 0 24000 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_9335
timestamp 1668089732
transform 1 0 24000 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_9336
timestamp 1668089732
transform 1 0 24000 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_9337
timestamp 1668089732
transform 1 0 24000 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_9338
timestamp 1668089732
transform 1 0 24000 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_9339
timestamp 1668089732
transform 1 0 24000 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_9340
timestamp 1668089732
transform 1 0 24000 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_9341
timestamp 1668089732
transform 1 0 24000 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_9342
timestamp 1668089732
transform 1 0 24000 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_9343
timestamp 1668089732
transform 1 0 24000 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_9344
timestamp 1668089732
transform 1 0 24000 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_9345
timestamp 1668089732
transform 1 0 24000 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_9346
timestamp 1668089732
transform 1 0 24000 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_9347
timestamp 1668089732
transform 1 0 24000 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_9348
timestamp 1668089732
transform 1 0 24000 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_9349
timestamp 1668089732
transform 1 0 24000 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_9350
timestamp 1668089732
transform 1 0 24000 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_9351
timestamp 1668089732
transform 1 0 24000 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_9352
timestamp 1668089732
transform 1 0 24000 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_9353
timestamp 1668089732
transform 1 0 24000 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_9354
timestamp 1668089732
transform 1 0 24000 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_9355
timestamp 1668089732
transform 1 0 24000 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_9356
timestamp 1668089732
transform 1 0 24000 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_9357
timestamp 1668089732
transform 1 0 24000 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_9358
timestamp 1668089732
transform 1 0 24000 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_9359
timestamp 1668089732
transform 1 0 24000 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_9360
timestamp 1668089732
transform 1 0 24000 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_9361
timestamp 1668089732
transform 1 0 24000 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_9362
timestamp 1668089732
transform 1 0 24160 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_9363
timestamp 1668089732
transform 1 0 24160 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_9364
timestamp 1668089732
transform 1 0 24160 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_9365
timestamp 1668089732
transform 1 0 24160 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_9366
timestamp 1668089732
transform 1 0 24160 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_9367
timestamp 1668089732
transform 1 0 24160 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_9368
timestamp 1668089732
transform 1 0 24160 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_9369
timestamp 1668089732
transform 1 0 24160 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_9370
timestamp 1668089732
transform 1 0 24160 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_9371
timestamp 1668089732
transform 1 0 24160 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_9372
timestamp 1668089732
transform 1 0 24160 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_9373
timestamp 1668089732
transform 1 0 24160 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_9374
timestamp 1668089732
transform 1 0 24160 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_9375
timestamp 1668089732
transform 1 0 24160 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_9376
timestamp 1668089732
transform 1 0 24160 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_9377
timestamp 1668089732
transform 1 0 24160 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_9378
timestamp 1668089732
transform 1 0 24160 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_9379
timestamp 1668089732
transform 1 0 24160 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_9380
timestamp 1668089732
transform 1 0 24160 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_9381
timestamp 1668089732
transform 1 0 24160 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_9382
timestamp 1668089732
transform 1 0 24160 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_9383
timestamp 1668089732
transform 1 0 24160 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_9384
timestamp 1668089732
transform 1 0 24160 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_9385
timestamp 1668089732
transform 1 0 24160 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_9386
timestamp 1668089732
transform 1 0 24160 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_9387
timestamp 1668089732
transform 1 0 24160 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_9388
timestamp 1668089732
transform 1 0 24160 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_9389
timestamp 1668089732
transform 1 0 24160 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_9390
timestamp 1668089732
transform 1 0 24160 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_9391
timestamp 1668089732
transform 1 0 24160 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_9392
timestamp 1668089732
transform 1 0 24160 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_9393
timestamp 1668089732
transform 1 0 24160 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_9394
timestamp 1668089732
transform 1 0 24160 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_9395
timestamp 1668089732
transform 1 0 24160 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_9396
timestamp 1668089732
transform 1 0 24160 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_9397
timestamp 1668089732
transform 1 0 24160 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_9398
timestamp 1668089732
transform 1 0 24160 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_9399
timestamp 1668089732
transform 1 0 24160 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_9400
timestamp 1668089732
transform 1 0 24160 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_9401
timestamp 1668089732
transform 1 0 24160 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_9402
timestamp 1668089732
transform 1 0 24160 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_9403
timestamp 1668089732
transform 1 0 24160 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_9404
timestamp 1668089732
transform 1 0 24160 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_9405
timestamp 1668089732
transform 1 0 24160 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_9406
timestamp 1668089732
transform 1 0 24160 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_9407
timestamp 1668089732
transform 1 0 24160 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_9408
timestamp 1668089732
transform 1 0 24160 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_9409
timestamp 1668089732
transform 1 0 24160 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_9410
timestamp 1668089732
transform 1 0 24160 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_9411
timestamp 1668089732
transform 1 0 24160 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_9412
timestamp 1668089732
transform 1 0 24160 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_9413
timestamp 1668089732
transform 1 0 24160 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_9414
timestamp 1668089732
transform 1 0 24160 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_9415
timestamp 1668089732
transform 1 0 24160 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_9416
timestamp 1668089732
transform 1 0 24160 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_9417
timestamp 1668089732
transform 1 0 24160 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_9418
timestamp 1668089732
transform 1 0 24160 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_9419
timestamp 1668089732
transform 1 0 24160 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_9420
timestamp 1668089732
transform 1 0 24160 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_9421
timestamp 1668089732
transform 1 0 24160 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_9422
timestamp 1668089732
transform 1 0 24160 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_9423
timestamp 1668089732
transform 1 0 24160 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_9424
timestamp 1668089732
transform 1 0 24320 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_9425
timestamp 1668089732
transform 1 0 24320 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_9426
timestamp 1668089732
transform 1 0 24320 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_9427
timestamp 1668089732
transform 1 0 24320 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_9428
timestamp 1668089732
transform 1 0 24320 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_9429
timestamp 1668089732
transform 1 0 24320 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_9430
timestamp 1668089732
transform 1 0 24320 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_9431
timestamp 1668089732
transform 1 0 24320 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_9432
timestamp 1668089732
transform 1 0 24320 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_9433
timestamp 1668089732
transform 1 0 24320 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_9434
timestamp 1668089732
transform 1 0 24320 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_9435
timestamp 1668089732
transform 1 0 24320 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_9436
timestamp 1668089732
transform 1 0 24320 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_9437
timestamp 1668089732
transform 1 0 24320 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_9438
timestamp 1668089732
transform 1 0 24320 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_9439
timestamp 1668089732
transform 1 0 24320 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_9440
timestamp 1668089732
transform 1 0 24320 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_9441
timestamp 1668089732
transform 1 0 24320 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_9442
timestamp 1668089732
transform 1 0 24320 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_9443
timestamp 1668089732
transform 1 0 24320 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_9444
timestamp 1668089732
transform 1 0 24320 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_9445
timestamp 1668089732
transform 1 0 24320 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_9446
timestamp 1668089732
transform 1 0 24320 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_9447
timestamp 1668089732
transform 1 0 24320 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_9448
timestamp 1668089732
transform 1 0 24320 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_9449
timestamp 1668089732
transform 1 0 24320 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_9450
timestamp 1668089732
transform 1 0 24320 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_9451
timestamp 1668089732
transform 1 0 24320 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_9452
timestamp 1668089732
transform 1 0 24320 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_9453
timestamp 1668089732
transform 1 0 24320 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_9454
timestamp 1668089732
transform 1 0 24320 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_9455
timestamp 1668089732
transform 1 0 24320 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_9456
timestamp 1668089732
transform 1 0 24320 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_9457
timestamp 1668089732
transform 1 0 24320 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_9458
timestamp 1668089732
transform 1 0 24320 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_9459
timestamp 1668089732
transform 1 0 24320 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_9460
timestamp 1668089732
transform 1 0 24320 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_9461
timestamp 1668089732
transform 1 0 24320 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_9462
timestamp 1668089732
transform 1 0 24320 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_9463
timestamp 1668089732
transform 1 0 24320 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_9464
timestamp 1668089732
transform 1 0 24320 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_9465
timestamp 1668089732
transform 1 0 24320 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_9466
timestamp 1668089732
transform 1 0 24320 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_9467
timestamp 1668089732
transform 1 0 24320 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_9468
timestamp 1668089732
transform 1 0 24320 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_9469
timestamp 1668089732
transform 1 0 24320 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_9470
timestamp 1668089732
transform 1 0 24320 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_9471
timestamp 1668089732
transform 1 0 24320 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_9472
timestamp 1668089732
transform 1 0 24320 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_9473
timestamp 1668089732
transform 1 0 24320 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_9474
timestamp 1668089732
transform 1 0 24320 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_9475
timestamp 1668089732
transform 1 0 24320 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_9476
timestamp 1668089732
transform 1 0 24320 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_9477
timestamp 1668089732
transform 1 0 24320 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_9478
timestamp 1668089732
transform 1 0 24320 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_9479
timestamp 1668089732
transform 1 0 24320 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_9480
timestamp 1668089732
transform 1 0 24320 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_9481
timestamp 1668089732
transform 1 0 24320 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_9482
timestamp 1668089732
transform 1 0 24320 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_9483
timestamp 1668089732
transform 1 0 24320 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_9484
timestamp 1668089732
transform 1 0 24320 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_9485
timestamp 1668089732
transform 1 0 24320 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_9486
timestamp 1668089732
transform 1 0 24480 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_9487
timestamp 1668089732
transform 1 0 24480 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_9488
timestamp 1668089732
transform 1 0 24480 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_9489
timestamp 1668089732
transform 1 0 24480 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_9490
timestamp 1668089732
transform 1 0 24480 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_9491
timestamp 1668089732
transform 1 0 24480 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_9492
timestamp 1668089732
transform 1 0 24480 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_9493
timestamp 1668089732
transform 1 0 24480 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_9494
timestamp 1668089732
transform 1 0 24480 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_9495
timestamp 1668089732
transform 1 0 24480 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_9496
timestamp 1668089732
transform 1 0 24480 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_9497
timestamp 1668089732
transform 1 0 24480 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_9498
timestamp 1668089732
transform 1 0 24480 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_9499
timestamp 1668089732
transform 1 0 24480 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_9500
timestamp 1668089732
transform 1 0 24480 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_9501
timestamp 1668089732
transform 1 0 24480 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_9502
timestamp 1668089732
transform 1 0 24480 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_9503
timestamp 1668089732
transform 1 0 24480 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_9504
timestamp 1668089732
transform 1 0 24480 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_9505
timestamp 1668089732
transform 1 0 24480 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_9506
timestamp 1668089732
transform 1 0 24480 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_9507
timestamp 1668089732
transform 1 0 24480 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_9508
timestamp 1668089732
transform 1 0 24480 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_9509
timestamp 1668089732
transform 1 0 24480 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_9510
timestamp 1668089732
transform 1 0 24480 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_9511
timestamp 1668089732
transform 1 0 24480 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_9512
timestamp 1668089732
transform 1 0 24480 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_9513
timestamp 1668089732
transform 1 0 24480 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_9514
timestamp 1668089732
transform 1 0 24480 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_9515
timestamp 1668089732
transform 1 0 24480 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_9516
timestamp 1668089732
transform 1 0 24480 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_9517
timestamp 1668089732
transform 1 0 24480 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_9518
timestamp 1668089732
transform 1 0 24480 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_9519
timestamp 1668089732
transform 1 0 24480 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_9520
timestamp 1668089732
transform 1 0 24480 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_9521
timestamp 1668089732
transform 1 0 24480 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_9522
timestamp 1668089732
transform 1 0 24480 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_9523
timestamp 1668089732
transform 1 0 24480 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_9524
timestamp 1668089732
transform 1 0 24480 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_9525
timestamp 1668089732
transform 1 0 24480 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_9526
timestamp 1668089732
transform 1 0 24480 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_9527
timestamp 1668089732
transform 1 0 24480 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_9528
timestamp 1668089732
transform 1 0 24480 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_9529
timestamp 1668089732
transform 1 0 24480 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_9530
timestamp 1668089732
transform 1 0 24480 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_9531
timestamp 1668089732
transform 1 0 24480 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_9532
timestamp 1668089732
transform 1 0 24480 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_9533
timestamp 1668089732
transform 1 0 24480 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_9534
timestamp 1668089732
transform 1 0 24480 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_9535
timestamp 1668089732
transform 1 0 24480 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_9536
timestamp 1668089732
transform 1 0 24480 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_9537
timestamp 1668089732
transform 1 0 24480 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_9538
timestamp 1668089732
transform 1 0 24480 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_9539
timestamp 1668089732
transform 1 0 24480 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_9540
timestamp 1668089732
transform 1 0 24480 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_9541
timestamp 1668089732
transform 1 0 24480 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_9542
timestamp 1668089732
transform 1 0 24480 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_9543
timestamp 1668089732
transform 1 0 24480 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_9544
timestamp 1668089732
transform 1 0 24480 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_9545
timestamp 1668089732
transform 1 0 24480 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_9546
timestamp 1668089732
transform 1 0 24480 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_9547
timestamp 1668089732
transform 1 0 24480 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_9548
timestamp 1668089732
transform 1 0 24640 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_9549
timestamp 1668089732
transform 1 0 24640 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_9550
timestamp 1668089732
transform 1 0 24640 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_9551
timestamp 1668089732
transform 1 0 24640 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_9552
timestamp 1668089732
transform 1 0 24640 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_9553
timestamp 1668089732
transform 1 0 24640 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_9554
timestamp 1668089732
transform 1 0 24640 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_9555
timestamp 1668089732
transform 1 0 24640 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_9556
timestamp 1668089732
transform 1 0 24640 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_9557
timestamp 1668089732
transform 1 0 24640 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_9558
timestamp 1668089732
transform 1 0 24640 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_9559
timestamp 1668089732
transform 1 0 24640 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_9560
timestamp 1668089732
transform 1 0 24640 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_9561
timestamp 1668089732
transform 1 0 24640 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_9562
timestamp 1668089732
transform 1 0 24640 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_9563
timestamp 1668089732
transform 1 0 24640 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_9564
timestamp 1668089732
transform 1 0 24640 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_9565
timestamp 1668089732
transform 1 0 24640 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_9566
timestamp 1668089732
transform 1 0 24640 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_9567
timestamp 1668089732
transform 1 0 24640 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_9568
timestamp 1668089732
transform 1 0 24640 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_9569
timestamp 1668089732
transform 1 0 24640 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_9570
timestamp 1668089732
transform 1 0 24640 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_9571
timestamp 1668089732
transform 1 0 24640 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_9572
timestamp 1668089732
transform 1 0 24640 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_9573
timestamp 1668089732
transform 1 0 24640 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_9574
timestamp 1668089732
transform 1 0 24640 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_9575
timestamp 1668089732
transform 1 0 24640 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_9576
timestamp 1668089732
transform 1 0 24640 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_9577
timestamp 1668089732
transform 1 0 24640 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_9578
timestamp 1668089732
transform 1 0 24640 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_9579
timestamp 1668089732
transform 1 0 24640 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_9580
timestamp 1668089732
transform 1 0 24640 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_9581
timestamp 1668089732
transform 1 0 24640 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_9582
timestamp 1668089732
transform 1 0 24640 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_9583
timestamp 1668089732
transform 1 0 24640 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_9584
timestamp 1668089732
transform 1 0 24640 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_9585
timestamp 1668089732
transform 1 0 24640 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_9586
timestamp 1668089732
transform 1 0 24640 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_9587
timestamp 1668089732
transform 1 0 24640 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_9588
timestamp 1668089732
transform 1 0 24640 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_9589
timestamp 1668089732
transform 1 0 24640 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_9590
timestamp 1668089732
transform 1 0 24640 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_9591
timestamp 1668089732
transform 1 0 24640 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_9592
timestamp 1668089732
transform 1 0 24640 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_9593
timestamp 1668089732
transform 1 0 24640 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_9594
timestamp 1668089732
transform 1 0 24640 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_9595
timestamp 1668089732
transform 1 0 24640 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_9596
timestamp 1668089732
transform 1 0 24640 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_9597
timestamp 1668089732
transform 1 0 24640 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_9598
timestamp 1668089732
transform 1 0 24640 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_9599
timestamp 1668089732
transform 1 0 24640 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_9600
timestamp 1668089732
transform 1 0 24640 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_9601
timestamp 1668089732
transform 1 0 24640 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_9602
timestamp 1668089732
transform 1 0 24640 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_9603
timestamp 1668089732
transform 1 0 24640 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_9604
timestamp 1668089732
transform 1 0 24640 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_9605
timestamp 1668089732
transform 1 0 24640 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_9606
timestamp 1668089732
transform 1 0 24640 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_9607
timestamp 1668089732
transform 1 0 24640 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_9608
timestamp 1668089732
transform 1 0 24640 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_9609
timestamp 1668089732
transform 1 0 24640 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_9610
timestamp 1668089732
transform 1 0 24800 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_9611
timestamp 1668089732
transform 1 0 24800 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_9612
timestamp 1668089732
transform 1 0 24800 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_9613
timestamp 1668089732
transform 1 0 24800 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_9614
timestamp 1668089732
transform 1 0 24800 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_9615
timestamp 1668089732
transform 1 0 24800 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_9616
timestamp 1668089732
transform 1 0 24800 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_9617
timestamp 1668089732
transform 1 0 24800 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_9618
timestamp 1668089732
transform 1 0 24800 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_9619
timestamp 1668089732
transform 1 0 24800 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_9620
timestamp 1668089732
transform 1 0 24800 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_9621
timestamp 1668089732
transform 1 0 24800 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_9622
timestamp 1668089732
transform 1 0 24800 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_9623
timestamp 1668089732
transform 1 0 24800 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_9624
timestamp 1668089732
transform 1 0 24800 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_9625
timestamp 1668089732
transform 1 0 24800 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_9626
timestamp 1668089732
transform 1 0 24800 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_9627
timestamp 1668089732
transform 1 0 24800 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_9628
timestamp 1668089732
transform 1 0 24800 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_9629
timestamp 1668089732
transform 1 0 24800 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_9630
timestamp 1668089732
transform 1 0 24800 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_9631
timestamp 1668089732
transform 1 0 24800 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_9632
timestamp 1668089732
transform 1 0 24800 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_9633
timestamp 1668089732
transform 1 0 24800 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_9634
timestamp 1668089732
transform 1 0 24800 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_9635
timestamp 1668089732
transform 1 0 24800 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_9636
timestamp 1668089732
transform 1 0 24800 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_9637
timestamp 1668089732
transform 1 0 24800 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_9638
timestamp 1668089732
transform 1 0 24800 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_9639
timestamp 1668089732
transform 1 0 24800 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_9640
timestamp 1668089732
transform 1 0 24800 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_9641
timestamp 1668089732
transform 1 0 24800 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_9642
timestamp 1668089732
transform 1 0 24800 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_9643
timestamp 1668089732
transform 1 0 24800 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_9644
timestamp 1668089732
transform 1 0 24800 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_9645
timestamp 1668089732
transform 1 0 24800 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_9646
timestamp 1668089732
transform 1 0 24800 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_9647
timestamp 1668089732
transform 1 0 24800 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_9648
timestamp 1668089732
transform 1 0 24800 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_9649
timestamp 1668089732
transform 1 0 24800 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_9650
timestamp 1668089732
transform 1 0 24800 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_9651
timestamp 1668089732
transform 1 0 24800 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_9652
timestamp 1668089732
transform 1 0 24800 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_9653
timestamp 1668089732
transform 1 0 24800 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_9654
timestamp 1668089732
transform 1 0 24800 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_9655
timestamp 1668089732
transform 1 0 24800 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_9656
timestamp 1668089732
transform 1 0 24800 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_9657
timestamp 1668089732
transform 1 0 24800 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_9658
timestamp 1668089732
transform 1 0 24800 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_9659
timestamp 1668089732
transform 1 0 24800 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_9660
timestamp 1668089732
transform 1 0 24800 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_9661
timestamp 1668089732
transform 1 0 24800 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_9662
timestamp 1668089732
transform 1 0 24800 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_9663
timestamp 1668089732
transform 1 0 24800 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_9664
timestamp 1668089732
transform 1 0 24800 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_9665
timestamp 1668089732
transform 1 0 24800 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_9666
timestamp 1668089732
transform 1 0 24800 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_9667
timestamp 1668089732
transform 1 0 24800 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_9668
timestamp 1668089732
transform 1 0 24800 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_9669
timestamp 1668089732
transform 1 0 24800 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_9670
timestamp 1668089732
transform 1 0 24800 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_9671
timestamp 1668089732
transform 1 0 24800 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_9672
timestamp 1668089732
transform 1 0 24960 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_9673
timestamp 1668089732
transform 1 0 24960 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_9674
timestamp 1668089732
transform 1 0 24960 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_9675
timestamp 1668089732
transform 1 0 24960 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_9676
timestamp 1668089732
transform 1 0 24960 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_9677
timestamp 1668089732
transform 1 0 24960 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_9678
timestamp 1668089732
transform 1 0 24960 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_9679
timestamp 1668089732
transform 1 0 24960 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_9680
timestamp 1668089732
transform 1 0 24960 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_9681
timestamp 1668089732
transform 1 0 24960 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_9682
timestamp 1668089732
transform 1 0 24960 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_9683
timestamp 1668089732
transform 1 0 24960 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_9684
timestamp 1668089732
transform 1 0 24960 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_9685
timestamp 1668089732
transform 1 0 24960 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_9686
timestamp 1668089732
transform 1 0 24960 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_9687
timestamp 1668089732
transform 1 0 24960 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_9688
timestamp 1668089732
transform 1 0 24960 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_9689
timestamp 1668089732
transform 1 0 24960 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_9690
timestamp 1668089732
transform 1 0 24960 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_9691
timestamp 1668089732
transform 1 0 24960 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_9692
timestamp 1668089732
transform 1 0 24960 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_9693
timestamp 1668089732
transform 1 0 24960 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_9694
timestamp 1668089732
transform 1 0 24960 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_9695
timestamp 1668089732
transform 1 0 24960 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_9696
timestamp 1668089732
transform 1 0 24960 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_9697
timestamp 1668089732
transform 1 0 24960 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_9698
timestamp 1668089732
transform 1 0 24960 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_9699
timestamp 1668089732
transform 1 0 24960 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_9700
timestamp 1668089732
transform 1 0 24960 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_9701
timestamp 1668089732
transform 1 0 24960 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_9702
timestamp 1668089732
transform 1 0 24960 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_9703
timestamp 1668089732
transform 1 0 24960 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_9704
timestamp 1668089732
transform 1 0 24960 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_9705
timestamp 1668089732
transform 1 0 24960 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_9706
timestamp 1668089732
transform 1 0 24960 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_9707
timestamp 1668089732
transform 1 0 24960 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_9708
timestamp 1668089732
transform 1 0 24960 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_9709
timestamp 1668089732
transform 1 0 24960 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_9710
timestamp 1668089732
transform 1 0 24960 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_9711
timestamp 1668089732
transform 1 0 24960 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_9712
timestamp 1668089732
transform 1 0 24960 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_9713
timestamp 1668089732
transform 1 0 24960 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_9714
timestamp 1668089732
transform 1 0 24960 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_9715
timestamp 1668089732
transform 1 0 24960 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_9716
timestamp 1668089732
transform 1 0 24960 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_9717
timestamp 1668089732
transform 1 0 24960 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_9718
timestamp 1668089732
transform 1 0 24960 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_9719
timestamp 1668089732
transform 1 0 24960 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_9720
timestamp 1668089732
transform 1 0 24960 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_9721
timestamp 1668089732
transform 1 0 24960 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_9722
timestamp 1668089732
transform 1 0 24960 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_9723
timestamp 1668089732
transform 1 0 24960 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_9724
timestamp 1668089732
transform 1 0 24960 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_9725
timestamp 1668089732
transform 1 0 24960 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_9726
timestamp 1668089732
transform 1 0 24960 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_9727
timestamp 1668089732
transform 1 0 24960 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_9728
timestamp 1668089732
transform 1 0 24960 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_9729
timestamp 1668089732
transform 1 0 24960 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_9730
timestamp 1668089732
transform 1 0 24960 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_9731
timestamp 1668089732
transform 1 0 24960 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_9732
timestamp 1668089732
transform 1 0 24960 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_9733
timestamp 1668089732
transform 1 0 24960 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_9734
timestamp 1668089732
transform 1 0 25120 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_9735
timestamp 1668089732
transform 1 0 25120 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_9736
timestamp 1668089732
transform 1 0 25120 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_9737
timestamp 1668089732
transform 1 0 25120 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_9738
timestamp 1668089732
transform 1 0 25120 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_9739
timestamp 1668089732
transform 1 0 25120 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_9740
timestamp 1668089732
transform 1 0 25120 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_9741
timestamp 1668089732
transform 1 0 25120 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_9742
timestamp 1668089732
transform 1 0 25120 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_9743
timestamp 1668089732
transform 1 0 25120 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_9744
timestamp 1668089732
transform 1 0 25120 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_9745
timestamp 1668089732
transform 1 0 25120 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_9746
timestamp 1668089732
transform 1 0 25120 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_9747
timestamp 1668089732
transform 1 0 25120 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_9748
timestamp 1668089732
transform 1 0 25120 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_9749
timestamp 1668089732
transform 1 0 25120 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_9750
timestamp 1668089732
transform 1 0 25120 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_9751
timestamp 1668089732
transform 1 0 25120 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_9752
timestamp 1668089732
transform 1 0 25120 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_9753
timestamp 1668089732
transform 1 0 25120 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_9754
timestamp 1668089732
transform 1 0 25120 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_9755
timestamp 1668089732
transform 1 0 25120 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_9756
timestamp 1668089732
transform 1 0 25120 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_9757
timestamp 1668089732
transform 1 0 25120 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_9758
timestamp 1668089732
transform 1 0 25120 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_9759
timestamp 1668089732
transform 1 0 25120 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_9760
timestamp 1668089732
transform 1 0 25120 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_9761
timestamp 1668089732
transform 1 0 25120 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_9762
timestamp 1668089732
transform 1 0 25120 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_9763
timestamp 1668089732
transform 1 0 25120 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_9764
timestamp 1668089732
transform 1 0 25120 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_9765
timestamp 1668089732
transform 1 0 25120 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_9766
timestamp 1668089732
transform 1 0 25120 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_9767
timestamp 1668089732
transform 1 0 25120 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_9768
timestamp 1668089732
transform 1 0 25120 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_9769
timestamp 1668089732
transform 1 0 25120 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_9770
timestamp 1668089732
transform 1 0 25120 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_9771
timestamp 1668089732
transform 1 0 25120 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_9772
timestamp 1668089732
transform 1 0 25120 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_9773
timestamp 1668089732
transform 1 0 25120 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_9774
timestamp 1668089732
transform 1 0 25120 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_9775
timestamp 1668089732
transform 1 0 25120 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_9776
timestamp 1668089732
transform 1 0 25120 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_9777
timestamp 1668089732
transform 1 0 25120 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_9778
timestamp 1668089732
transform 1 0 25120 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_9779
timestamp 1668089732
transform 1 0 25120 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_9780
timestamp 1668089732
transform 1 0 25120 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_9781
timestamp 1668089732
transform 1 0 25120 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_9782
timestamp 1668089732
transform 1 0 25120 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_9783
timestamp 1668089732
transform 1 0 25120 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_9784
timestamp 1668089732
transform 1 0 25120 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_9785
timestamp 1668089732
transform 1 0 25120 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_9786
timestamp 1668089732
transform 1 0 25120 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_9787
timestamp 1668089732
transform 1 0 25120 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_9788
timestamp 1668089732
transform 1 0 25120 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_9789
timestamp 1668089732
transform 1 0 25120 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_9790
timestamp 1668089732
transform 1 0 25120 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_9791
timestamp 1668089732
transform 1 0 25120 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_9792
timestamp 1668089732
transform 1 0 25120 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_9793
timestamp 1668089732
transform 1 0 25120 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_9794
timestamp 1668089732
transform 1 0 25120 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_9795
timestamp 1668089732
transform 1 0 25120 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_9796
timestamp 1668089732
transform 1 0 25280 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_9797
timestamp 1668089732
transform 1 0 25280 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_9798
timestamp 1668089732
transform 1 0 25280 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_9799
timestamp 1668089732
transform 1 0 25280 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_9800
timestamp 1668089732
transform 1 0 25280 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_9801
timestamp 1668089732
transform 1 0 25280 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_9802
timestamp 1668089732
transform 1 0 25280 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_9803
timestamp 1668089732
transform 1 0 25280 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_9804
timestamp 1668089732
transform 1 0 25280 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_9805
timestamp 1668089732
transform 1 0 25280 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_9806
timestamp 1668089732
transform 1 0 25280 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_9807
timestamp 1668089732
transform 1 0 25280 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_9808
timestamp 1668089732
transform 1 0 25280 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_9809
timestamp 1668089732
transform 1 0 25280 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_9810
timestamp 1668089732
transform 1 0 25280 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_9811
timestamp 1668089732
transform 1 0 25280 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_9812
timestamp 1668089732
transform 1 0 25280 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_9813
timestamp 1668089732
transform 1 0 25280 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_9814
timestamp 1668089732
transform 1 0 25280 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_9815
timestamp 1668089732
transform 1 0 25280 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_9816
timestamp 1668089732
transform 1 0 25280 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_9817
timestamp 1668089732
transform 1 0 25280 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_9818
timestamp 1668089732
transform 1 0 25280 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_9819
timestamp 1668089732
transform 1 0 25280 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_9820
timestamp 1668089732
transform 1 0 25280 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_9821
timestamp 1668089732
transform 1 0 25280 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_9822
timestamp 1668089732
transform 1 0 25280 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_9823
timestamp 1668089732
transform 1 0 25280 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_9824
timestamp 1668089732
transform 1 0 25280 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_9825
timestamp 1668089732
transform 1 0 25280 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_9826
timestamp 1668089732
transform 1 0 25280 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_9827
timestamp 1668089732
transform 1 0 25280 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_9828
timestamp 1668089732
transform 1 0 25280 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_9829
timestamp 1668089732
transform 1 0 25280 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_9830
timestamp 1668089732
transform 1 0 25280 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_9831
timestamp 1668089732
transform 1 0 25280 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_9832
timestamp 1668089732
transform 1 0 25280 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_9833
timestamp 1668089732
transform 1 0 25280 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_9834
timestamp 1668089732
transform 1 0 25280 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_9835
timestamp 1668089732
transform 1 0 25280 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_9836
timestamp 1668089732
transform 1 0 25280 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_9837
timestamp 1668089732
transform 1 0 25280 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_9838
timestamp 1668089732
transform 1 0 25280 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_9839
timestamp 1668089732
transform 1 0 25280 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_9840
timestamp 1668089732
transform 1 0 25280 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_9841
timestamp 1668089732
transform 1 0 25280 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_9842
timestamp 1668089732
transform 1 0 25280 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_9843
timestamp 1668089732
transform 1 0 25280 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_9844
timestamp 1668089732
transform 1 0 25280 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_9845
timestamp 1668089732
transform 1 0 25280 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_9846
timestamp 1668089732
transform 1 0 25280 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_9847
timestamp 1668089732
transform 1 0 25280 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_9848
timestamp 1668089732
transform 1 0 25280 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_9849
timestamp 1668089732
transform 1 0 25280 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_9850
timestamp 1668089732
transform 1 0 25280 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_9851
timestamp 1668089732
transform 1 0 25280 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_9852
timestamp 1668089732
transform 1 0 25280 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_9853
timestamp 1668089732
transform 1 0 25280 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_9854
timestamp 1668089732
transform 1 0 25280 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_9855
timestamp 1668089732
transform 1 0 25280 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_9856
timestamp 1668089732
transform 1 0 25280 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_9857
timestamp 1668089732
transform 1 0 25280 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_9858
timestamp 1668089732
transform 1 0 25440 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_9859
timestamp 1668089732
transform 1 0 25440 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_9860
timestamp 1668089732
transform 1 0 25440 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_9861
timestamp 1668089732
transform 1 0 25440 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_9862
timestamp 1668089732
transform 1 0 25440 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_9863
timestamp 1668089732
transform 1 0 25440 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_9864
timestamp 1668089732
transform 1 0 25440 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_9865
timestamp 1668089732
transform 1 0 25440 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_9866
timestamp 1668089732
transform 1 0 25440 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_9867
timestamp 1668089732
transform 1 0 25440 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_9868
timestamp 1668089732
transform 1 0 25440 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_9869
timestamp 1668089732
transform 1 0 25440 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_9870
timestamp 1668089732
transform 1 0 25440 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_9871
timestamp 1668089732
transform 1 0 25440 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_9872
timestamp 1668089732
transform 1 0 25440 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_9873
timestamp 1668089732
transform 1 0 25440 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_9874
timestamp 1668089732
transform 1 0 25440 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_9875
timestamp 1668089732
transform 1 0 25440 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_9876
timestamp 1668089732
transform 1 0 25440 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_9877
timestamp 1668089732
transform 1 0 25440 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_9878
timestamp 1668089732
transform 1 0 25440 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_9879
timestamp 1668089732
transform 1 0 25440 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_9880
timestamp 1668089732
transform 1 0 25440 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_9881
timestamp 1668089732
transform 1 0 25440 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_9882
timestamp 1668089732
transform 1 0 25440 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_9883
timestamp 1668089732
transform 1 0 25440 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_9884
timestamp 1668089732
transform 1 0 25440 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_9885
timestamp 1668089732
transform 1 0 25440 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_9886
timestamp 1668089732
transform 1 0 25440 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_9887
timestamp 1668089732
transform 1 0 25440 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_9888
timestamp 1668089732
transform 1 0 25440 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_9889
timestamp 1668089732
transform 1 0 25440 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_9890
timestamp 1668089732
transform 1 0 25440 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_9891
timestamp 1668089732
transform 1 0 25440 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_9892
timestamp 1668089732
transform 1 0 25440 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_9893
timestamp 1668089732
transform 1 0 25440 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_9894
timestamp 1668089732
transform 1 0 25440 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_9895
timestamp 1668089732
transform 1 0 25440 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_9896
timestamp 1668089732
transform 1 0 25440 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_9897
timestamp 1668089732
transform 1 0 25440 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_9898
timestamp 1668089732
transform 1 0 25440 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_9899
timestamp 1668089732
transform 1 0 25440 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_9900
timestamp 1668089732
transform 1 0 25440 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_9901
timestamp 1668089732
transform 1 0 25440 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_9902
timestamp 1668089732
transform 1 0 25440 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_9903
timestamp 1668089732
transform 1 0 25440 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_9904
timestamp 1668089732
transform 1 0 25440 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_9905
timestamp 1668089732
transform 1 0 25440 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_9906
timestamp 1668089732
transform 1 0 25440 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_9907
timestamp 1668089732
transform 1 0 25440 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_9908
timestamp 1668089732
transform 1 0 25440 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_9909
timestamp 1668089732
transform 1 0 25440 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_9910
timestamp 1668089732
transform 1 0 25440 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_9911
timestamp 1668089732
transform 1 0 25440 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_9912
timestamp 1668089732
transform 1 0 25440 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_9913
timestamp 1668089732
transform 1 0 25440 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_9914
timestamp 1668089732
transform 1 0 25440 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_9915
timestamp 1668089732
transform 1 0 25440 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_9916
timestamp 1668089732
transform 1 0 25440 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_9917
timestamp 1668089732
transform 1 0 25440 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_9918
timestamp 1668089732
transform 1 0 25440 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_9919
timestamp 1668089732
transform 1 0 25440 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_9920
timestamp 1668089732
transform 1 0 25600 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_9921
timestamp 1668089732
transform 1 0 25600 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_9922
timestamp 1668089732
transform 1 0 25600 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_9923
timestamp 1668089732
transform 1 0 25600 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_9924
timestamp 1668089732
transform 1 0 25600 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_9925
timestamp 1668089732
transform 1 0 25600 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_9926
timestamp 1668089732
transform 1 0 25600 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_9927
timestamp 1668089732
transform 1 0 25600 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_9928
timestamp 1668089732
transform 1 0 25600 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_9929
timestamp 1668089732
transform 1 0 25600 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_9930
timestamp 1668089732
transform 1 0 25600 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_9931
timestamp 1668089732
transform 1 0 25600 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_9932
timestamp 1668089732
transform 1 0 25600 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_9933
timestamp 1668089732
transform 1 0 25600 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_9934
timestamp 1668089732
transform 1 0 25600 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_9935
timestamp 1668089732
transform 1 0 25600 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_9936
timestamp 1668089732
transform 1 0 25600 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_9937
timestamp 1668089732
transform 1 0 25600 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_9938
timestamp 1668089732
transform 1 0 25600 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_9939
timestamp 1668089732
transform 1 0 25600 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_9940
timestamp 1668089732
transform 1 0 25600 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_9941
timestamp 1668089732
transform 1 0 25600 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_9942
timestamp 1668089732
transform 1 0 25600 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_9943
timestamp 1668089732
transform 1 0 25600 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_9944
timestamp 1668089732
transform 1 0 25600 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_9945
timestamp 1668089732
transform 1 0 25600 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_9946
timestamp 1668089732
transform 1 0 25600 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_9947
timestamp 1668089732
transform 1 0 25600 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_9948
timestamp 1668089732
transform 1 0 25600 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_9949
timestamp 1668089732
transform 1 0 25600 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_9950
timestamp 1668089732
transform 1 0 25600 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_9951
timestamp 1668089732
transform 1 0 25600 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_9952
timestamp 1668089732
transform 1 0 25600 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_9953
timestamp 1668089732
transform 1 0 25600 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_9954
timestamp 1668089732
transform 1 0 25600 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_9955
timestamp 1668089732
transform 1 0 25600 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_9956
timestamp 1668089732
transform 1 0 25600 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_9957
timestamp 1668089732
transform 1 0 25600 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_9958
timestamp 1668089732
transform 1 0 25600 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_9959
timestamp 1668089732
transform 1 0 25600 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_9960
timestamp 1668089732
transform 1 0 25600 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_9961
timestamp 1668089732
transform 1 0 25600 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_9962
timestamp 1668089732
transform 1 0 25600 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_9963
timestamp 1668089732
transform 1 0 25600 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_9964
timestamp 1668089732
transform 1 0 25600 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_9965
timestamp 1668089732
transform 1 0 25600 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_9966
timestamp 1668089732
transform 1 0 25600 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_9967
timestamp 1668089732
transform 1 0 25600 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_9968
timestamp 1668089732
transform 1 0 25600 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_9969
timestamp 1668089732
transform 1 0 25600 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_9970
timestamp 1668089732
transform 1 0 25600 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_9971
timestamp 1668089732
transform 1 0 25600 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_9972
timestamp 1668089732
transform 1 0 25600 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_9973
timestamp 1668089732
transform 1 0 25600 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_9974
timestamp 1668089732
transform 1 0 25600 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_9975
timestamp 1668089732
transform 1 0 25600 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_9976
timestamp 1668089732
transform 1 0 25600 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_9977
timestamp 1668089732
transform 1 0 25600 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_9978
timestamp 1668089732
transform 1 0 25600 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_9979
timestamp 1668089732
transform 1 0 25600 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_9980
timestamp 1668089732
transform 1 0 25600 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_9981
timestamp 1668089732
transform 1 0 25600 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_9982
timestamp 1668089732
transform 1 0 25760 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_9983
timestamp 1668089732
transform 1 0 25760 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_9984
timestamp 1668089732
transform 1 0 25760 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_9985
timestamp 1668089732
transform 1 0 25760 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_9986
timestamp 1668089732
transform 1 0 25760 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_9987
timestamp 1668089732
transform 1 0 25760 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_9988
timestamp 1668089732
transform 1 0 25760 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_9989
timestamp 1668089732
transform 1 0 25760 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_9990
timestamp 1668089732
transform 1 0 25760 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_9991
timestamp 1668089732
transform 1 0 25760 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_9992
timestamp 1668089732
transform 1 0 25760 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_9993
timestamp 1668089732
transform 1 0 25760 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_9994
timestamp 1668089732
transform 1 0 25760 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_9995
timestamp 1668089732
transform 1 0 25760 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_9996
timestamp 1668089732
transform 1 0 25760 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_9997
timestamp 1668089732
transform 1 0 25760 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_9998
timestamp 1668089732
transform 1 0 25760 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_9999
timestamp 1668089732
transform 1 0 25760 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_10000
timestamp 1668089732
transform 1 0 25760 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_10001
timestamp 1668089732
transform 1 0 25760 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_10002
timestamp 1668089732
transform 1 0 25760 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_10003
timestamp 1668089732
transform 1 0 25760 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_10004
timestamp 1668089732
transform 1 0 25760 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_10005
timestamp 1668089732
transform 1 0 25760 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_10006
timestamp 1668089732
transform 1 0 25760 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_10007
timestamp 1668089732
transform 1 0 25760 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_10008
timestamp 1668089732
transform 1 0 25760 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_10009
timestamp 1668089732
transform 1 0 25760 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_10010
timestamp 1668089732
transform 1 0 25760 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_10011
timestamp 1668089732
transform 1 0 25760 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_10012
timestamp 1668089732
transform 1 0 25760 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_10013
timestamp 1668089732
transform 1 0 25760 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_10014
timestamp 1668089732
transform 1 0 25760 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_10015
timestamp 1668089732
transform 1 0 25760 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_10016
timestamp 1668089732
transform 1 0 25760 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_10017
timestamp 1668089732
transform 1 0 25760 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_10018
timestamp 1668089732
transform 1 0 25760 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_10019
timestamp 1668089732
transform 1 0 25760 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_10020
timestamp 1668089732
transform 1 0 25760 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_10021
timestamp 1668089732
transform 1 0 25760 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_10022
timestamp 1668089732
transform 1 0 25760 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_10023
timestamp 1668089732
transform 1 0 25760 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_10024
timestamp 1668089732
transform 1 0 25760 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_10025
timestamp 1668089732
transform 1 0 25760 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_10026
timestamp 1668089732
transform 1 0 25760 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_10027
timestamp 1668089732
transform 1 0 25760 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_10028
timestamp 1668089732
transform 1 0 25760 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_10029
timestamp 1668089732
transform 1 0 25760 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_10030
timestamp 1668089732
transform 1 0 25760 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_10031
timestamp 1668089732
transform 1 0 25760 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_10032
timestamp 1668089732
transform 1 0 25760 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_10033
timestamp 1668089732
transform 1 0 25760 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_10034
timestamp 1668089732
transform 1 0 25760 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_10035
timestamp 1668089732
transform 1 0 25760 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_10036
timestamp 1668089732
transform 1 0 25760 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_10037
timestamp 1668089732
transform 1 0 25760 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_10038
timestamp 1668089732
transform 1 0 25760 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_10039
timestamp 1668089732
transform 1 0 25760 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_10040
timestamp 1668089732
transform 1 0 25760 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_10041
timestamp 1668089732
transform 1 0 25760 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_10042
timestamp 1668089732
transform 1 0 25760 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_10043
timestamp 1668089732
transform 1 0 25760 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_10044
timestamp 1668089732
transform 1 0 25920 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_10045
timestamp 1668089732
transform 1 0 25920 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_10046
timestamp 1668089732
transform 1 0 25920 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_10047
timestamp 1668089732
transform 1 0 25920 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_10048
timestamp 1668089732
transform 1 0 25920 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_10049
timestamp 1668089732
transform 1 0 25920 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_10050
timestamp 1668089732
transform 1 0 25920 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_10051
timestamp 1668089732
transform 1 0 25920 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_10052
timestamp 1668089732
transform 1 0 25920 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_10053
timestamp 1668089732
transform 1 0 25920 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_10054
timestamp 1668089732
transform 1 0 25920 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_10055
timestamp 1668089732
transform 1 0 25920 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_10056
timestamp 1668089732
transform 1 0 25920 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_10057
timestamp 1668089732
transform 1 0 25920 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_10058
timestamp 1668089732
transform 1 0 25920 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_10059
timestamp 1668089732
transform 1 0 25920 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_10060
timestamp 1668089732
transform 1 0 25920 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_10061
timestamp 1668089732
transform 1 0 25920 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_10062
timestamp 1668089732
transform 1 0 25920 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_10063
timestamp 1668089732
transform 1 0 25920 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_10064
timestamp 1668089732
transform 1 0 25920 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_10065
timestamp 1668089732
transform 1 0 25920 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_10066
timestamp 1668089732
transform 1 0 25920 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_10067
timestamp 1668089732
transform 1 0 25920 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_10068
timestamp 1668089732
transform 1 0 25920 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_10069
timestamp 1668089732
transform 1 0 25920 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_10070
timestamp 1668089732
transform 1 0 25920 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_10071
timestamp 1668089732
transform 1 0 25920 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_10072
timestamp 1668089732
transform 1 0 25920 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_10073
timestamp 1668089732
transform 1 0 25920 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_10074
timestamp 1668089732
transform 1 0 25920 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_10075
timestamp 1668089732
transform 1 0 25920 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_10076
timestamp 1668089732
transform 1 0 25920 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_10077
timestamp 1668089732
transform 1 0 25920 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_10078
timestamp 1668089732
transform 1 0 25920 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_10079
timestamp 1668089732
transform 1 0 25920 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_10080
timestamp 1668089732
transform 1 0 25920 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_10081
timestamp 1668089732
transform 1 0 25920 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_10082
timestamp 1668089732
transform 1 0 25920 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_10083
timestamp 1668089732
transform 1 0 25920 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_10084
timestamp 1668089732
transform 1 0 25920 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_10085
timestamp 1668089732
transform 1 0 25920 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_10086
timestamp 1668089732
transform 1 0 25920 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_10087
timestamp 1668089732
transform 1 0 25920 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_10088
timestamp 1668089732
transform 1 0 25920 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_10089
timestamp 1668089732
transform 1 0 25920 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_10090
timestamp 1668089732
transform 1 0 25920 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_10091
timestamp 1668089732
transform 1 0 25920 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_10092
timestamp 1668089732
transform 1 0 25920 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_10093
timestamp 1668089732
transform 1 0 25920 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_10094
timestamp 1668089732
transform 1 0 25920 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_10095
timestamp 1668089732
transform 1 0 25920 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_10096
timestamp 1668089732
transform 1 0 25920 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_10097
timestamp 1668089732
transform 1 0 25920 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_10098
timestamp 1668089732
transform 1 0 25920 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_10099
timestamp 1668089732
transform 1 0 25920 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_10100
timestamp 1668089732
transform 1 0 25920 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_10101
timestamp 1668089732
transform 1 0 25920 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_10102
timestamp 1668089732
transform 1 0 25920 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_10103
timestamp 1668089732
transform 1 0 25920 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_10104
timestamp 1668089732
transform 1 0 25920 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_10105
timestamp 1668089732
transform 1 0 25920 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_10106
timestamp 1668089732
transform 1 0 26080 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_10107
timestamp 1668089732
transform 1 0 26080 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_10108
timestamp 1668089732
transform 1 0 26080 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_10109
timestamp 1668089732
transform 1 0 26080 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_10110
timestamp 1668089732
transform 1 0 26080 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_10111
timestamp 1668089732
transform 1 0 26080 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_10112
timestamp 1668089732
transform 1 0 26080 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_10113
timestamp 1668089732
transform 1 0 26080 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_10114
timestamp 1668089732
transform 1 0 26080 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_10115
timestamp 1668089732
transform 1 0 26080 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_10116
timestamp 1668089732
transform 1 0 26080 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_10117
timestamp 1668089732
transform 1 0 26080 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_10118
timestamp 1668089732
transform 1 0 26080 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_10119
timestamp 1668089732
transform 1 0 26080 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_10120
timestamp 1668089732
transform 1 0 26080 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_10121
timestamp 1668089732
transform 1 0 26080 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_10122
timestamp 1668089732
transform 1 0 26080 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_10123
timestamp 1668089732
transform 1 0 26080 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_10124
timestamp 1668089732
transform 1 0 26080 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_10125
timestamp 1668089732
transform 1 0 26080 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_10126
timestamp 1668089732
transform 1 0 26080 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_10127
timestamp 1668089732
transform 1 0 26080 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_10128
timestamp 1668089732
transform 1 0 26080 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_10129
timestamp 1668089732
transform 1 0 26080 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_10130
timestamp 1668089732
transform 1 0 26080 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_10131
timestamp 1668089732
transform 1 0 26080 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_10132
timestamp 1668089732
transform 1 0 26080 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_10133
timestamp 1668089732
transform 1 0 26080 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_10134
timestamp 1668089732
transform 1 0 26080 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_10135
timestamp 1668089732
transform 1 0 26080 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_10136
timestamp 1668089732
transform 1 0 26080 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_10137
timestamp 1668089732
transform 1 0 26080 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_10138
timestamp 1668089732
transform 1 0 26080 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_10139
timestamp 1668089732
transform 1 0 26080 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_10140
timestamp 1668089732
transform 1 0 26080 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_10141
timestamp 1668089732
transform 1 0 26080 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_10142
timestamp 1668089732
transform 1 0 26080 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_10143
timestamp 1668089732
transform 1 0 26080 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_10144
timestamp 1668089732
transform 1 0 26080 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_10145
timestamp 1668089732
transform 1 0 26080 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_10146
timestamp 1668089732
transform 1 0 26080 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_10147
timestamp 1668089732
transform 1 0 26080 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_10148
timestamp 1668089732
transform 1 0 26080 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_10149
timestamp 1668089732
transform 1 0 26080 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_10150
timestamp 1668089732
transform 1 0 26080 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_10151
timestamp 1668089732
transform 1 0 26080 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_10152
timestamp 1668089732
transform 1 0 26080 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_10153
timestamp 1668089732
transform 1 0 26080 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_10154
timestamp 1668089732
transform 1 0 26080 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_10155
timestamp 1668089732
transform 1 0 26080 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_10156
timestamp 1668089732
transform 1 0 26080 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_10157
timestamp 1668089732
transform 1 0 26080 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_10158
timestamp 1668089732
transform 1 0 26080 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_10159
timestamp 1668089732
transform 1 0 26080 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_10160
timestamp 1668089732
transform 1 0 26080 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_10161
timestamp 1668089732
transform 1 0 26080 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_10162
timestamp 1668089732
transform 1 0 26080 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_10163
timestamp 1668089732
transform 1 0 26080 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_10164
timestamp 1668089732
transform 1 0 26080 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_10165
timestamp 1668089732
transform 1 0 26080 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_10166
timestamp 1668089732
transform 1 0 26080 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_10167
timestamp 1668089732
transform 1 0 26080 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_10168
timestamp 1668089732
transform 1 0 26240 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_10169
timestamp 1668089732
transform 1 0 26240 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_10170
timestamp 1668089732
transform 1 0 26240 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_10171
timestamp 1668089732
transform 1 0 26240 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_10172
timestamp 1668089732
transform 1 0 26240 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_10173
timestamp 1668089732
transform 1 0 26240 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_10174
timestamp 1668089732
transform 1 0 26240 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_10175
timestamp 1668089732
transform 1 0 26240 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_10176
timestamp 1668089732
transform 1 0 26240 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_10177
timestamp 1668089732
transform 1 0 26240 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_10178
timestamp 1668089732
transform 1 0 26240 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_10179
timestamp 1668089732
transform 1 0 26240 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_10180
timestamp 1668089732
transform 1 0 26240 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_10181
timestamp 1668089732
transform 1 0 26240 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_10182
timestamp 1668089732
transform 1 0 26240 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_10183
timestamp 1668089732
transform 1 0 26240 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_10184
timestamp 1668089732
transform 1 0 26240 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_10185
timestamp 1668089732
transform 1 0 26240 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_10186
timestamp 1668089732
transform 1 0 26240 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_10187
timestamp 1668089732
transform 1 0 26240 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_10188
timestamp 1668089732
transform 1 0 26240 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_10189
timestamp 1668089732
transform 1 0 26240 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_10190
timestamp 1668089732
transform 1 0 26240 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_10191
timestamp 1668089732
transform 1 0 26240 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_10192
timestamp 1668089732
transform 1 0 26240 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_10193
timestamp 1668089732
transform 1 0 26240 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_10194
timestamp 1668089732
transform 1 0 26240 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_10195
timestamp 1668089732
transform 1 0 26240 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_10196
timestamp 1668089732
transform 1 0 26240 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_10197
timestamp 1668089732
transform 1 0 26240 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_10198
timestamp 1668089732
transform 1 0 26240 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_10199
timestamp 1668089732
transform 1 0 26240 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_10200
timestamp 1668089732
transform 1 0 26240 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_10201
timestamp 1668089732
transform 1 0 26240 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_10202
timestamp 1668089732
transform 1 0 26240 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_10203
timestamp 1668089732
transform 1 0 26240 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_10204
timestamp 1668089732
transform 1 0 26240 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_10205
timestamp 1668089732
transform 1 0 26240 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_10206
timestamp 1668089732
transform 1 0 26240 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_10207
timestamp 1668089732
transform 1 0 26240 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_10208
timestamp 1668089732
transform 1 0 26240 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_10209
timestamp 1668089732
transform 1 0 26240 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_10210
timestamp 1668089732
transform 1 0 26240 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_10211
timestamp 1668089732
transform 1 0 26240 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_10212
timestamp 1668089732
transform 1 0 26240 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_10213
timestamp 1668089732
transform 1 0 26240 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_10214
timestamp 1668089732
transform 1 0 26240 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_10215
timestamp 1668089732
transform 1 0 26240 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_10216
timestamp 1668089732
transform 1 0 26240 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_10217
timestamp 1668089732
transform 1 0 26240 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_10218
timestamp 1668089732
transform 1 0 26240 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_10219
timestamp 1668089732
transform 1 0 26240 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_10220
timestamp 1668089732
transform 1 0 26240 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_10221
timestamp 1668089732
transform 1 0 26240 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_10222
timestamp 1668089732
transform 1 0 26240 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_10223
timestamp 1668089732
transform 1 0 26240 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_10224
timestamp 1668089732
transform 1 0 26240 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_10225
timestamp 1668089732
transform 1 0 26240 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_10226
timestamp 1668089732
transform 1 0 26240 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_10227
timestamp 1668089732
transform 1 0 26240 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_10228
timestamp 1668089732
transform 1 0 26240 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_10229
timestamp 1668089732
transform 1 0 26240 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_10230
timestamp 1668089732
transform 1 0 26400 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_10231
timestamp 1668089732
transform 1 0 26400 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_10232
timestamp 1668089732
transform 1 0 26400 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_10233
timestamp 1668089732
transform 1 0 26400 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_10234
timestamp 1668089732
transform 1 0 26400 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_10235
timestamp 1668089732
transform 1 0 26400 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_10236
timestamp 1668089732
transform 1 0 26400 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_10237
timestamp 1668089732
transform 1 0 26400 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_10238
timestamp 1668089732
transform 1 0 26400 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_10239
timestamp 1668089732
transform 1 0 26400 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_10240
timestamp 1668089732
transform 1 0 26400 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_10241
timestamp 1668089732
transform 1 0 26400 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_10242
timestamp 1668089732
transform 1 0 26400 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_10243
timestamp 1668089732
transform 1 0 26400 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_10244
timestamp 1668089732
transform 1 0 26400 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_10245
timestamp 1668089732
transform 1 0 26400 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_10246
timestamp 1668089732
transform 1 0 26400 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_10247
timestamp 1668089732
transform 1 0 26400 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_10248
timestamp 1668089732
transform 1 0 26400 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_10249
timestamp 1668089732
transform 1 0 26400 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_10250
timestamp 1668089732
transform 1 0 26400 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_10251
timestamp 1668089732
transform 1 0 26400 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_10252
timestamp 1668089732
transform 1 0 26400 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_10253
timestamp 1668089732
transform 1 0 26400 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_10254
timestamp 1668089732
transform 1 0 26400 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_10255
timestamp 1668089732
transform 1 0 26400 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_10256
timestamp 1668089732
transform 1 0 26400 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_10257
timestamp 1668089732
transform 1 0 26400 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_10258
timestamp 1668089732
transform 1 0 26400 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_10259
timestamp 1668089732
transform 1 0 26400 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_10260
timestamp 1668089732
transform 1 0 26400 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_10261
timestamp 1668089732
transform 1 0 26400 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_10262
timestamp 1668089732
transform 1 0 26400 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_10263
timestamp 1668089732
transform 1 0 26400 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_10264
timestamp 1668089732
transform 1 0 26400 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_10265
timestamp 1668089732
transform 1 0 26400 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_10266
timestamp 1668089732
transform 1 0 26400 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_10267
timestamp 1668089732
transform 1 0 26400 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_10268
timestamp 1668089732
transform 1 0 26400 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_10269
timestamp 1668089732
transform 1 0 26400 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_10270
timestamp 1668089732
transform 1 0 26400 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_10271
timestamp 1668089732
transform 1 0 26400 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_10272
timestamp 1668089732
transform 1 0 26400 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_10273
timestamp 1668089732
transform 1 0 26400 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_10274
timestamp 1668089732
transform 1 0 26400 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_10275
timestamp 1668089732
transform 1 0 26400 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_10276
timestamp 1668089732
transform 1 0 26400 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_10277
timestamp 1668089732
transform 1 0 26400 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_10278
timestamp 1668089732
transform 1 0 26400 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_10279
timestamp 1668089732
transform 1 0 26400 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_10280
timestamp 1668089732
transform 1 0 26400 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_10281
timestamp 1668089732
transform 1 0 26400 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_10282
timestamp 1668089732
transform 1 0 26400 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_10283
timestamp 1668089732
transform 1 0 26400 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_10284
timestamp 1668089732
transform 1 0 26400 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_10285
timestamp 1668089732
transform 1 0 26400 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_10286
timestamp 1668089732
transform 1 0 26400 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_10287
timestamp 1668089732
transform 1 0 26400 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_10288
timestamp 1668089732
transform 1 0 26400 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_10289
timestamp 1668089732
transform 1 0 26400 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_10290
timestamp 1668089732
transform 1 0 26400 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_10291
timestamp 1668089732
transform 1 0 26400 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_10292
timestamp 1668089732
transform 1 0 26560 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_10293
timestamp 1668089732
transform 1 0 26560 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_10294
timestamp 1668089732
transform 1 0 26560 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_10295
timestamp 1668089732
transform 1 0 26560 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_10296
timestamp 1668089732
transform 1 0 26560 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_10297
timestamp 1668089732
transform 1 0 26560 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_10298
timestamp 1668089732
transform 1 0 26560 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_10299
timestamp 1668089732
transform 1 0 26560 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_10300
timestamp 1668089732
transform 1 0 26560 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_10301
timestamp 1668089732
transform 1 0 26560 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_10302
timestamp 1668089732
transform 1 0 26560 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_10303
timestamp 1668089732
transform 1 0 26560 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_10304
timestamp 1668089732
transform 1 0 26560 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_10305
timestamp 1668089732
transform 1 0 26560 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_10306
timestamp 1668089732
transform 1 0 26560 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_10307
timestamp 1668089732
transform 1 0 26560 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_10308
timestamp 1668089732
transform 1 0 26560 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_10309
timestamp 1668089732
transform 1 0 26560 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_10310
timestamp 1668089732
transform 1 0 26560 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_10311
timestamp 1668089732
transform 1 0 26560 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_10312
timestamp 1668089732
transform 1 0 26560 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_10313
timestamp 1668089732
transform 1 0 26560 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_10314
timestamp 1668089732
transform 1 0 26560 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_10315
timestamp 1668089732
transform 1 0 26560 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_10316
timestamp 1668089732
transform 1 0 26560 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_10317
timestamp 1668089732
transform 1 0 26560 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_10318
timestamp 1668089732
transform 1 0 26560 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_10319
timestamp 1668089732
transform 1 0 26560 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_10320
timestamp 1668089732
transform 1 0 26560 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_10321
timestamp 1668089732
transform 1 0 26560 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_10322
timestamp 1668089732
transform 1 0 26560 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_10323
timestamp 1668089732
transform 1 0 26560 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_10324
timestamp 1668089732
transform 1 0 26560 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_10325
timestamp 1668089732
transform 1 0 26560 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_10326
timestamp 1668089732
transform 1 0 26560 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_10327
timestamp 1668089732
transform 1 0 26560 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_10328
timestamp 1668089732
transform 1 0 26560 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_10329
timestamp 1668089732
transform 1 0 26560 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_10330
timestamp 1668089732
transform 1 0 26560 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_10331
timestamp 1668089732
transform 1 0 26560 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_10332
timestamp 1668089732
transform 1 0 26560 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_10333
timestamp 1668089732
transform 1 0 26560 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_10334
timestamp 1668089732
transform 1 0 26560 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_10335
timestamp 1668089732
transform 1 0 26560 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_10336
timestamp 1668089732
transform 1 0 26560 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_10337
timestamp 1668089732
transform 1 0 26560 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_10338
timestamp 1668089732
transform 1 0 26560 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_10339
timestamp 1668089732
transform 1 0 26560 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_10340
timestamp 1668089732
transform 1 0 26560 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_10341
timestamp 1668089732
transform 1 0 26560 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_10342
timestamp 1668089732
transform 1 0 26560 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_10343
timestamp 1668089732
transform 1 0 26560 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_10344
timestamp 1668089732
transform 1 0 26560 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_10345
timestamp 1668089732
transform 1 0 26560 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_10346
timestamp 1668089732
transform 1 0 26560 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_10347
timestamp 1668089732
transform 1 0 26560 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_10348
timestamp 1668089732
transform 1 0 26560 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_10349
timestamp 1668089732
transform 1 0 26560 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_10350
timestamp 1668089732
transform 1 0 26560 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_10351
timestamp 1668089732
transform 1 0 26560 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_10352
timestamp 1668089732
transform 1 0 26560 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_10353
timestamp 1668089732
transform 1 0 26560 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_10354
timestamp 1668089732
transform 1 0 26720 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_10355
timestamp 1668089732
transform 1 0 26720 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_10356
timestamp 1668089732
transform 1 0 26720 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_10357
timestamp 1668089732
transform 1 0 26720 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_10358
timestamp 1668089732
transform 1 0 26720 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_10359
timestamp 1668089732
transform 1 0 26720 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_10360
timestamp 1668089732
transform 1 0 26720 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_10361
timestamp 1668089732
transform 1 0 26720 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_10362
timestamp 1668089732
transform 1 0 26720 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_10363
timestamp 1668089732
transform 1 0 26720 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_10364
timestamp 1668089732
transform 1 0 26720 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_10365
timestamp 1668089732
transform 1 0 26720 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_10366
timestamp 1668089732
transform 1 0 26720 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_10367
timestamp 1668089732
transform 1 0 26720 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_10368
timestamp 1668089732
transform 1 0 26720 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_10369
timestamp 1668089732
transform 1 0 26720 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_10370
timestamp 1668089732
transform 1 0 26720 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_10371
timestamp 1668089732
transform 1 0 26720 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_10372
timestamp 1668089732
transform 1 0 26720 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_10373
timestamp 1668089732
transform 1 0 26720 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_10374
timestamp 1668089732
transform 1 0 26720 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_10375
timestamp 1668089732
transform 1 0 26720 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_10376
timestamp 1668089732
transform 1 0 26720 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_10377
timestamp 1668089732
transform 1 0 26720 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_10378
timestamp 1668089732
transform 1 0 26720 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_10379
timestamp 1668089732
transform 1 0 26720 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_10380
timestamp 1668089732
transform 1 0 26720 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_10381
timestamp 1668089732
transform 1 0 26720 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_10382
timestamp 1668089732
transform 1 0 26720 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_10383
timestamp 1668089732
transform 1 0 26720 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_10384
timestamp 1668089732
transform 1 0 26720 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_10385
timestamp 1668089732
transform 1 0 26720 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_10386
timestamp 1668089732
transform 1 0 26720 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_10387
timestamp 1668089732
transform 1 0 26720 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_10388
timestamp 1668089732
transform 1 0 26720 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_10389
timestamp 1668089732
transform 1 0 26720 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_10390
timestamp 1668089732
transform 1 0 26720 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_10391
timestamp 1668089732
transform 1 0 26720 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_10392
timestamp 1668089732
transform 1 0 26720 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_10393
timestamp 1668089732
transform 1 0 26720 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_10394
timestamp 1668089732
transform 1 0 26720 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_10395
timestamp 1668089732
transform 1 0 26720 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_10396
timestamp 1668089732
transform 1 0 26720 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_10397
timestamp 1668089732
transform 1 0 26720 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_10398
timestamp 1668089732
transform 1 0 26720 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_10399
timestamp 1668089732
transform 1 0 26720 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_10400
timestamp 1668089732
transform 1 0 26720 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_10401
timestamp 1668089732
transform 1 0 26720 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_10402
timestamp 1668089732
transform 1 0 26720 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_10403
timestamp 1668089732
transform 1 0 26720 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_10404
timestamp 1668089732
transform 1 0 26720 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_10405
timestamp 1668089732
transform 1 0 26720 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_10406
timestamp 1668089732
transform 1 0 26720 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_10407
timestamp 1668089732
transform 1 0 26720 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_10408
timestamp 1668089732
transform 1 0 26720 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_10409
timestamp 1668089732
transform 1 0 26720 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_10410
timestamp 1668089732
transform 1 0 26720 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_10411
timestamp 1668089732
transform 1 0 26720 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_10412
timestamp 1668089732
transform 1 0 26720 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_10413
timestamp 1668089732
transform 1 0 26720 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_10414
timestamp 1668089732
transform 1 0 26720 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_10415
timestamp 1668089732
transform 1 0 26720 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_10416
timestamp 1668089732
transform 1 0 26880 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_10417
timestamp 1668089732
transform 1 0 26880 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_10418
timestamp 1668089732
transform 1 0 26880 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_10419
timestamp 1668089732
transform 1 0 26880 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_10420
timestamp 1668089732
transform 1 0 26880 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_10421
timestamp 1668089732
transform 1 0 26880 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_10422
timestamp 1668089732
transform 1 0 26880 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_10423
timestamp 1668089732
transform 1 0 26880 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_10424
timestamp 1668089732
transform 1 0 26880 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_10425
timestamp 1668089732
transform 1 0 26880 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_10426
timestamp 1668089732
transform 1 0 26880 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_10427
timestamp 1668089732
transform 1 0 26880 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_10428
timestamp 1668089732
transform 1 0 26880 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_10429
timestamp 1668089732
transform 1 0 26880 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_10430
timestamp 1668089732
transform 1 0 26880 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_10431
timestamp 1668089732
transform 1 0 26880 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_10432
timestamp 1668089732
transform 1 0 26880 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_10433
timestamp 1668089732
transform 1 0 26880 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_10434
timestamp 1668089732
transform 1 0 26880 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_10435
timestamp 1668089732
transform 1 0 26880 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_10436
timestamp 1668089732
transform 1 0 26880 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_10437
timestamp 1668089732
transform 1 0 26880 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_10438
timestamp 1668089732
transform 1 0 26880 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_10439
timestamp 1668089732
transform 1 0 26880 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_10440
timestamp 1668089732
transform 1 0 26880 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_10441
timestamp 1668089732
transform 1 0 26880 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_10442
timestamp 1668089732
transform 1 0 26880 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_10443
timestamp 1668089732
transform 1 0 26880 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_10444
timestamp 1668089732
transform 1 0 26880 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_10445
timestamp 1668089732
transform 1 0 26880 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_10446
timestamp 1668089732
transform 1 0 26880 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_10447
timestamp 1668089732
transform 1 0 26880 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_10448
timestamp 1668089732
transform 1 0 26880 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_10449
timestamp 1668089732
transform 1 0 26880 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_10450
timestamp 1668089732
transform 1 0 26880 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_10451
timestamp 1668089732
transform 1 0 26880 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_10452
timestamp 1668089732
transform 1 0 26880 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_10453
timestamp 1668089732
transform 1 0 26880 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_10454
timestamp 1668089732
transform 1 0 26880 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_10455
timestamp 1668089732
transform 1 0 26880 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_10456
timestamp 1668089732
transform 1 0 26880 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_10457
timestamp 1668089732
transform 1 0 26880 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_10458
timestamp 1668089732
transform 1 0 26880 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_10459
timestamp 1668089732
transform 1 0 26880 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_10460
timestamp 1668089732
transform 1 0 26880 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_10461
timestamp 1668089732
transform 1 0 26880 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_10462
timestamp 1668089732
transform 1 0 26880 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_10463
timestamp 1668089732
transform 1 0 26880 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_10464
timestamp 1668089732
transform 1 0 26880 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_10465
timestamp 1668089732
transform 1 0 26880 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_10466
timestamp 1668089732
transform 1 0 26880 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_10467
timestamp 1668089732
transform 1 0 26880 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_10468
timestamp 1668089732
transform 1 0 26880 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_10469
timestamp 1668089732
transform 1 0 26880 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_10470
timestamp 1668089732
transform 1 0 26880 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_10471
timestamp 1668089732
transform 1 0 26880 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_10472
timestamp 1668089732
transform 1 0 26880 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_10473
timestamp 1668089732
transform 1 0 26880 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_10474
timestamp 1668089732
transform 1 0 26880 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_10475
timestamp 1668089732
transform 1 0 26880 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_10476
timestamp 1668089732
transform 1 0 26880 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_10477
timestamp 1668089732
transform 1 0 26880 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_10478
timestamp 1668089732
transform 1 0 27040 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_10479
timestamp 1668089732
transform 1 0 27040 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_10480
timestamp 1668089732
transform 1 0 27040 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_10481
timestamp 1668089732
transform 1 0 27040 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_10482
timestamp 1668089732
transform 1 0 27040 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_10483
timestamp 1668089732
transform 1 0 27040 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_10484
timestamp 1668089732
transform 1 0 27040 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_10485
timestamp 1668089732
transform 1 0 27040 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_10486
timestamp 1668089732
transform 1 0 27040 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_10487
timestamp 1668089732
transform 1 0 27040 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_10488
timestamp 1668089732
transform 1 0 27040 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_10489
timestamp 1668089732
transform 1 0 27040 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_10490
timestamp 1668089732
transform 1 0 27040 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_10491
timestamp 1668089732
transform 1 0 27040 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_10492
timestamp 1668089732
transform 1 0 27040 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_10493
timestamp 1668089732
transform 1 0 27040 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_10494
timestamp 1668089732
transform 1 0 27040 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_10495
timestamp 1668089732
transform 1 0 27040 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_10496
timestamp 1668089732
transform 1 0 27040 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_10497
timestamp 1668089732
transform 1 0 27040 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_10498
timestamp 1668089732
transform 1 0 27040 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_10499
timestamp 1668089732
transform 1 0 27040 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_10500
timestamp 1668089732
transform 1 0 27040 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_10501
timestamp 1668089732
transform 1 0 27040 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_10502
timestamp 1668089732
transform 1 0 27040 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_10503
timestamp 1668089732
transform 1 0 27040 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_10504
timestamp 1668089732
transform 1 0 27040 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_10505
timestamp 1668089732
transform 1 0 27040 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_10506
timestamp 1668089732
transform 1 0 27040 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_10507
timestamp 1668089732
transform 1 0 27040 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_10508
timestamp 1668089732
transform 1 0 27040 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_10509
timestamp 1668089732
transform 1 0 27040 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_10510
timestamp 1668089732
transform 1 0 27040 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_10511
timestamp 1668089732
transform 1 0 27040 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_10512
timestamp 1668089732
transform 1 0 27040 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_10513
timestamp 1668089732
transform 1 0 27040 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_10514
timestamp 1668089732
transform 1 0 27040 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_10515
timestamp 1668089732
transform 1 0 27040 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_10516
timestamp 1668089732
transform 1 0 27040 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_10517
timestamp 1668089732
transform 1 0 27040 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_10518
timestamp 1668089732
transform 1 0 27040 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_10519
timestamp 1668089732
transform 1 0 27040 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_10520
timestamp 1668089732
transform 1 0 27040 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_10521
timestamp 1668089732
transform 1 0 27040 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_10522
timestamp 1668089732
transform 1 0 27040 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_10523
timestamp 1668089732
transform 1 0 27040 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_10524
timestamp 1668089732
transform 1 0 27040 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_10525
timestamp 1668089732
transform 1 0 27040 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_10526
timestamp 1668089732
transform 1 0 27040 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_10527
timestamp 1668089732
transform 1 0 27040 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_10528
timestamp 1668089732
transform 1 0 27040 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_10529
timestamp 1668089732
transform 1 0 27040 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_10530
timestamp 1668089732
transform 1 0 27040 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_10531
timestamp 1668089732
transform 1 0 27040 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_10532
timestamp 1668089732
transform 1 0 27040 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_10533
timestamp 1668089732
transform 1 0 27040 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_10534
timestamp 1668089732
transform 1 0 27040 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_10535
timestamp 1668089732
transform 1 0 27040 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_10536
timestamp 1668089732
transform 1 0 27040 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_10537
timestamp 1668089732
transform 1 0 27040 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_10538
timestamp 1668089732
transform 1 0 27040 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_10539
timestamp 1668089732
transform 1 0 27040 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_10540
timestamp 1668089732
transform 1 0 27200 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_10541
timestamp 1668089732
transform 1 0 27200 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_10542
timestamp 1668089732
transform 1 0 27200 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_10543
timestamp 1668089732
transform 1 0 27200 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_10544
timestamp 1668089732
transform 1 0 27200 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_10545
timestamp 1668089732
transform 1 0 27200 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_10546
timestamp 1668089732
transform 1 0 27200 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_10547
timestamp 1668089732
transform 1 0 27200 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_10548
timestamp 1668089732
transform 1 0 27200 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_10549
timestamp 1668089732
transform 1 0 27200 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_10550
timestamp 1668089732
transform 1 0 27200 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_10551
timestamp 1668089732
transform 1 0 27200 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_10552
timestamp 1668089732
transform 1 0 27200 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_10553
timestamp 1668089732
transform 1 0 27200 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_10554
timestamp 1668089732
transform 1 0 27200 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_10555
timestamp 1668089732
transform 1 0 27200 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_10556
timestamp 1668089732
transform 1 0 27200 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_10557
timestamp 1668089732
transform 1 0 27200 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_10558
timestamp 1668089732
transform 1 0 27200 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_10559
timestamp 1668089732
transform 1 0 27200 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_10560
timestamp 1668089732
transform 1 0 27200 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_10561
timestamp 1668089732
transform 1 0 27200 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_10562
timestamp 1668089732
transform 1 0 27200 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_10563
timestamp 1668089732
transform 1 0 27200 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_10564
timestamp 1668089732
transform 1 0 27200 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_10565
timestamp 1668089732
transform 1 0 27200 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_10566
timestamp 1668089732
transform 1 0 27200 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_10567
timestamp 1668089732
transform 1 0 27200 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_10568
timestamp 1668089732
transform 1 0 27200 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_10569
timestamp 1668089732
transform 1 0 27200 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_10570
timestamp 1668089732
transform 1 0 27200 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_10571
timestamp 1668089732
transform 1 0 27200 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_10572
timestamp 1668089732
transform 1 0 27200 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_10573
timestamp 1668089732
transform 1 0 27200 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_10574
timestamp 1668089732
transform 1 0 27200 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_10575
timestamp 1668089732
transform 1 0 27200 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_10576
timestamp 1668089732
transform 1 0 27200 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_10577
timestamp 1668089732
transform 1 0 27200 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_10578
timestamp 1668089732
transform 1 0 27200 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_10579
timestamp 1668089732
transform 1 0 27200 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_10580
timestamp 1668089732
transform 1 0 27200 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_10581
timestamp 1668089732
transform 1 0 27200 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_10582
timestamp 1668089732
transform 1 0 27200 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_10583
timestamp 1668089732
transform 1 0 27200 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_10584
timestamp 1668089732
transform 1 0 27200 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_10585
timestamp 1668089732
transform 1 0 27200 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_10586
timestamp 1668089732
transform 1 0 27200 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_10587
timestamp 1668089732
transform 1 0 27200 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_10588
timestamp 1668089732
transform 1 0 27200 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_10589
timestamp 1668089732
transform 1 0 27200 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_10590
timestamp 1668089732
transform 1 0 27200 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_10591
timestamp 1668089732
transform 1 0 27200 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_10592
timestamp 1668089732
transform 1 0 27200 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_10593
timestamp 1668089732
transform 1 0 27200 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_10594
timestamp 1668089732
transform 1 0 27200 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_10595
timestamp 1668089732
transform 1 0 27200 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_10596
timestamp 1668089732
transform 1 0 27200 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_10597
timestamp 1668089732
transform 1 0 27200 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_10598
timestamp 1668089732
transform 1 0 27200 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_10599
timestamp 1668089732
transform 1 0 27200 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_10600
timestamp 1668089732
transform 1 0 27200 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_10601
timestamp 1668089732
transform 1 0 27200 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_10602
timestamp 1668089732
transform 1 0 27360 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_10603
timestamp 1668089732
transform 1 0 27360 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_10604
timestamp 1668089732
transform 1 0 27360 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_10605
timestamp 1668089732
transform 1 0 27360 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_10606
timestamp 1668089732
transform 1 0 27360 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_10607
timestamp 1668089732
transform 1 0 27360 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_10608
timestamp 1668089732
transform 1 0 27360 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_10609
timestamp 1668089732
transform 1 0 27360 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_10610
timestamp 1668089732
transform 1 0 27360 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_10611
timestamp 1668089732
transform 1 0 27360 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_10612
timestamp 1668089732
transform 1 0 27360 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_10613
timestamp 1668089732
transform 1 0 27360 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_10614
timestamp 1668089732
transform 1 0 27360 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_10615
timestamp 1668089732
transform 1 0 27360 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_10616
timestamp 1668089732
transform 1 0 27360 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_10617
timestamp 1668089732
transform 1 0 27360 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_10618
timestamp 1668089732
transform 1 0 27360 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_10619
timestamp 1668089732
transform 1 0 27360 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_10620
timestamp 1668089732
transform 1 0 27360 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_10621
timestamp 1668089732
transform 1 0 27360 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_10622
timestamp 1668089732
transform 1 0 27360 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_10623
timestamp 1668089732
transform 1 0 27360 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_10624
timestamp 1668089732
transform 1 0 27360 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_10625
timestamp 1668089732
transform 1 0 27360 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_10626
timestamp 1668089732
transform 1 0 27360 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_10627
timestamp 1668089732
transform 1 0 27360 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_10628
timestamp 1668089732
transform 1 0 27360 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_10629
timestamp 1668089732
transform 1 0 27360 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_10630
timestamp 1668089732
transform 1 0 27360 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_10631
timestamp 1668089732
transform 1 0 27360 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_10632
timestamp 1668089732
transform 1 0 27360 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_10633
timestamp 1668089732
transform 1 0 27360 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_10634
timestamp 1668089732
transform 1 0 27360 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_10635
timestamp 1668089732
transform 1 0 27360 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_10636
timestamp 1668089732
transform 1 0 27360 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_10637
timestamp 1668089732
transform 1 0 27360 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_10638
timestamp 1668089732
transform 1 0 27360 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_10639
timestamp 1668089732
transform 1 0 27360 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_10640
timestamp 1668089732
transform 1 0 27360 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_10641
timestamp 1668089732
transform 1 0 27360 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_10642
timestamp 1668089732
transform 1 0 27360 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_10643
timestamp 1668089732
transform 1 0 27360 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_10644
timestamp 1668089732
transform 1 0 27360 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_10645
timestamp 1668089732
transform 1 0 27360 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_10646
timestamp 1668089732
transform 1 0 27360 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_10647
timestamp 1668089732
transform 1 0 27360 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_10648
timestamp 1668089732
transform 1 0 27360 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_10649
timestamp 1668089732
transform 1 0 27360 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_10650
timestamp 1668089732
transform 1 0 27360 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_10651
timestamp 1668089732
transform 1 0 27360 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_10652
timestamp 1668089732
transform 1 0 27360 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_10653
timestamp 1668089732
transform 1 0 27360 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_10654
timestamp 1668089732
transform 1 0 27360 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_10655
timestamp 1668089732
transform 1 0 27360 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_10656
timestamp 1668089732
transform 1 0 27360 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_10657
timestamp 1668089732
transform 1 0 27360 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_10658
timestamp 1668089732
transform 1 0 27360 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_10659
timestamp 1668089732
transform 1 0 27360 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_10660
timestamp 1668089732
transform 1 0 27360 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_10661
timestamp 1668089732
transform 1 0 27360 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_10662
timestamp 1668089732
transform 1 0 27360 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_10663
timestamp 1668089732
transform 1 0 27360 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_10664
timestamp 1668089732
transform 1 0 27520 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_10665
timestamp 1668089732
transform 1 0 27520 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_10666
timestamp 1668089732
transform 1 0 27520 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_10667
timestamp 1668089732
transform 1 0 27520 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_10668
timestamp 1668089732
transform 1 0 27520 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_10669
timestamp 1668089732
transform 1 0 27520 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_10670
timestamp 1668089732
transform 1 0 27520 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_10671
timestamp 1668089732
transform 1 0 27520 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_10672
timestamp 1668089732
transform 1 0 27520 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_10673
timestamp 1668089732
transform 1 0 27520 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_10674
timestamp 1668089732
transform 1 0 27520 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_10675
timestamp 1668089732
transform 1 0 27520 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_10676
timestamp 1668089732
transform 1 0 27520 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_10677
timestamp 1668089732
transform 1 0 27520 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_10678
timestamp 1668089732
transform 1 0 27520 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_10679
timestamp 1668089732
transform 1 0 27520 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_10680
timestamp 1668089732
transform 1 0 27520 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_10681
timestamp 1668089732
transform 1 0 27520 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_10682
timestamp 1668089732
transform 1 0 27520 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_10683
timestamp 1668089732
transform 1 0 27520 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_10684
timestamp 1668089732
transform 1 0 27520 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_10685
timestamp 1668089732
transform 1 0 27520 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_10686
timestamp 1668089732
transform 1 0 27520 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_10687
timestamp 1668089732
transform 1 0 27520 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_10688
timestamp 1668089732
transform 1 0 27520 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_10689
timestamp 1668089732
transform 1 0 27520 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_10690
timestamp 1668089732
transform 1 0 27520 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_10691
timestamp 1668089732
transform 1 0 27520 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_10692
timestamp 1668089732
transform 1 0 27520 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_10693
timestamp 1668089732
transform 1 0 27520 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_10694
timestamp 1668089732
transform 1 0 27520 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_10695
timestamp 1668089732
transform 1 0 27520 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_10696
timestamp 1668089732
transform 1 0 27520 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_10697
timestamp 1668089732
transform 1 0 27520 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_10698
timestamp 1668089732
transform 1 0 27520 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_10699
timestamp 1668089732
transform 1 0 27520 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_10700
timestamp 1668089732
transform 1 0 27520 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_10701
timestamp 1668089732
transform 1 0 27520 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_10702
timestamp 1668089732
transform 1 0 27520 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_10703
timestamp 1668089732
transform 1 0 27520 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_10704
timestamp 1668089732
transform 1 0 27520 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_10705
timestamp 1668089732
transform 1 0 27520 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_10706
timestamp 1668089732
transform 1 0 27520 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_10707
timestamp 1668089732
transform 1 0 27520 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_10708
timestamp 1668089732
transform 1 0 27520 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_10709
timestamp 1668089732
transform 1 0 27520 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_10710
timestamp 1668089732
transform 1 0 27520 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_10711
timestamp 1668089732
transform 1 0 27520 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_10712
timestamp 1668089732
transform 1 0 27520 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_10713
timestamp 1668089732
transform 1 0 27520 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_10714
timestamp 1668089732
transform 1 0 27520 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_10715
timestamp 1668089732
transform 1 0 27520 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_10716
timestamp 1668089732
transform 1 0 27520 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_10717
timestamp 1668089732
transform 1 0 27520 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_10718
timestamp 1668089732
transform 1 0 27520 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_10719
timestamp 1668089732
transform 1 0 27520 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_10720
timestamp 1668089732
transform 1 0 27520 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_10721
timestamp 1668089732
transform 1 0 27520 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_10722
timestamp 1668089732
transform 1 0 27520 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_10723
timestamp 1668089732
transform 1 0 27520 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_10724
timestamp 1668089732
transform 1 0 27520 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_10725
timestamp 1668089732
transform 1 0 27520 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_10726
timestamp 1668089732
transform 1 0 27680 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_10727
timestamp 1668089732
transform 1 0 27680 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_10728
timestamp 1668089732
transform 1 0 27680 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_10729
timestamp 1668089732
transform 1 0 27680 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_10730
timestamp 1668089732
transform 1 0 27680 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_10731
timestamp 1668089732
transform 1 0 27680 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_10732
timestamp 1668089732
transform 1 0 27680 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_10733
timestamp 1668089732
transform 1 0 27680 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_10734
timestamp 1668089732
transform 1 0 27680 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_10735
timestamp 1668089732
transform 1 0 27680 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_10736
timestamp 1668089732
transform 1 0 27680 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_10737
timestamp 1668089732
transform 1 0 27680 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_10738
timestamp 1668089732
transform 1 0 27680 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_10739
timestamp 1668089732
transform 1 0 27680 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_10740
timestamp 1668089732
transform 1 0 27680 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_10741
timestamp 1668089732
transform 1 0 27680 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_10742
timestamp 1668089732
transform 1 0 27680 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_10743
timestamp 1668089732
transform 1 0 27680 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_10744
timestamp 1668089732
transform 1 0 27680 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_10745
timestamp 1668089732
transform 1 0 27680 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_10746
timestamp 1668089732
transform 1 0 27680 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_10747
timestamp 1668089732
transform 1 0 27680 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_10748
timestamp 1668089732
transform 1 0 27680 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_10749
timestamp 1668089732
transform 1 0 27680 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_10750
timestamp 1668089732
transform 1 0 27680 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_10751
timestamp 1668089732
transform 1 0 27680 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_10752
timestamp 1668089732
transform 1 0 27680 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_10753
timestamp 1668089732
transform 1 0 27680 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_10754
timestamp 1668089732
transform 1 0 27680 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_10755
timestamp 1668089732
transform 1 0 27680 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_10756
timestamp 1668089732
transform 1 0 27680 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_10757
timestamp 1668089732
transform 1 0 27680 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_10758
timestamp 1668089732
transform 1 0 27680 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_10759
timestamp 1668089732
transform 1 0 27680 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_10760
timestamp 1668089732
transform 1 0 27680 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_10761
timestamp 1668089732
transform 1 0 27680 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_10762
timestamp 1668089732
transform 1 0 27680 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_10763
timestamp 1668089732
transform 1 0 27680 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_10764
timestamp 1668089732
transform 1 0 27680 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_10765
timestamp 1668089732
transform 1 0 27680 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_10766
timestamp 1668089732
transform 1 0 27680 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_10767
timestamp 1668089732
transform 1 0 27680 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_10768
timestamp 1668089732
transform 1 0 27680 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_10769
timestamp 1668089732
transform 1 0 27680 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_10770
timestamp 1668089732
transform 1 0 27680 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_10771
timestamp 1668089732
transform 1 0 27680 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_10772
timestamp 1668089732
transform 1 0 27680 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_10773
timestamp 1668089732
transform 1 0 27680 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_10774
timestamp 1668089732
transform 1 0 27680 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_10775
timestamp 1668089732
transform 1 0 27680 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_10776
timestamp 1668089732
transform 1 0 27680 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_10777
timestamp 1668089732
transform 1 0 27680 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_10778
timestamp 1668089732
transform 1 0 27680 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_10779
timestamp 1668089732
transform 1 0 27680 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_10780
timestamp 1668089732
transform 1 0 27680 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_10781
timestamp 1668089732
transform 1 0 27680 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_10782
timestamp 1668089732
transform 1 0 27680 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_10783
timestamp 1668089732
transform 1 0 27680 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_10784
timestamp 1668089732
transform 1 0 27680 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_10785
timestamp 1668089732
transform 1 0 27680 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_10786
timestamp 1668089732
transform 1 0 27680 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_10787
timestamp 1668089732
transform 1 0 27680 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_10788
timestamp 1668089732
transform 1 0 27840 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_10789
timestamp 1668089732
transform 1 0 27840 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_10790
timestamp 1668089732
transform 1 0 27840 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_10791
timestamp 1668089732
transform 1 0 27840 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_10792
timestamp 1668089732
transform 1 0 27840 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_10793
timestamp 1668089732
transform 1 0 27840 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_10794
timestamp 1668089732
transform 1 0 27840 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_10795
timestamp 1668089732
transform 1 0 27840 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_10796
timestamp 1668089732
transform 1 0 27840 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_10797
timestamp 1668089732
transform 1 0 27840 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_10798
timestamp 1668089732
transform 1 0 27840 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_10799
timestamp 1668089732
transform 1 0 27840 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_10800
timestamp 1668089732
transform 1 0 27840 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_10801
timestamp 1668089732
transform 1 0 27840 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_10802
timestamp 1668089732
transform 1 0 27840 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_10803
timestamp 1668089732
transform 1 0 27840 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_10804
timestamp 1668089732
transform 1 0 27840 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_10805
timestamp 1668089732
transform 1 0 27840 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_10806
timestamp 1668089732
transform 1 0 27840 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_10807
timestamp 1668089732
transform 1 0 27840 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_10808
timestamp 1668089732
transform 1 0 27840 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_10809
timestamp 1668089732
transform 1 0 27840 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_10810
timestamp 1668089732
transform 1 0 27840 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_10811
timestamp 1668089732
transform 1 0 27840 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_10812
timestamp 1668089732
transform 1 0 27840 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_10813
timestamp 1668089732
transform 1 0 27840 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_10814
timestamp 1668089732
transform 1 0 27840 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_10815
timestamp 1668089732
transform 1 0 27840 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_10816
timestamp 1668089732
transform 1 0 27840 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_10817
timestamp 1668089732
transform 1 0 27840 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_10818
timestamp 1668089732
transform 1 0 27840 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_10819
timestamp 1668089732
transform 1 0 27840 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_10820
timestamp 1668089732
transform 1 0 27840 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_10821
timestamp 1668089732
transform 1 0 27840 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_10822
timestamp 1668089732
transform 1 0 27840 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_10823
timestamp 1668089732
transform 1 0 27840 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_10824
timestamp 1668089732
transform 1 0 27840 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_10825
timestamp 1668089732
transform 1 0 27840 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_10826
timestamp 1668089732
transform 1 0 27840 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_10827
timestamp 1668089732
transform 1 0 27840 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_10828
timestamp 1668089732
transform 1 0 27840 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_10829
timestamp 1668089732
transform 1 0 27840 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_10830
timestamp 1668089732
transform 1 0 27840 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_10831
timestamp 1668089732
transform 1 0 27840 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_10832
timestamp 1668089732
transform 1 0 27840 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_10833
timestamp 1668089732
transform 1 0 27840 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_10834
timestamp 1668089732
transform 1 0 27840 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_10835
timestamp 1668089732
transform 1 0 27840 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_10836
timestamp 1668089732
transform 1 0 27840 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_10837
timestamp 1668089732
transform 1 0 27840 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_10838
timestamp 1668089732
transform 1 0 27840 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_10839
timestamp 1668089732
transform 1 0 27840 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_10840
timestamp 1668089732
transform 1 0 27840 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_10841
timestamp 1668089732
transform 1 0 27840 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_10842
timestamp 1668089732
transform 1 0 27840 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_10843
timestamp 1668089732
transform 1 0 27840 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_10844
timestamp 1668089732
transform 1 0 27840 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_10845
timestamp 1668089732
transform 1 0 27840 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_10846
timestamp 1668089732
transform 1 0 27840 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_10847
timestamp 1668089732
transform 1 0 27840 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_10848
timestamp 1668089732
transform 1 0 27840 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_10849
timestamp 1668089732
transform 1 0 27840 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_10850
timestamp 1668089732
transform 1 0 28000 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_10851
timestamp 1668089732
transform 1 0 28000 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_10852
timestamp 1668089732
transform 1 0 28000 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_10853
timestamp 1668089732
transform 1 0 28000 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_10854
timestamp 1668089732
transform 1 0 28000 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_10855
timestamp 1668089732
transform 1 0 28000 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_10856
timestamp 1668089732
transform 1 0 28000 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_10857
timestamp 1668089732
transform 1 0 28000 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_10858
timestamp 1668089732
transform 1 0 28000 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_10859
timestamp 1668089732
transform 1 0 28000 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_10860
timestamp 1668089732
transform 1 0 28000 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_10861
timestamp 1668089732
transform 1 0 28000 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_10862
timestamp 1668089732
transform 1 0 28000 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_10863
timestamp 1668089732
transform 1 0 28000 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_10864
timestamp 1668089732
transform 1 0 28000 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_10865
timestamp 1668089732
transform 1 0 28000 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_10866
timestamp 1668089732
transform 1 0 28000 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_10867
timestamp 1668089732
transform 1 0 28000 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_10868
timestamp 1668089732
transform 1 0 28000 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_10869
timestamp 1668089732
transform 1 0 28000 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_10870
timestamp 1668089732
transform 1 0 28000 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_10871
timestamp 1668089732
transform 1 0 28000 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_10872
timestamp 1668089732
transform 1 0 28000 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_10873
timestamp 1668089732
transform 1 0 28000 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_10874
timestamp 1668089732
transform 1 0 28000 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_10875
timestamp 1668089732
transform 1 0 28000 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_10876
timestamp 1668089732
transform 1 0 28000 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_10877
timestamp 1668089732
transform 1 0 28000 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_10878
timestamp 1668089732
transform 1 0 28000 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_10879
timestamp 1668089732
transform 1 0 28000 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_10880
timestamp 1668089732
transform 1 0 28000 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_10881
timestamp 1668089732
transform 1 0 28000 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_10882
timestamp 1668089732
transform 1 0 28000 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_10883
timestamp 1668089732
transform 1 0 28000 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_10884
timestamp 1668089732
transform 1 0 28000 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_10885
timestamp 1668089732
transform 1 0 28000 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_10886
timestamp 1668089732
transform 1 0 28000 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_10887
timestamp 1668089732
transform 1 0 28000 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_10888
timestamp 1668089732
transform 1 0 28000 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_10889
timestamp 1668089732
transform 1 0 28000 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_10890
timestamp 1668089732
transform 1 0 28000 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_10891
timestamp 1668089732
transform 1 0 28000 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_10892
timestamp 1668089732
transform 1 0 28000 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_10893
timestamp 1668089732
transform 1 0 28000 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_10894
timestamp 1668089732
transform 1 0 28000 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_10895
timestamp 1668089732
transform 1 0 28000 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_10896
timestamp 1668089732
transform 1 0 28000 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_10897
timestamp 1668089732
transform 1 0 28000 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_10898
timestamp 1668089732
transform 1 0 28000 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_10899
timestamp 1668089732
transform 1 0 28000 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_10900
timestamp 1668089732
transform 1 0 28000 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_10901
timestamp 1668089732
transform 1 0 28000 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_10902
timestamp 1668089732
transform 1 0 28000 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_10903
timestamp 1668089732
transform 1 0 28000 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_10904
timestamp 1668089732
transform 1 0 28000 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_10905
timestamp 1668089732
transform 1 0 28000 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_10906
timestamp 1668089732
transform 1 0 28000 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_10907
timestamp 1668089732
transform 1 0 28000 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_10908
timestamp 1668089732
transform 1 0 28000 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_10909
timestamp 1668089732
transform 1 0 28000 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_10910
timestamp 1668089732
transform 1 0 28000 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_10911
timestamp 1668089732
transform 1 0 28000 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_10912
timestamp 1668089732
transform 1 0 28160 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_10913
timestamp 1668089732
transform 1 0 28160 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_10914
timestamp 1668089732
transform 1 0 28160 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_10915
timestamp 1668089732
transform 1 0 28160 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_10916
timestamp 1668089732
transform 1 0 28160 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_10917
timestamp 1668089732
transform 1 0 28160 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_10918
timestamp 1668089732
transform 1 0 28160 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_10919
timestamp 1668089732
transform 1 0 28160 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_10920
timestamp 1668089732
transform 1 0 28160 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_10921
timestamp 1668089732
transform 1 0 28160 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_10922
timestamp 1668089732
transform 1 0 28160 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_10923
timestamp 1668089732
transform 1 0 28160 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_10924
timestamp 1668089732
transform 1 0 28160 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_10925
timestamp 1668089732
transform 1 0 28160 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_10926
timestamp 1668089732
transform 1 0 28160 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_10927
timestamp 1668089732
transform 1 0 28160 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_10928
timestamp 1668089732
transform 1 0 28160 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_10929
timestamp 1668089732
transform 1 0 28160 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_10930
timestamp 1668089732
transform 1 0 28160 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_10931
timestamp 1668089732
transform 1 0 28160 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_10932
timestamp 1668089732
transform 1 0 28160 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_10933
timestamp 1668089732
transform 1 0 28160 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_10934
timestamp 1668089732
transform 1 0 28160 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_10935
timestamp 1668089732
transform 1 0 28160 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_10936
timestamp 1668089732
transform 1 0 28160 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_10937
timestamp 1668089732
transform 1 0 28160 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_10938
timestamp 1668089732
transform 1 0 28160 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_10939
timestamp 1668089732
transform 1 0 28160 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_10940
timestamp 1668089732
transform 1 0 28160 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_10941
timestamp 1668089732
transform 1 0 28160 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_10942
timestamp 1668089732
transform 1 0 28160 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_10943
timestamp 1668089732
transform 1 0 28160 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_10944
timestamp 1668089732
transform 1 0 28160 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_10945
timestamp 1668089732
transform 1 0 28160 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_10946
timestamp 1668089732
transform 1 0 28160 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_10947
timestamp 1668089732
transform 1 0 28160 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_10948
timestamp 1668089732
transform 1 0 28160 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_10949
timestamp 1668089732
transform 1 0 28160 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_10950
timestamp 1668089732
transform 1 0 28160 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_10951
timestamp 1668089732
transform 1 0 28160 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_10952
timestamp 1668089732
transform 1 0 28160 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_10953
timestamp 1668089732
transform 1 0 28160 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_10954
timestamp 1668089732
transform 1 0 28160 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_10955
timestamp 1668089732
transform 1 0 28160 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_10956
timestamp 1668089732
transform 1 0 28160 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_10957
timestamp 1668089732
transform 1 0 28160 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_10958
timestamp 1668089732
transform 1 0 28160 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_10959
timestamp 1668089732
transform 1 0 28160 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_10960
timestamp 1668089732
transform 1 0 28160 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_10961
timestamp 1668089732
transform 1 0 28160 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_10962
timestamp 1668089732
transform 1 0 28160 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_10963
timestamp 1668089732
transform 1 0 28160 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_10964
timestamp 1668089732
transform 1 0 28160 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_10965
timestamp 1668089732
transform 1 0 28160 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_10966
timestamp 1668089732
transform 1 0 28160 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_10967
timestamp 1668089732
transform 1 0 28160 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_10968
timestamp 1668089732
transform 1 0 28160 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_10969
timestamp 1668089732
transform 1 0 28160 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_10970
timestamp 1668089732
transform 1 0 28160 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_10971
timestamp 1668089732
transform 1 0 28160 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_10972
timestamp 1668089732
transform 1 0 28160 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_10973
timestamp 1668089732
transform 1 0 28160 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_10974
timestamp 1668089732
transform 1 0 28320 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_10975
timestamp 1668089732
transform 1 0 28320 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_10976
timestamp 1668089732
transform 1 0 28320 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_10977
timestamp 1668089732
transform 1 0 28320 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_10978
timestamp 1668089732
transform 1 0 28320 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_10979
timestamp 1668089732
transform 1 0 28320 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_10980
timestamp 1668089732
transform 1 0 28320 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_10981
timestamp 1668089732
transform 1 0 28320 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_10982
timestamp 1668089732
transform 1 0 28320 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_10983
timestamp 1668089732
transform 1 0 28320 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_10984
timestamp 1668089732
transform 1 0 28320 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_10985
timestamp 1668089732
transform 1 0 28320 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_10986
timestamp 1668089732
transform 1 0 28320 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_10987
timestamp 1668089732
transform 1 0 28320 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_10988
timestamp 1668089732
transform 1 0 28320 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_10989
timestamp 1668089732
transform 1 0 28320 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_10990
timestamp 1668089732
transform 1 0 28320 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_10991
timestamp 1668089732
transform 1 0 28320 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_10992
timestamp 1668089732
transform 1 0 28320 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_10993
timestamp 1668089732
transform 1 0 28320 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_10994
timestamp 1668089732
transform 1 0 28320 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_10995
timestamp 1668089732
transform 1 0 28320 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_10996
timestamp 1668089732
transform 1 0 28320 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_10997
timestamp 1668089732
transform 1 0 28320 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_10998
timestamp 1668089732
transform 1 0 28320 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_10999
timestamp 1668089732
transform 1 0 28320 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_11000
timestamp 1668089732
transform 1 0 28320 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_11001
timestamp 1668089732
transform 1 0 28320 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_11002
timestamp 1668089732
transform 1 0 28320 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_11003
timestamp 1668089732
transform 1 0 28320 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_11004
timestamp 1668089732
transform 1 0 28320 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_11005
timestamp 1668089732
transform 1 0 28320 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_11006
timestamp 1668089732
transform 1 0 28320 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_11007
timestamp 1668089732
transform 1 0 28320 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_11008
timestamp 1668089732
transform 1 0 28320 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_11009
timestamp 1668089732
transform 1 0 28320 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_11010
timestamp 1668089732
transform 1 0 28320 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_11011
timestamp 1668089732
transform 1 0 28320 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_11012
timestamp 1668089732
transform 1 0 28320 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_11013
timestamp 1668089732
transform 1 0 28320 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_11014
timestamp 1668089732
transform 1 0 28320 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_11015
timestamp 1668089732
transform 1 0 28320 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_11016
timestamp 1668089732
transform 1 0 28320 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_11017
timestamp 1668089732
transform 1 0 28320 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_11018
timestamp 1668089732
transform 1 0 28320 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_11019
timestamp 1668089732
transform 1 0 28320 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_11020
timestamp 1668089732
transform 1 0 28320 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_11021
timestamp 1668089732
transform 1 0 28320 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_11022
timestamp 1668089732
transform 1 0 28320 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_11023
timestamp 1668089732
transform 1 0 28320 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_11024
timestamp 1668089732
transform 1 0 28320 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_11025
timestamp 1668089732
transform 1 0 28320 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_11026
timestamp 1668089732
transform 1 0 28320 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_11027
timestamp 1668089732
transform 1 0 28320 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_11028
timestamp 1668089732
transform 1 0 28320 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_11029
timestamp 1668089732
transform 1 0 28320 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_11030
timestamp 1668089732
transform 1 0 28320 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_11031
timestamp 1668089732
transform 1 0 28320 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_11032
timestamp 1668089732
transform 1 0 28320 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_11033
timestamp 1668089732
transform 1 0 28320 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_11034
timestamp 1668089732
transform 1 0 28320 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_11035
timestamp 1668089732
transform 1 0 28320 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_11036
timestamp 1668089732
transform 1 0 28480 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_11037
timestamp 1668089732
transform 1 0 28480 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_11038
timestamp 1668089732
transform 1 0 28480 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_11039
timestamp 1668089732
transform 1 0 28480 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_11040
timestamp 1668089732
transform 1 0 28480 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_11041
timestamp 1668089732
transform 1 0 28480 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_11042
timestamp 1668089732
transform 1 0 28480 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_11043
timestamp 1668089732
transform 1 0 28480 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_11044
timestamp 1668089732
transform 1 0 28480 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_11045
timestamp 1668089732
transform 1 0 28480 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_11046
timestamp 1668089732
transform 1 0 28480 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_11047
timestamp 1668089732
transform 1 0 28480 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_11048
timestamp 1668089732
transform 1 0 28480 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_11049
timestamp 1668089732
transform 1 0 28480 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_11050
timestamp 1668089732
transform 1 0 28480 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_11051
timestamp 1668089732
transform 1 0 28480 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_11052
timestamp 1668089732
transform 1 0 28480 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_11053
timestamp 1668089732
transform 1 0 28480 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_11054
timestamp 1668089732
transform 1 0 28480 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_11055
timestamp 1668089732
transform 1 0 28480 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_11056
timestamp 1668089732
transform 1 0 28480 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_11057
timestamp 1668089732
transform 1 0 28480 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_11058
timestamp 1668089732
transform 1 0 28480 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_11059
timestamp 1668089732
transform 1 0 28480 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_11060
timestamp 1668089732
transform 1 0 28480 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_11061
timestamp 1668089732
transform 1 0 28480 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_11062
timestamp 1668089732
transform 1 0 28480 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_11063
timestamp 1668089732
transform 1 0 28480 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_11064
timestamp 1668089732
transform 1 0 28480 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_11065
timestamp 1668089732
transform 1 0 28480 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_11066
timestamp 1668089732
transform 1 0 28480 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_11067
timestamp 1668089732
transform 1 0 28480 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_11068
timestamp 1668089732
transform 1 0 28480 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_11069
timestamp 1668089732
transform 1 0 28480 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_11070
timestamp 1668089732
transform 1 0 28480 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_11071
timestamp 1668089732
transform 1 0 28480 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_11072
timestamp 1668089732
transform 1 0 28480 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_11073
timestamp 1668089732
transform 1 0 28480 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_11074
timestamp 1668089732
transform 1 0 28480 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_11075
timestamp 1668089732
transform 1 0 28480 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_11076
timestamp 1668089732
transform 1 0 28480 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_11077
timestamp 1668089732
transform 1 0 28480 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_11078
timestamp 1668089732
transform 1 0 28480 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_11079
timestamp 1668089732
transform 1 0 28480 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_11080
timestamp 1668089732
transform 1 0 28480 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_11081
timestamp 1668089732
transform 1 0 28480 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_11082
timestamp 1668089732
transform 1 0 28480 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_11083
timestamp 1668089732
transform 1 0 28480 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_11084
timestamp 1668089732
transform 1 0 28480 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_11085
timestamp 1668089732
transform 1 0 28480 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_11086
timestamp 1668089732
transform 1 0 28480 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_11087
timestamp 1668089732
transform 1 0 28480 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_11088
timestamp 1668089732
transform 1 0 28480 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_11089
timestamp 1668089732
transform 1 0 28480 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_11090
timestamp 1668089732
transform 1 0 28480 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_11091
timestamp 1668089732
transform 1 0 28480 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_11092
timestamp 1668089732
transform 1 0 28480 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_11093
timestamp 1668089732
transform 1 0 28480 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_11094
timestamp 1668089732
transform 1 0 28480 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_11095
timestamp 1668089732
transform 1 0 28480 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_11096
timestamp 1668089732
transform 1 0 28480 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_11097
timestamp 1668089732
transform 1 0 28480 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_11098
timestamp 1668089732
transform 1 0 28640 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_11099
timestamp 1668089732
transform 1 0 28640 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_11100
timestamp 1668089732
transform 1 0 28640 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_11101
timestamp 1668089732
transform 1 0 28640 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_11102
timestamp 1668089732
transform 1 0 28640 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_11103
timestamp 1668089732
transform 1 0 28640 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_11104
timestamp 1668089732
transform 1 0 28640 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_11105
timestamp 1668089732
transform 1 0 28640 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_11106
timestamp 1668089732
transform 1 0 28640 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_11107
timestamp 1668089732
transform 1 0 28640 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_11108
timestamp 1668089732
transform 1 0 28640 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_11109
timestamp 1668089732
transform 1 0 28640 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_11110
timestamp 1668089732
transform 1 0 28640 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_11111
timestamp 1668089732
transform 1 0 28640 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_11112
timestamp 1668089732
transform 1 0 28640 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_11113
timestamp 1668089732
transform 1 0 28640 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_11114
timestamp 1668089732
transform 1 0 28640 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_11115
timestamp 1668089732
transform 1 0 28640 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_11116
timestamp 1668089732
transform 1 0 28640 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_11117
timestamp 1668089732
transform 1 0 28640 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_11118
timestamp 1668089732
transform 1 0 28640 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_11119
timestamp 1668089732
transform 1 0 28640 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_11120
timestamp 1668089732
transform 1 0 28640 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_11121
timestamp 1668089732
transform 1 0 28640 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_11122
timestamp 1668089732
transform 1 0 28640 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_11123
timestamp 1668089732
transform 1 0 28640 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_11124
timestamp 1668089732
transform 1 0 28640 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_11125
timestamp 1668089732
transform 1 0 28640 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_11126
timestamp 1668089732
transform 1 0 28640 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_11127
timestamp 1668089732
transform 1 0 28640 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_11128
timestamp 1668089732
transform 1 0 28640 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_11129
timestamp 1668089732
transform 1 0 28640 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_11130
timestamp 1668089732
transform 1 0 28640 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_11131
timestamp 1668089732
transform 1 0 28640 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_11132
timestamp 1668089732
transform 1 0 28640 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_11133
timestamp 1668089732
transform 1 0 28640 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_11134
timestamp 1668089732
transform 1 0 28640 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_11135
timestamp 1668089732
transform 1 0 28640 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_11136
timestamp 1668089732
transform 1 0 28640 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_11137
timestamp 1668089732
transform 1 0 28640 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_11138
timestamp 1668089732
transform 1 0 28640 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_11139
timestamp 1668089732
transform 1 0 28640 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_11140
timestamp 1668089732
transform 1 0 28640 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_11141
timestamp 1668089732
transform 1 0 28640 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_11142
timestamp 1668089732
transform 1 0 28640 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_11143
timestamp 1668089732
transform 1 0 28640 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_11144
timestamp 1668089732
transform 1 0 28640 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_11145
timestamp 1668089732
transform 1 0 28640 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_11146
timestamp 1668089732
transform 1 0 28640 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_11147
timestamp 1668089732
transform 1 0 28640 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_11148
timestamp 1668089732
transform 1 0 28640 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_11149
timestamp 1668089732
transform 1 0 28640 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_11150
timestamp 1668089732
transform 1 0 28640 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_11151
timestamp 1668089732
transform 1 0 28640 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_11152
timestamp 1668089732
transform 1 0 28640 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_11153
timestamp 1668089732
transform 1 0 28640 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_11154
timestamp 1668089732
transform 1 0 28640 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_11155
timestamp 1668089732
transform 1 0 28640 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_11156
timestamp 1668089732
transform 1 0 28640 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_11157
timestamp 1668089732
transform 1 0 28640 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_11158
timestamp 1668089732
transform 1 0 28640 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_11159
timestamp 1668089732
transform 1 0 28640 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_11160
timestamp 1668089732
transform 1 0 28800 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_11161
timestamp 1668089732
transform 1 0 28800 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_11162
timestamp 1668089732
transform 1 0 28800 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_11163
timestamp 1668089732
transform 1 0 28800 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_11164
timestamp 1668089732
transform 1 0 28800 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_11165
timestamp 1668089732
transform 1 0 28800 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_11166
timestamp 1668089732
transform 1 0 28800 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_11167
timestamp 1668089732
transform 1 0 28800 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_11168
timestamp 1668089732
transform 1 0 28800 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_11169
timestamp 1668089732
transform 1 0 28800 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_11170
timestamp 1668089732
transform 1 0 28800 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_11171
timestamp 1668089732
transform 1 0 28800 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_11172
timestamp 1668089732
transform 1 0 28800 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_11173
timestamp 1668089732
transform 1 0 28800 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_11174
timestamp 1668089732
transform 1 0 28800 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_11175
timestamp 1668089732
transform 1 0 28800 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_11176
timestamp 1668089732
transform 1 0 28800 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_11177
timestamp 1668089732
transform 1 0 28800 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_11178
timestamp 1668089732
transform 1 0 28800 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_11179
timestamp 1668089732
transform 1 0 28800 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_11180
timestamp 1668089732
transform 1 0 28800 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_11181
timestamp 1668089732
transform 1 0 28800 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_11182
timestamp 1668089732
transform 1 0 28800 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_11183
timestamp 1668089732
transform 1 0 28800 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_11184
timestamp 1668089732
transform 1 0 28800 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_11185
timestamp 1668089732
transform 1 0 28800 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_11186
timestamp 1668089732
transform 1 0 28800 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_11187
timestamp 1668089732
transform 1 0 28800 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_11188
timestamp 1668089732
transform 1 0 28800 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_11189
timestamp 1668089732
transform 1 0 28800 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_11190
timestamp 1668089732
transform 1 0 28800 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_11191
timestamp 1668089732
transform 1 0 28800 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_11192
timestamp 1668089732
transform 1 0 28800 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_11193
timestamp 1668089732
transform 1 0 28800 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_11194
timestamp 1668089732
transform 1 0 28800 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_11195
timestamp 1668089732
transform 1 0 28800 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_11196
timestamp 1668089732
transform 1 0 28800 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_11197
timestamp 1668089732
transform 1 0 28800 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_11198
timestamp 1668089732
transform 1 0 28800 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_11199
timestamp 1668089732
transform 1 0 28800 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_11200
timestamp 1668089732
transform 1 0 28800 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_11201
timestamp 1668089732
transform 1 0 28800 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_11202
timestamp 1668089732
transform 1 0 28800 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_11203
timestamp 1668089732
transform 1 0 28800 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_11204
timestamp 1668089732
transform 1 0 28800 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_11205
timestamp 1668089732
transform 1 0 28800 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_11206
timestamp 1668089732
transform 1 0 28800 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_11207
timestamp 1668089732
transform 1 0 28800 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_11208
timestamp 1668089732
transform 1 0 28800 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_11209
timestamp 1668089732
transform 1 0 28800 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_11210
timestamp 1668089732
transform 1 0 28800 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_11211
timestamp 1668089732
transform 1 0 28800 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_11212
timestamp 1668089732
transform 1 0 28800 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_11213
timestamp 1668089732
transform 1 0 28800 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_11214
timestamp 1668089732
transform 1 0 28800 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_11215
timestamp 1668089732
transform 1 0 28800 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_11216
timestamp 1668089732
transform 1 0 28800 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_11217
timestamp 1668089732
transform 1 0 28800 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_11218
timestamp 1668089732
transform 1 0 28800 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_11219
timestamp 1668089732
transform 1 0 28800 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_11220
timestamp 1668089732
transform 1 0 28800 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_11221
timestamp 1668089732
transform 1 0 28800 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_11222
timestamp 1668089732
transform 1 0 28960 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_11223
timestamp 1668089732
transform 1 0 28960 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_11224
timestamp 1668089732
transform 1 0 28960 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_11225
timestamp 1668089732
transform 1 0 28960 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_11226
timestamp 1668089732
transform 1 0 28960 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_11227
timestamp 1668089732
transform 1 0 28960 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_11228
timestamp 1668089732
transform 1 0 28960 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_11229
timestamp 1668089732
transform 1 0 28960 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_11230
timestamp 1668089732
transform 1 0 28960 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_11231
timestamp 1668089732
transform 1 0 28960 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_11232
timestamp 1668089732
transform 1 0 28960 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_11233
timestamp 1668089732
transform 1 0 28960 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_11234
timestamp 1668089732
transform 1 0 28960 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_11235
timestamp 1668089732
transform 1 0 28960 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_11236
timestamp 1668089732
transform 1 0 28960 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_11237
timestamp 1668089732
transform 1 0 28960 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_11238
timestamp 1668089732
transform 1 0 28960 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_11239
timestamp 1668089732
transform 1 0 28960 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_11240
timestamp 1668089732
transform 1 0 28960 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_11241
timestamp 1668089732
transform 1 0 28960 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_11242
timestamp 1668089732
transform 1 0 28960 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_11243
timestamp 1668089732
transform 1 0 28960 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_11244
timestamp 1668089732
transform 1 0 28960 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_11245
timestamp 1668089732
transform 1 0 28960 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_11246
timestamp 1668089732
transform 1 0 28960 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_11247
timestamp 1668089732
transform 1 0 28960 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_11248
timestamp 1668089732
transform 1 0 28960 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_11249
timestamp 1668089732
transform 1 0 28960 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_11250
timestamp 1668089732
transform 1 0 28960 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_11251
timestamp 1668089732
transform 1 0 28960 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_11252
timestamp 1668089732
transform 1 0 28960 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_11253
timestamp 1668089732
transform 1 0 28960 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_11254
timestamp 1668089732
transform 1 0 28960 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_11255
timestamp 1668089732
transform 1 0 28960 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_11256
timestamp 1668089732
transform 1 0 28960 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_11257
timestamp 1668089732
transform 1 0 28960 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_11258
timestamp 1668089732
transform 1 0 28960 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_11259
timestamp 1668089732
transform 1 0 28960 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_11260
timestamp 1668089732
transform 1 0 28960 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_11261
timestamp 1668089732
transform 1 0 28960 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_11262
timestamp 1668089732
transform 1 0 28960 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_11263
timestamp 1668089732
transform 1 0 28960 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_11264
timestamp 1668089732
transform 1 0 28960 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_11265
timestamp 1668089732
transform 1 0 28960 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_11266
timestamp 1668089732
transform 1 0 28960 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_11267
timestamp 1668089732
transform 1 0 28960 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_11268
timestamp 1668089732
transform 1 0 28960 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_11269
timestamp 1668089732
transform 1 0 28960 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_11270
timestamp 1668089732
transform 1 0 28960 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_11271
timestamp 1668089732
transform 1 0 28960 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_11272
timestamp 1668089732
transform 1 0 28960 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_11273
timestamp 1668089732
transform 1 0 28960 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_11274
timestamp 1668089732
transform 1 0 28960 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_11275
timestamp 1668089732
transform 1 0 28960 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_11276
timestamp 1668089732
transform 1 0 28960 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_11277
timestamp 1668089732
transform 1 0 28960 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_11278
timestamp 1668089732
transform 1 0 28960 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_11279
timestamp 1668089732
transform 1 0 28960 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_11280
timestamp 1668089732
transform 1 0 28960 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_11281
timestamp 1668089732
transform 1 0 28960 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_11282
timestamp 1668089732
transform 1 0 28960 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_11283
timestamp 1668089732
transform 1 0 28960 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_11284
timestamp 1668089732
transform 1 0 29120 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_11285
timestamp 1668089732
transform 1 0 29120 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_11286
timestamp 1668089732
transform 1 0 29120 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_11287
timestamp 1668089732
transform 1 0 29120 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_11288
timestamp 1668089732
transform 1 0 29120 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_11289
timestamp 1668089732
transform 1 0 29120 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_11290
timestamp 1668089732
transform 1 0 29120 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_11291
timestamp 1668089732
transform 1 0 29120 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_11292
timestamp 1668089732
transform 1 0 29120 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_11293
timestamp 1668089732
transform 1 0 29120 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_11294
timestamp 1668089732
transform 1 0 29120 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_11295
timestamp 1668089732
transform 1 0 29120 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_11296
timestamp 1668089732
transform 1 0 29120 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_11297
timestamp 1668089732
transform 1 0 29120 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_11298
timestamp 1668089732
transform 1 0 29120 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_11299
timestamp 1668089732
transform 1 0 29120 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_11300
timestamp 1668089732
transform 1 0 29120 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_11301
timestamp 1668089732
transform 1 0 29120 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_11302
timestamp 1668089732
transform 1 0 29120 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_11303
timestamp 1668089732
transform 1 0 29120 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_11304
timestamp 1668089732
transform 1 0 29120 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_11305
timestamp 1668089732
transform 1 0 29120 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_11306
timestamp 1668089732
transform 1 0 29120 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_11307
timestamp 1668089732
transform 1 0 29120 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_11308
timestamp 1668089732
transform 1 0 29120 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_11309
timestamp 1668089732
transform 1 0 29120 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_11310
timestamp 1668089732
transform 1 0 29120 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_11311
timestamp 1668089732
transform 1 0 29120 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_11312
timestamp 1668089732
transform 1 0 29120 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_11313
timestamp 1668089732
transform 1 0 29120 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_11314
timestamp 1668089732
transform 1 0 29120 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_11315
timestamp 1668089732
transform 1 0 29120 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_11316
timestamp 1668089732
transform 1 0 29120 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_11317
timestamp 1668089732
transform 1 0 29120 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_11318
timestamp 1668089732
transform 1 0 29120 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_11319
timestamp 1668089732
transform 1 0 29120 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_11320
timestamp 1668089732
transform 1 0 29120 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_11321
timestamp 1668089732
transform 1 0 29120 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_11322
timestamp 1668089732
transform 1 0 29120 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_11323
timestamp 1668089732
transform 1 0 29120 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_11324
timestamp 1668089732
transform 1 0 29120 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_11325
timestamp 1668089732
transform 1 0 29120 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_11326
timestamp 1668089732
transform 1 0 29120 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_11327
timestamp 1668089732
transform 1 0 29120 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_11328
timestamp 1668089732
transform 1 0 29120 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_11329
timestamp 1668089732
transform 1 0 29120 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_11330
timestamp 1668089732
transform 1 0 29120 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_11331
timestamp 1668089732
transform 1 0 29120 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_11332
timestamp 1668089732
transform 1 0 29120 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_11333
timestamp 1668089732
transform 1 0 29120 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_11334
timestamp 1668089732
transform 1 0 29120 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_11335
timestamp 1668089732
transform 1 0 29120 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_11336
timestamp 1668089732
transform 1 0 29120 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_11337
timestamp 1668089732
transform 1 0 29120 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_11338
timestamp 1668089732
transform 1 0 29120 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_11339
timestamp 1668089732
transform 1 0 29120 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_11340
timestamp 1668089732
transform 1 0 29120 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_11341
timestamp 1668089732
transform 1 0 29120 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_11342
timestamp 1668089732
transform 1 0 29120 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_11343
timestamp 1668089732
transform 1 0 29120 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_11344
timestamp 1668089732
transform 1 0 29120 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_11345
timestamp 1668089732
transform 1 0 29120 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_11346
timestamp 1668089732
transform 1 0 29280 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_11347
timestamp 1668089732
transform 1 0 29280 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_11348
timestamp 1668089732
transform 1 0 29280 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_11349
timestamp 1668089732
transform 1 0 29280 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_11350
timestamp 1668089732
transform 1 0 29280 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_11351
timestamp 1668089732
transform 1 0 29280 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_11352
timestamp 1668089732
transform 1 0 29280 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_11353
timestamp 1668089732
transform 1 0 29280 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_11354
timestamp 1668089732
transform 1 0 29280 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_11355
timestamp 1668089732
transform 1 0 29280 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_11356
timestamp 1668089732
transform 1 0 29280 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_11357
timestamp 1668089732
transform 1 0 29280 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_11358
timestamp 1668089732
transform 1 0 29280 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_11359
timestamp 1668089732
transform 1 0 29280 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_11360
timestamp 1668089732
transform 1 0 29280 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_11361
timestamp 1668089732
transform 1 0 29280 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_11362
timestamp 1668089732
transform 1 0 29280 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_11363
timestamp 1668089732
transform 1 0 29280 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_11364
timestamp 1668089732
transform 1 0 29280 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_11365
timestamp 1668089732
transform 1 0 29280 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_11366
timestamp 1668089732
transform 1 0 29280 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_11367
timestamp 1668089732
transform 1 0 29280 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_11368
timestamp 1668089732
transform 1 0 29280 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_11369
timestamp 1668089732
transform 1 0 29280 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_11370
timestamp 1668089732
transform 1 0 29280 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_11371
timestamp 1668089732
transform 1 0 29280 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_11372
timestamp 1668089732
transform 1 0 29280 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_11373
timestamp 1668089732
transform 1 0 29280 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_11374
timestamp 1668089732
transform 1 0 29280 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_11375
timestamp 1668089732
transform 1 0 29280 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_11376
timestamp 1668089732
transform 1 0 29280 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_11377
timestamp 1668089732
transform 1 0 29280 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_11378
timestamp 1668089732
transform 1 0 29280 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_11379
timestamp 1668089732
transform 1 0 29280 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_11380
timestamp 1668089732
transform 1 0 29280 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_11381
timestamp 1668089732
transform 1 0 29280 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_11382
timestamp 1668089732
transform 1 0 29280 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_11383
timestamp 1668089732
transform 1 0 29280 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_11384
timestamp 1668089732
transform 1 0 29280 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_11385
timestamp 1668089732
transform 1 0 29280 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_11386
timestamp 1668089732
transform 1 0 29280 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_11387
timestamp 1668089732
transform 1 0 29280 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_11388
timestamp 1668089732
transform 1 0 29280 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_11389
timestamp 1668089732
transform 1 0 29280 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_11390
timestamp 1668089732
transform 1 0 29280 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_11391
timestamp 1668089732
transform 1 0 29280 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_11392
timestamp 1668089732
transform 1 0 29280 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_11393
timestamp 1668089732
transform 1 0 29280 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_11394
timestamp 1668089732
transform 1 0 29280 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_11395
timestamp 1668089732
transform 1 0 29280 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_11396
timestamp 1668089732
transform 1 0 29280 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_11397
timestamp 1668089732
transform 1 0 29280 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_11398
timestamp 1668089732
transform 1 0 29280 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_11399
timestamp 1668089732
transform 1 0 29280 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_11400
timestamp 1668089732
transform 1 0 29280 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_11401
timestamp 1668089732
transform 1 0 29280 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_11402
timestamp 1668089732
transform 1 0 29280 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_11403
timestamp 1668089732
transform 1 0 29280 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_11404
timestamp 1668089732
transform 1 0 29280 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_11405
timestamp 1668089732
transform 1 0 29280 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_11406
timestamp 1668089732
transform 1 0 29280 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_11407
timestamp 1668089732
transform 1 0 29280 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_11408
timestamp 1668089732
transform 1 0 29440 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_11409
timestamp 1668089732
transform 1 0 29440 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_11410
timestamp 1668089732
transform 1 0 29440 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_11411
timestamp 1668089732
transform 1 0 29440 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_11412
timestamp 1668089732
transform 1 0 29440 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_11413
timestamp 1668089732
transform 1 0 29440 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_11414
timestamp 1668089732
transform 1 0 29440 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_11415
timestamp 1668089732
transform 1 0 29440 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_11416
timestamp 1668089732
transform 1 0 29440 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_11417
timestamp 1668089732
transform 1 0 29440 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_11418
timestamp 1668089732
transform 1 0 29440 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_11419
timestamp 1668089732
transform 1 0 29440 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_11420
timestamp 1668089732
transform 1 0 29440 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_11421
timestamp 1668089732
transform 1 0 29440 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_11422
timestamp 1668089732
transform 1 0 29440 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_11423
timestamp 1668089732
transform 1 0 29440 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_11424
timestamp 1668089732
transform 1 0 29440 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_11425
timestamp 1668089732
transform 1 0 29440 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_11426
timestamp 1668089732
transform 1 0 29440 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_11427
timestamp 1668089732
transform 1 0 29440 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_11428
timestamp 1668089732
transform 1 0 29440 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_11429
timestamp 1668089732
transform 1 0 29440 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_11430
timestamp 1668089732
transform 1 0 29440 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_11431
timestamp 1668089732
transform 1 0 29440 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_11432
timestamp 1668089732
transform 1 0 29440 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_11433
timestamp 1668089732
transform 1 0 29440 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_11434
timestamp 1668089732
transform 1 0 29440 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_11435
timestamp 1668089732
transform 1 0 29440 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_11436
timestamp 1668089732
transform 1 0 29440 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_11437
timestamp 1668089732
transform 1 0 29440 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_11438
timestamp 1668089732
transform 1 0 29440 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_11439
timestamp 1668089732
transform 1 0 29440 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_11440
timestamp 1668089732
transform 1 0 29440 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_11441
timestamp 1668089732
transform 1 0 29440 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_11442
timestamp 1668089732
transform 1 0 29440 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_11443
timestamp 1668089732
transform 1 0 29440 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_11444
timestamp 1668089732
transform 1 0 29440 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_11445
timestamp 1668089732
transform 1 0 29440 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_11446
timestamp 1668089732
transform 1 0 29440 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_11447
timestamp 1668089732
transform 1 0 29440 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_11448
timestamp 1668089732
transform 1 0 29440 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_11449
timestamp 1668089732
transform 1 0 29440 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_11450
timestamp 1668089732
transform 1 0 29440 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_11451
timestamp 1668089732
transform 1 0 29440 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_11452
timestamp 1668089732
transform 1 0 29440 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_11453
timestamp 1668089732
transform 1 0 29440 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_11454
timestamp 1668089732
transform 1 0 29440 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_11455
timestamp 1668089732
transform 1 0 29440 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_11456
timestamp 1668089732
transform 1 0 29440 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_11457
timestamp 1668089732
transform 1 0 29440 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_11458
timestamp 1668089732
transform 1 0 29440 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_11459
timestamp 1668089732
transform 1 0 29440 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_11460
timestamp 1668089732
transform 1 0 29440 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_11461
timestamp 1668089732
transform 1 0 29440 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_11462
timestamp 1668089732
transform 1 0 29440 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_11463
timestamp 1668089732
transform 1 0 29440 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_11464
timestamp 1668089732
transform 1 0 29440 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_11465
timestamp 1668089732
transform 1 0 29440 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_11466
timestamp 1668089732
transform 1 0 29440 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_11467
timestamp 1668089732
transform 1 0 29440 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_11468
timestamp 1668089732
transform 1 0 29440 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_11469
timestamp 1668089732
transform 1 0 29440 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_11470
timestamp 1668089732
transform 1 0 29600 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_11471
timestamp 1668089732
transform 1 0 29600 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_11472
timestamp 1668089732
transform 1 0 29600 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_11473
timestamp 1668089732
transform 1 0 29600 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_11474
timestamp 1668089732
transform 1 0 29600 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_11475
timestamp 1668089732
transform 1 0 29600 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_11476
timestamp 1668089732
transform 1 0 29600 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_11477
timestamp 1668089732
transform 1 0 29600 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_11478
timestamp 1668089732
transform 1 0 29600 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_11479
timestamp 1668089732
transform 1 0 29600 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_11480
timestamp 1668089732
transform 1 0 29600 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_11481
timestamp 1668089732
transform 1 0 29600 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_11482
timestamp 1668089732
transform 1 0 29600 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_11483
timestamp 1668089732
transform 1 0 29600 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_11484
timestamp 1668089732
transform 1 0 29600 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_11485
timestamp 1668089732
transform 1 0 29600 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_11486
timestamp 1668089732
transform 1 0 29600 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_11487
timestamp 1668089732
transform 1 0 29600 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_11488
timestamp 1668089732
transform 1 0 29600 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_11489
timestamp 1668089732
transform 1 0 29600 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_11490
timestamp 1668089732
transform 1 0 29600 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_11491
timestamp 1668089732
transform 1 0 29600 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_11492
timestamp 1668089732
transform 1 0 29600 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_11493
timestamp 1668089732
transform 1 0 29600 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_11494
timestamp 1668089732
transform 1 0 29600 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_11495
timestamp 1668089732
transform 1 0 29600 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_11496
timestamp 1668089732
transform 1 0 29600 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_11497
timestamp 1668089732
transform 1 0 29600 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_11498
timestamp 1668089732
transform 1 0 29600 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_11499
timestamp 1668089732
transform 1 0 29600 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_11500
timestamp 1668089732
transform 1 0 29600 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_11501
timestamp 1668089732
transform 1 0 29600 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_11502
timestamp 1668089732
transform 1 0 29600 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_11503
timestamp 1668089732
transform 1 0 29600 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_11504
timestamp 1668089732
transform 1 0 29600 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_11505
timestamp 1668089732
transform 1 0 29600 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_11506
timestamp 1668089732
transform 1 0 29600 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_11507
timestamp 1668089732
transform 1 0 29600 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_11508
timestamp 1668089732
transform 1 0 29600 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_11509
timestamp 1668089732
transform 1 0 29600 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_11510
timestamp 1668089732
transform 1 0 29600 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_11511
timestamp 1668089732
transform 1 0 29600 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_11512
timestamp 1668089732
transform 1 0 29600 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_11513
timestamp 1668089732
transform 1 0 29600 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_11514
timestamp 1668089732
transform 1 0 29600 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_11515
timestamp 1668089732
transform 1 0 29600 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_11516
timestamp 1668089732
transform 1 0 29600 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_11517
timestamp 1668089732
transform 1 0 29600 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_11518
timestamp 1668089732
transform 1 0 29600 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_11519
timestamp 1668089732
transform 1 0 29600 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_11520
timestamp 1668089732
transform 1 0 29600 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_11521
timestamp 1668089732
transform 1 0 29600 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_11522
timestamp 1668089732
transform 1 0 29600 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_11523
timestamp 1668089732
transform 1 0 29600 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_11524
timestamp 1668089732
transform 1 0 29600 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_11525
timestamp 1668089732
transform 1 0 29600 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_11526
timestamp 1668089732
transform 1 0 29600 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_11527
timestamp 1668089732
transform 1 0 29600 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_11528
timestamp 1668089732
transform 1 0 29600 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_11529
timestamp 1668089732
transform 1 0 29600 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_11530
timestamp 1668089732
transform 1 0 29600 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_11531
timestamp 1668089732
transform 1 0 29600 0 1 9760
box 0 0 200 200
use unit_pad  unit_pad_11532
timestamp 1668089732
transform 1 0 29760 0 1 0
box 0 0 200 200
use unit_pad  unit_pad_11533
timestamp 1668089732
transform 1 0 29760 0 1 160
box 0 0 200 200
use unit_pad  unit_pad_11534
timestamp 1668089732
transform 1 0 29760 0 1 320
box 0 0 200 200
use unit_pad  unit_pad_11535
timestamp 1668089732
transform 1 0 29760 0 1 480
box 0 0 200 200
use unit_pad  unit_pad_11536
timestamp 1668089732
transform 1 0 29760 0 1 640
box 0 0 200 200
use unit_pad  unit_pad_11537
timestamp 1668089732
transform 1 0 29760 0 1 800
box 0 0 200 200
use unit_pad  unit_pad_11538
timestamp 1668089732
transform 1 0 29760 0 1 960
box 0 0 200 200
use unit_pad  unit_pad_11539
timestamp 1668089732
transform 1 0 29760 0 1 1120
box 0 0 200 200
use unit_pad  unit_pad_11540
timestamp 1668089732
transform 1 0 29760 0 1 1280
box 0 0 200 200
use unit_pad  unit_pad_11541
timestamp 1668089732
transform 1 0 29760 0 1 1440
box 0 0 200 200
use unit_pad  unit_pad_11542
timestamp 1668089732
transform 1 0 29760 0 1 1600
box 0 0 200 200
use unit_pad  unit_pad_11543
timestamp 1668089732
transform 1 0 29760 0 1 1760
box 0 0 200 200
use unit_pad  unit_pad_11544
timestamp 1668089732
transform 1 0 29760 0 1 1920
box 0 0 200 200
use unit_pad  unit_pad_11545
timestamp 1668089732
transform 1 0 29760 0 1 2080
box 0 0 200 200
use unit_pad  unit_pad_11546
timestamp 1668089732
transform 1 0 29760 0 1 2240
box 0 0 200 200
use unit_pad  unit_pad_11547
timestamp 1668089732
transform 1 0 29760 0 1 2400
box 0 0 200 200
use unit_pad  unit_pad_11548
timestamp 1668089732
transform 1 0 29760 0 1 2560
box 0 0 200 200
use unit_pad  unit_pad_11549
timestamp 1668089732
transform 1 0 29760 0 1 2720
box 0 0 200 200
use unit_pad  unit_pad_11550
timestamp 1668089732
transform 1 0 29760 0 1 2880
box 0 0 200 200
use unit_pad  unit_pad_11551
timestamp 1668089732
transform 1 0 29760 0 1 3040
box 0 0 200 200
use unit_pad  unit_pad_11552
timestamp 1668089732
transform 1 0 29760 0 1 3200
box 0 0 200 200
use unit_pad  unit_pad_11553
timestamp 1668089732
transform 1 0 29760 0 1 3360
box 0 0 200 200
use unit_pad  unit_pad_11554
timestamp 1668089732
transform 1 0 29760 0 1 3520
box 0 0 200 200
use unit_pad  unit_pad_11555
timestamp 1668089732
transform 1 0 29760 0 1 3680
box 0 0 200 200
use unit_pad  unit_pad_11556
timestamp 1668089732
transform 1 0 29760 0 1 3840
box 0 0 200 200
use unit_pad  unit_pad_11557
timestamp 1668089732
transform 1 0 29760 0 1 4000
box 0 0 200 200
use unit_pad  unit_pad_11558
timestamp 1668089732
transform 1 0 29760 0 1 4160
box 0 0 200 200
use unit_pad  unit_pad_11559
timestamp 1668089732
transform 1 0 29760 0 1 4320
box 0 0 200 200
use unit_pad  unit_pad_11560
timestamp 1668089732
transform 1 0 29760 0 1 4480
box 0 0 200 200
use unit_pad  unit_pad_11561
timestamp 1668089732
transform 1 0 29760 0 1 4640
box 0 0 200 200
use unit_pad  unit_pad_11562
timestamp 1668089732
transform 1 0 29760 0 1 4800
box 0 0 200 200
use unit_pad  unit_pad_11563
timestamp 1668089732
transform 1 0 29760 0 1 4960
box 0 0 200 200
use unit_pad  unit_pad_11564
timestamp 1668089732
transform 1 0 29760 0 1 5120
box 0 0 200 200
use unit_pad  unit_pad_11565
timestamp 1668089732
transform 1 0 29760 0 1 5280
box 0 0 200 200
use unit_pad  unit_pad_11566
timestamp 1668089732
transform 1 0 29760 0 1 5440
box 0 0 200 200
use unit_pad  unit_pad_11567
timestamp 1668089732
transform 1 0 29760 0 1 5600
box 0 0 200 200
use unit_pad  unit_pad_11568
timestamp 1668089732
transform 1 0 29760 0 1 5760
box 0 0 200 200
use unit_pad  unit_pad_11569
timestamp 1668089732
transform 1 0 29760 0 1 5920
box 0 0 200 200
use unit_pad  unit_pad_11570
timestamp 1668089732
transform 1 0 29760 0 1 6080
box 0 0 200 200
use unit_pad  unit_pad_11571
timestamp 1668089732
transform 1 0 29760 0 1 6240
box 0 0 200 200
use unit_pad  unit_pad_11572
timestamp 1668089732
transform 1 0 29760 0 1 6400
box 0 0 200 200
use unit_pad  unit_pad_11573
timestamp 1668089732
transform 1 0 29760 0 1 6560
box 0 0 200 200
use unit_pad  unit_pad_11574
timestamp 1668089732
transform 1 0 29760 0 1 6720
box 0 0 200 200
use unit_pad  unit_pad_11575
timestamp 1668089732
transform 1 0 29760 0 1 6880
box 0 0 200 200
use unit_pad  unit_pad_11576
timestamp 1668089732
transform 1 0 29760 0 1 7040
box 0 0 200 200
use unit_pad  unit_pad_11577
timestamp 1668089732
transform 1 0 29760 0 1 7200
box 0 0 200 200
use unit_pad  unit_pad_11578
timestamp 1668089732
transform 1 0 29760 0 1 7360
box 0 0 200 200
use unit_pad  unit_pad_11579
timestamp 1668089732
transform 1 0 29760 0 1 7520
box 0 0 200 200
use unit_pad  unit_pad_11580
timestamp 1668089732
transform 1 0 29760 0 1 7680
box 0 0 200 200
use unit_pad  unit_pad_11581
timestamp 1668089732
transform 1 0 29760 0 1 7840
box 0 0 200 200
use unit_pad  unit_pad_11582
timestamp 1668089732
transform 1 0 29760 0 1 8000
box 0 0 200 200
use unit_pad  unit_pad_11583
timestamp 1668089732
transform 1 0 29760 0 1 8160
box 0 0 200 200
use unit_pad  unit_pad_11584
timestamp 1668089732
transform 1 0 29760 0 1 8320
box 0 0 200 200
use unit_pad  unit_pad_11585
timestamp 1668089732
transform 1 0 29760 0 1 8480
box 0 0 200 200
use unit_pad  unit_pad_11586
timestamp 1668089732
transform 1 0 29760 0 1 8640
box 0 0 200 200
use unit_pad  unit_pad_11587
timestamp 1668089732
transform 1 0 29760 0 1 8800
box 0 0 200 200
use unit_pad  unit_pad_11588
timestamp 1668089732
transform 1 0 29760 0 1 8960
box 0 0 200 200
use unit_pad  unit_pad_11589
timestamp 1668089732
transform 1 0 29760 0 1 9120
box 0 0 200 200
use unit_pad  unit_pad_11590
timestamp 1668089732
transform 1 0 29760 0 1 9280
box 0 0 200 200
use unit_pad  unit_pad_11591
timestamp 1668089732
transform 1 0 29760 0 1 9440
box 0 0 200 200
use unit_pad  unit_pad_11592
timestamp 1668089732
transform 1 0 29760 0 1 9600
box 0 0 200 200
use unit_pad  unit_pad_11593
timestamp 1668089732
transform 1 0 29760 0 1 9760
box 0 0 200 200
<< end >>
