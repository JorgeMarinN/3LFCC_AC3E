magic
tech sky130A
timestamp 1666629273
<< error_p >>
rect 48350 45532 48361 48361
rect 54857 45532 54868 52039
rect 48350 45521 54868 45532
<< metal4 >>
rect 48349 52039 54869 52040
rect 48349 45521 48350 52039
rect 54868 45521 54869 52039
rect 48349 18479 54869 45521
<< via4 >>
rect 48350 45521 54868 52039
<< metal5 >>
rect 25000 68869 75389 75389
rect 25000 62029 68549 68549
rect 25000 31520 31520 62029
rect 31840 55189 61709 61709
rect 31840 38360 38360 55189
rect 38680 52039 54869 54869
rect 38680 48349 48350 52039
rect 38680 45200 45200 48349
rect 48349 45521 48350 48349
rect 54868 45521 54869 52039
rect 48349 45520 54869 45521
rect 55189 45200 61709 55189
rect 38680 38680 61709 45200
rect 62029 38360 68549 62029
rect 31840 31840 68549 38360
rect 68869 31520 75389 68869
rect 25000 25000 75389 31520
<< end >>
