magic
tech sky130A
timestamp 1668199884
<< error_p >>
rect 25 550 75 557
rect 2 112 4 538
rect 265 373 385 385
rect 265 277 277 373
rect 373 277 385 373
rect 265 265 385 277
rect 550 25 557 75
rect 0 2 2 17
rect 112 2 538 4
rect 0 0 17 2
<< dnwell >>
rect 0 0 550 550
<< pwell >>
rect 0 0 550 550
<< mvnmos >>
rect 25 106 75 544
rect 106 25 544 75
<< mvndiff >>
rect 106 546 544 550
rect 104 544 546 546
rect 0 538 25 544
rect 0 112 2 538
rect 19 112 25 538
rect 0 106 25 112
rect 75 538 550 544
rect 75 112 81 538
rect 98 490 550 538
rect 98 160 160 490
rect 490 160 550 490
rect 98 112 550 160
rect 75 106 550 112
rect 104 104 546 106
rect 106 98 544 104
rect 106 81 112 98
rect 538 81 544 98
rect 106 75 544 81
rect 106 19 544 25
rect 106 2 112 19
rect 538 2 544 19
rect 106 0 544 2
<< mvndiffc >>
rect 2 112 19 538
rect 81 112 98 538
rect 112 81 538 98
rect 112 2 538 19
<< mvpsubdiff >>
rect 160 478 490 490
rect 160 172 172 478
rect 478 172 490 478
rect 160 160 490 172
<< mvpsubdiffcont >>
rect 172 172 478 478
<< poly >>
rect 25 544 75 550
rect 25 75 75 106
rect 0 67 106 75
rect 0 33 33 67
rect 67 33 106 67
rect 0 25 106 33
rect 544 25 550 75
rect 25 0 75 25
<< polycont >>
rect 33 33 67 67
<< locali >>
rect 98 546 550 550
rect 0 538 19 546
rect 0 511 2 538
rect 0 112 2 139
rect 0 104 19 112
rect 81 538 550 546
rect 98 490 550 538
rect 98 160 160 490
rect 490 160 550 490
rect 98 112 550 160
rect 81 104 550 112
rect 98 98 550 104
rect 104 81 112 98
rect 538 81 546 98
rect 25 67 75 75
rect 25 33 33 67
rect 67 33 75 67
rect 25 25 75 33
rect 104 2 112 19
rect 538 2 546 19
rect 0 0 2 2
rect 104 0 139 2
rect 511 0 546 2
<< viali >>
rect 2 112 19 538
rect 81 112 98 538
rect 160 478 490 490
rect 160 172 172 478
rect 172 172 478 478
rect 478 172 490 478
rect 160 160 490 172
rect 112 81 538 98
rect 33 33 67 67
rect 112 2 538 19
<< metal1 >>
rect 106 549 544 550
rect 101 544 549 549
rect 0 538 22 544
rect 0 112 2 538
rect 19 112 22 538
rect 0 106 22 112
rect 78 538 550 544
rect 78 112 81 538
rect 98 490 550 538
rect 98 160 160 490
rect 490 160 550 490
rect 98 112 550 160
rect 78 106 550 112
rect 101 101 549 106
rect 106 98 544 101
rect 106 81 112 98
rect 538 81 544 98
rect 106 78 544 81
rect 25 67 75 75
rect 25 33 33 67
rect 67 33 75 67
rect 25 25 75 33
rect 106 19 544 22
rect 106 2 112 19
rect 538 2 544 19
rect 106 0 544 2
<< via1 >>
rect 160 160 490 490
rect 33 33 67 67
<< metal2 >>
rect 25 75 75 550
rect 150 490 500 500
rect 150 160 160 490
rect 490 160 500 490
rect 150 150 500 160
rect 0 67 550 75
rect 0 33 33 67
rect 67 33 550 67
rect 0 25 550 33
rect 25 0 75 25
<< via2 >>
rect 265 265 385 385
<< via3 >>
rect 265 265 385 385
<< via4 >>
rect 265 265 385 385
<< properties >>
string MASKHINTS_HVI 0 0 300 300
string MASKHINTS_HVNTM 0 0 300 300
<< end >>
