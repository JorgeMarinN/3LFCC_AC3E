magic
tech sky130A
timestamp 1661199807
<< checkpaint >>
rect 170 61370 38630 137830
rect 6770 -630 38630 61370
<< metal2 >>
rect 4000 131460 6000 132000
rect 4000 131270 5760 131460
rect 4000 130400 6000 131270
rect 4000 66960 6540 67200
rect 6730 66960 7600 67200
rect 4000 65600 7600 66960
rect 10000 56640 14200 58000
rect 10000 56400 13140 56640
rect 13330 56400 14200 56640
rect 10000 5925 12700 6800
rect 10000 5749 12362 5925
rect 10000 5200 12700 5749
<< metal3 >>
rect 7000 133000 38000 136000
rect 4200 131000 5200 131039
rect 2000 130100 5200 131000
rect 2000 104000 5000 130100
rect 34000 106000 38000 133000
rect 2000 95000 32000 104000
rect 2000 68000 5000 95000
rect 6961 66000 7900 66400
rect 34000 66000 38000 93000
rect 6961 65400 38000 66000
rect 7000 63000 38000 65400
rect 14000 58200 38000 63000
rect 13561 58000 38000 58200
rect 13561 57200 14500 58000
rect 8000 35000 11000 56000
rect 34000 37000 38000 58000
rect 8000 27000 32000 35000
rect 8000 7100 11000 27000
rect 8000 7000 11800 7100
rect 10800 6161 11800 7000
rect 34000 4000 38000 25000
rect 13000 1000 38000 4000
<< metal4 >>
rect 7000 133000 38000 136000
rect 4200 131000 5200 131039
rect 2000 130100 5200 131000
rect 2000 104000 5000 130100
rect 34000 106000 38000 133000
rect 2000 95000 32000 104000
rect 2000 68000 5000 95000
rect 6961 66000 7900 66400
rect 34000 66000 38000 93000
rect 6961 65400 38000 66000
rect 7000 63000 38000 65400
rect 14000 58200 38000 63000
rect 13561 58000 38000 58200
rect 13561 57200 14500 58000
rect 8000 35000 11000 56000
rect 34000 37000 38000 58000
rect 8000 27000 32000 35000
rect 8000 7100 11000 27000
rect 8000 7000 11800 7100
rect 10800 6161 11800 7000
rect 34000 4000 38000 25000
rect 13000 1000 38000 4000
<< metal5 >>
rect 7000 133000 38000 136000
rect 4200 131000 5200 131039
rect 2000 130100 5200 131000
rect 2000 104000 5000 130100
rect 34000 106000 38000 133000
rect 2000 95000 32000 104000
rect 2000 68000 5000 95000
rect 6961 66000 7900 66400
rect 34000 66000 38000 93000
rect 6961 65400 38000 66000
rect 7000 63000 38000 65400
rect 14000 58200 38000 63000
rect 13561 58000 38000 58200
rect 13561 57200 14500 58000
rect 8000 35000 11000 56000
rect 34000 37000 38000 58000
rect 8000 27000 32000 35000
rect 8000 7100 11000 27000
rect 8000 7000 11800 7100
rect 10800 6161 11800 7000
rect 34000 4000 38000 25000
rect 13000 1000 38000 4000
use nmos_waffle_36x36  nmos_waffle_36x36_0
timestamp 1624430562
transform 1 0 12800 0 1 5400
box -5400 -5400 25200 25200
use nmos_waffle_36x36  nmos_waffle_36x36_1
timestamp 1624430562
transform 0 1 12800 -1 0 56200
box -5400 -5400 25200 25200
use pmos_waffle_48x48  pmos_waffle_48x48_0
timestamp 1624430562
transform 0 1 6200 1 0 67400
box -5400 -5400 31800 31800
use pmos_waffle_48x48  pmos_waffle_48x48_1
timestamp 1624430562
transform 1 0 6200 0 -1 131800
box -5400 -5400 31800 31800
<< labels >>
rlabel metal2 4168 131219 4797 131806 1 S1
rlabel metal2 4225 66197 4854 66784 1 S2
rlabel metal2 10261 57177 10890 57764 1 S3
rlabel metal2 10064 5384 10693 5971 1 S4
rlabel metal5 13240 2292 13869 2879 1 Vss
rlabel metal5 8350 30451 8979 31038 1 fc2
rlabel metal5 37352 61196 37981 61783 1 Vout
rlabel metal5 7310 134235 7939 134822 1 Vdd
rlabel metal5 2366 99271 2995 99858 1 fc1
<< end >>
