magic
tech sky130A
timestamp 1666025761
<< metal1 >>
rect 2000 169795 2500 169800
rect 2000 169305 2005 169795
rect 2495 169305 2500 169795
rect 2000 166800 2500 169305
rect 136500 169795 137000 169800
rect 136500 169305 136505 169795
rect 136995 169305 137000 169795
rect 2000 166600 136400 166800
rect 136500 166550 137000 169305
rect 2000 166545 137000 166550
rect 2000 166355 6345 166545
rect 6435 166355 71345 166545
rect 71435 166355 80345 166545
rect 80435 166355 132345 166545
rect 132435 166355 137000 166545
rect 2000 166350 137000 166355
rect 1000 166245 137000 166300
rect 1000 166105 6840 166245
rect 6870 166105 71840 166245
rect 71870 166105 80840 166245
rect 80870 166105 132840 166245
rect 132870 166105 137000 166245
rect 1000 166100 137000 166105
<< via1 >>
rect 2005 169305 2495 169795
rect 136505 169305 136995 169795
rect 6345 167015 6435 167205
rect 6840 167015 6870 167205
rect 71345 167015 71435 167205
rect 71840 167015 71870 167205
rect 80345 167015 80435 167205
rect 80840 167015 80870 167205
rect 132345 167015 132435 167205
rect 132840 167015 132870 167205
rect 6345 166355 6435 166545
rect 71345 166355 71435 166545
rect 80345 166355 80435 166545
rect 132345 166355 132435 166545
rect 6840 166105 6870 166245
rect 71840 166105 71870 166245
rect 80840 166105 80870 166245
rect 132840 166105 132870 166245
<< metal2 >>
rect 2000 169795 2500 169800
rect 2000 169305 2005 169795
rect 2495 169305 2500 169795
rect 6250 169600 6350 173100
rect 71250 169600 71350 173100
rect 80250 169600 80350 173100
rect 132250 169600 132350 173100
rect 136500 169795 137000 169800
rect 2000 169300 2500 169305
rect 136500 169305 136505 169795
rect 136995 169305 137000 169795
rect 136500 169300 137000 169305
rect 6340 167205 6440 167210
rect 6340 167015 6345 167205
rect 6435 167015 6440 167205
rect 6340 166545 6440 167015
rect 6835 167205 6875 167210
rect 6835 167015 6840 167205
rect 6870 167015 6875 167205
rect 6340 166355 6345 166545
rect 6435 166355 6440 166545
rect 6340 166350 6440 166355
rect 6600 166050 6700 166890
rect 6835 166245 6875 167015
rect 71340 167205 71440 167210
rect 71340 167015 71345 167205
rect 71435 167015 71440 167205
rect 71340 166545 71440 167015
rect 71835 167205 71875 167210
rect 71835 167015 71840 167205
rect 71870 167015 71875 167205
rect 71340 166355 71345 166545
rect 71435 166355 71440 166545
rect 71340 166350 71440 166355
rect 6835 166105 6840 166245
rect 6870 166105 6875 166245
rect 6835 166100 6875 166105
rect 1000 165950 6700 166050
rect 71600 165900 71700 166890
rect 71835 166245 71875 167015
rect 80340 167205 80440 167210
rect 80340 167015 80345 167205
rect 80435 167015 80440 167205
rect 80340 166545 80440 167015
rect 80835 167205 80875 167210
rect 80835 167015 80840 167205
rect 80870 167015 80875 167205
rect 80340 166355 80345 166545
rect 80435 166355 80440 166545
rect 80340 166350 80440 166355
rect 71835 166105 71840 166245
rect 71870 166105 71875 166245
rect 71835 166100 71875 166105
rect 1200 165800 71700 165900
rect 80600 165750 80700 166890
rect 80835 166245 80875 167015
rect 132340 167205 132440 167210
rect 132340 167015 132345 167205
rect 132435 167015 132440 167205
rect 132340 166545 132440 167015
rect 132835 167205 132875 167210
rect 132835 167015 132840 167205
rect 132870 167015 132875 167205
rect 132340 166355 132345 166545
rect 132435 166355 132440 166545
rect 132340 166350 132440 166355
rect 80835 166105 80840 166245
rect 80870 166105 80875 166245
rect 80835 166100 80875 166105
rect 1400 165650 80700 165750
rect 132600 165600 132700 166890
rect 132835 166245 132875 167015
rect 132835 166105 132840 166245
rect 132870 166105 132875 166245
rect 132835 166100 132875 166105
rect 1600 165500 132700 165600
<< via2 >>
rect 2005 169305 2495 169795
rect 136505 169305 136995 169795
<< metal3 >>
rect 2000 169795 2500 176500
rect 2000 169305 2005 169795
rect 2495 169305 2500 169795
rect 2000 169300 2500 169305
rect 136500 169795 137000 176500
rect 136500 169305 136505 169795
rect 136995 169305 137000 169795
rect 136500 169300 137000 169305
use converter  converter_0
timestamp 1665354016
transform 1 0 800 0 1 0
box 0 0 137200 207200
use level_shifter  level_shifter_0
timestamp 1665425771
transform 0 -1 8468 1 0 167947
box -1223 0 1802 4468
use level_shifter  level_shifter_1
timestamp 1665425771
transform 0 -1 73468 1 0 167947
box -1223 0 1802 4468
use level_shifter  level_shifter_2
timestamp 1665425771
transform 0 -1 82468 1 0 167947
box -1223 0 1802 4468
use level_shifter  level_shifter_3
timestamp 1665425771
transform 0 -1 134468 1 0 167947
box -1223 0 1802 4468
<< labels >>
rlabel metal1 1000 166100 1200 166300 7 VDD
rlabel metal2 1000 165950 1100 166050 7 D1
rlabel metal2 1200 165800 1300 165900 7 D2
rlabel metal2 1400 165650 1500 165750 7 D3
rlabel metal2 1600 165500 1700 165600 7 D4
<< end >>
