magic
tech sky130A
timestamp 1668373927
<< metal5 >>
rect 19700 16900 40300 17000
rect 19600 16800 40400 16900
rect 19500 16700 40500 16800
rect 19400 16600 40600 16700
rect 19300 16500 40700 16600
rect 1600 16400 6000 16500
rect 7000 16400 8000 16500
rect 19200 16400 40800 16500
rect 1500 16300 6100 16400
rect 7000 16300 8100 16400
rect 19100 16300 40900 16400
rect 1400 16200 6200 16300
rect 7000 16200 8200 16300
rect 1300 16100 6300 16200
rect 7000 16100 8300 16200
rect 1200 16000 6400 16100
rect 7000 16000 8400 16100
rect 19000 16000 41000 16300
rect 1100 15900 6500 16000
rect 1000 15800 6500 15900
rect 900 15700 6500 15800
rect 800 15600 6500 15700
rect 700 15500 6500 15600
rect 600 15400 6500 15500
rect 500 15300 6500 15400
rect 400 15200 6500 15300
rect 300 15100 6500 15200
rect 200 15000 6500 15100
rect 100 14900 2200 15000
rect 0 14800 2100 14900
rect 0 8200 2000 14800
rect 7000 12000 8500 16000
rect 19000 15000 19500 16000
rect 22100 15000 23700 16000
rect 26300 15900 27900 16000
rect 26300 15400 27800 15900
rect 28400 15500 28700 16000
rect 30700 15900 32400 16000
rect 34600 15900 38300 16000
rect 30800 15800 32400 15900
rect 34700 15800 38200 15900
rect 30900 15700 32400 15800
rect 34800 15700 38100 15800
rect 31000 15600 32400 15700
rect 34900 15600 38000 15700
rect 31100 15500 32400 15600
rect 35000 15500 37900 15600
rect 28360 15400 28700 15500
rect 31200 15400 32400 15500
rect 35100 15400 37800 15500
rect 26300 15300 27240 15400
rect 26300 15200 27170 15300
rect 26300 15000 27100 15200
rect 12000 14300 13500 14500
rect 12000 14100 12200 14300
rect 12450 14200 13050 14300
rect 12550 14100 12950 14200
rect 13300 14100 13500 14300
rect 12000 14000 12300 14100
rect 12650 14000 12850 14100
rect 13200 14000 13500 14100
rect 12000 13900 12400 14000
rect 13100 13900 13500 14000
rect 12000 13700 12500 13900
rect 13000 13700 13500 13900
rect 12000 13600 12400 13700
rect 13100 13600 13500 13700
rect 12000 13500 12300 13600
rect 12650 13500 12850 13600
rect 13200 13500 13500 13600
rect 12000 13200 12200 13500
rect 12550 13400 12950 13500
rect 12450 13300 13050 13400
rect 12400 13200 13100 13300
rect 13300 13200 13500 13500
rect 12000 13000 13500 13200
rect 7000 11900 11000 12000
rect 12000 11900 13000 12000
rect 14000 11900 17500 12000
rect 7000 11800 11100 11900
rect 12000 11800 13100 11900
rect 14000 11800 17600 11900
rect 7000 11700 11200 11800
rect 12000 11700 13200 11800
rect 14000 11700 17700 11800
rect 7000 11600 11300 11700
rect 12000 11600 13300 11700
rect 14000 11600 17800 11700
rect 7000 11500 11400 11600
rect 12000 11500 13400 11600
rect 14000 11500 17900 11600
rect 7000 10500 11500 11500
rect 0 8100 2100 8200
rect 100 8000 2200 8100
rect 200 7900 6500 8000
rect 300 7800 6500 7900
rect 400 7700 6500 7800
rect 500 7600 6500 7700
rect 600 7500 6500 7600
rect 700 7400 6500 7500
rect 800 7300 6500 7400
rect 900 7200 6500 7300
rect 1000 7100 6500 7200
rect 1100 7000 6500 7100
rect 7000 7000 8500 10500
rect 1200 6900 6500 7000
rect 7100 6900 8500 7000
rect 1300 6800 6500 6900
rect 7200 6800 8500 6900
rect 1400 6700 6500 6800
rect 7300 6700 8500 6800
rect 1500 6600 6500 6700
rect 7400 6600 8500 6700
rect 1600 6500 6500 6600
rect 7500 6500 8500 6600
rect 10000 6500 11500 10500
rect 12000 7000 13500 11500
rect 12100 6900 13500 7000
rect 12200 6800 13500 6900
rect 12300 6700 13500 6800
rect 12400 6600 13500 6700
rect 12500 6500 13500 6600
rect 14000 11400 18000 11500
rect 14000 11300 18100 11400
rect 14000 11200 18200 11300
rect 14000 11100 18300 11200
rect 14000 11000 18400 11100
rect 14000 10500 18500 11000
rect 14000 2000 15500 10500
rect 17000 8000 18500 10500
rect 16000 7500 18500 8000
rect 19000 8600 19800 15000
rect 21800 9100 24000 15000
rect 26000 14800 27100 15000
rect 26000 14700 26640 14800
rect 26000 14600 26570 14700
rect 26000 13500 26500 14600
rect 26800 13500 27100 14800
rect 26000 13100 27100 13500
rect 26000 12000 26500 13100
rect 26000 11900 26570 12000
rect 26000 11800 26640 11900
rect 26800 11800 27100 13100
rect 26000 11400 27100 11800
rect 27400 15000 27800 15400
rect 28260 15300 28700 15400
rect 31300 15300 32400 15400
rect 35200 15300 37700 15400
rect 28160 15200 28660 15300
rect 31400 15200 32400 15300
rect 35300 15200 37600 15300
rect 28060 15100 28560 15200
rect 31500 15100 32400 15200
rect 35400 15100 37500 15200
rect 27960 15000 28460 15100
rect 31600 15000 32400 15100
rect 35500 15000 37400 15100
rect 40500 15000 41000 16000
rect 27400 14900 28360 15000
rect 31700 14900 32700 15000
rect 35600 14900 37300 15000
rect 27400 14800 28260 14900
rect 31800 14800 32700 14900
rect 35700 14800 37200 14900
rect 27400 14700 28160 14800
rect 31900 14700 32700 14800
rect 35800 14700 37100 14800
rect 27400 14600 28060 14700
rect 32000 14600 32700 14700
rect 35900 14600 37000 14700
rect 27400 14500 27960 14600
rect 27400 14400 27860 14500
rect 27400 12100 27800 14400
rect 29300 14200 29500 14300
rect 29200 14100 29500 14200
rect 29100 14000 29500 14100
rect 29000 13900 30300 14000
rect 28900 13800 30400 13900
rect 28800 13700 30500 13800
rect 32100 13700 32700 14600
rect 36000 14500 36900 14600
rect 36100 14400 36800 14500
rect 36200 14300 36700 14400
rect 36300 14200 36600 14300
rect 28700 13600 32700 13700
rect 28600 13500 32700 13600
rect 28500 13400 32700 13500
rect 28400 13200 32700 13400
rect 28500 13100 32700 13200
rect 28600 13000 32700 13100
rect 28700 12900 32700 13000
rect 28800 12800 32700 12900
rect 28900 12700 32700 12800
rect 29000 12600 32700 12700
rect 29100 12500 32700 12600
rect 29200 12400 29500 12500
rect 30700 12400 32700 12500
rect 29300 12300 29500 12400
rect 30800 12300 32700 12400
rect 30900 12200 32700 12300
rect 31000 12100 32700 12200
rect 27400 12000 27960 12100
rect 31100 12000 32700 12100
rect 27400 11900 28060 12000
rect 31200 11900 32700 12000
rect 27400 11800 28160 11900
rect 31300 11800 32700 11900
rect 27400 11700 28260 11800
rect 31400 11700 32700 11800
rect 27400 11600 28360 11700
rect 31500 11600 32700 11700
rect 26000 11300 27170 11400
rect 26000 11200 27240 11300
rect 27400 11200 27800 11600
rect 27960 11500 28460 11600
rect 31600 11500 32700 11600
rect 28060 11400 28560 11500
rect 31700 11400 32700 11500
rect 28160 11300 28660 11400
rect 31800 11300 32700 11400
rect 28260 11200 28700 11300
rect 31900 11200 32700 11300
rect 26000 10700 27800 11200
rect 28360 11100 28700 11200
rect 32000 11100 32700 11200
rect 26000 10600 27900 10700
rect 28400 10600 28700 11100
rect 29400 10800 29600 10900
rect 29400 10700 29700 10800
rect 29400 10600 29800 10700
rect 26000 10500 29900 10600
rect 26000 10400 30000 10500
rect 26000 10300 30100 10400
rect 26000 10200 30200 10300
rect 26000 10100 30300 10200
rect 26000 10000 30400 10100
rect 32100 10000 32700 11100
rect 34700 12500 34900 12600
rect 38000 12500 38200 12600
rect 34700 12400 35000 12500
rect 37900 12400 38200 12500
rect 34700 12300 35100 12400
rect 37800 12300 38200 12400
rect 34700 12200 35200 12300
rect 37700 12200 38200 12300
rect 34700 12100 35300 12200
rect 37600 12100 38200 12200
rect 34700 12000 35400 12100
rect 37500 12000 38200 12100
rect 34700 11900 35500 12000
rect 37400 11900 38200 12000
rect 34700 11800 35600 11900
rect 37300 11800 38200 11900
rect 34700 11700 35700 11800
rect 37200 11700 38200 11800
rect 34700 11600 35800 11700
rect 37100 11600 38200 11700
rect 34700 11500 35900 11600
rect 37000 11500 38200 11600
rect 34700 11400 36000 11500
rect 36900 11400 38200 11500
rect 34700 11300 36100 11400
rect 36800 11300 38200 11400
rect 34700 11200 36200 11300
rect 36700 11200 38200 11300
rect 34700 11100 36300 11200
rect 36600 11100 38200 11200
rect 26000 9700 30500 10000
rect 32100 9700 33700 10000
rect 26000 9630 30400 9700
rect 25750 9620 30400 9630
rect 25740 9610 30400 9620
rect 25730 9600 30400 9610
rect 24830 9590 25120 9600
rect 25720 9590 30300 9600
rect 24820 9580 25130 9590
rect 25710 9580 30300 9590
rect 24810 9570 25140 9580
rect 25700 9570 30300 9580
rect 24800 9560 25150 9570
rect 25690 9560 30300 9570
rect 24790 9550 25160 9560
rect 25680 9550 30300 9560
rect 24790 9540 25170 9550
rect 25670 9540 30300 9550
rect 24790 9530 25180 9540
rect 25660 9530 30300 9540
rect 24790 9520 25190 9530
rect 25650 9520 30300 9530
rect 24790 9510 25200 9520
rect 25640 9510 30300 9520
rect 24790 9500 25210 9510
rect 25630 9500 30300 9510
rect 24790 9490 25220 9500
rect 25620 9490 30200 9500
rect 24790 9480 25230 9490
rect 25610 9480 30200 9490
rect 24790 9470 25240 9480
rect 25600 9470 30200 9480
rect 24790 9460 25250 9470
rect 25590 9460 30200 9470
rect 24790 9450 25260 9460
rect 25580 9450 25830 9460
rect 24790 9440 25270 9450
rect 25570 9440 25820 9450
rect 24790 9430 25280 9440
rect 25560 9430 25810 9440
rect 24790 9420 25290 9430
rect 25550 9420 25800 9430
rect 24790 9410 25300 9420
rect 25540 9410 25790 9420
rect 24790 9400 25310 9410
rect 25530 9400 25780 9410
rect 26000 9400 30200 9460
rect 24790 9390 25320 9400
rect 25520 9390 25770 9400
rect 24790 9380 25330 9390
rect 25510 9380 25760 9390
rect 24790 9370 25340 9380
rect 25500 9370 25750 9380
rect 24790 9210 24950 9370
rect 25110 9360 25740 9370
rect 25120 9350 25730 9360
rect 25130 9340 25720 9350
rect 25140 9330 25710 9340
rect 25150 9320 25700 9330
rect 25160 9310 25690 9320
rect 25170 9300 25680 9310
rect 25180 9290 25670 9300
rect 25190 9280 25660 9290
rect 25200 9270 25650 9280
rect 25210 9260 25640 9270
rect 25220 9250 25630 9260
rect 25230 9240 25620 9250
rect 25240 9230 25610 9240
rect 25250 9220 25600 9230
rect 25260 9210 25590 9220
rect 24790 9180 24960 9210
rect 25270 9200 25580 9210
rect 25280 9190 25570 9200
rect 25290 9180 25560 9190
rect 24790 9150 24970 9180
rect 25300 9170 25550 9180
rect 25310 9160 25540 9170
rect 25320 9150 25530 9160
rect 24800 9120 24980 9150
rect 25330 9140 25520 9150
rect 25340 9130 25510 9140
rect 21900 9000 23900 9100
rect 24810 9090 24990 9120
rect 24820 9060 25000 9090
rect 24830 9030 25010 9060
rect 24840 9000 25020 9030
rect 22000 8900 23800 9000
rect 24850 8970 25030 9000
rect 24860 8940 25040 8970
rect 24870 8910 25050 8940
rect 22100 8800 23700 8900
rect 24880 8880 25060 8910
rect 24170 8870 24460 8880
rect 24160 8860 24470 8870
rect 24150 8850 24480 8860
rect 24890 8850 25070 8880
rect 24140 8840 24490 8850
rect 24130 8830 24500 8840
rect 24130 8820 24510 8830
rect 24900 8820 25080 8850
rect 24130 8810 24520 8820
rect 24130 8800 24530 8810
rect 22200 8700 23600 8800
rect 24130 8790 24540 8800
rect 24910 8790 25090 8820
rect 24130 8780 24550 8790
rect 24130 8770 24560 8780
rect 24130 8760 24570 8770
rect 24920 8760 25100 8790
rect 24130 8750 24580 8760
rect 24130 8740 24590 8750
rect 24130 8730 24600 8740
rect 24930 8730 25110 8760
rect 24130 8720 24610 8730
rect 24130 8710 24620 8720
rect 24130 8700 24630 8710
rect 24940 8700 25120 8730
rect 22300 8600 23500 8700
rect 24130 8690 24640 8700
rect 24130 8680 24650 8690
rect 24130 8670 24660 8680
rect 24130 8660 24670 8670
rect 24130 8650 24680 8660
rect 19000 8500 19900 8600
rect 22400 8500 23400 8600
rect 19000 8400 20000 8500
rect 24130 8490 24290 8650
rect 24450 8640 24690 8650
rect 24460 8630 24700 8640
rect 24470 8620 24710 8630
rect 24480 8610 24720 8620
rect 24490 8600 24730 8610
rect 24500 8590 24740 8600
rect 24510 8580 24750 8590
rect 24520 8570 24760 8580
rect 24530 8560 24770 8570
rect 24540 8550 24780 8560
rect 24550 8540 24790 8550
rect 24950 8540 25130 8700
rect 26000 8600 26500 9400
rect 28000 9300 30100 9400
rect 28100 9200 30000 9300
rect 28200 9100 29900 9200
rect 29400 9000 29800 9100
rect 29400 8900 29700 9000
rect 29400 8800 29600 8900
rect 24560 8530 25130 8540
rect 24570 8520 25130 8530
rect 24580 8510 25130 8520
rect 24590 8500 25130 8510
rect 25900 8500 26500 8600
rect 24600 8490 25130 8500
rect 24130 8460 24300 8490
rect 24610 8480 25130 8490
rect 24620 8470 25130 8480
rect 24630 8460 25130 8470
rect 24130 8430 24310 8460
rect 24640 8450 25130 8460
rect 24650 8440 25130 8450
rect 24660 8430 25130 8440
rect 24140 8400 24320 8430
rect 24670 8420 25130 8430
rect 24680 8410 25130 8420
rect 24690 8400 25130 8410
rect 25800 8400 26500 8500
rect 32100 8400 32700 9700
rect 19000 8300 20100 8400
rect 24150 8370 24330 8400
rect 24700 8390 25130 8400
rect 24710 8380 25130 8390
rect 24720 8370 25130 8380
rect 24160 8340 24340 8370
rect 24730 8360 25130 8370
rect 24740 8350 25130 8360
rect 24750 8340 25130 8350
rect 24170 8310 24350 8340
rect 24760 8330 25130 8340
rect 24770 8320 25130 8330
rect 24780 8310 25130 8320
rect 19000 8200 20200 8300
rect 24180 8280 24360 8310
rect 25700 8300 26600 8400
rect 32000 8300 32700 8400
rect 33400 8300 33700 9700
rect 24190 8250 24370 8280
rect 23400 8220 23720 8230
rect 24200 8220 24380 8250
rect 23390 8210 23730 8220
rect 23380 8200 23740 8210
rect 19000 8100 20300 8200
rect 23370 8190 23750 8200
rect 24210 8190 24390 8220
rect 25600 8200 26700 8300
rect 31900 8200 34400 8300
rect 23360 8180 23760 8190
rect 23360 8170 23770 8180
rect 23360 8160 23780 8170
rect 24220 8160 24400 8190
rect 23360 8150 23790 8160
rect 23360 8140 23800 8150
rect 23360 8130 23810 8140
rect 24230 8130 24410 8160
rect 23360 8120 23820 8130
rect 23360 8110 23830 8120
rect 23360 8100 23840 8110
rect 24240 8100 24420 8130
rect 25500 8100 26800 8200
rect 31800 8140 34400 8200
rect 31800 8100 32700 8140
rect 19000 8000 20400 8100
rect 23360 8090 23850 8100
rect 23360 8080 23860 8090
rect 23360 8070 23870 8080
rect 24250 8070 24430 8100
rect 23360 8060 23880 8070
rect 23360 8050 23890 8060
rect 23360 8040 23900 8050
rect 24260 8040 24440 8070
rect 23360 8030 23910 8040
rect 19000 7900 20500 8000
rect 19000 7800 20600 7900
rect 23360 7870 23520 8030
rect 23680 8020 23920 8030
rect 23690 8010 23930 8020
rect 24270 8010 24450 8040
rect 23700 8000 23940 8010
rect 23710 7990 23950 8000
rect 23720 7980 23960 7990
rect 24280 7980 24450 8010
rect 25400 8000 26900 8100
rect 31700 8000 32700 8100
rect 34700 8000 38200 11100
rect 40200 8000 41000 15000
rect 23730 7970 23970 7980
rect 23740 7960 23980 7970
rect 23750 7950 23990 7960
rect 23760 7940 24000 7950
rect 23770 7930 24010 7940
rect 23780 7920 24020 7930
rect 23790 7910 24030 7920
rect 23800 7900 24040 7910
rect 23810 7890 24050 7900
rect 23820 7880 24060 7890
rect 23830 7870 24070 7880
rect 23360 7840 23530 7870
rect 23840 7860 24080 7870
rect 23850 7850 24090 7860
rect 23860 7840 24100 7850
rect 23360 7810 23540 7840
rect 23870 7830 24110 7840
rect 23880 7820 24120 7830
rect 24290 7820 24450 7980
rect 25300 7900 27000 8000
rect 31600 7900 32400 8000
rect 23890 7810 24450 7820
rect 19000 7700 20700 7800
rect 23370 7780 23550 7810
rect 23900 7800 24450 7810
rect 25200 7800 27100 7900
rect 31500 7800 32400 7900
rect 32920 7820 34180 7980
rect 23910 7790 24450 7800
rect 23920 7780 24450 7790
rect 23380 7750 23560 7780
rect 23930 7770 24450 7780
rect 23940 7760 24450 7770
rect 23950 7750 24450 7760
rect 23390 7720 23570 7750
rect 23960 7740 24450 7750
rect 23970 7730 24450 7740
rect 23980 7720 24450 7730
rect 19000 7600 20800 7700
rect 23400 7690 23580 7720
rect 23990 7710 24450 7720
rect 24000 7700 24450 7710
rect 25100 7700 27200 7800
rect 31400 7700 32400 7800
rect 24010 7690 24450 7700
rect 23410 7660 23590 7690
rect 24020 7680 24450 7690
rect 24030 7670 24450 7680
rect 24040 7660 24450 7670
rect 23420 7630 23600 7660
rect 24050 7650 24450 7660
rect 24060 7640 24450 7650
rect 24070 7630 24450 7640
rect 23430 7600 23610 7630
rect 24080 7620 24450 7630
rect 24090 7610 24450 7620
rect 24100 7600 24450 7610
rect 25000 7600 27300 7700
rect 31300 7600 32400 7700
rect 19000 7500 20900 7600
rect 23440 7570 23620 7600
rect 24110 7590 24450 7600
rect 23440 7540 23630 7570
rect 16000 7400 18400 7500
rect 19000 7400 21000 7500
rect 23440 7420 23640 7540
rect 24900 7500 27400 7600
rect 31200 7500 32400 7600
rect 33160 7500 33940 7660
rect 23430 7410 23640 7420
rect 23420 7400 23640 7410
rect 24800 7400 27500 7500
rect 31100 7400 32400 7500
rect 16000 7300 18300 7400
rect 19000 7300 21100 7400
rect 23410 7390 23640 7400
rect 23400 7380 23640 7390
rect 23390 7370 23630 7380
rect 23380 7360 23620 7370
rect 23370 7350 23610 7360
rect 23360 7340 23600 7350
rect 23350 7330 23590 7340
rect 23340 7320 23580 7330
rect 23330 7310 23570 7320
rect 23320 7300 23560 7310
rect 24700 7300 27600 7400
rect 31000 7300 32400 7400
rect 16000 7200 18200 7300
rect 19000 7200 21200 7300
rect 23310 7290 23550 7300
rect 23300 7280 23540 7290
rect 23290 7270 23530 7280
rect 23280 7260 23520 7270
rect 23270 7250 23510 7260
rect 23260 7240 23500 7250
rect 23250 7230 23490 7240
rect 23250 7220 23480 7230
rect 23250 7210 23470 7220
rect 23250 7200 23460 7210
rect 24600 7200 27700 7300
rect 30900 7200 32400 7300
rect 16000 7100 18100 7200
rect 19000 7100 21300 7200
rect 23250 7190 23450 7200
rect 23250 7180 23440 7190
rect 23250 7170 23430 7180
rect 23250 7160 23420 7170
rect 16000 7000 18000 7100
rect 19000 7000 21400 7100
rect 23250 7000 23410 7160
rect 24500 7100 27800 7200
rect 30800 7100 32400 7200
rect 33400 7180 33700 7340
rect 24400 7000 27900 7100
rect 30700 7000 32400 7100
rect 35000 7000 37900 8000
rect 40500 7000 41000 8000
rect 16000 6900 17900 7000
rect 16000 6800 17800 6900
rect 16000 6700 17700 6800
rect 19000 6700 41000 7000
rect 16000 6600 17600 6700
rect 19100 6600 40900 6700
rect 16000 6500 17500 6600
rect 19200 6500 40800 6600
rect 19300 6400 40700 6500
rect 19400 6300 40600 6400
rect 19500 6200 40500 6300
rect 19600 6100 40400 6200
rect 19700 6000 40300 6100
<< comment >>
rect -100 21000 41100 21100
rect -100 0 0 21000
rect 41000 0 41100 21000
rect -100 -100 41100 0
<< end >>
