magic
tech sky130A
timestamp 1668218559
<< metal5 >>
rect 3500 13500 16000 16500
rect 3500 10000 6500 13500
rect 0 0 10000 10000
<< end >>
