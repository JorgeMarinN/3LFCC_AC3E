magic
tech sky130A
timestamp 1667487468
<< metal1 >>
rect 1000 41895 137200 41900
rect 1000 41605 1005 41895
rect 137195 41605 137200 41895
rect 1000 41600 137200 41605
rect 5050 41545 137200 41550
rect 5050 41455 5055 41545
rect 5145 41455 137200 41545
rect 5050 41450 137200 41455
rect 56750 41395 137200 41400
rect 56750 41305 56755 41395
rect 56845 41305 137200 41395
rect 56750 41300 137200 41305
rect 65750 41245 137200 41250
rect 65750 41155 65755 41245
rect 65845 41155 137200 41245
rect 65750 41150 137200 41155
rect 130950 41095 137200 41100
rect 130950 41005 130955 41095
rect 131045 41005 137200 41095
rect 130950 41000 137200 41005
rect 1000 40945 137200 40950
rect 1000 40705 4897 40945
rect 4930 40705 56597 40945
rect 56630 40705 65597 40945
rect 65630 40705 130797 40945
rect 130830 40705 137200 40945
rect 1000 40700 137200 40705
rect 1000 40350 137200 40650
rect 8000 40295 56000 40300
rect 8000 40005 8005 40295
rect 55995 40005 56000 40295
rect 60000 40295 65000 40300
rect 8000 40000 56000 40005
rect 60000 40005 60005 40295
rect 64995 40005 65000 40295
rect 69000 40295 130000 40300
rect 60000 40000 65000 40005
rect 69000 40005 69005 40295
rect 129995 40005 130000 40295
rect 69000 40000 130000 40005
<< via1 >>
rect 1005 41605 137195 41895
rect 5055 41455 5145 41545
rect 56755 41305 56845 41395
rect 65755 41155 65845 41245
rect 130955 41005 131045 41095
rect 4897 40705 4930 40945
rect 56597 40705 56630 40945
rect 65597 40705 65630 40945
rect 130797 40705 130830 40945
rect 4897 39906 4930 40136
rect 5335 39806 5425 40096
rect 8005 40005 55995 40295
rect 56597 39906 56630 40136
rect 57035 39806 57125 40096
rect 60005 40005 64995 40295
rect 65597 39906 65630 40136
rect 66035 39806 66125 40096
rect 69005 40005 129995 40295
rect 130797 39906 130830 40136
rect 131235 39806 131325 40096
<< metal2 >>
rect 1000 41895 137200 41900
rect 1000 41605 1005 41895
rect 137195 41605 137200 41895
rect 1000 41600 137200 41605
rect 2500 37995 3000 41600
rect 5050 41545 5150 41550
rect 5050 41455 5055 41545
rect 5145 41455 5150 41545
rect 4892 40945 4935 40950
rect 4892 40705 4897 40945
rect 4930 40705 4935 40945
rect 4892 40136 4935 40705
rect 5050 40266 5150 41455
rect 4892 39906 4897 40136
rect 4930 39906 4935 40136
rect 4892 39901 4935 39906
rect 5330 40096 5430 41600
rect 5330 39806 5335 40096
rect 5425 39806 5430 40096
rect 8000 40295 56000 41600
rect 56750 41395 56850 41400
rect 56750 41305 56755 41395
rect 56845 41305 56850 41395
rect 8000 40005 8005 40295
rect 55995 40005 56000 40295
rect 8000 40000 56000 40005
rect 56592 40945 56635 40950
rect 56592 40705 56597 40945
rect 56630 40705 56635 40945
rect 56592 40136 56635 40705
rect 56750 40266 56850 41305
rect 56592 39906 56597 40136
rect 56630 39906 56635 40136
rect 56592 39901 56635 39906
rect 57030 40096 57130 41600
rect 5330 39801 5430 39806
rect 57030 39806 57035 40096
rect 57125 39806 57130 40096
rect 60000 40295 65000 41600
rect 65750 41245 65850 41250
rect 65750 41155 65755 41245
rect 65845 41155 65850 41245
rect 60000 40005 60005 40295
rect 64995 40005 65000 40295
rect 60000 40000 65000 40005
rect 65592 40945 65635 40950
rect 65592 40705 65597 40945
rect 65630 40705 65635 40945
rect 65592 40136 65635 40705
rect 65750 40266 65850 41155
rect 65592 39906 65597 40136
rect 65630 39906 65635 40136
rect 65592 39901 65635 39906
rect 66030 40096 66130 41600
rect 57030 39801 57130 39806
rect 66030 39806 66035 40096
rect 66125 39806 66130 40096
rect 69000 40295 130000 41600
rect 130950 41095 131050 41100
rect 130950 41005 130955 41095
rect 131045 41005 131050 41095
rect 69000 40005 69005 40295
rect 129995 40005 130000 40295
rect 69000 40000 130000 40005
rect 130792 40945 130835 40950
rect 130792 40705 130797 40945
rect 130830 40705 130835 40945
rect 130792 40136 130835 40705
rect 130950 40266 131050 41005
rect 130792 39906 130797 40136
rect 130830 39906 130835 40136
rect 130792 39901 130835 39906
rect 131230 40096 131330 41600
rect 66030 39801 66130 39806
rect 131230 39806 131235 40096
rect 131325 39806 131330 40096
rect 131230 39801 131330 39806
rect 2500 37505 2505 37995
rect 2995 37505 3000 37995
rect 2500 37500 3000 37505
rect 5347 34185 5647 37451
rect 5347 33515 5362 34185
rect 5632 33515 5647 34185
rect 5347 33500 5647 33515
rect 57047 34185 57347 37451
rect 57047 33515 57062 34185
rect 57332 33515 57347 34185
rect 57047 33500 57347 33515
rect 66047 34185 66347 37451
rect 66047 33515 66062 34185
rect 66332 33515 66347 34185
rect 66047 33500 66347 33515
rect 131247 34185 131547 37451
rect 131247 33515 131262 34185
rect 131532 33515 131547 34185
rect 131247 33500 131547 33515
<< via2 >>
rect 2505 37505 2995 37995
rect 5362 33515 5632 34185
rect 57062 33515 57332 34185
rect 66062 33515 66332 34185
rect 131262 33515 131532 34185
<< metal3 >>
rect 2500 37995 3000 38000
rect 2500 37505 2505 37995
rect 2995 37505 3000 37995
rect 2500 31000 3000 37505
rect 5347 34185 5647 37451
rect 5347 33515 5362 34185
rect 5632 33515 5647 34185
rect 5347 33500 5647 33515
rect 57047 34185 57347 37451
rect 57047 33515 57062 34185
rect 57332 33515 57347 34185
rect 57047 33500 57347 33515
rect 66047 34185 66347 37451
rect 66047 33515 66062 34185
rect 66332 33515 66347 34185
rect 66047 33500 66347 33515
rect 131247 34185 131547 37451
rect 131247 33515 131262 34185
rect 131532 33515 131547 34185
rect 131247 33500 131547 33515
<< via3 >>
rect 5362 33515 5632 34185
rect 57062 33515 57332 34185
rect 66062 33515 66332 34185
rect 131262 33515 131532 34185
<< metal4 >>
rect 5347 34185 5647 37451
rect 5347 33515 5362 34185
rect 5632 33515 5647 34185
rect 5347 33500 5647 33515
rect 57047 34185 57347 37451
rect 57047 33515 57062 34185
rect 57332 33515 57347 34185
rect 57047 33500 57347 33515
rect 66047 34185 66347 37451
rect 66047 33515 66062 34185
rect 66332 33515 66347 34185
rect 66047 33500 66347 33515
rect 131247 34185 131547 37451
rect 131247 33515 131262 34185
rect 131532 33515 131547 34185
rect 131247 33500 131547 33515
<< via4 >>
rect 5362 33515 5632 34185
rect 57062 33515 57332 34185
rect 66062 33515 66332 34185
rect 131262 33515 131532 34185
<< metal5 >>
rect 5347 34185 5647 37451
rect 5347 33515 5362 34185
rect 5632 33515 5647 34185
rect 5347 33500 5647 33515
rect 57047 34185 57347 37451
rect 57047 33515 57062 34185
rect 57332 33515 57347 34185
rect 57047 33500 57347 33515
rect 66047 34185 66347 37451
rect 66047 33515 66062 34185
rect 66332 33515 66347 34185
rect 66047 33500 66347 33515
rect 131247 34185 131547 37451
rect 131247 33515 131262 34185
rect 131532 33515 131547 34185
rect 131247 33500 131547 33515
use converter  converter_0
timestamp 1667484097
transform 1 0 0 0 1 0
box 0 0 137760 209000
use level_shifter  level_shifter_0
timestamp 1666543010
transform 0 1 129200 -1 0 40426
box 0 0 3025 4468
use level_shifter  level_shifter_1
timestamp 1666543010
transform 0 1 64000 -1 0 40426
box 0 0 3025 4468
use level_shifter  level_shifter_2
timestamp 1666543010
transform 0 1 55000 -1 0 40426
box 0 0 3025 4468
use level_shifter  level_shifter_3
timestamp 1666543010
transform 0 1 3300 -1 0 40426
box 0 0 3025 4468
<< labels >>
rlabel metal1 137000 40350 137200 40650 3 VLS
rlabel metal1 137000 40700 137200 40950 7 VDD
rlabel metal1 137100 41000 137200 41100 7 D1
rlabel metal1 137100 41150 137200 41250 7 D2
rlabel metal1 137100 41300 137200 41400 7 D3
rlabel metal1 137100 41450 137200 41550 7 D4
<< end >>
