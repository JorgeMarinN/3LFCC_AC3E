magic
tech sky130A
timestamp 1668389896
<< metal1 >>
rect -51720 222600 -47200 225600
rect -51720 222400 -50400 222600
rect -50200 222400 -47200 222600
rect -51720 219400 -47200 222400
rect -51720 215600 -50400 219400
rect -72600 209000 -69600 215600
rect -69400 209000 -66400 215600
rect -66200 209000 -63200 215600
rect -63000 209000 -60000 215600
rect -59800 209000 -56800 215600
rect -56600 209000 -53600 215600
rect -53400 209000 -50400 215600
rect -50200 209000 -47200 219400
rect 48280 222600 59000 225600
rect 48280 222400 49400 222600
rect 49600 222400 52600 222600
rect 52800 222400 55800 222600
rect 56000 222400 59000 222600
rect 48280 219400 59000 222400
rect 48280 215600 49400 219400
rect -72600 208985 -47200 209000
rect -72600 207815 -72585 208985
rect -63215 207815 -47200 208985
rect -72600 207800 -47200 207815
rect -63000 207300 -60000 207800
rect -59800 207300 -56800 207800
rect -56600 207300 -53600 207800
rect -53400 207300 -50400 207800
rect -50200 207300 -47200 207800
rect -27400 207300 -24400 215600
rect -24200 207300 -21200 215600
rect -21000 207300 -18000 215600
rect -17800 207300 -14800 215600
rect -14600 207300 -11600 215600
rect -11400 207300 -8400 215600
rect -8200 207300 -5200 215600
rect -5000 207300 -2000 215600
rect 33600 207300 36600 215600
rect 36800 207300 39800 215600
rect 40000 207300 43000 215600
rect 43200 207300 46200 215600
rect 46400 207300 49400 215600
rect 49600 207300 52600 219400
rect 52800 207300 55800 219400
rect 56000 207300 59000 219400
rect 99000 225585 106000 225600
rect 99000 224115 99015 225585
rect 105985 224115 106000 225585
rect 99000 208985 106000 224115
rect 99000 207815 99015 208985
rect 105985 207815 106000 208985
rect 99000 207800 106000 207815
rect -3000 167050 3000 167300
rect -2000 166395 2000 166400
rect -2000 166105 -1795 166395
rect 1795 166105 2000 166395
rect -2000 166100 2000 166105
<< via1 >>
rect -72585 207815 -63215 208985
rect 99015 224115 105985 225585
rect 99015 207815 105985 208985
rect -1795 166105 1795 166395
<< metal2 >>
rect -51720 222600 -47200 225600
rect -51720 222400 -50400 222600
rect -50200 222400 -47200 222600
rect -51720 219400 -47200 222400
rect -51720 215600 -50400 219400
rect -72600 209000 -69600 215600
rect -69400 209000 -66400 215600
rect -66200 209000 -63200 215600
rect -63000 209000 -60000 215600
rect -59800 209000 -56800 215600
rect -56600 209000 -53600 215600
rect -53400 209000 -50400 215600
rect -50200 209000 -47200 219400
rect 48280 222600 59000 225600
rect 48280 222400 49400 222600
rect 49600 222400 52600 222600
rect 52800 222400 55800 222600
rect 56000 222400 59000 222600
rect 48280 219400 59000 222400
rect 48280 215600 49400 219400
rect -72600 208985 -47200 209000
rect -72600 207815 -72585 208985
rect -63215 207815 -47200 208985
rect -72600 207800 -47200 207815
rect -63000 207300 -60000 207800
rect -59800 207300 -56800 207800
rect -56600 207300 -53600 207800
rect -53400 207300 -50400 207800
rect -50200 207300 -47200 207800
rect -32500 215385 -30500 215400
rect -32500 212415 -31985 215385
rect -31005 212415 -30500 215385
rect -32500 212185 -30500 212415
rect -32500 209215 -31985 212185
rect -31005 209215 -30500 212185
rect -63000 204100 -60000 204300
rect -59800 204100 -56800 204300
rect -56600 204100 -53600 204300
rect -53400 204100 -50400 204300
rect -50200 204100 -47200 204300
rect -32500 197000 -30500 209215
rect -27400 207300 -24400 215600
rect -24200 207300 -21200 215600
rect -21000 207300 -18000 215600
rect -17800 207300 -14800 215600
rect -14600 207300 -11600 215600
rect -11400 207300 -8400 215600
rect -8200 207300 -5200 215600
rect -5000 207300 -2000 215600
rect 30500 215385 32500 215400
rect 30500 212415 31015 215385
rect 31985 212415 32500 215385
rect 30500 212185 32500 212415
rect 30500 209215 31015 212185
rect 31985 209215 32500 212185
rect -27400 204100 -24400 204300
rect -24200 204100 -21200 204300
rect -21000 204100 -18000 204300
rect -17800 204100 -14800 204300
rect -14600 204100 -11600 204300
rect -11400 204100 -8400 204300
rect -8200 204100 -5200 204300
rect -5000 204100 -2000 204300
rect 30500 197000 32500 209215
rect 33600 207300 36600 215600
rect 36800 207300 39800 215600
rect 40000 207300 43000 215600
rect 43200 207300 46200 215600
rect 46400 207300 49400 215600
rect 49600 207300 52600 219400
rect 52800 207300 55800 219400
rect 56000 207300 59000 219400
rect 99000 225585 106000 225600
rect 99000 224115 99015 225585
rect 105985 224115 106000 225585
rect 99000 208985 106000 224115
rect 99000 207815 99015 208985
rect 105985 207815 106000 208985
rect 99000 207800 106000 207815
rect 33600 204100 36600 204300
rect 36800 204100 39800 204300
rect 40000 204100 43000 204300
rect 43200 204100 46200 204300
rect 46400 204100 49400 204300
rect 49600 204100 52600 204300
rect 52800 204100 55800 204300
rect 56000 204100 59000 204300
rect -129000 167000 -70000 172000
rect -2000 169995 2000 170500
rect -2000 168505 -1495 169995
rect 1495 168505 2000 169995
rect -2000 166395 2000 168505
rect 70000 167000 129000 172000
rect -2000 166105 -1795 166395
rect 1795 166105 2000 166395
rect -2000 166100 2000 166105
<< via2 >>
rect -72585 207815 -63215 208985
rect -31985 212415 -31005 215385
rect -31985 209215 -31005 212185
rect 31015 212415 31985 215385
rect 31015 209215 31985 212185
rect 99015 224115 105985 225585
rect 99015 207815 105985 208985
rect -1495 168505 1495 169995
<< metal3 >>
rect -101720 222600 -83000 225600
rect -51720 222600 -47200 225600
rect 48280 222600 59000 225600
rect -132000 215400 -129000 215600
rect -110000 215400 -107000 215600
rect -105000 215400 -102000 215600
rect -86000 215400 -83000 222600
rect -50200 222400 -47200 222600
rect 56000 222400 59000 222600
rect -51720 219400 -47200 222400
rect 48280 219400 59000 222400
rect 60000 222600 68280 225600
rect 99000 225585 106000 225600
rect 99000 224115 99015 225585
rect 105985 224115 106000 225585
rect 99000 224100 106000 224115
rect 60000 215400 63000 222600
rect 68000 215400 71000 215600
rect 82000 215400 85000 215600
rect 95000 215400 98000 215600
rect -132000 215385 123200 215400
rect -132000 212415 -31985 215385
rect -31005 212415 31015 215385
rect 31985 212415 123200 215385
rect -132000 212400 123200 212415
rect -132000 212200 -129000 212400
rect -110000 212200 -107000 212400
rect -105000 212200 -102000 212400
rect -86000 212200 -83000 212400
rect 60000 212200 63000 212400
rect 68000 212200 71000 212400
rect 82000 212200 85000 212400
rect 95000 212200 98000 212400
rect 107000 212200 110000 212400
rect 120200 212200 123200 212400
rect -136800 212185 136800 212200
rect -136800 209215 -31985 212185
rect -31005 209215 31015 212185
rect 31985 209215 136800 212185
rect -136800 209200 136800 209215
rect -136800 206000 -133800 209200
rect -132000 206000 -129000 209200
rect -110000 206000 -107000 209200
rect -72600 208985 -47200 209000
rect -72600 207815 -72585 208985
rect -63215 207815 -47200 208985
rect -72600 207500 -47200 207815
rect -72600 207300 -69600 207500
rect -59800 207300 -56800 207500
rect -50200 207300 -47200 207500
rect 31800 208985 106000 209000
rect 31800 207815 99015 208985
rect 105985 207815 106000 208985
rect 31800 207500 106000 207815
rect -72600 204300 -47200 207300
rect -59800 204100 -56800 204300
rect -50200 204100 -47200 204300
rect -65000 201100 -47200 204100
rect -59800 200900 -56800 201100
rect -50200 200900 -47200 201100
rect -27400 204300 -2000 207300
rect -27400 204100 -24400 204300
rect -16000 204100 -13000 204300
rect -5000 204100 -2000 204300
rect -27400 201100 -2000 204100
rect 31800 202600 33400 207500
rect -27400 200900 -24400 201100
rect -16000 200900 -13000 201100
rect -5000 200900 -2000 201100
rect 23000 201100 33400 202600
rect 33600 204300 93000 207300
rect 107000 206000 110000 209200
rect 120200 206000 123200 209200
rect 133800 206000 136800 209200
rect 33600 204100 36600 204300
rect 43200 204100 46200 204300
rect 52800 204100 55800 204300
rect 33600 201100 65000 204100
rect 23000 200900 25000 201100
rect -65000 198000 -38000 200900
rect -27400 198000 25000 200900
rect 33600 200900 36600 201100
rect 43200 200900 46200 201100
rect 52800 200900 55800 201100
rect 33600 198000 65000 200900
rect -3000 180000 3000 198000
rect -2000 169995 2000 180000
rect -2000 168505 -1495 169995
rect 1495 168505 2000 169995
rect -2000 168000 2000 168505
<< via3 >>
rect 99015 224115 105985 225585
rect -31985 212415 -31005 215385
rect 31015 212415 31985 215385
rect -31985 209215 -31005 212185
rect 31015 209215 31985 212185
rect -72585 207815 -63215 208985
rect 99015 207815 105985 208985
<< metal4 >>
rect -101720 222600 -83000 225600
rect -51720 222600 -47200 225600
rect 48280 222600 59000 225600
rect -132000 215400 -129000 215600
rect -110000 215400 -107000 215600
rect -105000 215400 -102000 215600
rect -86000 215400 -83000 222600
rect -50200 222400 -47200 222600
rect 56000 222400 59000 222600
rect -51720 219400 -47200 222400
rect 48280 219400 59000 222400
rect 60000 222600 68280 225600
rect 99000 225585 106000 225600
rect 99000 224115 99015 225585
rect 105985 224115 106000 225585
rect 99000 224100 106000 224115
rect 60000 215400 63000 222600
rect 68000 215400 71000 215600
rect 82000 215400 85000 215600
rect 95000 215400 98000 215600
rect -132000 215385 123200 215400
rect -132000 212415 -31985 215385
rect -31005 212415 31015 215385
rect 31985 212415 123200 215385
rect -132000 212400 123200 212415
rect -132000 212200 -129000 212400
rect -110000 212200 -107000 212400
rect -105000 212200 -102000 212400
rect -86000 212200 -83000 212400
rect 60000 212200 63000 212400
rect 68000 212200 71000 212400
rect 82000 212200 85000 212400
rect 95000 212200 98000 212400
rect 107000 212200 110000 212400
rect 120200 212200 123200 212400
rect -136800 212185 136800 212200
rect -136800 209215 -31985 212185
rect -31005 209215 31015 212185
rect 31985 209215 136800 212185
rect -136800 209200 136800 209215
rect -136800 206000 -133800 209200
rect -132000 206000 -129000 209200
rect -110000 206000 -107000 209200
rect -72600 208985 -47200 209000
rect -72600 207815 -72585 208985
rect -63215 207815 -47200 208985
rect -72600 207500 -47200 207815
rect -72600 207300 -69600 207500
rect -59800 207300 -56800 207500
rect -50200 207300 -47200 207500
rect 31800 208985 106000 209000
rect 31800 207815 99015 208985
rect 105985 207815 106000 208985
rect 31800 207500 106000 207815
rect -72600 204300 -47200 207300
rect -59800 204100 -56800 204300
rect -50200 204100 -47200 204300
rect -65000 201100 -47200 204100
rect -59800 200900 -56800 201100
rect -50200 200900 -47200 201100
rect -27400 204300 -2000 207300
rect -27400 204100 -24400 204300
rect -16000 204100 -13000 204300
rect -5000 204100 -2000 204300
rect -27400 201100 -2000 204100
rect 31800 202600 33400 207500
rect -27400 200900 -24400 201100
rect -16000 200900 -13000 201100
rect -5000 200900 -2000 201100
rect 23000 201100 33400 202600
rect 33600 204300 93000 207300
rect 107000 206000 110000 209200
rect 120200 206000 123200 209200
rect 133800 206000 136800 209200
rect 33600 204100 36600 204300
rect 43200 204100 46200 204300
rect 52800 204100 55800 204300
rect 33600 201100 65000 204100
rect 23000 200900 25000 201100
rect -65000 198000 -38000 200900
rect -27400 198000 25000 200900
rect 33600 200900 36600 201100
rect 43200 200900 46200 201100
rect 52800 200900 55800 201100
rect 33600 198000 65000 200900
rect -3000 180000 3000 198000
<< via4 >>
rect 99015 224115 105985 225585
rect -31985 212415 -31005 215385
rect 31015 212415 31985 215385
rect -31985 209215 -31005 212185
rect 31015 209215 31985 212185
rect -72585 207815 -63215 208985
rect 99015 207815 105985 208985
<< metal5 >>
rect -101720 222600 -83000 225600
rect -51720 222600 -47200 225600
rect 48280 222600 59000 225600
rect -132000 215400 -129000 215600
rect -110000 215400 -107000 215600
rect -105000 215400 -102000 215600
rect -86000 215400 -83000 222600
rect -50200 222400 -47200 222600
rect 56000 222400 59000 222600
rect -51720 219400 -47200 222400
rect 48280 219400 59000 222400
rect 60000 222600 68280 225600
rect 99000 225585 106000 225600
rect 99000 224115 99015 225585
rect 105985 224115 106000 225585
rect 99000 224100 106000 224115
rect 60000 215400 63000 222600
rect 68000 215400 71000 215600
rect 82000 215400 85000 215600
rect 95000 215400 98000 215600
rect -132000 215385 123200 215400
rect -132000 212415 -31985 215385
rect -31005 212415 31015 215385
rect 31985 212415 123200 215385
rect -132000 212400 123200 212415
rect -132000 212200 -129000 212400
rect -110000 212200 -107000 212400
rect -105000 212200 -102000 212400
rect -86000 212200 -83000 212400
rect 60000 212200 63000 212400
rect 68000 212200 71000 212400
rect 82000 212200 85000 212400
rect 95000 212200 98000 212400
rect 107000 212200 110000 212400
rect 120200 212200 123200 212400
rect -136800 212185 136800 212200
rect -136800 209215 -31985 212185
rect -31005 209215 31015 212185
rect 31985 209215 136800 212185
rect -136800 209200 136800 209215
rect -136800 206000 -133800 209200
rect -132000 206000 -129000 209200
rect -110000 206000 -107000 209200
rect -72600 208985 -47200 209000
rect -72600 207815 -72585 208985
rect -63215 207815 -47200 208985
rect -72600 207500 -47200 207815
rect -72600 207300 -69600 207500
rect -59800 207300 -56800 207500
rect -50200 207300 -47200 207500
rect 31800 208985 106000 209000
rect 31800 207815 99015 208985
rect 105985 207815 106000 208985
rect 31800 207500 106000 207815
rect -72600 204300 -47200 207300
rect -59800 204100 -56800 204300
rect -50200 204100 -47200 204300
rect -65000 201100 -47200 204100
rect -59800 200900 -56800 201100
rect -50200 200900 -47200 201100
rect -27400 204300 -2000 207300
rect -27400 204100 -24400 204300
rect -16000 204100 -13000 204300
rect -5000 204100 -2000 204300
rect -27400 201100 -2000 204100
rect 31800 202600 33400 207500
rect -27400 200900 -24400 201100
rect -16000 200900 -13000 201100
rect -5000 200900 -2000 201100
rect 23000 201100 33400 202600
rect 33600 204300 93000 207300
rect 107000 206000 110000 209200
rect 120200 206000 123200 209200
rect 133800 206000 136800 209200
rect 33600 204100 36600 204300
rect 43200 204100 46200 204300
rect 52800 204100 55800 204300
rect 33600 201100 65000 204100
rect 23000 200900 25000 201100
rect -65000 198000 -38000 200900
rect -27400 198000 25000 200900
rect 33600 200900 36600 201100
rect 43200 200900 46200 201100
rect 52800 200900 55800 201100
rect 33600 198000 65000 200900
rect -3000 180000 3000 198000
use core  core_0
timestamp 1667487468
transform -1 0 -800 0 -1 208000
box 0 0 137760 209000
use core  core_1
timestamp 1667487468
transform 1 0 800 0 -1 208000
box 0 0 137760 209000
use power_pad_1_5  power_pad_1_5_0
timestamp 1668387596
transform 1 0 -31720 0 1 215600
box 0 0 30000 10000
use power_pad_1_5  power_pad_1_5_1
timestamp 1668387596
transform 1 0 -81720 0 1 215600
box 0 0 30000 10000
use power_pad_1_5  power_pad_1_5_2
timestamp 1668387596
transform 1 0 18280 0 1 215600
box 0 0 30000 10000
use power_pad_3_5  power_pad_3_5_0
timestamp 1668387625
transform 1 0 -131720 0 1 215600
box 0 0 30000 10000
use power_pad_3_5  power_pad_3_5_1
timestamp 1668387625
transform 1 0 68280 0 1 215600
box 0 0 30000 10000
use stack30um_1_5  stack30um_1_5_0
timestamp 1668366526
transform 1 0 -27400 0 1 201100
box 0 0 3000 3000
use stack30um_1_5  stack30um_1_5_1
timestamp 1668366526
transform 1 0 -24200 0 1 201100
box 0 0 3000 3000
use stack30um_1_5  stack30um_1_5_2
timestamp 1668366526
transform 1 0 -21000 0 1 201100
box 0 0 3000 3000
use stack30um_1_5  stack30um_1_5_3
timestamp 1668366526
transform 1 0 -17800 0 1 201100
box 0 0 3000 3000
use stack30um_1_5  stack30um_1_5_4
timestamp 1668366526
transform 1 0 -14600 0 1 201100
box 0 0 3000 3000
use stack30um_1_5  stack30um_1_5_5
timestamp 1668366526
transform 1 0 -11400 0 1 201100
box 0 0 3000 3000
use stack30um_1_5  stack30um_1_5_6
timestamp 1668366526
transform 1 0 -8200 0 1 201100
box 0 0 3000 3000
use stack30um_1_5  stack30um_1_5_7
timestamp 1668366526
transform 1 0 -5000 0 1 201100
box 0 0 3000 3000
use stack30um_1_5  stack30um_1_5_8
timestamp 1668366526
transform 1 0 -27400 0 1 204300
box 0 0 3000 3000
use stack30um_1_5  stack30um_1_5_9
timestamp 1668366526
transform 1 0 -24200 0 1 204300
box 0 0 3000 3000
use stack30um_1_5  stack30um_1_5_10
timestamp 1668366526
transform 1 0 -21000 0 1 204300
box 0 0 3000 3000
use stack30um_1_5  stack30um_1_5_11
timestamp 1668366526
transform 1 0 -17800 0 1 204300
box 0 0 3000 3000
use stack30um_1_5  stack30um_1_5_12
timestamp 1668366526
transform 1 0 -14600 0 1 204300
box 0 0 3000 3000
use stack30um_1_5  stack30um_1_5_13
timestamp 1668366526
transform 1 0 -11400 0 1 204300
box 0 0 3000 3000
use stack30um_1_5  stack30um_1_5_14
timestamp 1668366526
transform 1 0 -8200 0 1 204300
box 0 0 3000 3000
use stack30um_1_5  stack30um_1_5_15
timestamp 1668366526
transform 1 0 -5000 0 1 204300
box 0 0 3000 3000
use stack30um_1_5  stack30um_1_5_16
timestamp 1668366526
transform 1 0 -63000 0 1 201100
box 0 0 3000 3000
use stack30um_1_5  stack30um_1_5_17
timestamp 1668366526
transform 1 0 -59800 0 1 201100
box 0 0 3000 3000
use stack30um_1_5  stack30um_1_5_18
timestamp 1668366526
transform 1 0 -56600 0 1 201100
box 0 0 3000 3000
use stack30um_1_5  stack30um_1_5_19
timestamp 1668366526
transform 1 0 -53400 0 1 201100
box 0 0 3000 3000
use stack30um_1_5  stack30um_1_5_20
timestamp 1668366526
transform 1 0 -50200 0 1 201100
box 0 0 3000 3000
use stack30um_1_5  stack30um_1_5_21
timestamp 1668366526
transform 1 0 -63000 0 1 204300
box 0 0 3000 3000
use stack30um_1_5  stack30um_1_5_22
timestamp 1668366526
transform 1 0 -59800 0 1 204300
box 0 0 3000 3000
use stack30um_1_5  stack30um_1_5_23
timestamp 1668366526
transform 1 0 -56600 0 1 204300
box 0 0 3000 3000
use stack30um_1_5  stack30um_1_5_24
timestamp 1668366526
transform 1 0 -53400 0 1 204300
box 0 0 3000 3000
use stack30um_1_5  stack30um_1_5_25
timestamp 1668366526
transform 1 0 -50200 0 1 204300
box 0 0 3000 3000
use stack30um_1_5  stack30um_1_5_26
timestamp 1668366526
transform 1 0 33600 0 1 201100
box 0 0 3000 3000
use stack30um_1_5  stack30um_1_5_27
timestamp 1668366526
transform 1 0 36800 0 1 201100
box 0 0 3000 3000
use stack30um_1_5  stack30um_1_5_28
timestamp 1668366526
transform 1 0 40000 0 1 201100
box 0 0 3000 3000
use stack30um_1_5  stack30um_1_5_29
timestamp 1668366526
transform 1 0 43200 0 1 201100
box 0 0 3000 3000
use stack30um_1_5  stack30um_1_5_30
timestamp 1668366526
transform 1 0 46400 0 1 201100
box 0 0 3000 3000
use stack30um_1_5  stack30um_1_5_31
timestamp 1668366526
transform 1 0 49600 0 1 201100
box 0 0 3000 3000
use stack30um_1_5  stack30um_1_5_32
timestamp 1668366526
transform 1 0 52800 0 1 201100
box 0 0 3000 3000
use stack30um_1_5  stack30um_1_5_33
timestamp 1668366526
transform 1 0 56000 0 1 201100
box 0 0 3000 3000
use stack30um_1_5  stack30um_1_5_34
timestamp 1668366526
transform 1 0 33600 0 1 204300
box 0 0 3000 3000
use stack30um_1_5  stack30um_1_5_35
timestamp 1668366526
transform 1 0 36800 0 1 204300
box 0 0 3000 3000
use stack30um_1_5  stack30um_1_5_36
timestamp 1668366526
transform 1 0 40000 0 1 204300
box 0 0 3000 3000
use stack30um_1_5  stack30um_1_5_37
timestamp 1668366526
transform 1 0 43200 0 1 204300
box 0 0 3000 3000
use stack30um_1_5  stack30um_1_5_38
timestamp 1668366526
transform 1 0 46400 0 1 204300
box 0 0 3000 3000
use stack30um_1_5  stack30um_1_5_39
timestamp 1668366526
transform 1 0 49600 0 1 204300
box 0 0 3000 3000
use stack30um_1_5  stack30um_1_5_40
timestamp 1668366526
transform 1 0 52800 0 1 204300
box 0 0 3000 3000
use stack30um_1_5  stack30um_1_5_41
timestamp 1668366526
transform 1 0 56000 0 1 204300
box 0 0 3000 3000
<< labels >>
rlabel metal5 -27400 204300 -2000 207300 3 GND
rlabel metal5 -51720 222600 -47200 225600 3 Vout1
rlabel metal5 48280 222600 59000 225600 3 Vout2
rlabel metal5 -132000 206000 -129000 215600 3 VH
<< end >>
