magic
tech sky130A
timestamp 1668309370
<< poly >>
rect 100 49900 200 50000
rect 300 49700 400 50000
rect 0 49500 200 49600
rect 500 49500 600 50000
rect 0 49300 400 49400
rect 700 49300 800 50000
rect 0 49100 600 49200
rect 900 49100 1000 50000
rect 0 48900 800 49000
rect 1100 48900 1200 50000
rect 0 48700 1000 48800
rect 1300 48700 1400 50000
rect 0 48500 1200 48600
rect 1500 48500 1600 50000
rect 0 48300 1400 48400
rect 1700 48300 1800 50000
rect 0 48100 1600 48200
rect 1900 48100 2000 50000
rect 0 47900 1800 48000
rect 2100 47900 2200 50000
rect 0 47700 2000 47800
rect 2300 47700 2400 50000
rect 0 47500 2200 47600
rect 2500 47500 2600 50000
rect 0 47300 2400 47400
rect 2700 47300 2800 50000
rect 0 47100 2600 47200
rect 2900 47100 3000 50000
rect 0 46900 2800 47000
rect 3100 46900 3200 50000
rect 0 46700 3000 46800
rect 3300 46700 3400 50000
rect 0 46500 3200 46600
rect 3500 46500 3600 50000
rect 0 46300 3400 46400
rect 3700 46300 3800 50000
rect 0 46100 3600 46200
rect 3900 46100 4000 50000
rect 0 45900 3800 46000
rect 4100 45900 4200 50000
rect 0 45700 4000 45800
rect 4300 45700 4400 50000
rect 0 45500 4200 45600
rect 4500 45500 4600 50000
rect 0 45300 4400 45400
rect 4700 45300 4800 50000
rect 0 45100 4600 45200
rect 4900 45100 5000 50000
rect 0 44900 4800 45000
rect 5100 44900 5200 50000
rect 0 44700 5000 44800
rect 5300 44700 5400 50000
rect 0 44500 5200 44600
rect 5500 44500 5600 50000
rect 0 44300 5400 44400
rect 5700 44300 5800 50000
rect 0 44100 5600 44200
rect 5900 44100 6000 50000
rect 0 43900 5800 44000
rect 6100 43900 6200 50000
rect 0 43700 6000 43800
rect 6300 43700 6400 50000
rect 0 43500 6200 43600
rect 6500 43500 6600 50000
rect 0 43300 6400 43400
rect 6700 43300 6800 50000
rect 0 43100 6600 43200
rect 6900 43100 7000 50000
rect 0 42900 6800 43000
rect 7100 42900 7200 50000
rect 0 42700 7000 42800
rect 7300 42700 7400 50000
rect 0 42500 7200 42600
rect 7500 42500 7600 50000
rect 0 42300 7400 42400
rect 7700 42300 7800 50000
rect 0 42100 7600 42200
rect 7900 42100 8000 50000
rect 0 41900 7800 42000
rect 8100 41900 8200 50000
rect 0 41700 8000 41800
rect 8300 41700 8400 50000
rect 0 41500 8200 41600
rect 8500 41500 8600 50000
rect 0 41300 8400 41400
rect 8700 41300 8800 50000
rect 0 41100 8600 41200
rect 8900 41100 9000 50000
rect 0 40900 8800 41000
rect 9100 40900 9200 50000
rect 0 40700 9000 40800
rect 9300 40700 9400 50000
rect 0 40500 9200 40600
rect 9500 40500 9600 50000
rect 0 40300 9400 40400
rect 9700 40300 9800 50000
rect 0 40100 9600 40200
rect 9900 40100 10000 50000
rect 0 39900 9800 40000
rect 10100 39900 10200 50000
rect 0 39700 10000 39800
rect 10300 39700 10400 50000
rect 0 39500 10200 39600
rect 10500 39500 10600 50000
rect 0 39300 10400 39400
rect 10700 39300 10800 50000
rect 0 39100 10600 39200
rect 10900 39100 11000 50000
rect 0 38900 10800 39000
rect 11100 38900 11200 50000
rect 0 38700 11000 38800
rect 11300 38700 11400 50000
rect 0 38500 11200 38600
rect 11500 38500 11600 50000
rect 0 38300 11400 38400
rect 11700 38300 11800 50000
rect 0 38100 11600 38200
rect 11900 38100 12000 50000
rect 0 37900 11800 38000
rect 12100 37900 12200 50000
rect 0 37700 12000 37800
rect 12300 37700 12400 50000
rect 0 37500 12200 37600
rect 12500 37500 12600 50000
rect 0 37300 12400 37400
rect 12700 37300 12800 50000
rect 0 37100 12600 37200
rect 12900 37100 13000 50000
rect 0 36900 12800 37000
rect 13100 36900 13200 50000
rect 0 36700 13000 36800
rect 13300 36700 13400 50000
rect 0 36500 13200 36600
rect 13500 36500 13600 50000
rect 0 36300 13400 36400
rect 13700 36300 13800 50000
rect 0 36100 13600 36200
rect 13900 36100 14000 50000
rect 0 35900 13800 36000
rect 14100 35900 14200 50000
rect 0 35700 14000 35800
rect 14300 35700 14400 50000
rect 0 35500 14200 35600
rect 14500 35500 14600 50000
rect 0 35300 14400 35400
rect 14700 35300 14800 50000
rect 0 35100 14600 35200
rect 14900 35100 15000 50000
rect 0 34900 14800 35000
rect 15100 34900 15200 50000
rect 0 34700 15000 34800
rect 15300 34700 15400 50000
rect 0 34500 15200 34600
rect 15500 34500 15600 50000
rect 0 34300 15400 34400
rect 15700 34300 15800 50000
rect 0 34100 15600 34200
rect 15900 34100 16000 50000
rect 0 33900 15800 34000
rect 16100 33900 16200 50000
rect 0 33700 16000 33800
rect 16300 33700 16400 50000
rect 0 33500 16200 33600
rect 16500 33500 16600 50000
rect 0 33300 16400 33400
rect 16700 33300 16800 50000
rect 0 33100 16600 33200
rect 16900 33100 17000 50000
rect 0 32900 16800 33000
rect 17100 32900 17200 50000
rect 0 32700 17000 32800
rect 17300 32700 17400 50000
rect 0 32500 17200 32600
rect 17500 32500 17600 50000
rect 0 32300 17400 32400
rect 17700 32300 17800 50000
rect 0 32100 17600 32200
rect 17900 32100 18000 50000
rect 0 31900 17800 32000
rect 18100 31900 18200 50000
rect 0 31700 18000 31800
rect 18300 31700 18400 50000
rect 0 31500 18200 31600
rect 18500 31500 18600 50000
rect 0 31300 18400 31400
rect 18700 31300 18800 50000
rect 0 31100 18600 31200
rect 18900 31100 19000 50000
rect 0 30900 18800 31000
rect 19100 30900 19200 50000
rect 0 30700 19000 30800
rect 19300 30700 19400 50000
rect 0 30500 19200 30600
rect 19500 30500 19600 50000
rect 0 30300 19400 30400
rect 19700 30300 19800 50000
rect 0 30100 19600 30200
rect 19900 30100 20000 50000
rect 0 29900 19800 30000
rect 20100 29900 20200 50000
rect 0 29700 20000 29800
rect 20300 29700 20400 50000
rect 0 29500 20200 29600
rect 20500 29500 20600 50000
rect 0 29300 20400 29400
rect 20700 29300 20800 50000
rect 0 29100 20600 29200
rect 20900 29100 21000 50000
rect 0 28900 20800 29000
rect 21100 28900 21200 50000
rect 0 28700 21000 28800
rect 21300 28700 21400 50000
rect 0 28500 21200 28600
rect 21500 28500 21600 50000
rect 0 28300 21400 28400
rect 21700 28300 21800 50000
rect 0 28100 21600 28200
rect 21900 28100 22000 50000
rect 0 27900 21800 28000
rect 22100 27900 22200 50000
rect 0 27700 22000 27800
rect 22300 27700 22400 50000
rect 0 27500 22200 27600
rect 22500 27500 22600 50000
rect 0 27300 22400 27400
rect 22700 27300 22800 50000
rect 0 27100 22600 27200
rect 22900 27100 23000 50000
rect 0 26900 22800 27000
rect 23100 26900 23200 50000
rect 0 26700 23000 26800
rect 23300 26700 23400 50000
rect 0 26500 23200 26600
rect 23500 26500 23600 50000
rect 0 26300 23400 26400
rect 23700 26300 23800 50000
rect 0 26100 23600 26200
rect 23900 26100 24000 50000
rect 0 25900 23800 26000
rect 24100 25900 24200 50000
rect 0 25700 24000 25800
rect 24300 25700 24400 50000
rect 0 25500 24200 25600
rect 24500 25500 24600 50000
rect 0 25300 24400 25400
rect 24700 25300 24800 50000
rect 0 25100 24600 25200
rect 24900 25100 25000 50000
rect 25100 25300 25200 50000
rect 25300 25500 25400 50000
rect 25500 25700 25600 50000
rect 25700 25900 25800 50000
rect 25900 26100 26000 50000
rect 26100 26300 26200 50000
rect 26300 26500 26400 50000
rect 26500 26700 26600 50000
rect 26700 26900 26800 50000
rect 26900 27100 27000 50000
rect 27100 27300 27200 50000
rect 27300 27500 27400 50000
rect 27500 27700 27600 50000
rect 27700 27900 27800 50000
rect 27900 28100 28000 50000
rect 28100 28300 28200 50000
rect 28300 28500 28400 50000
rect 28500 28700 28600 50000
rect 28700 28900 28800 50000
rect 28900 29100 29000 50000
rect 29100 29300 29200 50000
rect 29300 29500 29400 50000
rect 29500 29700 29600 50000
rect 29700 29900 29800 50000
rect 29900 30100 30000 50000
rect 30100 30300 30200 50000
rect 30300 30500 30400 50000
rect 30500 30700 30600 50000
rect 30700 30900 30800 50000
rect 30900 31100 31000 50000
rect 31100 31300 31200 50000
rect 31300 31500 31400 50000
rect 31500 31700 31600 50000
rect 31700 31900 31800 50000
rect 31900 32100 32000 50000
rect 32100 32300 32200 50000
rect 32300 32500 32400 50000
rect 32500 32700 32600 50000
rect 32700 32900 32800 50000
rect 32900 33100 33000 50000
rect 33100 33300 33200 50000
rect 33300 33500 33400 50000
rect 33500 33700 33600 50000
rect 33700 33900 33800 50000
rect 33900 34100 34000 50000
rect 34100 34300 34200 50000
rect 34300 34500 34400 50000
rect 34500 34700 34600 50000
rect 34700 34900 34800 50000
rect 34900 35100 35000 50000
rect 35100 35300 35200 50000
rect 35300 35500 35400 50000
rect 35500 35700 35600 50000
rect 35700 35900 35800 50000
rect 35900 36100 36000 50000
rect 36100 36300 36200 50000
rect 36300 36500 36400 50000
rect 36500 36700 36600 50000
rect 36700 36900 36800 50000
rect 36900 37100 37000 50000
rect 37100 37300 37200 50000
rect 37300 37500 37400 50000
rect 37500 37700 37600 50000
rect 37700 37900 37800 50000
rect 37900 38100 38000 50000
rect 38100 38300 38200 50000
rect 38300 38500 38400 50000
rect 38500 38700 38600 50000
rect 38700 38900 38800 50000
rect 38900 39100 39000 50000
rect 39100 39300 39200 50000
rect 39300 39500 39400 50000
rect 39500 39700 39600 50000
rect 39700 39900 39800 50000
rect 39900 40100 40000 50000
rect 40100 40300 40200 50000
rect 40300 40500 40400 50000
rect 40500 40700 40600 50000
rect 40700 40900 40800 50000
rect 40900 41100 41000 50000
rect 41100 41300 41200 50000
rect 41300 41500 41400 50000
rect 41500 41700 41600 50000
rect 41700 41900 41800 50000
rect 41900 42100 42000 50000
rect 42100 42300 42200 50000
rect 42300 42500 42400 50000
rect 42500 42700 42600 50000
rect 42700 42900 42800 50000
rect 42900 43100 43000 50000
rect 43100 43300 43200 50000
rect 43300 43500 43400 50000
rect 43500 43700 43600 50000
rect 43700 43900 43800 50000
rect 43900 44100 44000 50000
rect 44100 44300 44200 50000
rect 44300 44500 44400 50000
rect 44500 44700 44600 50000
rect 44700 44900 44800 50000
rect 44900 45100 45000 50000
rect 45100 45300 45200 50000
rect 45300 45500 45400 50000
rect 45500 45700 45600 50000
rect 45700 45900 45800 50000
rect 45900 46100 46000 50000
rect 46100 46300 46200 50000
rect 46300 46500 46400 50000
rect 46500 46700 46600 50000
rect 46700 46900 46800 50000
rect 46900 47100 47000 50000
rect 47100 47300 47200 50000
rect 47300 47500 47400 50000
rect 47500 47700 47600 50000
rect 47700 47900 47800 50000
rect 47900 48100 48000 50000
rect 48100 48300 48200 50000
rect 48300 48500 48400 50000
rect 48500 48700 48600 50000
rect 48700 48900 48800 50000
rect 48900 49100 49000 50000
rect 49100 49300 49200 50000
rect 49300 49500 49400 50000
rect 49500 49700 49600 50000
rect 49700 49900 49800 50000
rect 49900 49700 50000 49800
rect 49700 49500 50000 49600
rect 49500 49300 50000 49400
rect 49300 49100 50000 49200
rect 49100 48900 50000 49000
rect 48900 48700 50000 48800
rect 48700 48500 50000 48600
rect 48500 48300 50000 48400
rect 48300 48100 50000 48200
rect 48100 47900 50000 48000
rect 47900 47700 50000 47800
rect 47700 47500 50000 47600
rect 47500 47300 50000 47400
rect 47300 47100 50000 47200
rect 47100 46900 50000 47000
rect 46900 46700 50000 46800
rect 46700 46500 50000 46600
rect 46500 46300 50000 46400
rect 46300 46100 50000 46200
rect 46100 45900 50000 46000
rect 45900 45700 50000 45800
rect 45700 45500 50000 45600
rect 45500 45300 50000 45400
rect 45300 45100 50000 45200
rect 45100 44900 50000 45000
rect 44900 44700 50000 44800
rect 44700 44500 50000 44600
rect 44500 44300 50000 44400
rect 44300 44100 50000 44200
rect 44100 43900 50000 44000
rect 43900 43700 50000 43800
rect 43700 43500 50000 43600
rect 43500 43300 50000 43400
rect 43300 43100 50000 43200
rect 43100 42900 50000 43000
rect 42900 42700 50000 42800
rect 42700 42500 50000 42600
rect 42500 42300 50000 42400
rect 42300 42100 50000 42200
rect 42100 41900 50000 42000
rect 41900 41700 50000 41800
rect 41700 41500 50000 41600
rect 41500 41300 50000 41400
rect 41300 41100 50000 41200
rect 41100 40900 50000 41000
rect 40900 40700 50000 40800
rect 40700 40500 50000 40600
rect 40500 40300 50000 40400
rect 40300 40100 50000 40200
rect 40100 39900 50000 40000
rect 39900 39700 50000 39800
rect 39700 39500 50000 39600
rect 39500 39300 50000 39400
rect 39300 39100 50000 39200
rect 39100 38900 50000 39000
rect 38900 38700 50000 38800
rect 38700 38500 50000 38600
rect 38500 38300 50000 38400
rect 38300 38100 50000 38200
rect 38100 37900 50000 38000
rect 37900 37700 50000 37800
rect 37700 37500 50000 37600
rect 37500 37300 50000 37400
rect 37300 37100 50000 37200
rect 37100 36900 50000 37000
rect 36900 36700 50000 36800
rect 36700 36500 50000 36600
rect 36500 36300 50000 36400
rect 36300 36100 50000 36200
rect 36100 35900 50000 36000
rect 35900 35700 50000 35800
rect 35700 35500 50000 35600
rect 35500 35300 50000 35400
rect 35300 35100 50000 35200
rect 35100 34900 50000 35000
rect 34900 34700 50000 34800
rect 34700 34500 50000 34600
rect 34500 34300 50000 34400
rect 34300 34100 50000 34200
rect 34100 33900 50000 34000
rect 33900 33700 50000 33800
rect 33700 33500 50000 33600
rect 33500 33300 50000 33400
rect 33300 33100 50000 33200
rect 33100 32900 50000 33000
rect 32900 32700 50000 32800
rect 32700 32500 50000 32600
rect 32500 32300 50000 32400
rect 32300 32100 50000 32200
rect 32100 31900 50000 32000
rect 31900 31700 50000 31800
rect 31700 31500 50000 31600
rect 31500 31300 50000 31400
rect 31300 31100 50000 31200
rect 31100 30900 50000 31000
rect 30900 30700 50000 30800
rect 30700 30500 50000 30600
rect 30500 30300 50000 30400
rect 30300 30100 50000 30200
rect 30100 29900 50000 30000
rect 29900 29700 50000 29800
rect 29700 29500 50000 29600
rect 29500 29300 50000 29400
rect 29300 29100 50000 29200
rect 29100 28900 50000 29000
rect 28900 28700 50000 28800
rect 28700 28500 50000 28600
rect 28500 28300 50000 28400
rect 28300 28100 50000 28200
rect 28100 27900 50000 28000
rect 27900 27700 50000 27800
rect 27700 27500 50000 27600
rect 27500 27300 50000 27400
rect 27300 27100 50000 27200
rect 27100 26900 50000 27000
rect 26900 26700 50000 26800
rect 26700 26500 50000 26600
rect 26500 26300 50000 26400
rect 26300 26100 50000 26200
rect 26100 25900 50000 26000
rect 25900 25700 50000 25800
rect 25700 25500 50000 25600
rect 25500 25300 50000 25400
rect 25300 25100 50000 25200
rect 0 24900 24800 25000
rect 25100 24900 50000 25000
rect 0 24700 24600 24800
rect 0 24500 24400 24600
rect 0 24300 24200 24400
rect 0 24100 24000 24200
rect 0 23900 23800 24000
rect 0 23700 23600 23800
rect 0 23500 23400 23600
rect 0 23300 23200 23400
rect 0 23100 23000 23200
rect 0 22900 22800 23000
rect 0 22700 22600 22800
rect 0 22500 22400 22600
rect 0 22300 22200 22400
rect 0 22100 22000 22200
rect 0 21900 21800 22000
rect 0 21700 21600 21800
rect 0 21500 21400 21600
rect 0 21300 21200 21400
rect 0 21100 21000 21200
rect 0 20900 20800 21000
rect 0 20700 20600 20800
rect 0 20500 20400 20600
rect 0 20300 20200 20400
rect 0 20100 20000 20200
rect 0 19900 19800 20000
rect 0 19700 19600 19800
rect 0 19500 19400 19600
rect 0 19300 19200 19400
rect 0 19100 19000 19200
rect 0 18900 18800 19000
rect 0 18700 18600 18800
rect 0 18500 18400 18600
rect 0 18300 18200 18400
rect 0 18100 18000 18200
rect 0 17900 17800 18000
rect 0 17700 17600 17800
rect 0 17500 17400 17600
rect 0 17300 17200 17400
rect 0 17100 17000 17200
rect 0 16900 16800 17000
rect 0 16700 16600 16800
rect 0 16500 16400 16600
rect 0 16300 16200 16400
rect 0 16100 16000 16200
rect 0 15900 15800 16000
rect 0 15700 15600 15800
rect 0 15500 15400 15600
rect 0 15300 15200 15400
rect 0 15100 15000 15200
rect 0 14900 14800 15000
rect 0 14700 14600 14800
rect 0 14500 14400 14600
rect 0 14300 14200 14400
rect 0 14100 14000 14200
rect 0 13900 13800 14000
rect 0 13700 13600 13800
rect 0 13500 13400 13600
rect 0 13300 13200 13400
rect 0 13100 13000 13200
rect 0 12900 12800 13000
rect 0 12700 12600 12800
rect 0 12500 12400 12600
rect 0 12300 12200 12400
rect 0 12100 12000 12200
rect 0 11900 11800 12000
rect 0 11700 11600 11800
rect 0 11500 11400 11600
rect 0 11300 11200 11400
rect 0 11100 11000 11200
rect 0 10900 10800 11000
rect 0 10700 10600 10800
rect 0 10500 10400 10600
rect 0 10300 10200 10400
rect 0 10100 10000 10200
rect 0 9900 9800 10000
rect 0 9700 9600 9800
rect 0 9500 9400 9600
rect 0 9300 9200 9400
rect 0 9100 9000 9200
rect 0 8900 8800 9000
rect 0 8700 8600 8800
rect 0 8500 8400 8600
rect 0 8300 8200 8400
rect 0 8100 8000 8200
rect 0 7900 7800 8000
rect 0 7700 7600 7800
rect 0 7500 7400 7600
rect 0 7300 7200 7400
rect 0 7100 7000 7200
rect 0 6900 6800 7000
rect 0 6700 6600 6800
rect 0 6500 6400 6600
rect 0 6300 6200 6400
rect 0 6100 6000 6200
rect 0 5900 5800 6000
rect 0 5700 5600 5800
rect 0 5500 5400 5600
rect 0 5300 5200 5400
rect 0 5100 5000 5200
rect 0 4900 4800 5000
rect 0 4700 4600 4800
rect 0 4500 4400 4600
rect 0 4300 4200 4400
rect 0 4100 4000 4200
rect 0 3900 3800 4000
rect 0 3700 3600 3800
rect 0 3500 3400 3600
rect 0 3300 3200 3400
rect 0 3100 3000 3200
rect 0 2900 2800 3000
rect 0 2700 2600 2800
rect 0 2500 2400 2600
rect 0 2300 2200 2400
rect 0 2100 2000 2200
rect 0 1900 1800 2000
rect 0 1700 1600 1800
rect 0 1500 1400 1600
rect 0 1300 1200 1400
rect 0 1100 1000 1200
rect 0 900 800 1000
rect 0 700 600 800
rect 0 500 400 600
rect 0 300 200 400
rect 300 0 400 200
rect 500 0 600 400
rect 700 0 800 600
rect 900 0 1000 800
rect 1100 0 1200 1000
rect 1300 0 1400 1200
rect 1500 0 1600 1400
rect 1700 0 1800 1600
rect 1900 0 2000 1800
rect 2100 0 2200 2000
rect 2300 0 2400 2200
rect 2500 0 2600 2400
rect 2700 0 2800 2600
rect 2900 0 3000 2800
rect 3100 0 3200 3000
rect 3300 0 3400 3200
rect 3500 0 3600 3400
rect 3700 0 3800 3600
rect 3900 0 4000 3800
rect 4100 0 4200 4000
rect 4300 0 4400 4200
rect 4500 0 4600 4400
rect 4700 0 4800 4600
rect 4900 0 5000 4800
rect 5100 0 5200 5000
rect 5300 0 5400 5200
rect 5500 0 5600 5400
rect 5700 0 5800 5600
rect 5900 0 6000 5800
rect 6100 0 6200 6000
rect 6300 0 6400 6200
rect 6500 0 6600 6400
rect 6700 0 6800 6600
rect 6900 0 7000 6800
rect 7100 0 7200 7000
rect 7300 0 7400 7200
rect 7500 0 7600 7400
rect 7700 0 7800 7600
rect 7900 0 8000 7800
rect 8100 0 8200 8000
rect 8300 0 8400 8200
rect 8500 0 8600 8400
rect 8700 0 8800 8600
rect 8900 0 9000 8800
rect 9100 0 9200 9000
rect 9300 0 9400 9200
rect 9500 0 9600 9400
rect 9700 0 9800 9600
rect 9900 0 10000 9800
rect 10100 0 10200 10000
rect 10300 0 10400 10200
rect 10500 0 10600 10400
rect 10700 0 10800 10600
rect 10900 0 11000 10800
rect 11100 0 11200 11000
rect 11300 0 11400 11200
rect 11500 0 11600 11400
rect 11700 0 11800 11600
rect 11900 0 12000 11800
rect 12100 0 12200 12000
rect 12300 0 12400 12200
rect 12500 0 12600 12400
rect 12700 0 12800 12600
rect 12900 0 13000 12800
rect 13100 0 13200 13000
rect 13300 0 13400 13200
rect 13500 0 13600 13400
rect 13700 0 13800 13600
rect 13900 0 14000 13800
rect 14100 0 14200 14000
rect 14300 0 14400 14200
rect 14500 0 14600 14400
rect 14700 0 14800 14600
rect 14900 0 15000 14800
rect 15100 0 15200 15000
rect 15300 0 15400 15200
rect 15500 0 15600 15400
rect 15700 0 15800 15600
rect 15900 0 16000 15800
rect 16100 0 16200 16000
rect 16300 0 16400 16200
rect 16500 0 16600 16400
rect 16700 0 16800 16600
rect 16900 0 17000 16800
rect 17100 0 17200 17000
rect 17300 0 17400 17200
rect 17500 0 17600 17400
rect 17700 0 17800 17600
rect 17900 0 18000 17800
rect 18100 0 18200 18000
rect 18300 0 18400 18200
rect 18500 0 18600 18400
rect 18700 0 18800 18600
rect 18900 0 19000 18800
rect 19100 0 19200 19000
rect 19300 0 19400 19200
rect 19500 0 19600 19400
rect 19700 0 19800 19600
rect 19900 0 20000 19800
rect 20100 0 20200 20000
rect 20300 0 20400 20200
rect 20500 0 20600 20400
rect 20700 0 20800 20600
rect 20900 0 21000 20800
rect 21100 0 21200 21000
rect 21300 0 21400 21200
rect 21500 0 21600 21400
rect 21700 0 21800 21600
rect 21900 0 22000 21800
rect 22100 0 22200 22000
rect 22300 0 22400 22200
rect 22500 0 22600 22400
rect 22700 0 22800 22600
rect 22900 0 23000 22800
rect 23100 0 23200 23000
rect 23300 0 23400 23200
rect 23500 0 23600 23400
rect 23700 0 23800 23600
rect 23900 0 24000 23800
rect 24100 0 24200 24000
rect 24300 0 24400 24200
rect 24500 0 24600 24400
rect 24700 0 24800 24600
rect 24900 0 25000 24800
rect 25300 24700 50000 24800
rect 25100 0 25200 24600
rect 25500 24500 50000 24600
rect 25300 0 25400 24400
rect 25700 24300 50000 24400
rect 25500 0 25600 24200
rect 25900 24100 50000 24200
rect 25700 0 25800 24000
rect 26100 23900 50000 24000
rect 25900 0 26000 23800
rect 26300 23700 50000 23800
rect 26100 0 26200 23600
rect 26500 23500 50000 23600
rect 26300 0 26400 23400
rect 26700 23300 50000 23400
rect 26500 0 26600 23200
rect 26900 23100 50000 23200
rect 26700 0 26800 23000
rect 27100 22900 50000 23000
rect 26900 0 27000 22800
rect 27300 22700 50000 22800
rect 27100 0 27200 22600
rect 27500 22500 50000 22600
rect 27300 0 27400 22400
rect 27700 22300 50000 22400
rect 27500 0 27600 22200
rect 27900 22100 50000 22200
rect 27700 0 27800 22000
rect 28100 21900 50000 22000
rect 27900 0 28000 21800
rect 28300 21700 50000 21800
rect 28100 0 28200 21600
rect 28500 21500 50000 21600
rect 28300 0 28400 21400
rect 28700 21300 50000 21400
rect 28500 0 28600 21200
rect 28900 21100 50000 21200
rect 28700 0 28800 21000
rect 29100 20900 50000 21000
rect 28900 0 29000 20800
rect 29300 20700 50000 20800
rect 29100 0 29200 20600
rect 29500 20500 50000 20600
rect 29300 0 29400 20400
rect 29700 20300 50000 20400
rect 29500 0 29600 20200
rect 29900 20100 50000 20200
rect 29700 0 29800 20000
rect 30100 19900 50000 20000
rect 29900 0 30000 19800
rect 30300 19700 50000 19800
rect 30100 0 30200 19600
rect 30500 19500 50000 19600
rect 30300 0 30400 19400
rect 30700 19300 50000 19400
rect 30500 0 30600 19200
rect 30900 19100 50000 19200
rect 30700 0 30800 19000
rect 31100 18900 50000 19000
rect 30900 0 31000 18800
rect 31300 18700 50000 18800
rect 31100 0 31200 18600
rect 31500 18500 50000 18600
rect 31300 0 31400 18400
rect 31700 18300 50000 18400
rect 31500 0 31600 18200
rect 31900 18100 50000 18200
rect 31700 0 31800 18000
rect 32100 17900 50000 18000
rect 31900 0 32000 17800
rect 32300 17700 50000 17800
rect 32100 0 32200 17600
rect 32500 17500 50000 17600
rect 32300 0 32400 17400
rect 32700 17300 50000 17400
rect 32500 0 32600 17200
rect 32900 17100 50000 17200
rect 32700 0 32800 17000
rect 33100 16900 50000 17000
rect 32900 0 33000 16800
rect 33300 16700 50000 16800
rect 33100 0 33200 16600
rect 33500 16500 50000 16600
rect 33300 0 33400 16400
rect 33700 16300 50000 16400
rect 33500 0 33600 16200
rect 33900 16100 50000 16200
rect 33700 0 33800 16000
rect 34100 15900 50000 16000
rect 33900 0 34000 15800
rect 34300 15700 50000 15800
rect 34100 0 34200 15600
rect 34500 15500 50000 15600
rect 34300 0 34400 15400
rect 34700 15300 50000 15400
rect 34500 0 34600 15200
rect 34900 15100 50000 15200
rect 34700 0 34800 15000
rect 35100 14900 50000 15000
rect 34900 0 35000 14800
rect 35300 14700 50000 14800
rect 35100 0 35200 14600
rect 35500 14500 50000 14600
rect 35300 0 35400 14400
rect 35700 14300 50000 14400
rect 35500 0 35600 14200
rect 35900 14100 50000 14200
rect 35700 0 35800 14000
rect 36100 13900 50000 14000
rect 35900 0 36000 13800
rect 36300 13700 50000 13800
rect 36100 0 36200 13600
rect 36500 13500 50000 13600
rect 36300 0 36400 13400
rect 36700 13300 50000 13400
rect 36500 0 36600 13200
rect 36900 13100 50000 13200
rect 36700 0 36800 13000
rect 37100 12900 50000 13000
rect 36900 0 37000 12800
rect 37300 12700 50000 12800
rect 37100 0 37200 12600
rect 37500 12500 50000 12600
rect 37300 0 37400 12400
rect 37700 12300 50000 12400
rect 37500 0 37600 12200
rect 37900 12100 50000 12200
rect 37700 0 37800 12000
rect 38100 11900 50000 12000
rect 37900 0 38000 11800
rect 38300 11700 50000 11800
rect 38100 0 38200 11600
rect 38500 11500 50000 11600
rect 38300 0 38400 11400
rect 38700 11300 50000 11400
rect 38500 0 38600 11200
rect 38900 11100 50000 11200
rect 38700 0 38800 11000
rect 39100 10900 50000 11000
rect 38900 0 39000 10800
rect 39300 10700 50000 10800
rect 39100 0 39200 10600
rect 39500 10500 50000 10600
rect 39300 0 39400 10400
rect 39700 10300 50000 10400
rect 39500 0 39600 10200
rect 39900 10100 50000 10200
rect 39700 0 39800 10000
rect 40100 9900 50000 10000
rect 39900 0 40000 9800
rect 40300 9700 50000 9800
rect 40100 0 40200 9600
rect 40500 9500 50000 9600
rect 40300 0 40400 9400
rect 40700 9300 50000 9400
rect 40500 0 40600 9200
rect 40900 9100 50000 9200
rect 40700 0 40800 9000
rect 41100 8900 50000 9000
rect 40900 0 41000 8800
rect 41300 8700 50000 8800
rect 41100 0 41200 8600
rect 41500 8500 50000 8600
rect 41300 0 41400 8400
rect 41700 8300 50000 8400
rect 41500 0 41600 8200
rect 41900 8100 50000 8200
rect 41700 0 41800 8000
rect 42100 7900 50000 8000
rect 41900 0 42000 7800
rect 42300 7700 50000 7800
rect 42100 0 42200 7600
rect 42500 7500 50000 7600
rect 42300 0 42400 7400
rect 42700 7300 50000 7400
rect 42500 0 42600 7200
rect 42900 7100 50000 7200
rect 42700 0 42800 7000
rect 43100 6900 50000 7000
rect 42900 0 43000 6800
rect 43300 6700 50000 6800
rect 43100 0 43200 6600
rect 43500 6500 50000 6600
rect 43300 0 43400 6400
rect 43700 6300 50000 6400
rect 43500 0 43600 6200
rect 43900 6100 50000 6200
rect 43700 0 43800 6000
rect 44100 5900 50000 6000
rect 43900 0 44000 5800
rect 44300 5700 50000 5800
rect 44100 0 44200 5600
rect 44500 5500 50000 5600
rect 44300 0 44400 5400
rect 44700 5300 50000 5400
rect 44500 0 44600 5200
rect 44900 5100 50000 5200
rect 44700 0 44800 5000
rect 45100 4900 50000 5000
rect 44900 0 45000 4800
rect 45300 4700 50000 4800
rect 45100 0 45200 4600
rect 45500 4500 50000 4600
rect 45300 0 45400 4400
rect 45700 4300 50000 4400
rect 45500 0 45600 4200
rect 45900 4100 50000 4200
rect 45700 0 45800 4000
rect 46100 3900 50000 4000
rect 45900 0 46000 3800
rect 46300 3700 50000 3800
rect 46100 0 46200 3600
rect 46500 3500 50000 3600
rect 46300 0 46400 3400
rect 46700 3300 50000 3400
rect 46500 0 46600 3200
rect 46900 3100 50000 3200
rect 46700 0 46800 3000
rect 47100 2900 50000 3000
rect 46900 0 47000 2800
rect 47300 2700 50000 2800
rect 47100 0 47200 2600
rect 47500 2500 50000 2600
rect 47300 0 47400 2400
rect 47700 2300 50000 2400
rect 47500 0 47600 2200
rect 47900 2100 50000 2200
rect 47700 0 47800 2000
rect 48100 1900 50000 2000
rect 47900 0 48000 1800
rect 48300 1700 50000 1800
rect 48100 0 48200 1600
rect 48500 1500 50000 1600
rect 48300 0 48400 1400
rect 48700 1300 50000 1400
rect 48500 0 48600 1200
rect 48900 1100 50000 1200
rect 48700 0 48800 1000
rect 49100 900 50000 1000
rect 48900 0 49000 800
rect 49300 700 50000 800
rect 49100 0 49200 600
rect 49500 500 50000 600
rect 49300 0 49400 400
rect 49700 300 50000 400
rect 49500 0 49600 200
rect 49900 100 50000 200
<< end >>
