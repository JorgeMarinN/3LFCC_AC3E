magic
tech sky130A
timestamp 1669823032
<< metal1 >>
rect 203500 23500 206500 23700
<< metal3 >>
rect 66000 99000 71000 99500
rect 500 98500 66500 99000
rect 70500 98500 71000 99000
rect 500 98000 71000 98500
rect 500 81000 1500 98000
rect 0 61600 800 62100
rect 900 61600 1100 62100
rect 500 47480 1500 47500
rect 500 47020 1020 47480
rect 1480 47020 1500 47480
rect 500 47000 1500 47020
rect 500 40500 1000 47000
rect 0 40000 1000 40500
rect 0 18400 800 18900
rect 900 18400 1100 18900
rect 0 8080 1500 8100
rect 0 7620 1020 8080
rect 1480 7620 1500 8080
rect 0 7600 1500 7620
<< rmetal3 >>
rect 800 61600 900 62100
rect 800 18400 900 18900
<< via3 >>
rect 66500 98500 70500 99000
rect 1020 47020 1480 47480
rect 1020 7620 1480 8080
<< metal4 >>
rect 66000 118000 131000 122000
rect 66000 99000 70000 118000
rect 70500 117000 126500 117500
rect 66000 98500 66500 99000
rect 66000 85500 70000 98500
rect 70500 85500 71000 117000
rect 66000 79500 71000 85500
rect 66000 71500 70000 79500
rect 70500 71500 71000 79500
rect 66000 64500 71000 71500
rect 66000 60000 70000 64500
rect 70500 61000 71000 64500
rect 126000 61000 126500 117000
rect 70500 60500 126500 61000
rect 127000 60000 131000 118000
rect 66000 56000 131000 60000
rect 1000 47480 1500 47500
rect 1000 47020 1020 47480
rect 1480 47020 1500 47480
rect 1000 47000 1500 47020
rect 1000 8080 1500 8100
rect 1000 7620 1020 8080
rect 1480 7620 1500 8080
rect 1000 7600 1500 7620
<< via4 >>
rect 70000 117500 127000 118000
rect 70000 99000 70500 117500
rect 70000 98500 70500 99000
rect 70000 85500 70500 98500
rect 70000 71500 70500 79500
rect 70000 60500 70500 64500
rect 126500 60500 127000 117500
rect 70000 60000 127000 60500
rect 1020 47020 1480 47480
rect 1020 7620 1480 8080
<< metal5 >>
rect 66000 118000 131000 122000
rect 66000 85500 70000 118000
rect 70500 117000 126500 117500
rect 70500 85500 71000 117000
rect 66000 85000 71000 85500
rect 66000 79500 71000 80000
rect 66000 71500 70000 79500
rect 70500 71500 71000 79500
rect 66000 71000 71000 71500
rect 66000 64500 71000 65000
rect 66000 60000 70000 64500
rect 70500 61000 71000 64500
rect 126000 61000 126500 117000
rect 70500 60500 126500 61000
rect 127000 60000 131000 118000
rect 66000 56000 131000 60000
<< fillblock >>
rect 1819 122000 288920 122455
rect 1819 121980 170530 122000
rect 1819 112020 132020 121980
rect 141980 112020 170530 121980
rect 1819 112000 170530 112020
rect 180530 112000 240000 122000
rect 250000 121980 288920 122000
rect 250000 112020 278550 121980
rect 288510 112020 288920 121980
rect 250000 112000 288920 112020
rect 1819 97700 288920 112000
rect 1819 97680 166000 97700
rect 1819 87720 55020 97680
rect 64980 87720 166000 97680
rect 1819 87700 166000 87720
rect 176000 87700 288920 97700
rect 1819 63100 288920 87700
rect 1819 53100 55000 63100
rect 65000 63080 288920 63100
rect 65000 53120 166020 63080
rect 175980 53120 288920 63080
rect 65000 53100 288920 53120
rect 1819 46200 288920 53100
rect 1819 45500 200000 46200
rect 1819 35500 53000 45500
rect 63000 40800 200000 45500
rect 63000 35500 110000 40800
rect 1819 31000 110000 35500
rect 1819 21000 95000 31000
rect 105000 30800 110000 31000
rect 120000 36200 200000 40800
rect 210000 45680 288920 46200
rect 210000 36200 212020 45680
rect 120000 35720 212020 36200
rect 221980 35720 288920 45680
rect 120000 30800 288920 35720
rect 105000 21000 288920 30800
rect 1819 11080 288920 21000
rect 1819 10980 110020 11080
rect 1819 1480 53020 10980
rect 62980 1480 73020 10980
rect 82980 1480 110020 10980
rect 119980 11000 212020 11080
rect 119980 1480 200000 11000
rect 210000 1480 212020 11000
rect 221980 1480 288920 11080
<< comment >>
rect 0 0 1000 1000
use ac3e  ac3e_0
timestamp 1668294652
transform 1 0 132100 0 1 79100
box -100 -100 32100 32100
use calibration  calibration_0
timestamp 1668451787
transform 1 0 132000 0 1 112000
box 0 0 48530 10000
use calibration  calibration_1
timestamp 1668451787
transform 1 0 240000 0 1 112000
box 0 0 48530 10000
use calibration_pad  calibration_pad_0
timestamp 1668450285
transform 1 0 200000 0 1 1000
box 0 0 10000 22500
use calibration_pad  calibration_pad_1
timestamp 1668450285
transform 1 0 200000 0 -1 46200
box 0 0 10000 22500
use ind2  ind2_0
timestamp 1668216304
transform 1 0 1000 0 -1 92160
box 0 0 50020 45160
use ind2  ind2_1
timestamp 1668216304
transform 1 0 71000 0 -1 111660
box 0 0 50020 45160
use ind2  ind2_2
timestamp 1668216304
transform 1 0 182000 0 -1 111660
box 0 0 50020 45160
use ind2  ind2_3
timestamp 1668216304
transform 1 0 228000 0 -1 59660
box 0 0 50020 45160
use ind3  ind3_0
timestamp 1668216541
transform 1 0 1000 0 -1 41439
box 0 0 40299 35439
use ind3  ind3_1
timestamp 1668216541
transform 1 0 126000 0 -1 49939
box 0 0 40299 35439
use ind_pad  ind_pad_0
timestamp 1668309265
transform 1 0 55000 0 1 53100
box 0 0 16000 16500
use ind_pad  ind_pad_1
timestamp 1668309265
transform 1 0 55000 0 -1 97700
box 0 0 16000 16500
use ind_pad  ind_pad_2
timestamp 1668309265
transform 1 0 110000 0 1 1100
box 0 0 16000 16500
use ind_pad  ind_pad_3
timestamp 1668309265
transform 1 0 110000 0 -1 40800
box 0 0 16000 16500
use ind_pad  ind_pad_4
timestamp 1668309265
transform 1 0 166000 0 1 53100
box 0 0 16000 16500
use ind_pad  ind_pad_5
timestamp 1668309265
transform 1 0 166000 0 -1 97700
box 0 0 16000 16500
use ind_pad  ind_pad_6
timestamp 1668309265
transform 1 0 212000 0 1 1100
box 0 0 16000 16500
use ind_pad  ind_pad_7
timestamp 1668309265
transform 1 0 212000 0 -1 45700
box 0 0 16000 16500
use ind_pad  ind_pad_8
timestamp 1668309265
transform 1 0 73000 0 1 1000
box 0 0 16000 16500
use ind_pad  ind_pad_9
timestamp 1668309265
transform -1 0 105000 0 -1 31000
box 0 0 16000 16500
use ind_pad  ind_pad_10
timestamp 1668309265
transform 1 0 53000 0 1 1000
box 0 0 16000 16500
use ind_pad  ind_pad_11
timestamp 1668309265
transform 1 0 53000 0 -1 45500
box 0 0 16000 16500
use ucu  ucu_0
timestamp 1668296084
transform 1 0 257100 0 1 94100
box -100 -100 32100 17100
use uns  uns_0
timestamp 1668297044
transform 1 0 257100 0 1 81100
box -100 -100 32100 17100
use utfsm  utfsm_0
timestamp 1668455399
transform 1 0 1100 0 1 97100
box -100 -100 49100 26100
<< end >>
