magic
tech sky130A
timestamp 1660620067
<< metal2 >>
rect 5200 57300 5500 64300
rect -1500 5200 5300 5500
<< via2 >>
rect 7600 58400 25800 59000
rect 3600 7100 4100 26500
<< metal4 >>
rect 6100 58200 7100 64300
rect 1100 7100 4400 57200
rect -1500 6100 4400 7100
rect -1500 3400 5400 4400
use nmos_waffle_36x36  nmos_waffle_36x36_0
timestamp 1624430562
transform 1 0 5400 0 1 5400
box -5400 -5400 25200 25200
use nmos_waffle_36x36  nmos_waffle_36x36_1
timestamp 1624430562
transform 0 1 5400 -1 0 57200
box -5400 -5400 25200 25200
<< labels >>
rlabel metal4 6300 63400 6900 64100 1 Vout
rlabel metal2 5200 63500 5500 64100 1 S2
rlabel metal4 -1400 6300 -900 6900 1 V1
rlabel metal4 -1300 3600 -800 4200 1 GND
rlabel metal2 -1400 5200 -900 5500 1 S1
<< end >>
