magic
tech sky130A
timestamp 1669842011
<< checkpaint >>
rect -1966 -966 51966 51966
rect -966 -1966 51966 -966
<< poly >>
rect 3000 48000 4000 50000
rect 0 47000 2000 48000
rect 5000 46000 6000 50000
rect 0 45000 4000 46000
rect 7000 44000 8000 50000
rect 0 43000 6000 44000
rect 9000 42000 10000 50000
rect 0 41000 8000 42000
rect 11000 40000 12000 50000
rect 0 39000 10000 40000
rect 13000 38000 14000 50000
rect 0 37000 12000 38000
rect 15000 36000 16000 50000
rect 0 35000 14000 36000
rect 17000 34000 18000 50000
rect 0 33000 16000 34000
rect 19000 32000 20000 50000
rect 0 31000 18000 32000
rect 21000 30000 22000 50000
rect 0 29000 20000 30000
rect 23000 28000 24000 50000
rect 0 27000 22000 28000
rect 25000 26000 26000 50000
rect 27000 28000 28000 50000
rect 29000 30000 30000 50000
rect 31000 32000 32000 50000
rect 33000 34000 34000 50000
rect 35000 36000 36000 50000
rect 37000 38000 38000 50000
rect 39000 40000 40000 50000
rect 41000 42000 42000 50000
rect 43000 44000 44000 50000
rect 45000 46000 46000 50000
rect 47000 48000 48000 50000
rect 49000 47000 50000 48000
rect 47000 45000 50000 46000
rect 45000 43000 50000 44000
rect 43000 41000 50000 42000
rect 41000 39000 50000 40000
rect 39000 37000 50000 38000
rect 37000 35000 50000 36000
rect 35000 33000 50000 34000
rect 33000 31000 50000 32000
rect 31000 29000 50000 30000
rect 29000 27000 50000 28000
rect 0 25000 24000 26000
rect 27000 25000 50000 26000
rect 0 23000 22000 24000
rect 0 21000 20000 22000
rect 0 19000 18000 20000
rect 0 17000 16000 18000
rect 0 15000 14000 16000
rect 0 13000 12000 14000
rect 0 11000 10000 12000
rect 0 9000 8000 10000
rect 0 7000 6000 8000
rect 0 5000 4000 6000
rect 0 3000 2000 4000
rect 3000 0 4000 2000
rect 5000 0 6000 4000
rect 7000 0 8000 6000
rect 9000 0 10000 8000
rect 11000 0 12000 10000
rect 13000 0 14000 12000
rect 15000 0 16000 14000
rect 17000 0 18000 16000
rect 19000 0 20000 18000
rect 21000 0 22000 20000
rect 23000 0 24000 22000
rect 25000 0 26000 24000
rect 28000 23000 50000 24000
rect 27000 0 28000 22000
rect 30000 21000 50000 22000
rect 29000 0 30000 20000
rect 32000 19000 50000 20000
rect 31000 0 32000 18000
rect 34000 17000 50000 18000
rect 33000 0 34000 16000
rect 36000 15000 50000 16000
rect 35000 0 36000 14000
rect 38000 13000 50000 14000
rect 37000 0 38000 12000
rect 40000 11000 50000 12000
rect 39000 0 40000 10000
rect 42000 9000 50000 10000
rect 41000 0 42000 8000
rect 44000 7000 50000 8000
rect 43000 0 44000 6000
rect 46000 5000 50000 6000
rect 45000 0 46000 4000
rect 48000 3000 50000 4000
rect 47000 0 48000 2000
<< end >>
