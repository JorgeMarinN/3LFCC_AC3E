magic
tech sky130A
timestamp 1668387755
<< metal1 >>
rect 0 21500 10000 22010
rect 0 500 500 21500
rect 9500 500 10000 21500
rect 0 0 10000 500
<< metal2 >>
rect 0 0 10000 22010
<< metal3 >>
rect 0 0 10000 22010
<< metal4 >>
rect 0 0 10000 22010
<< metal5 >>
rect 0 0 10000 22010
use stack30um_1_5  stack30um_1_5_0
timestamp 1668366526
transform 1 0 500 0 1 500
box 0 0 3000 3000
use stack30um_1_5  stack30um_1_5_1
timestamp 1668366526
transform 1 0 500 0 1 3500
box 0 0 3000 3000
use stack30um_1_5  stack30um_1_5_2
timestamp 1668366526
transform 1 0 500 0 1 6500
box 0 0 3000 3000
use stack30um_1_5  stack30um_1_5_3
timestamp 1668366526
transform 1 0 500 0 1 9500
box 0 0 3000 3000
use stack30um_1_5  stack30um_1_5_4
timestamp 1668366526
transform 1 0 500 0 1 12500
box 0 0 3000 3000
use stack30um_1_5  stack30um_1_5_5
timestamp 1668366526
transform 1 0 500 0 1 15500
box 0 0 3000 3000
use stack30um_1_5  stack30um_1_5_6
timestamp 1668366526
transform 1 0 500 0 1 18500
box 0 0 3000 3000
use stack30um_1_5  stack30um_1_5_7
timestamp 1668366526
transform 1 0 3500 0 1 500
box 0 0 3000 3000
use stack30um_1_5  stack30um_1_5_8
timestamp 1668366526
transform 1 0 3500 0 1 3500
box 0 0 3000 3000
use stack30um_1_5  stack30um_1_5_9
timestamp 1668366526
transform 1 0 3500 0 1 6500
box 0 0 3000 3000
use stack30um_1_5  stack30um_1_5_10
timestamp 1668366526
transform 1 0 3500 0 1 9500
box 0 0 3000 3000
use stack30um_1_5  stack30um_1_5_11
timestamp 1668366526
transform 1 0 3500 0 1 12500
box 0 0 3000 3000
use stack30um_1_5  stack30um_1_5_12
timestamp 1668366526
transform 1 0 3500 0 1 15500
box 0 0 3000 3000
use stack30um_1_5  stack30um_1_5_13
timestamp 1668366526
transform 1 0 3500 0 1 18500
box 0 0 3000 3000
use stack30um_1_5  stack30um_1_5_14
timestamp 1668366526
transform 1 0 6500 0 1 500
box 0 0 3000 3000
use stack30um_1_5  stack30um_1_5_15
timestamp 1668366526
transform 1 0 6500 0 1 3500
box 0 0 3000 3000
use stack30um_1_5  stack30um_1_5_16
timestamp 1668366526
transform 1 0 6500 0 1 6500
box 0 0 3000 3000
use stack30um_1_5  stack30um_1_5_17
timestamp 1668366526
transform 1 0 6500 0 1 9500
box 0 0 3000 3000
use stack30um_1_5  stack30um_1_5_18
timestamp 1668366526
transform 1 0 6500 0 1 12500
box 0 0 3000 3000
use stack30um_1_5  stack30um_1_5_19
timestamp 1668366526
transform 1 0 6500 0 1 15500
box 0 0 3000 3000
use stack30um_1_5  stack30um_1_5_20
timestamp 1668366526
transform 1 0 6500 0 1 18500
box 0 0 3000 3000
<< end >>
