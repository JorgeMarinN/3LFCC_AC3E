magic
tech sky130A
timestamp 1663434635
<< metal3 >>
rect 8000 150000 69000 154000
rect 8000 148300 8100 150000
rect 68900 148300 69000 150000
rect 8000 148200 69000 148300
rect 82000 150000 130000 154000
rect 82000 148300 82100 150000
rect 129900 148300 130000 150000
rect 82000 147000 130000 148300
<< via3 >>
rect 8100 148300 68900 150000
rect 82100 148300 129900 150000
<< metal4 >>
rect 8000 150000 69000 154000
rect 8000 148300 8100 150000
rect 68900 148300 69000 150000
rect 8000 147000 69000 148300
rect 82000 150000 130000 154000
rect 82000 148300 82100 150000
rect 129900 148300 130000 150000
rect 82000 148200 130000 148300
<< via4 >>
rect 8100 148300 68900 150000
rect 82100 148300 129900 150000
<< metal5 >>
rect 8000 150000 69000 154000
rect 8000 148300 8100 150000
rect 68900 148300 69000 150000
rect 8000 148200 69000 148300
rect 82000 150000 130000 154000
rect 82000 148300 82100 150000
rect 129900 148300 130000 150000
rect 82000 147000 130000 148300
use flying_cap  flying_cap_0
timestamp 1663424981
transform 1 0 30 0 1 0
box 0 0 137170 148000
use power_stage  power_stage_0
timestamp 1663434482
transform 0 -1 137200 1 0 150000
box 0 0 37200 137200
<< end >>
