magic
tech sky130A
timestamp 1660060145
<< metal2 >>
rect -771 5206 5230 5419
<< metal4 >>
rect -578 26326 3934 27131
rect 3389 6628 4360 7097
rect 3389 6614 4791 6628
rect 3386 6176 4791 6614
rect 3386 6167 4542 6176
rect 26273 3507 30785 4312
use nmos_waffle_36x36  nmos_waffle_36x36_0
timestamp 1624430562
transform 1 0 5374 0 1 5407
box -5400 -5400 25200 25200
<< labels >>
rlabel metal2 -739 5222 -336 5385 7 G
rlabel metal4 -457 26414 83 26978 7 D
rlabel metal4 30259 3665 30692 4164 3 S
<< end >>
