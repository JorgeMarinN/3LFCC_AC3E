magic
tech sky130A
timestamp 1669080206
<< error_s >>
rect 400 136794 36800 136800
rect 400 100400 415 136794
rect 400 98794 36800 98800
rect 400 62400 415 98794
rect 400 61194 30200 61200
rect 400 31400 415 61194
rect 400 30194 30200 30200
rect 400 400 415 30194
<< obsactive >>
rect -9585 136794 46815 146794
rect -9585 135000 415 136794
rect -9585 128000 -4000 135000
rect 0 128000 415 135000
rect -9585 100394 415 128000
rect 36815 100394 46815 136794
rect -9585 98794 46815 100394
rect -9585 70000 415 98794
rect -9585 63000 -4000 70000
rect 0 63000 415 70000
rect -9585 62394 415 63000
rect 36815 62394 46815 98794
rect -9585 61194 46815 62394
rect -9585 61000 415 61194
rect -9585 54000 -4000 61000
rect 0 54000 415 61000
rect -9585 31394 415 54000
rect 30215 52394 46815 61194
rect 30215 31394 40215 52394
rect -9585 30194 40215 31394
rect -9585 9000 415 30194
rect -9585 2000 -4000 9000
rect 0 2000 415 9000
rect -9585 394 415 2000
rect 30215 394 40215 30194
rect -9585 -1000 40215 394
use power_stage  power_stage_0
timestamp 1663434482
transform 1 0 0 0 1 0
box 0 0 37200 137200
<< end >>
