magic
tech sky130A
timestamp 1666495176
<< metal1 >>
rect -13000 221385 13000 221400
rect -13000 218415 -12985 221385
rect 12985 218415 13000 221385
rect -13000 218400 13000 218415
rect -12700 218200 -9700 218400
rect -9500 218200 -6500 218400
rect -6300 218200 -3300 218400
rect -3100 218200 -100 218400
rect 100 218200 3100 218400
rect 3300 218200 6300 218400
rect 6500 218200 9500 218400
rect 9700 218200 12700 218400
rect -13000 218185 13000 218200
rect -13000 215215 -12985 218185
rect 12985 215215 13000 218185
rect -13000 215200 13000 215215
rect -12700 202200 -9700 215200
rect -9500 202200 -6500 215200
rect -6300 202200 -3300 215200
rect -3100 202200 -100 215200
rect 100 202200 3100 215200
rect 3300 202200 6300 215200
rect 6500 202200 9500 215200
rect 9700 202200 12700 215200
rect -13000 202185 13000 202200
rect -13000 201215 -12985 202185
rect 12985 201215 13000 202185
rect -13000 201200 13000 201215
rect -2000 166950 2000 167150
<< via1 >>
rect -12985 218415 12985 221385
rect -12985 215215 12985 218185
rect -12985 201215 12985 202185
<< metal2 >>
rect -13000 221385 13000 221400
rect -13000 218415 -12985 221385
rect 12985 218415 13000 221385
rect -13000 218400 13000 218415
rect -12700 218200 -9700 218400
rect -9500 218200 -6500 218400
rect -6300 218200 -3300 218400
rect -3100 218200 -100 218400
rect 100 218200 3100 218400
rect 3300 218200 6300 218400
rect 6500 218200 9500 218400
rect 9700 218200 12700 218400
rect -13000 218185 13000 218200
rect -13000 215215 -12985 218185
rect 12985 215215 13000 218185
rect -13000 215200 13000 215215
rect -12700 202200 -9700 215200
rect -9500 202200 -6500 215200
rect -6300 202200 -3300 215200
rect -3100 202200 -100 215200
rect 100 202200 3100 215200
rect 3300 202200 6300 215200
rect 6500 202200 9500 215200
rect 9700 202200 12700 215200
rect -13000 202185 13000 202200
rect -13000 201215 -12985 202185
rect 12985 201215 13000 202185
rect -13000 201200 13000 201215
<< via2 >>
rect -12985 218415 12985 221385
rect -12985 215215 12985 218185
rect -12985 201215 12985 202185
<< metal3 >>
rect -13000 221385 13000 221400
rect -13000 218415 -12985 221385
rect 12985 218415 13000 221385
rect -13000 218400 13000 218415
rect -13000 218185 13000 218200
rect -13000 215215 -12985 218185
rect 12985 215215 13000 218185
rect -13000 215200 13000 215215
rect -136000 212000 136000 215000
rect -136000 211800 -133000 212000
rect -132800 211800 -129800 212000
rect 129800 211800 132800 212000
rect 133000 211800 136000 212000
rect -136000 208800 136000 211800
rect -136000 206000 -133000 208800
rect -132800 206000 -129800 208800
rect -93000 205600 93000 208600
rect 129800 206000 132800 208800
rect 133000 206000 136000 208800
rect -61000 205400 -58000 205600
rect -57800 205400 -54800 205600
rect 54800 205400 57800 205600
rect 58000 205400 61000 205600
rect -65000 202400 65000 205400
rect -61000 200000 -58000 202400
rect -57800 200000 -54800 202400
rect -13000 202185 13000 202200
rect -13000 201215 -12985 202185
rect 12985 201215 13000 202185
rect -13000 200000 13000 201215
rect 54800 200000 57800 202400
rect 58000 200000 61000 202400
rect -4000 177000 4000 200000
<< via3 >>
rect -12985 218415 12985 221385
rect -12985 215215 12985 218185
rect -12985 201215 12985 202185
<< metal4 >>
rect -13000 221385 13000 221400
rect -13000 218415 -12985 221385
rect 12985 218415 13000 221385
rect -13000 218400 13000 218415
rect -13000 218185 13000 218200
rect -13000 215215 -12985 218185
rect 12985 215215 13000 218185
rect -13000 215200 13000 215215
rect -136000 212000 136000 215000
rect -136000 211800 -133000 212000
rect -132800 211800 -129800 212000
rect 129800 211800 132800 212000
rect 133000 211800 136000 212000
rect -136000 208800 136000 211800
rect -136000 206000 -133000 208800
rect -132800 206000 -129800 208800
rect -93000 205600 93000 208600
rect 129800 206000 132800 208800
rect 133000 206000 136000 208800
rect -61000 205400 -58000 205600
rect -57800 205400 -54800 205600
rect 54800 205400 57800 205600
rect 58000 205400 61000 205600
rect -65000 202400 65000 205400
rect -61000 200000 -58000 202400
rect -57800 200000 -54800 202400
rect -13000 202185 13000 202200
rect -13000 201215 -12985 202185
rect 12985 201215 13000 202185
rect -13000 200000 13000 201215
rect 54800 200000 57800 202400
rect 58000 200000 61000 202400
rect -4000 177000 4000 200000
<< via4 >>
rect -12985 218415 12985 221385
rect -12985 215215 12985 218185
rect -12985 201215 12985 202185
<< metal5 >>
rect -13000 221385 13000 221400
rect -13000 218415 -12985 221385
rect 12985 218415 13000 221385
rect -13000 218400 13000 218415
rect -13000 218185 13000 218200
rect -13000 215215 -12985 218185
rect 12985 215215 13000 218185
rect -13000 215200 13000 215215
rect -136000 212000 136000 215000
rect -136000 211800 -133000 212000
rect -132800 211800 -129800 212000
rect 129800 211800 132800 212000
rect 133000 211800 136000 212000
rect -136000 208800 136000 211800
rect -136000 206000 -133000 208800
rect -132800 206000 -129800 208800
rect -93000 205600 93000 208600
rect 129800 206000 132800 208800
rect 133000 206000 136000 208800
rect -61000 205400 -58000 205600
rect -57800 205400 -54800 205600
rect 54800 205400 57800 205600
rect 58000 205400 61000 205600
rect -65000 202400 65000 205400
rect -61000 200000 -58000 202400
rect -57800 200000 -54800 202400
rect -13000 202185 13000 202200
rect -13000 201215 -12985 202185
rect 12985 201215 13000 202185
rect -13000 200000 13000 201215
rect 54800 200000 57800 202400
rect 58000 200000 61000 202400
rect -4000 177000 4000 200000
use core  core_0
timestamp 1666382007
transform -1 0 -800 0 -1 208000
box 0 0 137200 208000
use core  core_1
timestamp 1666382007
transform 1 0 800 0 -1 208000
box 0 0 137200 208000
<< labels >>
rlabel metal5 -1500 218400 1500 221400 7 GND
rlabel metal5 -1500 212000 1500 215000 7 VH
rlabel metal5 -1500 205600 1500 208600 7 Vout
<< end >>
