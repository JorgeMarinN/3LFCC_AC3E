magic
tech sky130A
timestamp 1667308578
<< metal1 >>
rect 900 292395 8000 292400
rect 900 292305 905 292395
rect 995 292305 8000 292395
rect 900 292300 8000 292305
rect 283000 292395 291100 292400
rect 283000 292305 291005 292395
rect 291095 292305 291100 292395
rect 283000 292300 291100 292305
rect 1050 292245 8200 292250
rect 1050 292155 1055 292245
rect 1145 292155 8200 292245
rect 1050 292150 8200 292155
rect 283000 292245 290950 292250
rect 283000 292155 290855 292245
rect 290945 292155 290950 292245
rect 283000 292150 290950 292155
rect 1200 292095 8400 292100
rect 1200 292005 1205 292095
rect 1295 292005 8400 292095
rect 1200 292000 8400 292005
rect 283000 292095 290800 292100
rect 283000 292005 290705 292095
rect 290795 292005 290800 292095
rect 283000 292000 290800 292005
rect 1350 291945 8600 291950
rect 1350 291855 1355 291945
rect 1445 291855 8600 291945
rect 1350 291850 8600 291855
rect 283000 291945 290650 291950
rect 283000 291855 290555 291945
rect 290645 291855 290650 291945
rect 283000 291850 290650 291855
<< via1 >>
rect 905 292305 995 292395
rect 291005 292305 291095 292395
rect 1055 292155 1145 292245
rect 290855 292155 290945 292245
rect 1205 292005 1295 292095
rect 290705 292005 290795 292095
rect 1355 291855 1445 291945
rect 290555 291855 290645 291945
<< metal2 >>
rect 900 292395 1000 292400
rect 900 292305 905 292395
rect 995 292305 1000 292395
rect 900 124495 1000 292305
rect 291000 292395 291100 292400
rect 291000 292305 291005 292395
rect 291095 292305 291100 292395
rect 1050 292245 1150 292250
rect 1050 292155 1055 292245
rect 1145 292155 1150 292245
rect 1050 146045 1150 292155
rect 290850 292245 290950 292250
rect 290850 292155 290855 292245
rect 290945 292155 290950 292245
rect 1200 292095 1300 292100
rect 1200 292005 1205 292095
rect 1295 292005 1300 292095
rect 1200 167595 1300 292005
rect 290700 292095 290800 292100
rect 290700 292005 290705 292095
rect 290795 292005 290800 292095
rect 1350 291945 1450 291950
rect 1350 291855 1355 291945
rect 1445 291855 1450 291945
rect 1350 189195 1450 291855
rect 290550 291945 290650 291950
rect 290550 291855 290555 291945
rect 290645 291855 290650 291945
rect 290550 204495 290650 291855
rect 290550 204405 290555 204495
rect 290645 204405 290650 204495
rect 290550 204400 290650 204405
rect 1350 189105 1355 189195
rect 1445 189105 1450 189195
rect 1350 189100 1450 189105
rect 290700 181295 290800 292005
rect 290700 181205 290705 181295
rect 290795 181205 290800 181295
rect 290700 181200 290800 181205
rect 1200 167505 1205 167595
rect 1295 167505 1300 167595
rect 1200 167500 1300 167505
rect 290850 158695 290950 292155
rect 290850 158605 290855 158695
rect 290945 158605 290950 158695
rect 290850 158600 290950 158605
rect 1050 145955 1055 146045
rect 1145 145955 1150 146045
rect 1050 145950 1150 145955
rect 291000 136495 291100 292305
rect 291000 136405 291005 136495
rect 291095 136405 291100 136495
rect 291000 136400 291100 136405
rect 900 124405 905 124495
rect 995 124405 1000 124495
rect 900 124400 1000 124405
<< via2 >>
rect 290555 204405 290645 204495
rect 1355 189105 1445 189195
rect 290705 181205 290795 181295
rect 1205 167505 1295 167595
rect 290855 158605 290945 158695
rect 1055 145955 1145 146045
rect 291005 136405 291095 136495
rect 905 124405 995 124495
<< metal3 >>
rect 4500 246000 5500 343000
rect 6000 291000 7000 351000
rect 34000 350000 62597 351150
rect 73000 351000 85300 351150
rect 87947 351000 90500 351150
rect 73000 350000 90500 351000
rect 108647 351000 111147 351150
rect 113797 351000 119000 351150
rect 108647 350000 119000 351000
rect 159497 351000 161997 351150
rect 164647 351000 181000 351150
rect 159497 350000 181000 351000
rect 206697 350000 236000 351150
rect 285000 291000 286000 351000
rect 6000 290000 8000 291000
rect 283000 290000 286000 291000
rect 286500 246000 287500 342000
rect 4500 245000 8000 246000
rect 283000 245000 287500 246000
rect 290550 204495 292000 204700
rect 290550 204405 290555 204495
rect 290645 204405 292000 204495
rect 290550 204200 292000 204405
rect 0 189195 1450 189400
rect 0 189105 1355 189195
rect 1445 189105 1450 189195
rect 0 188900 1450 189105
rect 290700 181295 292000 181500
rect 290700 181205 290705 181295
rect 290795 181205 292000 181295
rect 290700 181000 292000 181205
rect 0 167595 1300 167800
rect 0 167505 1205 167595
rect 1295 167505 1300 167595
rect 0 167300 1300 167505
rect 290850 158695 292000 158900
rect 290850 158605 290855 158695
rect 290945 158605 292000 158695
rect 290850 158400 292000 158605
rect 0 146045 1150 146200
rect 0 145955 1055 146045
rect 1145 145955 1150 146045
rect 0 145700 1150 145955
rect 291000 136495 292000 136700
rect 291000 136405 291005 136495
rect 291095 136405 292000 136495
rect 291000 136200 292000 136405
rect 0 124495 1000 124700
rect 0 124405 905 124495
rect 995 124405 1000 124495
rect 0 124200 1000 124405
<< metal4 >>
rect 34000 350000 62597 351150
rect 73000 351000 85300 351150
rect 87947 351000 90500 351150
rect 73000 350000 90500 351000
rect 108647 351000 111147 351150
rect 113797 351000 119000 351150
rect 108647 350000 119000 351000
rect 159497 351000 161997 351150
rect 164647 351000 181000 351150
rect 159497 350000 181000 351000
rect 206697 350000 236000 351150
<< metal5 >>
rect 34000 350000 62597 351150
rect 73000 351000 85300 351150
rect 87947 351000 90500 351150
rect 73000 350000 90500 351000
rect 108647 351000 111147 351150
rect 113797 351000 119000 351150
rect 108647 350000 119000 351000
rect 159497 351000 161997 351150
rect 164647 351000 181000 351150
rect 159497 350000 181000 351000
rect 206697 350000 236000 351150
<< comment >>
rect 14280 341100 44280 351100
rect 64280 341100 94280 351100
rect 114280 341100 144280 351100
rect 164280 341100 194280 351100
rect 214280 341100 244280 351100
rect 0 0 1000 1000
use interleaved  interleaved_0
timestamp 1667308048
transform 1 0 146280 0 1 125500
box -139120 0 138560 225600
<< labels >>
rlabel metal3 0 124200 1000 124700 7 D1
rlabel metal3 0 145700 1150 146200 7 D2
rlabel metal3 0 167300 1300 167800 7 D3
rlabel metal3 0 188900 1450 189400 7 D4
rlabel metal3 291000 136200 292000 136700 3 D5
rlabel metal3 290850 158400 292000 158900 3 D6
rlabel metal3 290700 181000 292000 181500 3 D7
rlabel metal3 290550 204200 292000 204700 3 D8
<< end >>
