magic
tech sky130A
timestamp 1667308048
<< metal1 >>
rect -72600 225585 -47200 225600
rect -72600 222615 -72585 225585
rect -47215 222615 -47200 225585
rect -72600 222600 -47200 222615
rect -72600 222400 -69600 222600
rect -69400 222400 -66400 222600
rect -66200 222400 -63200 222600
rect -63000 222400 -60000 222600
rect -59800 222400 -56800 222600
rect -56600 222400 -53600 222600
rect -53400 222400 -50400 222600
rect -50200 222400 -47200 222600
rect -72600 222385 -47200 222400
rect -72600 219415 -72585 222385
rect -47215 219415 -47200 222385
rect -72600 219400 -47200 219415
rect -72600 209000 -69600 219400
rect -69400 209000 -66400 219400
rect -66200 209000 -63200 219400
rect -63000 209000 -60000 219400
rect -59800 209000 -56800 219400
rect -56600 209000 -53600 219400
rect -53400 209000 -50400 219400
rect -50200 209000 -47200 219400
rect -72600 208985 -47200 209000
rect -72600 207815 -72585 208985
rect -47215 207815 -47200 208985
rect -72600 207800 -47200 207815
rect -63000 207300 -60000 207800
rect -59800 207300 -56800 207800
rect -56600 207300 -53600 207800
rect -53400 207300 -50400 207800
rect -50200 207300 -47200 207800
rect -63000 207285 -47200 207300
rect -63000 204315 -62985 207285
rect -47215 204315 -47200 207285
rect -63000 204300 -47200 204315
rect -63000 204100 -60000 204300
rect -59800 204100 -56800 204300
rect -56600 204100 -53600 204300
rect -53400 204100 -50400 204300
rect -50200 204100 -47200 204300
rect -63000 204085 -47200 204100
rect -63000 201115 -62985 204085
rect -47215 201115 -47200 204085
rect -63000 201100 -47200 201115
rect -27600 225585 -2000 225600
rect -27600 222615 -27585 225585
rect -2015 222615 -2000 225585
rect -27600 222600 -2000 222615
rect -27600 222400 -24400 222600
rect -24200 222400 -21200 222600
rect -21000 222400 -18000 222600
rect -17800 222400 -14800 222600
rect -14600 222400 -11600 222600
rect -11400 222400 -8400 222600
rect -8200 222400 -5200 222600
rect -5000 222400 -2000 222600
rect -27600 222385 -2000 222400
rect -27600 219415 -27585 222385
rect -2015 219415 -2000 222385
rect -27600 219400 -2000 219415
rect -27600 207300 -24400 219400
rect -24200 207300 -21200 219400
rect -21000 207300 -18000 219400
rect -17800 207300 -14800 219400
rect -14600 207300 -11600 219400
rect -11400 207300 -8400 219400
rect -8200 207300 -5200 219400
rect -5000 207300 -2000 219400
rect -27600 207285 -2000 207300
rect -27600 204315 -27585 207285
rect -2015 204315 -2000 207285
rect -27600 204300 -2000 204315
rect -27600 204100 -24400 204300
rect -24200 204100 -21200 204300
rect -21000 204100 -18000 204300
rect -17800 204100 -14800 204300
rect -14600 204100 -11600 204300
rect -11400 204100 -8400 204300
rect -8200 204100 -5200 204300
rect -5000 204100 -2000 204300
rect -27600 204085 -2000 204100
rect -27600 201115 -27585 204085
rect -2015 201115 -2000 204085
rect -27600 201100 -2000 201115
rect 33600 225585 59000 225600
rect 33600 222615 33615 225585
rect 58985 222615 59000 225585
rect 33600 222600 59000 222615
rect 33600 222400 36600 222600
rect 36800 222400 39800 222600
rect 40000 222400 43000 222600
rect 43200 222400 46200 222600
rect 46400 222400 49400 222600
rect 49600 222400 52600 222600
rect 52800 222400 55800 222600
rect 56000 222400 59000 222600
rect 33600 222385 59000 222400
rect 33600 219415 33615 222385
rect 58985 219415 59000 222385
rect 33600 219400 59000 219415
rect 33600 207300 36600 219400
rect 36800 207300 39800 219400
rect 40000 207300 43000 219400
rect 43200 207300 46200 219400
rect 46400 207300 49400 219400
rect 49600 207300 52600 219400
rect 52800 207300 55800 219400
rect 56000 207300 59000 219400
rect 99000 225585 106000 225600
rect 99000 224115 99015 225585
rect 105985 224115 106000 225585
rect 99000 208985 106000 224115
rect 99000 207815 99015 208985
rect 105985 207815 106000 208985
rect 99000 207800 106000 207815
rect 33600 207285 59000 207300
rect 33600 204315 33615 207285
rect 58985 204315 59000 207285
rect 33600 204300 59000 204315
rect 33600 204100 36600 204300
rect 36800 204100 39800 204300
rect 40000 204100 43000 204300
rect 43200 204100 46200 204300
rect 46400 204100 49400 204300
rect 49600 204100 52600 204300
rect 52800 204100 55800 204300
rect 56000 204100 59000 204300
rect 33600 204085 59000 204100
rect 33600 201115 33615 204085
rect 58985 201115 59000 204085
rect 33600 201100 59000 201115
rect -3000 166950 3000 167150
<< via1 >>
rect -72585 222615 -47215 225585
rect -72585 219415 -47215 222385
rect -72585 207815 -47215 208985
rect -62985 204315 -47215 207285
rect -62985 201115 -47215 204085
rect -27585 222615 -2015 225585
rect -27585 219415 -2015 222385
rect -27585 204315 -2015 207285
rect -27585 201115 -2015 204085
rect 33615 222615 58985 225585
rect 33615 219415 58985 222385
rect 99015 224115 105985 225585
rect 99015 207815 105985 208985
rect 33615 204315 58985 207285
rect 33615 201115 58985 204085
<< metal2 >>
rect -72600 225585 -47200 225600
rect -72600 222615 -72585 225585
rect -47215 222615 -47200 225585
rect -72600 222600 -47200 222615
rect -72600 222400 -69600 222600
rect -69400 222400 -66400 222600
rect -66200 222400 -63200 222600
rect -63000 222400 -60000 222600
rect -59800 222400 -56800 222600
rect -56600 222400 -53600 222600
rect -53400 222400 -50400 222600
rect -50200 222400 -47200 222600
rect -72600 222385 -47200 222400
rect -72600 219415 -72585 222385
rect -47215 219415 -47200 222385
rect -72600 219400 -47200 219415
rect -72600 209000 -69600 219400
rect -69400 209000 -66400 219400
rect -66200 209000 -63200 219400
rect -63000 209000 -60000 219400
rect -59800 209000 -56800 219400
rect -56600 209000 -53600 219400
rect -53400 209000 -50400 219400
rect -50200 209000 -47200 219400
rect -27600 225585 -2000 225600
rect -27600 222615 -27585 225585
rect -2015 222615 -2000 225585
rect -27600 222600 -2000 222615
rect -27600 222400 -24400 222600
rect -24200 222400 -21200 222600
rect -21000 222400 -18000 222600
rect -17800 222400 -14800 222600
rect -14600 222400 -11600 222600
rect -11400 222400 -8400 222600
rect -8200 222400 -5200 222600
rect -5000 222400 -2000 222600
rect -27600 222385 -2000 222400
rect -27600 219415 -27585 222385
rect -2015 219415 -2000 222385
rect -27600 219400 -2000 219415
rect -72600 208985 -47200 209000
rect -72600 207815 -72585 208985
rect -47215 207815 -47200 208985
rect -72600 207800 -47200 207815
rect -63000 207300 -60000 207800
rect -59800 207300 -56800 207800
rect -56600 207300 -53600 207800
rect -53400 207300 -50400 207800
rect -50200 207300 -47200 207800
rect -63000 207285 -47200 207300
rect -63000 204315 -62985 207285
rect -47215 204315 -47200 207285
rect -63000 204300 -47200 204315
rect -63000 204100 -60000 204300
rect -59800 204100 -56800 204300
rect -56600 204100 -53600 204300
rect -53400 204100 -50400 204300
rect -50200 204100 -47200 204300
rect -63000 204085 -47200 204100
rect -63000 201115 -62985 204085
rect -47215 201115 -47200 204085
rect -63000 201100 -47200 201115
rect -32500 215385 -30500 215400
rect -32500 212415 -32485 215385
rect -30505 212415 -30500 215385
rect -32500 212185 -30500 212415
rect -32500 209215 -32485 212185
rect -30505 209215 -30500 212185
rect -32500 197000 -30500 209215
rect -27600 207300 -24400 219400
rect -24200 207300 -21200 219400
rect -21000 207300 -18000 219400
rect -17800 207300 -14800 219400
rect -14600 207300 -11600 219400
rect -11400 207300 -8400 219400
rect -8200 207300 -5200 219400
rect -5000 207300 -2000 219400
rect 33600 225585 59000 225600
rect 33600 222615 33615 225585
rect 58985 222615 59000 225585
rect 33600 222600 59000 222615
rect 33600 222400 36600 222600
rect 36800 222400 39800 222600
rect 40000 222400 43000 222600
rect 43200 222400 46200 222600
rect 46400 222400 49400 222600
rect 49600 222400 52600 222600
rect 52800 222400 55800 222600
rect 56000 222400 59000 222600
rect 33600 222385 59000 222400
rect 33600 219415 33615 222385
rect 58985 219415 59000 222385
rect 33600 219400 59000 219415
rect -27600 207285 -2000 207300
rect -27600 204315 -27585 207285
rect -2015 204315 -2000 207285
rect -27600 204300 -2000 204315
rect -27600 204100 -24400 204300
rect -24200 204100 -21200 204300
rect -21000 204100 -18000 204300
rect -17800 204100 -14800 204300
rect -14600 204100 -11600 204300
rect -11400 204100 -8400 204300
rect -8200 204100 -5200 204300
rect -5000 204100 -2000 204300
rect -27600 204085 -2000 204100
rect -27600 201115 -27585 204085
rect -2015 201115 -2000 204085
rect -27600 201100 -2000 201115
rect 30500 215385 32500 215400
rect 30500 212415 30515 215385
rect 32485 212415 32500 215385
rect 30500 212185 32500 212415
rect 30500 209215 30515 212185
rect 32485 209215 32500 212185
rect 30500 197000 32500 209215
rect 33600 207300 36600 219400
rect 36800 207300 39800 219400
rect 40000 207300 43000 219400
rect 43200 207300 46200 219400
rect 46400 207300 49400 219400
rect 49600 207300 52600 219400
rect 52800 207300 55800 219400
rect 56000 207300 59000 219400
rect 99000 225585 106000 225600
rect 99000 224115 99015 225585
rect 105985 224115 106000 225585
rect 99000 208985 106000 224115
rect 99000 207815 99015 208985
rect 105985 207815 106000 208985
rect 99000 207800 106000 207815
rect 33600 207285 59000 207300
rect 33600 204315 33615 207285
rect 58985 204315 59000 207285
rect 33600 204300 59000 204315
rect 33600 204100 36600 204300
rect 36800 204100 39800 204300
rect 40000 204100 43000 204300
rect 43200 204100 46200 204300
rect 46400 204100 49400 204300
rect 49600 204100 52600 204300
rect 52800 204100 55800 204300
rect 56000 204100 59000 204300
rect 33600 204085 59000 204100
rect 33600 201115 33615 204085
rect 58985 201115 59000 204085
rect 33600 201100 59000 201115
<< via2 >>
rect -72585 222615 -47215 225585
rect -72585 219415 -47215 222385
rect -27585 222615 -2015 225585
rect -27585 219415 -2015 222385
rect -72585 207815 -47215 208985
rect -62985 204315 -47215 207285
rect -62985 201115 -47215 204085
rect -32485 212415 -30505 215385
rect -32485 209215 -30505 212185
rect 33615 222615 58985 225585
rect 33615 219415 58985 222385
rect -27585 204315 -2015 207285
rect -27585 201115 -2015 204085
rect 30515 212415 32485 215385
rect 30515 209215 32485 212185
rect 99015 224115 105985 225585
rect 99015 207815 105985 208985
rect 33615 204315 58985 207285
rect 33615 201115 58985 204085
<< metal3 >>
rect -132000 222600 -102000 225600
rect -132000 215400 -129000 222600
rect -110000 215400 -107000 222600
rect -105000 215400 -102000 222600
rect -72600 225585 -47200 225600
rect -72600 222615 -72585 225585
rect -47215 222615 -47200 225585
rect -72600 222600 -47200 222615
rect -72600 222400 -69600 222600
rect -50200 222400 -47200 222600
rect -72600 222385 -47200 222400
rect -72600 219415 -72585 222385
rect -47215 219415 -47200 222385
rect -72600 219400 -47200 219415
rect -27600 225585 -2000 225600
rect -27600 222615 -27585 225585
rect -2015 222615 -2000 225585
rect -27600 222600 -2000 222615
rect -27600 222400 -24600 222600
rect -5000 222400 -2000 222600
rect -27600 222385 -2000 222400
rect -27600 219415 -27585 222385
rect -2015 219415 -2000 222385
rect -27600 219400 -2000 219415
rect 33600 225585 59000 225600
rect 33600 222615 33615 225585
rect 58985 222615 59000 225585
rect 33600 222600 59000 222615
rect 33600 222400 36600 222600
rect 56000 222400 59000 222600
rect 33600 222385 59000 222400
rect 33600 219415 33615 222385
rect 58985 219415 59000 222385
rect 33600 219400 59000 219415
rect 60000 222600 98000 225600
rect 99000 225585 106000 225600
rect 99000 224115 99015 225585
rect 105985 224115 106000 225585
rect 99000 224100 106000 224115
rect 60000 215400 63000 222600
rect 68000 215400 71000 222600
rect 95000 215400 98000 222600
rect -132000 215385 123200 215400
rect -132000 212415 -32485 215385
rect -30505 212415 30515 215385
rect 32485 212415 123200 215385
rect -132000 212400 123200 212415
rect -132000 212200 -129000 212400
rect -110000 212200 -107000 212400
rect -105000 212200 -102000 212400
rect 60000 212200 63000 212400
rect 68000 212200 71000 212400
rect 95000 212200 98000 212400
rect 107000 212200 110000 212400
rect 120200 212200 123200 212400
rect -136800 212185 136800 212200
rect -136800 209215 -32485 212185
rect -30505 209215 30515 212185
rect 32485 209215 136800 212185
rect -136800 209200 136800 209215
rect -136800 206000 -133800 209200
rect -132000 206000 -129000 209200
rect -110000 206000 -107000 209200
rect -72600 208985 -47200 209000
rect -72600 207815 -72585 208985
rect -47215 207815 -47200 208985
rect -72600 207500 -47200 207815
rect -72600 207300 -69600 207500
rect -59800 207300 -56800 207500
rect -50200 207300 -47200 207500
rect 31800 208985 106000 209000
rect 31800 207815 99015 208985
rect 105985 207815 106000 208985
rect 31800 207500 106000 207815
rect -72600 207285 -47200 207300
rect -72600 204315 -62985 207285
rect -47215 204315 -47200 207285
rect -72600 204300 -47200 204315
rect -59800 204100 -56800 204300
rect -50200 204100 -47200 204300
rect -65000 204085 -47200 204100
rect -65000 201115 -62985 204085
rect -47215 201115 -47200 204085
rect -65000 201100 -47200 201115
rect -59800 200900 -56800 201100
rect -50200 200900 -47200 201100
rect -27600 207285 -2000 207300
rect -27600 204315 -27585 207285
rect -2015 204315 -2000 207285
rect -27600 204300 -2000 204315
rect -27600 204100 -24400 204300
rect -16000 204100 -13000 204300
rect -5000 204100 -2000 204300
rect -27600 204085 -2000 204100
rect -27600 201115 -27585 204085
rect -2015 201115 -2000 204085
rect 31800 202600 33400 207500
rect -27600 201100 -2000 201115
rect -27600 200900 -24400 201100
rect -16000 200900 -13000 201100
rect -5000 200900 -2000 201100
rect 23000 201100 33400 202600
rect 33600 207285 93000 207300
rect 33600 204315 33615 207285
rect 58985 204315 93000 207285
rect 107000 206000 110000 209200
rect 120200 206000 123200 209200
rect 133800 206000 136800 209200
rect 33600 204300 93000 204315
rect 33600 204100 36600 204300
rect 43200 204100 46200 204300
rect 52800 204100 55800 204300
rect 33600 204085 65000 204100
rect 33600 201115 33615 204085
rect 58985 201115 65000 204085
rect 33600 201100 65000 201115
rect 23000 200900 25000 201100
rect -65000 198000 -38000 200900
rect -27600 198000 25000 200900
rect 33600 200900 36600 201100
rect 43200 200900 46200 201100
rect 52800 200900 55800 201100
rect 33600 198000 65000 200900
rect -3000 180000 3000 198000
<< via3 >>
rect -72585 222615 -47215 225585
rect -72585 219415 -47215 222385
rect -27585 222615 -2015 225585
rect -27585 219415 -2015 222385
rect 33615 222615 58985 225585
rect 33615 219415 58985 222385
rect 99015 224115 105985 225585
rect -32485 212415 -30505 215385
rect 30515 212415 32485 215385
rect -32485 209215 -30505 212185
rect 30515 209215 32485 212185
rect -72585 207815 -47215 208985
rect 99015 207815 105985 208985
rect -62985 204315 -47215 207285
rect -62985 201115 -47215 204085
rect -27585 204315 -2015 207285
rect -27585 201115 -2015 204085
rect 33615 204315 58985 207285
rect 33615 201115 58985 204085
<< metal4 >>
rect -132000 222600 -102000 225600
rect -132000 215400 -129000 222600
rect -110000 215400 -107000 222600
rect -105000 215400 -102000 222600
rect -72600 225585 -47200 225600
rect -72600 222615 -72585 225585
rect -47215 222615 -47200 225585
rect -72600 222600 -47200 222615
rect -72600 222400 -69600 222600
rect -50200 222400 -47200 222600
rect -72600 222385 -47200 222400
rect -72600 219415 -72585 222385
rect -47215 219415 -47200 222385
rect -72600 219400 -47200 219415
rect -27600 225585 -2000 225600
rect -27600 222615 -27585 225585
rect -2015 222615 -2000 225585
rect -27600 222600 -2000 222615
rect -27600 222400 -24600 222600
rect -5000 222400 -2000 222600
rect -27600 222385 -2000 222400
rect -27600 219415 -27585 222385
rect -2015 219415 -2000 222385
rect -27600 219400 -2000 219415
rect 33600 225585 59000 225600
rect 33600 222615 33615 225585
rect 58985 222615 59000 225585
rect 33600 222600 59000 222615
rect 33600 222400 36600 222600
rect 56000 222400 59000 222600
rect 33600 222385 59000 222400
rect 33600 219415 33615 222385
rect 58985 219415 59000 222385
rect 33600 219400 59000 219415
rect 60000 222600 98000 225600
rect 99000 225585 106000 225600
rect 99000 224115 99015 225585
rect 105985 224115 106000 225585
rect 99000 224100 106000 224115
rect 60000 215400 63000 222600
rect 68000 215400 71000 222600
rect 95000 215400 98000 222600
rect -132000 215385 123200 215400
rect -132000 212415 -32485 215385
rect -30505 212415 30515 215385
rect 32485 212415 123200 215385
rect -132000 212400 123200 212415
rect -132000 212200 -129000 212400
rect -110000 212200 -107000 212400
rect -105000 212200 -102000 212400
rect 60000 212200 63000 212400
rect 68000 212200 71000 212400
rect 95000 212200 98000 212400
rect 107000 212200 110000 212400
rect 120200 212200 123200 212400
rect -136800 212185 136800 212200
rect -136800 209215 -32485 212185
rect -30505 209215 30515 212185
rect 32485 209215 136800 212185
rect -136800 209200 136800 209215
rect -136800 206000 -133800 209200
rect -132000 206000 -129000 209200
rect -110000 206000 -107000 209200
rect -72600 208985 -47200 209000
rect -72600 207815 -72585 208985
rect -47215 207815 -47200 208985
rect -72600 207500 -47200 207815
rect -72600 207300 -69600 207500
rect -59800 207300 -56800 207500
rect -50200 207300 -47200 207500
rect 31800 208985 106000 209000
rect 31800 207815 99015 208985
rect 105985 207815 106000 208985
rect 31800 207500 106000 207815
rect -72600 207285 -47200 207300
rect -72600 204315 -62985 207285
rect -47215 204315 -47200 207285
rect -72600 204300 -47200 204315
rect -59800 204100 -56800 204300
rect -50200 204100 -47200 204300
rect -65000 204085 -47200 204100
rect -65000 201115 -62985 204085
rect -47215 201115 -47200 204085
rect -65000 201100 -47200 201115
rect -59800 200900 -56800 201100
rect -50200 200900 -47200 201100
rect -27600 207285 -2000 207300
rect -27600 204315 -27585 207285
rect -2015 204315 -2000 207285
rect -27600 204300 -2000 204315
rect -27600 204100 -24400 204300
rect -16000 204100 -13000 204300
rect -5000 204100 -2000 204300
rect -27600 204085 -2000 204100
rect -27600 201115 -27585 204085
rect -2015 201115 -2000 204085
rect 31800 202600 33400 207500
rect -27600 201100 -2000 201115
rect -27600 200900 -24400 201100
rect -16000 200900 -13000 201100
rect -5000 200900 -2000 201100
rect 23000 201100 33400 202600
rect 33600 207285 93000 207300
rect 33600 204315 33615 207285
rect 58985 204315 93000 207285
rect 107000 206000 110000 209200
rect 120200 206000 123200 209200
rect 133800 206000 136800 209200
rect 33600 204300 93000 204315
rect 33600 204100 36600 204300
rect 43200 204100 46200 204300
rect 52800 204100 55800 204300
rect 33600 204085 65000 204100
rect 33600 201115 33615 204085
rect 58985 201115 65000 204085
rect 33600 201100 65000 201115
rect 23000 200900 25000 201100
rect -65000 198000 -38000 200900
rect -27600 198000 25000 200900
rect 33600 200900 36600 201100
rect 43200 200900 46200 201100
rect 52800 200900 55800 201100
rect 33600 198000 65000 200900
rect -3000 180000 3000 198000
<< via4 >>
rect -72585 222615 -47215 225585
rect -72585 219415 -47215 222385
rect -27585 222615 -2015 225585
rect -27585 219415 -2015 222385
rect 33615 222615 58985 225585
rect 33615 219415 58985 222385
rect 99015 224115 105985 225585
rect -32485 212415 -30505 215385
rect 30515 212415 32485 215385
rect -32485 209215 -30505 212185
rect 30515 209215 32485 212185
rect -72585 207815 -47215 208985
rect 99015 207815 105985 208985
rect -62985 204315 -47215 207285
rect -62985 201115 -47215 204085
rect -27585 204315 -2015 207285
rect -27585 201115 -2015 204085
rect 33615 204315 58985 207285
rect 33615 201115 58985 204085
<< metal5 >>
rect -132000 222600 -102000 225600
rect -132000 215400 -129000 222600
rect -110000 215400 -107000 222600
rect -105000 215400 -102000 222600
rect -72600 225585 -47200 225600
rect -72600 222615 -72585 225585
rect -47215 222615 -47200 225585
rect -72600 222600 -47200 222615
rect -72600 222400 -69600 222600
rect -50200 222400 -47200 222600
rect -72600 222385 -47200 222400
rect -72600 219415 -72585 222385
rect -47215 219415 -47200 222385
rect -72600 219400 -47200 219415
rect -27600 225585 -2000 225600
rect -27600 222615 -27585 225585
rect -2015 222615 -2000 225585
rect -27600 222600 -2000 222615
rect -27600 222400 -24600 222600
rect -5000 222400 -2000 222600
rect -27600 222385 -2000 222400
rect -27600 219415 -27585 222385
rect -2015 219415 -2000 222385
rect -27600 219400 -2000 219415
rect 33600 225585 59000 225600
rect 33600 222615 33615 225585
rect 58985 222615 59000 225585
rect 33600 222600 59000 222615
rect 33600 222400 36600 222600
rect 56000 222400 59000 222600
rect 33600 222385 59000 222400
rect 33600 219415 33615 222385
rect 58985 219415 59000 222385
rect 33600 219400 59000 219415
rect 60000 222600 98000 225600
rect 99000 225585 106000 225600
rect 99000 224115 99015 225585
rect 105985 224115 106000 225585
rect 99000 224100 106000 224115
rect 60000 215400 63000 222600
rect 68000 215400 71000 222600
rect 95000 215400 98000 222600
rect -132000 215385 123200 215400
rect -132000 212415 -32485 215385
rect -30505 212415 30515 215385
rect 32485 212415 123200 215385
rect -132000 212400 123200 212415
rect -132000 212200 -129000 212400
rect -110000 212200 -107000 212400
rect -105000 212200 -102000 212400
rect 60000 212200 63000 212400
rect 68000 212200 71000 212400
rect 95000 212200 98000 212400
rect 107000 212200 110000 212400
rect 120200 212200 123200 212400
rect -136800 212185 136800 212200
rect -136800 209215 -32485 212185
rect -30505 209215 30515 212185
rect 32485 209215 136800 212185
rect -136800 209200 136800 209215
rect -136800 206000 -133800 209200
rect -132000 206000 -129000 209200
rect -110000 206000 -107000 209200
rect -72600 208985 -47200 209000
rect -72600 207815 -72585 208985
rect -47215 207815 -47200 208985
rect -72600 207500 -47200 207815
rect -72600 207300 -69600 207500
rect -59800 207300 -56800 207500
rect -50200 207300 -47200 207500
rect 31800 208985 106000 209000
rect 31800 207815 99015 208985
rect 105985 207815 106000 208985
rect 31800 207500 106000 207815
rect -72600 207285 -47200 207300
rect -72600 204315 -62985 207285
rect -47215 204315 -47200 207285
rect -72600 204300 -47200 204315
rect -59800 204100 -56800 204300
rect -50200 204100 -47200 204300
rect -65000 204085 -47200 204100
rect -65000 201115 -62985 204085
rect -47215 201115 -47200 204085
rect -65000 201100 -47200 201115
rect -59800 200900 -56800 201100
rect -50200 200900 -47200 201100
rect -27600 207285 -2000 207300
rect -27600 204315 -27585 207285
rect -2015 204315 -2000 207285
rect -27600 204300 -2000 204315
rect -27600 204100 -24400 204300
rect -16000 204100 -13000 204300
rect -5000 204100 -2000 204300
rect -27600 204085 -2000 204100
rect -27600 201115 -27585 204085
rect -2015 201115 -2000 204085
rect 31800 202600 33400 207500
rect -27600 201100 -2000 201115
rect -27600 200900 -24400 201100
rect -16000 200900 -13000 201100
rect -5000 200900 -2000 201100
rect 23000 201100 33400 202600
rect 33600 207285 93000 207300
rect 33600 204315 33615 207285
rect 58985 204315 93000 207285
rect 107000 206000 110000 209200
rect 120200 206000 123200 209200
rect 133800 206000 136800 209200
rect 33600 204300 93000 204315
rect 33600 204100 36600 204300
rect 43200 204100 46200 204300
rect 52800 204100 55800 204300
rect 33600 204085 65000 204100
rect 33600 201115 33615 204085
rect 58985 201115 65000 204085
rect 33600 201100 65000 201115
rect 23000 200900 25000 201100
rect -65000 198000 -38000 200900
rect -27600 198000 25000 200900
rect 33600 200900 36600 201100
rect 43200 200900 46200 201100
rect 52800 200900 55800 201100
rect 33600 198000 65000 200900
rect -3000 180000 3000 198000
use core  core_0
timestamp 1667307464
transform -1 0 -1360 0 -1 208000
box 0 0 137760 208000
use core  core_1
timestamp 1667307464
transform 1 0 800 0 -1 208000
box 0 0 137760 208000
<< labels >>
rlabel metal5 -27600 222600 -2000 225600 3 GND
rlabel metal5 -132000 222600 -102000 225600 3 VH
rlabel metal5 -72600 222600 -47200 225600 3 Vout1
rlabel metal5 33600 222600 59000 225600 3 Vout2
<< end >>
