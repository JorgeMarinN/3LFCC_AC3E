** sch_path: /foss/designs/personal/converter/sim/converter.sch
**.subckt converter s1 s2 s3 s4 VP VN fc1_read fc2_read out
*.ipin s1
*.ipin s2
*.ipin s3
*.ipin s4
*.iopin VP
*.iopin VN
*.opin fc1_read
*.opin fc2_read
*.iopin out
X1v s1 s2 s3 s4 fc1_read fc2_read out VP VN power_stage
XC1 fc2_read fc1_read sky130_fd_pr__cap_mim_m3_1 W=30 L=30 MF=1978 m=1978
XC2 fc1_read fc2_read sky130_fd_pr__cap_mim_m3_2 W=30 L=30 VM=1978 m=1978
**.ends

* expanding   symbol:  power_stage.sym # of pins=9
** sym_path: /foss/designs/personal/converter/sim/power_stage.sym
** sch_path: /foss/designs/personal/converter/sim/power_stage.sch
.subckt power_stage  s1 s2 s3 s4 fc1 fc2 out VP VN
*.ipin s1
*.ipin s2
*.ipin s3
*.ipin s4
*.iopin VP
*.iopin VN
*.opin out
*.opin fc1
*.opin fc2
XM3 out s3 fc2 fc2 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=4.38 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2520 m=2520
XM2 out s2 fc1 fc1 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=4.38 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4512 m=4512
XM1 fc1 s1 VP VP sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=4.38 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4512 m=4512
XM4 fc2 s4 VN VN sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=4.38 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2520 m=2520
.ends

.end
