magic
tech sky130A
timestamp 1660617642
<< metal2 >>
rect -771 5206 5230 5419
<< via2 >>
rect 3400 7850 3850 26300
<< metal4 >>
rect 2800 27131 4350 27150
rect -578 26326 4350 27131
rect 2800 7097 4350 26326
rect 2800 6628 4360 7097
rect 2800 6176 4791 6628
rect 2800 6167 4542 6176
rect 2800 6150 4350 6167
rect 26273 3507 30785 4312
use nmos_waffle_36x36  nmos_waffle_36x36_0
timestamp 1624430562
transform 1 0 5374 0 1 5407
box -5400 -5400 25200 25200
<< labels >>
rlabel metal2 -739 5222 -336 5385 7 G
rlabel metal4 -457 26414 83 26978 7 D
rlabel metal4 30259 3665 30692 4164 3 S
<< end >>
