magic
tech sky130A
magscale 1 2
timestamp 1666540277
<< metal2 >>
rect 2300 586800 16000 587000
rect 567796 586800 581496 587000
rect 2300 568890 2500 586800
rect 2300 568710 2310 568890
rect 2490 568710 2500 568890
rect 2300 568700 2500 568710
rect 4300 586500 16400 586700
rect 567396 586500 579496 586700
rect 4300 568890 4500 586500
rect 4300 568710 4310 568890
rect 4490 568710 4500 568890
rect 4300 568700 4500 568710
rect 6300 586200 16800 586400
rect 566996 586200 577496 586400
rect 6300 568890 6500 586200
rect 6300 568710 6310 568890
rect 6490 568710 6500 568890
rect 6300 568700 6500 568710
rect 8300 585900 17200 586100
rect 566596 585900 575496 586100
rect 8300 568890 8500 585900
rect 8300 568710 8310 568890
rect 8490 568710 8500 568890
rect 8300 568700 8500 568710
rect 575296 568890 575496 585900
rect 575296 568710 575306 568890
rect 575486 568710 575496 568890
rect 575296 568700 575496 568710
rect 577296 568890 577496 586200
rect 577296 568710 577306 568890
rect 577486 568710 577496 568890
rect 577296 568700 577496 568710
rect 579296 568890 579496 586500
rect 579296 568710 579306 568890
rect 579486 568710 579496 568890
rect 579296 568700 579496 568710
rect 581296 568890 581496 586800
rect 581296 568710 581306 568890
rect 581486 568710 581496 568890
rect 581296 568700 581496 568710
<< via2 >>
rect 2310 568710 2490 568890
rect 4310 568710 4490 568890
rect 6310 568710 6490 568890
rect 8310 568710 8490 568890
rect 575306 568710 575486 568890
rect 577306 568710 577486 568890
rect 579306 568710 579486 568890
rect 581306 568710 581486 568890
<< metal3 >>
rect 68000 702000 170600 702300
rect 175894 702000 181000 702300
rect 68000 700000 181000 702000
rect 217294 702000 222294 702300
rect 227594 702000 291400 702300
rect 217294 700000 291400 702000
rect 292600 702000 323994 702300
rect 329294 702000 470394 702300
rect 292600 700000 470394 702000
rect 2300 568890 2500 568900
rect 2300 568710 2310 568890
rect 2490 568710 2500 568890
rect 2300 379000 2500 568710
rect 4300 568890 4500 568900
rect 4300 568710 4310 568890
rect 4490 568710 4500 568890
rect 0 377800 4000 379000
rect 0 335300 4000 335758
rect 4300 335300 4500 568710
rect 0 335100 4500 335300
rect 6300 568890 6500 568900
rect 6300 568710 6310 568890
rect 6490 568710 6500 568890
rect 0 334558 4000 335100
rect 0 292100 4000 292536
rect 6300 292100 6500 568710
rect 0 291900 6500 292100
rect 8300 568890 8500 568900
rect 8300 568710 8310 568890
rect 8490 568710 8500 568890
rect 0 291336 4000 291900
rect 0 249000 4000 249514
rect 8300 249000 8500 568710
rect 575296 568890 575496 568900
rect 575296 568710 575306 568890
rect 575486 568710 575496 568890
rect 575296 273000 575496 568710
rect 577296 568890 577496 568900
rect 577296 568710 577306 568890
rect 577486 568710 577496 568890
rect 577296 317400 577496 568710
rect 579296 568890 579496 568900
rect 579296 568710 579306 568890
rect 579486 568710 579496 568890
rect 579296 362600 579496 568710
rect 581296 568890 581496 568900
rect 581296 568710 581306 568890
rect 581486 568710 581496 568890
rect 581296 409524 581496 568710
rect 580000 408324 584000 409524
rect 580000 362600 584000 363101
rect 579296 362400 584000 362600
rect 580000 361901 584000 362400
rect 580000 317400 584000 317880
rect 577296 317200 584000 317400
rect 580000 316680 584000 317200
rect 580000 273000 584000 273458
rect 575296 272800 584000 273000
rect 580000 272258 584000 272800
rect 0 248800 8500 249000
rect 0 248314 4000 248800
<< metal4 >>
rect 68000 702000 170600 702300
rect 175894 702000 181000 702300
rect 68000 700000 181000 702000
rect 217294 702000 222294 702300
rect 227594 702000 291400 702300
rect 217294 700000 291400 702000
rect 292600 702000 323994 702300
rect 329294 702000 470394 702300
rect 292600 700000 470394 702000
<< metal5 >>
rect 68000 702000 170600 702300
rect 175894 702000 181000 702300
rect 68000 700000 181000 702000
rect 217294 702000 222294 702300
rect 227594 702000 291400 702300
rect 217294 700000 291400 702000
rect 292600 702000 323994 702300
rect 329294 702000 470394 702300
rect 292600 700000 470394 702000
<< comment >>
rect 16146 668718 75266 686998
rect 114158 669884 173278 688164
rect 232978 684470 292098 702750
rect 358410 657244 417530 675524
rect 506012 669496 565132 687776
use interleaved  interleaved_0
timestamp 1666538287
transform 1 0 292000 0 1 253200
box -276000 0 276000 448800
<< end >>
