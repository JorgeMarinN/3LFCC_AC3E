magic
tech sky130A
timestamp 1668349622
<< metal3 >>
rect 0 196 200 200
rect 0 4 4 196
rect 196 4 200 196
rect 0 0 200 4
<< rmetal3 >>
rect 80 80 120 120
<< via3 >>
rect 4 120 196 196
rect 4 80 80 120
rect 120 80 196 120
rect 4 4 196 80
<< metal4 >>
rect 0 196 200 200
rect 0 4 4 196
rect 196 4 200 196
rect 0 0 200 4
<< via4 >>
rect 21 120 179 179
rect 21 80 80 120
rect 80 80 120 120
rect 120 80 179 120
rect 21 21 179 80
<< metal5 >>
rect 0 179 200 200
rect 0 21 21 179
rect 179 21 200 179
rect 0 0 200 21
<< end >>
