magic
tech sky130A
timestamp 1668216541
<< metal3 >>
rect 0 25699 12980 25719
rect 0 22479 20 25699
rect 3240 25668 12980 25699
rect 3240 22510 9771 25668
rect 12929 22510 12980 25668
rect 3240 22479 12980 22510
rect 0 22459 12980 22479
<< via3 >>
rect 20 22479 3240 25699
rect 9771 22510 12929 25668
<< metal4 >>
rect 0 25699 3260 25719
rect 0 22479 20 25699
rect 3240 22479 3260 25699
rect 0 22459 3260 22479
rect 9751 25668 12980 25719
rect 9751 22510 9771 25668
rect 12929 22510 12980 25668
rect 9751 22459 12980 22510
<< via4 >>
rect 20 22479 3240 25699
rect 9771 22510 12929 25668
<< metal5 >>
rect 0 32179 40299 35439
rect 4860 27319 35439 30579
rect 0 25699 3260 25719
rect 0 22479 20 25699
rect 3240 22479 3260 25699
rect 0 22459 3260 22479
rect 4860 3260 8120 27319
rect 9720 25668 12980 25719
rect 9720 22510 9771 25668
rect 12929 22510 12980 25668
rect 9720 8120 12980 22510
rect 32179 8120 35439 27319
rect 9720 4860 35439 8120
rect 37039 3260 40299 32179
rect 4860 0 40299 3260
<< end >>
