magic
tech sky130A
magscale 1 2
timestamp 1663460437
<< error_p >>
rect -1675 2062 1675 2066
rect -1675 -2062 -1645 2062
rect -1609 1996 1609 2000
rect -1609 -1996 -1579 1996
rect 1579 -1996 1609 1996
rect -1609 -2000 1609 -1996
rect 1645 -2062 1675 2062
rect -1675 -2066 1675 -2062
<< nwell >>
rect -1645 -2062 1645 2062
<< mvpmos >>
rect -1551 -2000 -1451 2000
rect -1393 -2000 -1293 2000
rect -1235 -2000 -1135 2000
rect -1077 -2000 -977 2000
rect -919 -2000 -819 2000
rect -761 -2000 -661 2000
rect -603 -2000 -503 2000
rect -445 -2000 -345 2000
rect -287 -2000 -187 2000
rect -129 -2000 -29 2000
rect 29 -2000 129 2000
rect 187 -2000 287 2000
rect 345 -2000 445 2000
rect 503 -2000 603 2000
rect 661 -2000 761 2000
rect 819 -2000 919 2000
rect 977 -2000 1077 2000
rect 1135 -2000 1235 2000
rect 1293 -2000 1393 2000
rect 1451 -2000 1551 2000
<< mvpdiff >>
rect -1609 1988 -1551 2000
rect -1609 -1988 -1597 1988
rect -1563 -1988 -1551 1988
rect -1609 -2000 -1551 -1988
rect -1451 1988 -1393 2000
rect -1451 -1988 -1439 1988
rect -1405 -1988 -1393 1988
rect -1451 -2000 -1393 -1988
rect -1293 1988 -1235 2000
rect -1293 -1988 -1281 1988
rect -1247 -1988 -1235 1988
rect -1293 -2000 -1235 -1988
rect -1135 1988 -1077 2000
rect -1135 -1988 -1123 1988
rect -1089 -1988 -1077 1988
rect -1135 -2000 -1077 -1988
rect -977 1988 -919 2000
rect -977 -1988 -965 1988
rect -931 -1988 -919 1988
rect -977 -2000 -919 -1988
rect -819 1988 -761 2000
rect -819 -1988 -807 1988
rect -773 -1988 -761 1988
rect -819 -2000 -761 -1988
rect -661 1988 -603 2000
rect -661 -1988 -649 1988
rect -615 -1988 -603 1988
rect -661 -2000 -603 -1988
rect -503 1988 -445 2000
rect -503 -1988 -491 1988
rect -457 -1988 -445 1988
rect -503 -2000 -445 -1988
rect -345 1988 -287 2000
rect -345 -1988 -333 1988
rect -299 -1988 -287 1988
rect -345 -2000 -287 -1988
rect -187 1988 -129 2000
rect -187 -1988 -175 1988
rect -141 -1988 -129 1988
rect -187 -2000 -129 -1988
rect -29 1988 29 2000
rect -29 -1988 -17 1988
rect 17 -1988 29 1988
rect -29 -2000 29 -1988
rect 129 1988 187 2000
rect 129 -1988 141 1988
rect 175 -1988 187 1988
rect 129 -2000 187 -1988
rect 287 1988 345 2000
rect 287 -1988 299 1988
rect 333 -1988 345 1988
rect 287 -2000 345 -1988
rect 445 1988 503 2000
rect 445 -1988 457 1988
rect 491 -1988 503 1988
rect 445 -2000 503 -1988
rect 603 1988 661 2000
rect 603 -1988 615 1988
rect 649 -1988 661 1988
rect 603 -2000 661 -1988
rect 761 1988 819 2000
rect 761 -1988 773 1988
rect 807 -1988 819 1988
rect 761 -2000 819 -1988
rect 919 1988 977 2000
rect 919 -1988 931 1988
rect 965 -1988 977 1988
rect 919 -2000 977 -1988
rect 1077 1988 1135 2000
rect 1077 -1988 1089 1988
rect 1123 -1988 1135 1988
rect 1077 -2000 1135 -1988
rect 1235 1988 1293 2000
rect 1235 -1988 1247 1988
rect 1281 -1988 1293 1988
rect 1235 -2000 1293 -1988
rect 1393 1988 1451 2000
rect 1393 -1988 1405 1988
rect 1439 -1988 1451 1988
rect 1393 -2000 1451 -1988
rect 1551 1988 1609 2000
rect 1551 -1988 1563 1988
rect 1597 -1988 1609 1988
rect 1551 -2000 1609 -1988
<< mvpdiffc >>
rect -1597 -1988 -1563 1988
rect -1439 -1988 -1405 1988
rect -1281 -1988 -1247 1988
rect -1123 -1988 -1089 1988
rect -965 -1988 -931 1988
rect -807 -1988 -773 1988
rect -649 -1988 -615 1988
rect -491 -1988 -457 1988
rect -333 -1988 -299 1988
rect -175 -1988 -141 1988
rect -17 -1988 17 1988
rect 141 -1988 175 1988
rect 299 -1988 333 1988
rect 457 -1988 491 1988
rect 615 -1988 649 1988
rect 773 -1988 807 1988
rect 931 -1988 965 1988
rect 1089 -1988 1123 1988
rect 1247 -1988 1281 1988
rect 1405 -1988 1439 1988
rect 1563 -1988 1597 1988
<< poly >>
rect -1551 2000 -1451 2026
rect -1393 2000 -1293 2026
rect -1235 2000 -1135 2026
rect -1077 2000 -977 2026
rect -919 2000 -819 2026
rect -761 2000 -661 2026
rect -603 2000 -503 2026
rect -445 2000 -345 2026
rect -287 2000 -187 2026
rect -129 2000 -29 2026
rect 29 2000 129 2026
rect 187 2000 287 2026
rect 345 2000 445 2026
rect 503 2000 603 2026
rect 661 2000 761 2026
rect 819 2000 919 2026
rect 977 2000 1077 2026
rect 1135 2000 1235 2026
rect 1293 2000 1393 2026
rect 1451 2000 1551 2026
rect -1551 -2026 -1451 -2000
rect -1393 -2026 -1293 -2000
rect -1235 -2026 -1135 -2000
rect -1077 -2026 -977 -2000
rect -919 -2026 -819 -2000
rect -761 -2026 -661 -2000
rect -603 -2026 -503 -2000
rect -445 -2026 -345 -2000
rect -287 -2026 -187 -2000
rect -129 -2026 -29 -2000
rect 29 -2026 129 -2000
rect 187 -2026 287 -2000
rect 345 -2026 445 -2000
rect 503 -2026 603 -2000
rect 661 -2026 761 -2000
rect 819 -2026 919 -2000
rect 977 -2026 1077 -2000
rect 1135 -2026 1235 -2000
rect 1293 -2026 1393 -2000
rect 1451 -2026 1551 -2000
<< locali >>
rect -1597 1988 -1563 2004
rect -1597 -2004 -1563 -1988
rect -1439 1988 -1405 2004
rect -1439 -2004 -1405 -1988
rect -1281 1988 -1247 2004
rect -1281 -2004 -1247 -1988
rect -1123 1988 -1089 2004
rect -1123 -2004 -1089 -1988
rect -965 1988 -931 2004
rect -965 -2004 -931 -1988
rect -807 1988 -773 2004
rect -807 -2004 -773 -1988
rect -649 1988 -615 2004
rect -649 -2004 -615 -1988
rect -491 1988 -457 2004
rect -491 -2004 -457 -1988
rect -333 1988 -299 2004
rect -333 -2004 -299 -1988
rect -175 1988 -141 2004
rect -175 -2004 -141 -1988
rect -17 1988 17 2004
rect -17 -2004 17 -1988
rect 141 1988 175 2004
rect 141 -2004 175 -1988
rect 299 1988 333 2004
rect 299 -2004 333 -1988
rect 457 1988 491 2004
rect 457 -2004 491 -1988
rect 615 1988 649 2004
rect 615 -2004 649 -1988
rect 773 1988 807 2004
rect 773 -2004 807 -1988
rect 931 1988 965 2004
rect 931 -2004 965 -1988
rect 1089 1988 1123 2004
rect 1089 -2004 1123 -1988
rect 1247 1988 1281 2004
rect 1247 -2004 1281 -1988
rect 1405 1988 1439 2004
rect 1405 -2004 1439 -1988
rect 1563 1988 1597 2004
rect 1563 -2004 1597 -1988
<< viali >>
rect -1597 -1988 -1563 1988
rect -1439 -1988 -1405 1988
rect -1281 -1988 -1247 1988
rect -1123 -1988 -1089 1988
rect -965 -1988 -931 1988
rect -807 -1988 -773 1988
rect -649 -1988 -615 1988
rect -491 -1988 -457 1988
rect -333 -1988 -299 1988
rect -175 -1988 -141 1988
rect -17 -1988 17 1988
rect 141 -1988 175 1988
rect 299 -1988 333 1988
rect 457 -1988 491 1988
rect 615 -1988 649 1988
rect 773 -1988 807 1988
rect 931 -1988 965 1988
rect 1089 -1988 1123 1988
rect 1247 -1988 1281 1988
rect 1405 -1988 1439 1988
rect 1563 -1988 1597 1988
<< metal1 >>
rect -1603 1988 -1557 2000
rect -1603 -1988 -1597 1988
rect -1563 -1988 -1557 1988
rect -1603 -2000 -1557 -1988
rect -1445 1988 -1399 2000
rect -1445 -1988 -1439 1988
rect -1405 -1988 -1399 1988
rect -1445 -2000 -1399 -1988
rect -1287 1988 -1241 2000
rect -1287 -1988 -1281 1988
rect -1247 -1988 -1241 1988
rect -1287 -2000 -1241 -1988
rect -1129 1988 -1083 2000
rect -1129 -1988 -1123 1988
rect -1089 -1988 -1083 1988
rect -1129 -2000 -1083 -1988
rect -971 1988 -925 2000
rect -971 -1988 -965 1988
rect -931 -1988 -925 1988
rect -971 -2000 -925 -1988
rect -813 1988 -767 2000
rect -813 -1988 -807 1988
rect -773 -1988 -767 1988
rect -813 -2000 -767 -1988
rect -655 1988 -609 2000
rect -655 -1988 -649 1988
rect -615 -1988 -609 1988
rect -655 -2000 -609 -1988
rect -497 1988 -451 2000
rect -497 -1988 -491 1988
rect -457 -1988 -451 1988
rect -497 -2000 -451 -1988
rect -339 1988 -293 2000
rect -339 -1988 -333 1988
rect -299 -1988 -293 1988
rect -339 -2000 -293 -1988
rect -181 1988 -135 2000
rect -181 -1988 -175 1988
rect -141 -1988 -135 1988
rect -181 -2000 -135 -1988
rect -23 1988 23 2000
rect -23 -1988 -17 1988
rect 17 -1988 23 1988
rect -23 -2000 23 -1988
rect 135 1988 181 2000
rect 135 -1988 141 1988
rect 175 -1988 181 1988
rect 135 -2000 181 -1988
rect 293 1988 339 2000
rect 293 -1988 299 1988
rect 333 -1988 339 1988
rect 293 -2000 339 -1988
rect 451 1988 497 2000
rect 451 -1988 457 1988
rect 491 -1988 497 1988
rect 451 -2000 497 -1988
rect 609 1988 655 2000
rect 609 -1988 615 1988
rect 649 -1988 655 1988
rect 609 -2000 655 -1988
rect 767 1988 813 2000
rect 767 -1988 773 1988
rect 807 -1988 813 1988
rect 767 -2000 813 -1988
rect 925 1988 971 2000
rect 925 -1988 931 1988
rect 965 -1988 971 1988
rect 925 -2000 971 -1988
rect 1083 1988 1129 2000
rect 1083 -1988 1089 1988
rect 1123 -1988 1129 1988
rect 1083 -2000 1129 -1988
rect 1241 1988 1287 2000
rect 1241 -1988 1247 1988
rect 1281 -1988 1287 1988
rect 1241 -2000 1287 -1988
rect 1399 1988 1445 2000
rect 1399 -1988 1405 1988
rect 1439 -1988 1445 1988
rect 1399 -2000 1445 -1988
rect 1557 1988 1603 2000
rect 1557 -1988 1563 1988
rect 1597 -1988 1603 1988
rect 1557 -2000 1603 -1988
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 20 l .5 m 1 nf 20 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
