magic
tech sky130A
timestamp 1666497650
<< checkpaint >>
rect -966 167866 137946 169966
rect -966 163914 137966 167866
rect 69034 163834 137966 163914
rect -1966 119094 11536 142326
rect -1966 77623 11536 100855
<< metal3 >>
rect 1000 166980 68990 167000
rect 1000 166020 1020 166980
rect 68970 166020 68990 166980
rect 1000 165880 68990 166020
rect 71180 166980 135980 168000
rect 71180 166020 71200 166980
rect 135960 166020 135980 166980
rect 71180 166000 135980 166020
rect 1000 165720 2000 165880
rect 4190 165720 5190 165880
rect 7380 165720 8380 165880
rect 10570 165720 11570 165880
rect 13760 165720 14760 165880
rect 16950 165720 17950 165880
rect 20140 165720 21140 165880
rect 23330 165720 24330 165880
rect 26520 165720 27520 165880
rect 29710 165720 30710 165880
rect 32900 165720 33900 165880
rect 36090 165720 37090 165880
rect 39280 165720 40280 165880
rect 42470 165720 43470 165880
rect 45660 165720 46660 165880
rect 48850 165720 49850 165880
rect 52040 165720 53040 165880
rect 55230 165720 56230 165880
rect 58420 165720 59420 165880
rect 61610 165720 62610 165880
rect 64800 165720 65800 165880
rect 67990 165720 68990 165880
rect 71180 165720 72180 165800
rect 74370 165720 75370 165800
rect 77560 165720 78560 165800
rect 80750 165720 81750 165800
rect 83940 165720 84940 165800
rect 87130 165720 88130 165800
rect 90320 165720 91320 165800
rect 93510 165720 94510 165800
rect 96700 165720 97700 165800
rect 99890 165720 100890 165800
rect 103080 165720 104080 165800
rect 106270 165720 107270 165800
rect 109460 165720 110460 165800
rect 112650 165720 113650 165800
rect 115840 165720 116840 165800
rect 119030 165720 120030 165800
rect 122220 165720 123220 165800
rect 125410 165720 126410 165800
rect 128600 165720 129600 165800
rect 131790 165720 132790 165800
rect 134980 165720 135980 165800
rect 0 164690 3030 165720
rect 3190 164690 6220 165720
rect 6380 164690 9410 165720
rect 9570 164690 12600 165720
rect 12760 164690 15790 165720
rect 15950 164690 18980 165720
rect 19140 164690 22170 165720
rect 22330 164690 25360 165720
rect 25520 164690 28550 165720
rect 28710 164690 31740 165720
rect 31900 164690 34930 165720
rect 35090 164690 38120 165720
rect 38280 164690 41310 165720
rect 41470 164690 44500 165720
rect 44660 164690 47690 165720
rect 47850 164690 50880 165720
rect 51040 164690 54070 165720
rect 54230 164690 57260 165720
rect 57420 164690 60450 165720
rect 60610 164690 63640 165720
rect 63800 164690 66830 165720
rect 66990 164690 70020 165720
rect 70180 164690 73210 165720
rect 73370 164690 76400 165720
rect 76560 164690 79590 165720
rect 79750 164690 82780 165720
rect 82940 164690 85970 165720
rect 86130 164690 89160 165720
rect 89320 164690 92350 165720
rect 92510 164690 95540 165720
rect 95700 164690 98730 165720
rect 98890 164690 101920 165720
rect 102080 164690 105110 165720
rect 105270 164690 108300 165720
rect 108460 164690 111490 165720
rect 111650 164690 114680 165720
rect 114840 164690 117870 165720
rect 118030 164690 121060 165720
rect 121220 164690 124250 165720
rect 124410 164690 127440 165720
rect 127600 164690 130630 165720
rect 130790 164690 133820 165720
rect 133980 164690 137010 165720
rect 0 163690 137170 164690
rect 0 162690 3030 163690
rect 3190 162690 6220 163690
rect 6380 162690 9410 163690
rect 9570 162690 12600 163690
rect 12760 162690 15790 163690
rect 15950 162690 18980 163690
rect 19140 162690 22170 163690
rect 22330 162690 25360 163690
rect 25520 162690 28550 163690
rect 28710 162690 31740 163690
rect 31900 162690 34930 163690
rect 35090 162690 38120 163690
rect 38280 162690 41310 163690
rect 41470 162690 44500 163690
rect 44660 162690 47690 163690
rect 47850 162690 50880 163690
rect 51040 162690 54070 163690
rect 54230 162690 57260 163690
rect 57420 162690 60450 163690
rect 60610 162690 63640 163690
rect 63800 162690 66830 163690
rect 66990 162690 70020 163690
rect 70180 162690 73210 163690
rect 73370 162690 76400 163690
rect 76560 162690 79590 163690
rect 79750 162690 82780 163690
rect 82940 162690 85970 163690
rect 86130 162690 89160 163690
rect 89320 162690 92350 163690
rect 92510 162690 95540 163690
rect 95700 162690 98730 163690
rect 98890 162690 101920 163690
rect 102080 162690 105110 163690
rect 105270 162690 108300 163690
rect 108460 162690 111490 163690
rect 111650 162690 114680 163690
rect 114840 162690 117870 163690
rect 118030 162690 121060 163690
rect 121220 162690 124250 163690
rect 124410 162690 127440 163690
rect 127600 162690 130630 163690
rect 130790 162690 133820 163690
rect 133980 162690 137010 163690
rect 1000 162530 2000 162690
rect 4190 162530 5190 162690
rect 7380 162530 8380 162690
rect 10570 162530 11570 162690
rect 13760 162530 14760 162690
rect 16950 162530 17950 162690
rect 20140 162530 21140 162690
rect 23330 162530 24330 162690
rect 26520 162530 27520 162690
rect 29710 162530 30710 162690
rect 32900 162530 33900 162690
rect 36090 162530 37090 162690
rect 39280 162530 40280 162690
rect 42470 162530 43470 162690
rect 45660 162530 46660 162690
rect 48850 162530 49850 162690
rect 52040 162530 53040 162690
rect 55230 162530 56230 162690
rect 58420 162530 59420 162690
rect 61610 162530 62610 162690
rect 64800 162530 65800 162690
rect 67990 162530 68990 162690
rect 71180 162530 72180 162690
rect 74370 162530 75370 162690
rect 77560 162530 78560 162690
rect 80750 162530 81750 162690
rect 83940 162530 84940 162690
rect 87130 162530 88130 162690
rect 90320 162530 91320 162690
rect 93510 162530 94510 162690
rect 96700 162530 97700 162690
rect 99890 162530 100890 162690
rect 103080 162530 104080 162690
rect 106270 162530 107270 162690
rect 109460 162530 110460 162690
rect 112650 162530 113650 162690
rect 115840 162530 116840 162690
rect 119030 162530 120030 162690
rect 122220 162530 123220 162690
rect 125410 162530 126410 162690
rect 128600 162530 129600 162690
rect 131790 162530 132790 162690
rect 134980 162530 135980 162690
rect 0 161500 3030 162530
rect 3190 161500 6220 162530
rect 6380 161500 9410 162530
rect 9570 161500 12600 162530
rect 12760 161500 15790 162530
rect 15950 161500 18980 162530
rect 19140 161500 22170 162530
rect 22330 161500 25360 162530
rect 25520 161500 28550 162530
rect 28710 161500 31740 162530
rect 31900 161500 34930 162530
rect 35090 161500 38120 162530
rect 38280 161500 41310 162530
rect 41470 161500 44500 162530
rect 44660 161500 47690 162530
rect 47850 161500 50880 162530
rect 51040 161500 54070 162530
rect 54230 161500 57260 162530
rect 57420 161500 60450 162530
rect 60610 161500 63640 162530
rect 63800 161500 66830 162530
rect 66990 161500 70020 162530
rect 70180 161500 73210 162530
rect 73370 161500 76400 162530
rect 76560 161500 79590 162530
rect 79750 161500 82780 162530
rect 82940 161500 85970 162530
rect 86130 161500 89160 162530
rect 89320 161500 92350 162530
rect 92510 161500 95540 162530
rect 95700 161500 98730 162530
rect 98890 161500 101920 162530
rect 102080 161500 105110 162530
rect 105270 161500 108300 162530
rect 108460 161500 111490 162530
rect 111650 161500 114680 162530
rect 114840 161500 117870 162530
rect 118030 161500 121060 162530
rect 121220 161500 124250 162530
rect 124410 161500 127440 162530
rect 127600 161500 130630 162530
rect 130790 161500 133820 162530
rect 133980 161500 137010 162530
rect 0 160500 137170 161500
rect 0 159500 3030 160500
rect 3190 159500 6220 160500
rect 6380 159500 9410 160500
rect 9570 159500 12600 160500
rect 12760 159500 15790 160500
rect 15950 159500 18980 160500
rect 19140 159500 22170 160500
rect 22330 159500 25360 160500
rect 25520 159500 28550 160500
rect 28710 159500 31740 160500
rect 31900 159500 34930 160500
rect 35090 159500 38120 160500
rect 38280 159500 41310 160500
rect 41470 159500 44500 160500
rect 44660 159500 47690 160500
rect 47850 159500 50880 160500
rect 51040 159500 54070 160500
rect 54230 159500 57260 160500
rect 57420 159500 60450 160500
rect 60610 159500 63640 160500
rect 63800 159500 66830 160500
rect 66990 159500 70020 160500
rect 70180 159500 73210 160500
rect 73370 159500 76400 160500
rect 76560 159500 79590 160500
rect 79750 159500 82780 160500
rect 82940 159500 85970 160500
rect 86130 159500 89160 160500
rect 89320 159500 92350 160500
rect 92510 159500 95540 160500
rect 95700 159500 98730 160500
rect 98890 159500 101920 160500
rect 102080 159500 105110 160500
rect 105270 159500 108300 160500
rect 108460 159500 111490 160500
rect 111650 159500 114680 160500
rect 114840 159500 117870 160500
rect 118030 159500 121060 160500
rect 121220 159500 124250 160500
rect 124410 159500 127440 160500
rect 127600 159500 130630 160500
rect 130790 159500 133820 160500
rect 133980 159500 137010 160500
rect 1000 159340 2000 159500
rect 4190 159340 5190 159500
rect 7380 159340 8380 159500
rect 10570 159340 11570 159500
rect 13760 159340 14760 159500
rect 16950 159340 17950 159500
rect 20140 159340 21140 159500
rect 23330 159340 24330 159500
rect 26520 159340 27520 159500
rect 29710 159340 30710 159500
rect 32900 159340 33900 159500
rect 36090 159340 37090 159500
rect 39280 159340 40280 159500
rect 42470 159340 43470 159500
rect 45660 159340 46660 159500
rect 48850 159340 49850 159500
rect 52040 159340 53040 159500
rect 55230 159340 56230 159500
rect 58420 159340 59420 159500
rect 61610 159340 62610 159500
rect 64800 159340 65800 159500
rect 67990 159340 68990 159500
rect 71180 159340 72180 159500
rect 74370 159340 75370 159500
rect 77560 159340 78560 159500
rect 80750 159340 81750 159500
rect 83940 159340 84940 159500
rect 87130 159340 88130 159500
rect 90320 159340 91320 159500
rect 93510 159340 94510 159500
rect 96700 159340 97700 159500
rect 99890 159340 100890 159500
rect 103080 159340 104080 159500
rect 106270 159340 107270 159500
rect 109460 159340 110460 159500
rect 112650 159340 113650 159500
rect 115840 159340 116840 159500
rect 119030 159340 120030 159500
rect 122220 159340 123220 159500
rect 125410 159340 126410 159500
rect 128600 159340 129600 159500
rect 131790 159340 132790 159500
rect 134980 159340 135980 159500
rect 0 158310 3030 159340
rect 3190 158310 6220 159340
rect 6380 158310 9410 159340
rect 9570 158310 12600 159340
rect 12760 158310 15790 159340
rect 15950 158310 18980 159340
rect 19140 158310 22170 159340
rect 22330 158310 25360 159340
rect 25520 158310 28550 159340
rect 28710 158310 31740 159340
rect 31900 158310 34930 159340
rect 35090 158310 38120 159340
rect 38280 158310 41310 159340
rect 41470 158310 44500 159340
rect 44660 158310 47690 159340
rect 47850 158310 50880 159340
rect 51040 158310 54070 159340
rect 54230 158310 57260 159340
rect 57420 158310 60450 159340
rect 60610 158310 63640 159340
rect 63800 158310 66830 159340
rect 66990 158310 70020 159340
rect 70180 158310 73210 159340
rect 73370 158310 76400 159340
rect 76560 158310 79590 159340
rect 79750 158310 82780 159340
rect 82940 158310 85970 159340
rect 86130 158310 89160 159340
rect 89320 158310 92350 159340
rect 92510 158310 95540 159340
rect 95700 158310 98730 159340
rect 98890 158310 101920 159340
rect 102080 158310 105110 159340
rect 105270 158310 108300 159340
rect 108460 158310 111490 159340
rect 111650 158310 114680 159340
rect 114840 158310 117870 159340
rect 118030 158310 121060 159340
rect 121220 158310 124250 159340
rect 124410 158310 127440 159340
rect 127600 158310 130630 159340
rect 130790 158310 133820 159340
rect 133980 158310 137010 159340
rect 0 157310 137170 158310
rect 0 156310 3030 157310
rect 3190 156310 6220 157310
rect 6380 156310 9410 157310
rect 9570 156310 12600 157310
rect 12760 156310 15790 157310
rect 15950 156310 18980 157310
rect 19140 156310 22170 157310
rect 22330 156310 25360 157310
rect 25520 156310 28550 157310
rect 28710 156310 31740 157310
rect 31900 156310 34930 157310
rect 35090 156310 38120 157310
rect 38280 156310 41310 157310
rect 41470 156310 44500 157310
rect 44660 156310 47690 157310
rect 47850 156310 50880 157310
rect 51040 156310 54070 157310
rect 54230 156310 57260 157310
rect 57420 156310 60450 157310
rect 60610 156310 63640 157310
rect 63800 156310 66830 157310
rect 66990 156310 70020 157310
rect 70180 156310 73210 157310
rect 73370 156310 76400 157310
rect 76560 156310 79590 157310
rect 79750 156310 82780 157310
rect 82940 156310 85970 157310
rect 86130 156310 89160 157310
rect 89320 156310 92350 157310
rect 92510 156310 95540 157310
rect 95700 156310 98730 157310
rect 98890 156310 101920 157310
rect 102080 156310 105110 157310
rect 105270 156310 108300 157310
rect 108460 156310 111490 157310
rect 111650 156310 114680 157310
rect 114840 156310 117870 157310
rect 118030 156310 121060 157310
rect 121220 156310 124250 157310
rect 124410 156310 127440 157310
rect 127600 156310 130630 157310
rect 130790 156310 133820 157310
rect 133980 156310 137010 157310
rect 1000 156150 2000 156310
rect 4190 156150 5190 156310
rect 7380 156150 8380 156310
rect 10570 156150 11570 156310
rect 13760 156150 14760 156310
rect 16950 156150 17950 156310
rect 20140 156150 21140 156310
rect 23330 156150 24330 156310
rect 26520 156150 27520 156310
rect 29710 156150 30710 156310
rect 32900 156150 33900 156310
rect 36090 156150 37090 156310
rect 39280 156150 40280 156310
rect 42470 156150 43470 156310
rect 45660 156150 46660 156310
rect 48850 156150 49850 156310
rect 52040 156150 53040 156310
rect 55230 156150 56230 156310
rect 58420 156150 59420 156310
rect 61610 156150 62610 156310
rect 64800 156150 65800 156310
rect 67990 156150 68990 156310
rect 71180 156150 72180 156310
rect 74370 156150 75370 156310
rect 77560 156150 78560 156310
rect 80750 156150 81750 156310
rect 83940 156150 84940 156310
rect 87130 156150 88130 156310
rect 90320 156150 91320 156310
rect 93510 156150 94510 156310
rect 96700 156150 97700 156310
rect 99890 156150 100890 156310
rect 103080 156150 104080 156310
rect 106270 156150 107270 156310
rect 109460 156150 110460 156310
rect 112650 156150 113650 156310
rect 115840 156150 116840 156310
rect 119030 156150 120030 156310
rect 122220 156150 123220 156310
rect 125410 156150 126410 156310
rect 128600 156150 129600 156310
rect 131790 156150 132790 156310
rect 134980 156150 135980 156310
rect 0 155120 3030 156150
rect 3190 155120 6220 156150
rect 6380 155120 9410 156150
rect 9570 155120 12600 156150
rect 12760 155120 15790 156150
rect 15950 155120 18980 156150
rect 19140 155120 22170 156150
rect 22330 155120 25360 156150
rect 25520 155120 28550 156150
rect 28710 155120 31740 156150
rect 31900 155120 34930 156150
rect 35090 155120 38120 156150
rect 38280 155120 41310 156150
rect 41470 155120 44500 156150
rect 44660 155120 47690 156150
rect 47850 155120 50880 156150
rect 51040 155120 54070 156150
rect 54230 155120 57260 156150
rect 57420 155120 60450 156150
rect 60610 155120 63640 156150
rect 63800 155120 66830 156150
rect 66990 155120 70020 156150
rect 70180 155120 73210 156150
rect 73370 155120 76400 156150
rect 76560 155120 79590 156150
rect 79750 155120 82780 156150
rect 82940 155120 85970 156150
rect 86130 155120 89160 156150
rect 89320 155120 92350 156150
rect 92510 155120 95540 156150
rect 95700 155120 98730 156150
rect 98890 155120 101920 156150
rect 102080 155120 105110 156150
rect 105270 155120 108300 156150
rect 108460 155120 111490 156150
rect 111650 155120 114680 156150
rect 114840 155120 117870 156150
rect 118030 155120 121060 156150
rect 121220 155120 124250 156150
rect 124410 155120 127440 156150
rect 127600 155120 130630 156150
rect 130790 155120 133820 156150
rect 133980 155120 137010 156150
rect 0 154120 137170 155120
rect 0 153120 3030 154120
rect 3190 153120 6220 154120
rect 6380 153120 9410 154120
rect 9570 153120 12600 154120
rect 12760 153120 15790 154120
rect 15950 153120 18980 154120
rect 19140 153120 22170 154120
rect 22330 153120 25360 154120
rect 25520 153120 28550 154120
rect 28710 153120 31740 154120
rect 31900 153120 34930 154120
rect 35090 153120 38120 154120
rect 38280 153120 41310 154120
rect 41470 153120 44500 154120
rect 44660 153120 47690 154120
rect 47850 153120 50880 154120
rect 51040 153120 54070 154120
rect 54230 153120 57260 154120
rect 57420 153120 60450 154120
rect 60610 153120 63640 154120
rect 63800 153120 66830 154120
rect 66990 153120 70020 154120
rect 70180 153120 73210 154120
rect 73370 153120 76400 154120
rect 76560 153120 79590 154120
rect 79750 153120 82780 154120
rect 82940 153120 85970 154120
rect 86130 153120 89160 154120
rect 89320 153120 92350 154120
rect 92510 153120 95540 154120
rect 95700 153120 98730 154120
rect 98890 153120 101920 154120
rect 102080 153120 105110 154120
rect 105270 153120 108300 154120
rect 108460 153120 111490 154120
rect 111650 153120 114680 154120
rect 114840 153120 117870 154120
rect 118030 153120 121060 154120
rect 121220 153120 124250 154120
rect 124410 153120 127440 154120
rect 127600 153120 130630 154120
rect 130790 153120 133820 154120
rect 133980 153120 137010 154120
rect 1000 152960 2000 153120
rect 4190 152960 5190 153120
rect 7380 152960 8380 153120
rect 10570 152960 11570 153120
rect 13760 152960 14760 153120
rect 16950 152960 17950 153120
rect 20140 152960 21140 153120
rect 23330 152960 24330 153120
rect 26520 152960 27520 153120
rect 29710 152960 30710 153120
rect 32900 152960 33900 153120
rect 36090 152960 37090 153120
rect 39280 152960 40280 153120
rect 42470 152960 43470 153120
rect 45660 152960 46660 153120
rect 48850 152960 49850 153120
rect 52040 152960 53040 153120
rect 55230 152960 56230 153120
rect 58420 152960 59420 153120
rect 61610 152960 62610 153120
rect 64800 152960 65800 153120
rect 67990 152960 68990 153120
rect 71180 152960 72180 153120
rect 74370 152960 75370 153120
rect 77560 152960 78560 153120
rect 80750 152960 81750 153120
rect 83940 152960 84940 153120
rect 87130 152960 88130 153120
rect 90320 152960 91320 153120
rect 93510 152960 94510 153120
rect 96700 152960 97700 153120
rect 99890 152960 100890 153120
rect 103080 152960 104080 153120
rect 106270 152960 107270 153120
rect 109460 152960 110460 153120
rect 112650 152960 113650 153120
rect 115840 152960 116840 153120
rect 119030 152960 120030 153120
rect 122220 152960 123220 153120
rect 125410 152960 126410 153120
rect 128600 152960 129600 153120
rect 131790 152960 132790 153120
rect 134980 152960 135980 153120
rect 0 151930 3030 152960
rect 3190 151930 6220 152960
rect 6380 151930 9410 152960
rect 9570 151930 12600 152960
rect 12760 151930 15790 152960
rect 15950 151930 18980 152960
rect 19140 151930 22170 152960
rect 22330 151930 25360 152960
rect 25520 151930 28550 152960
rect 28710 151930 31740 152960
rect 31900 151930 34930 152960
rect 35090 151930 38120 152960
rect 38280 151930 41310 152960
rect 41470 151930 44500 152960
rect 44660 151930 47690 152960
rect 47850 151930 50880 152960
rect 51040 151930 54070 152960
rect 54230 151930 57260 152960
rect 57420 151930 60450 152960
rect 60610 151930 63640 152960
rect 63800 151930 66830 152960
rect 66990 151930 70020 152960
rect 70180 151930 73210 152960
rect 73370 151930 76400 152960
rect 76560 151930 79590 152960
rect 79750 151930 82780 152960
rect 82940 151930 85970 152960
rect 86130 151930 89160 152960
rect 89320 151930 92350 152960
rect 92510 151930 95540 152960
rect 95700 151930 98730 152960
rect 98890 151930 101920 152960
rect 102080 151930 105110 152960
rect 105270 151930 108300 152960
rect 108460 151930 111490 152960
rect 111650 151930 114680 152960
rect 114840 151930 117870 152960
rect 118030 151930 121060 152960
rect 121220 151930 124250 152960
rect 124410 151930 127440 152960
rect 127600 151930 130630 152960
rect 130790 151930 133820 152960
rect 133980 151930 137010 152960
rect 0 150930 137170 151930
rect 0 149930 3030 150930
rect 3190 149930 6220 150930
rect 6380 149930 9410 150930
rect 9570 149930 12600 150930
rect 12760 149930 15790 150930
rect 15950 149930 18980 150930
rect 19140 149930 22170 150930
rect 22330 149930 25360 150930
rect 25520 149930 28550 150930
rect 28710 149930 31740 150930
rect 31900 149930 34930 150930
rect 35090 149930 38120 150930
rect 38280 149930 41310 150930
rect 41470 149930 44500 150930
rect 44660 149930 47690 150930
rect 47850 149930 50880 150930
rect 51040 149930 54070 150930
rect 54230 149930 57260 150930
rect 57420 149930 60450 150930
rect 60610 149930 63640 150930
rect 63800 149930 66830 150930
rect 66990 149930 70020 150930
rect 70180 149930 73210 150930
rect 73370 149930 76400 150930
rect 76560 149930 79590 150930
rect 79750 149930 82780 150930
rect 82940 149930 85970 150930
rect 86130 149930 89160 150930
rect 89320 149930 92350 150930
rect 92510 149930 95540 150930
rect 95700 149930 98730 150930
rect 98890 149930 101920 150930
rect 102080 149930 105110 150930
rect 105270 149930 108300 150930
rect 108460 149930 111490 150930
rect 111650 149930 114680 150930
rect 114840 149930 117870 150930
rect 118030 149930 121060 150930
rect 121220 149930 124250 150930
rect 124410 149930 127440 150930
rect 127600 149930 130630 150930
rect 130790 149930 133820 150930
rect 133980 149930 137010 150930
rect 1000 149770 2000 149930
rect 4190 149770 5190 149930
rect 7380 149770 8380 149930
rect 10570 149770 11570 149930
rect 13760 149770 14760 149930
rect 16950 149770 17950 149930
rect 20140 149770 21140 149930
rect 23330 149770 24330 149930
rect 26520 149770 27520 149930
rect 29710 149770 30710 149930
rect 32900 149770 33900 149930
rect 36090 149770 37090 149930
rect 39280 149770 40280 149930
rect 42470 149770 43470 149930
rect 45660 149770 46660 149930
rect 48850 149770 49850 149930
rect 52040 149770 53040 149930
rect 55230 149770 56230 149930
rect 58420 149770 59420 149930
rect 61610 149770 62610 149930
rect 64800 149770 65800 149930
rect 67990 149770 68990 149930
rect 71180 149770 72180 149930
rect 74370 149770 75370 149930
rect 77560 149770 78560 149930
rect 80750 149770 81750 149930
rect 83940 149770 84940 149930
rect 87130 149770 88130 149930
rect 90320 149770 91320 149930
rect 93510 149770 94510 149930
rect 96700 149770 97700 149930
rect 99890 149770 100890 149930
rect 103080 149770 104080 149930
rect 106270 149770 107270 149930
rect 109460 149770 110460 149930
rect 112650 149770 113650 149930
rect 115840 149770 116840 149930
rect 119030 149770 120030 149930
rect 122220 149770 123220 149930
rect 125410 149770 126410 149930
rect 128600 149770 129600 149930
rect 131790 149770 132790 149930
rect 134980 149770 135980 149930
rect 0 148740 3030 149770
rect 3190 148740 6220 149770
rect 6380 148740 9410 149770
rect 9570 148740 12600 149770
rect 12760 148740 15790 149770
rect 15950 148740 18980 149770
rect 19140 148740 22170 149770
rect 22330 148740 25360 149770
rect 25520 148740 28550 149770
rect 28710 148740 31740 149770
rect 31900 148740 34930 149770
rect 35090 148740 38120 149770
rect 38280 148740 41310 149770
rect 41470 148740 44500 149770
rect 44660 148740 47690 149770
rect 47850 148740 50880 149770
rect 51040 148740 54070 149770
rect 54230 148740 57260 149770
rect 57420 148740 60450 149770
rect 60610 148740 63640 149770
rect 63800 148740 66830 149770
rect 66990 148740 70020 149770
rect 70180 148740 73210 149770
rect 73370 148740 76400 149770
rect 76560 148740 79590 149770
rect 79750 148740 82780 149770
rect 82940 148740 85970 149770
rect 86130 148740 89160 149770
rect 89320 148740 92350 149770
rect 92510 148740 95540 149770
rect 95700 148740 98730 149770
rect 98890 148740 101920 149770
rect 102080 148740 105110 149770
rect 105270 148740 108300 149770
rect 108460 148740 111490 149770
rect 111650 148740 114680 149770
rect 114840 148740 117870 149770
rect 118030 148740 121060 149770
rect 121220 148740 124250 149770
rect 124410 148740 127440 149770
rect 127600 148740 130630 149770
rect 130790 148740 133820 149770
rect 133980 148740 137010 149770
rect 0 147740 137170 148740
rect 0 146740 3030 147740
rect 3190 146740 6220 147740
rect 6380 146740 9410 147740
rect 9570 146740 12600 147740
rect 12760 146740 15790 147740
rect 15950 146740 18980 147740
rect 19140 146740 22170 147740
rect 22330 146740 25360 147740
rect 25520 146740 28550 147740
rect 28710 146740 31740 147740
rect 31900 146740 34930 147740
rect 35090 146740 38120 147740
rect 38280 146740 41310 147740
rect 41470 146740 44500 147740
rect 44660 146740 47690 147740
rect 47850 146740 50880 147740
rect 51040 146740 54070 147740
rect 54230 146740 57260 147740
rect 57420 146740 60450 147740
rect 60610 146740 63640 147740
rect 63800 146740 66830 147740
rect 66990 146740 70020 147740
rect 70180 146740 73210 147740
rect 73370 146740 76400 147740
rect 76560 146740 79590 147740
rect 79750 146740 82780 147740
rect 82940 146740 85970 147740
rect 86130 146740 89160 147740
rect 89320 146740 92350 147740
rect 92510 146740 95540 147740
rect 95700 146740 98730 147740
rect 98890 146740 101920 147740
rect 102080 146740 105110 147740
rect 105270 146740 108300 147740
rect 108460 146740 111490 147740
rect 111650 146740 114680 147740
rect 114840 146740 117870 147740
rect 118030 146740 121060 147740
rect 121220 146740 124250 147740
rect 124410 146740 127440 147740
rect 127600 146740 130630 147740
rect 130790 146740 133820 147740
rect 133980 146740 137010 147740
rect 1000 146580 2000 146740
rect 4190 146580 5190 146740
rect 7380 146580 8380 146740
rect 10570 146580 11570 146740
rect 13760 146580 14760 146740
rect 16950 146580 17950 146740
rect 20140 146580 21140 146740
rect 23330 146580 24330 146740
rect 26520 146580 27520 146740
rect 29710 146580 30710 146740
rect 32900 146580 33900 146740
rect 36090 146580 37090 146740
rect 39280 146580 40280 146740
rect 42470 146580 43470 146740
rect 45660 146580 46660 146740
rect 48850 146580 49850 146740
rect 52040 146580 53040 146740
rect 55230 146580 56230 146740
rect 58420 146580 59420 146740
rect 61610 146580 62610 146740
rect 64800 146580 65800 146740
rect 67990 146580 68990 146740
rect 71180 146580 72180 146740
rect 74370 146580 75370 146740
rect 77560 146580 78560 146740
rect 80750 146580 81750 146740
rect 83940 146580 84940 146740
rect 87130 146580 88130 146740
rect 90320 146580 91320 146740
rect 93510 146580 94510 146740
rect 96700 146580 97700 146740
rect 99890 146580 100890 146740
rect 103080 146580 104080 146740
rect 106270 146580 107270 146740
rect 109460 146580 110460 146740
rect 112650 146580 113650 146740
rect 115840 146580 116840 146740
rect 119030 146580 120030 146740
rect 122220 146580 123220 146740
rect 125410 146580 126410 146740
rect 128600 146580 129600 146740
rect 131790 146580 132790 146740
rect 134980 146580 135980 146740
rect 0 145550 3030 146580
rect 3190 145550 6220 146580
rect 6380 145550 9410 146580
rect 9570 145550 12600 146580
rect 12760 145550 15790 146580
rect 15950 145550 18980 146580
rect 19140 145550 22170 146580
rect 22330 145550 25360 146580
rect 25520 145550 28550 146580
rect 28710 145550 31740 146580
rect 31900 145550 34930 146580
rect 35090 145550 38120 146580
rect 38280 145550 41310 146580
rect 41470 145550 44500 146580
rect 44660 145550 47690 146580
rect 47850 145550 50880 146580
rect 51040 145550 54070 146580
rect 54230 145550 57260 146580
rect 57420 145550 60450 146580
rect 60610 145550 63640 146580
rect 63800 145550 66830 146580
rect 66990 145550 70020 146580
rect 70180 145550 73210 146580
rect 73370 145550 76400 146580
rect 76560 145550 79590 146580
rect 79750 145550 82780 146580
rect 82940 145550 85970 146580
rect 86130 145550 89160 146580
rect 89320 145550 92350 146580
rect 92510 145550 95540 146580
rect 95700 145550 98730 146580
rect 98890 145550 101920 146580
rect 102080 145550 105110 146580
rect 105270 145550 108300 146580
rect 108460 145550 111490 146580
rect 111650 145550 114680 146580
rect 114840 145550 117870 146580
rect 118030 145550 121060 146580
rect 121220 145550 124250 146580
rect 124410 145550 127440 146580
rect 127600 145550 130630 146580
rect 130790 145550 133820 146580
rect 133980 145550 137010 146580
rect 0 144550 137170 145550
rect 0 143550 3030 144550
rect 3190 143550 6220 144550
rect 6380 143550 9410 144550
rect 9570 143550 12600 144550
rect 12760 143550 15790 144550
rect 15950 143550 18980 144550
rect 19140 143550 22170 144550
rect 22330 143550 25360 144550
rect 25520 143550 28550 144550
rect 28710 143550 31740 144550
rect 31900 143550 34930 144550
rect 35090 143550 38120 144550
rect 38280 143550 41310 144550
rect 41470 143550 44500 144550
rect 44660 143550 47690 144550
rect 47850 143550 50880 144550
rect 51040 143550 54070 144550
rect 54230 143550 57260 144550
rect 57420 143550 60450 144550
rect 60610 143550 63640 144550
rect 63800 143550 66830 144550
rect 66990 143550 70020 144550
rect 70180 143550 73210 144550
rect 73370 143550 76400 144550
rect 76560 143550 79590 144550
rect 79750 143550 82780 144550
rect 82940 143550 85970 144550
rect 86130 143550 89160 144550
rect 89320 143550 92350 144550
rect 92510 143550 95540 144550
rect 95700 143550 98730 144550
rect 98890 143550 101920 144550
rect 102080 143550 105110 144550
rect 105270 143550 108300 144550
rect 108460 143550 111490 144550
rect 111650 143550 114680 144550
rect 114840 143550 117870 144550
rect 118030 143550 121060 144550
rect 121220 143550 124250 144550
rect 124410 143550 127440 144550
rect 127600 143550 130630 144550
rect 130790 143550 133820 144550
rect 133980 143550 137010 144550
rect 1000 143390 2000 143550
rect 4190 143390 5190 143550
rect 7380 143390 8380 143550
rect 10570 143390 11570 143550
rect 13760 143390 14760 143550
rect 16950 143390 17950 143550
rect 20140 143390 21140 143550
rect 23330 143390 24330 143550
rect 26520 143390 27520 143550
rect 29710 143390 30710 143550
rect 32900 143390 33900 143550
rect 36090 143390 37090 143550
rect 39280 143390 40280 143550
rect 42470 143390 43470 143550
rect 45660 143390 46660 143550
rect 48850 143390 49850 143550
rect 52040 143390 53040 143550
rect 55230 143390 56230 143550
rect 58420 143390 59420 143550
rect 61610 143390 62610 143550
rect 64800 143390 65800 143550
rect 67990 143390 68990 143550
rect 71180 143390 72180 143550
rect 74370 143390 75370 143550
rect 77560 143390 78560 143550
rect 80750 143390 81750 143550
rect 83940 143390 84940 143550
rect 87130 143390 88130 143550
rect 90320 143390 91320 143550
rect 93510 143390 94510 143550
rect 96700 143390 97700 143550
rect 99890 143390 100890 143550
rect 103080 143390 104080 143550
rect 106270 143390 107270 143550
rect 109460 143390 110460 143550
rect 112650 143390 113650 143550
rect 115840 143390 116840 143550
rect 119030 143390 120030 143550
rect 122220 143390 123220 143550
rect 125410 143390 126410 143550
rect 128600 143390 129600 143550
rect 131790 143390 132790 143550
rect 134980 143390 135980 143550
rect 0 142360 3030 143390
rect 3190 142360 6220 143390
rect 6380 142360 9410 143390
rect 9570 142360 12600 143390
rect 12760 142360 15790 143390
rect 15950 142360 18980 143390
rect 19140 142360 22170 143390
rect 22330 142360 25360 143390
rect 25520 142360 28550 143390
rect 28710 142360 31740 143390
rect 31900 142360 34930 143390
rect 35090 142360 38120 143390
rect 38280 142360 41310 143390
rect 41470 142360 44500 143390
rect 44660 142360 47690 143390
rect 47850 142360 50880 143390
rect 51040 142360 54070 143390
rect 54230 142360 57260 143390
rect 57420 142360 60450 143390
rect 60610 142360 63640 143390
rect 63800 142360 66830 143390
rect 66990 142360 70020 143390
rect 70180 142360 73210 143390
rect 73370 142360 76400 143390
rect 76560 142360 79590 143390
rect 79750 142360 82780 143390
rect 82940 142360 85970 143390
rect 86130 142360 89160 143390
rect 89320 142360 92350 143390
rect 92510 142360 95540 143390
rect 95700 142360 98730 143390
rect 98890 142360 101920 143390
rect 102080 142360 105110 143390
rect 105270 142360 108300 143390
rect 108460 142360 111490 143390
rect 111650 142360 114680 143390
rect 114840 142360 117870 143390
rect 118030 142360 121060 143390
rect 121220 142360 124250 143390
rect 124410 142360 127440 143390
rect 127600 142360 130630 143390
rect 130790 142360 133820 143390
rect 133980 142360 137010 143390
rect 0 141360 137170 142360
rect 0 140360 3030 141360
rect 3190 140360 6220 141360
rect 6380 140360 9410 141360
rect 9570 140360 12600 141360
rect 12760 140360 15790 141360
rect 15950 140360 18980 141360
rect 19140 140360 22170 141360
rect 22330 140360 25360 141360
rect 25520 140360 28550 141360
rect 28710 140360 31740 141360
rect 31900 140360 34930 141360
rect 35090 140360 38120 141360
rect 38280 140360 41310 141360
rect 41470 140360 44500 141360
rect 44660 140360 47690 141360
rect 47850 140360 50880 141360
rect 51040 140360 54070 141360
rect 54230 140360 57260 141360
rect 57420 140360 60450 141360
rect 60610 140360 63640 141360
rect 63800 140360 66830 141360
rect 66990 140360 70020 141360
rect 70180 140360 73210 141360
rect 73370 140360 76400 141360
rect 76560 140360 79590 141360
rect 79750 140360 82780 141360
rect 82940 140360 85970 141360
rect 86130 140360 89160 141360
rect 89320 140360 92350 141360
rect 92510 140360 95540 141360
rect 95700 140360 98730 141360
rect 98890 140360 101920 141360
rect 102080 140360 105110 141360
rect 105270 140360 108300 141360
rect 108460 140360 111490 141360
rect 111650 140360 114680 141360
rect 114840 140360 117870 141360
rect 118030 140360 121060 141360
rect 121220 140360 124250 141360
rect 124410 140360 127440 141360
rect 127600 140360 130630 141360
rect 130790 140360 133820 141360
rect 133980 140360 137010 141360
rect 1000 140200 2000 140360
rect 4190 140200 5190 140360
rect 7380 140200 8380 140360
rect 10570 140200 11570 140360
rect 13760 140200 14760 140360
rect 16950 140200 17950 140360
rect 20140 140200 21140 140360
rect 23330 140200 24330 140360
rect 26520 140200 27520 140360
rect 29710 140200 30710 140360
rect 32900 140200 33900 140360
rect 36090 140200 37090 140360
rect 39280 140200 40280 140360
rect 42470 140200 43470 140360
rect 45660 140200 46660 140360
rect 48850 140200 49850 140360
rect 52040 140200 53040 140360
rect 55230 140200 56230 140360
rect 58420 140200 59420 140360
rect 61610 140200 62610 140360
rect 64800 140200 65800 140360
rect 67990 140200 68990 140360
rect 71180 140200 72180 140360
rect 74370 140200 75370 140360
rect 77560 140200 78560 140360
rect 80750 140200 81750 140360
rect 83940 140200 84940 140360
rect 87130 140200 88130 140360
rect 90320 140200 91320 140360
rect 93510 140200 94510 140360
rect 96700 140200 97700 140360
rect 99890 140200 100890 140360
rect 103080 140200 104080 140360
rect 106270 140200 107270 140360
rect 109460 140200 110460 140360
rect 112650 140200 113650 140360
rect 115840 140200 116840 140360
rect 119030 140200 120030 140360
rect 122220 140200 123220 140360
rect 125410 140200 126410 140360
rect 128600 140200 129600 140360
rect 131790 140200 132790 140360
rect 134980 140200 135980 140360
rect 0 140160 3030 140200
rect 3190 140160 6220 140200
rect 6380 140160 9410 140200
rect 0 140110 9410 140160
rect 0 121310 50 140110
rect 9320 139170 9410 140110
rect 9570 139170 12600 140200
rect 12760 139170 15790 140200
rect 15950 139170 18980 140200
rect 19140 139170 22170 140200
rect 22330 139170 25360 140200
rect 25520 139170 28550 140200
rect 28710 139170 31740 140200
rect 31900 139170 34930 140200
rect 35090 139170 38120 140200
rect 38280 139170 41310 140200
rect 41470 139170 44500 140200
rect 44660 139170 47690 140200
rect 47850 139170 50880 140200
rect 51040 139170 54070 140200
rect 54230 139170 57260 140200
rect 57420 139170 60450 140200
rect 60610 139170 63640 140200
rect 63800 139170 66830 140200
rect 66990 139170 70020 140200
rect 70180 139170 73210 140200
rect 73370 139170 76400 140200
rect 76560 139170 79590 140200
rect 79750 139170 82780 140200
rect 82940 139170 85970 140200
rect 86130 139170 89160 140200
rect 89320 139170 92350 140200
rect 92510 139170 95540 140200
rect 95700 139170 98730 140200
rect 98890 139170 101920 140200
rect 102080 139170 105110 140200
rect 105270 139170 108300 140200
rect 108460 139170 111490 140200
rect 111650 139170 114680 140200
rect 114840 139170 117870 140200
rect 118030 139170 121060 140200
rect 121220 139170 124250 140200
rect 124410 139170 127440 140200
rect 127600 139170 130630 140200
rect 130790 139170 133820 140200
rect 133980 139170 137010 140200
rect 9320 138170 137170 139170
rect 9320 137170 9410 138170
rect 9570 137170 12600 138170
rect 12760 137170 15790 138170
rect 15950 137170 18980 138170
rect 19140 137170 22170 138170
rect 22330 137170 25360 138170
rect 25520 137170 28550 138170
rect 28710 137170 31740 138170
rect 31900 137170 34930 138170
rect 35090 137170 38120 138170
rect 38280 137170 41310 138170
rect 41470 137170 44500 138170
rect 44660 137170 47690 138170
rect 47850 137170 50880 138170
rect 51040 137170 54070 138170
rect 54230 137170 57260 138170
rect 57420 137170 60450 138170
rect 60610 137170 63640 138170
rect 63800 137170 66830 138170
rect 66990 137170 70020 138170
rect 70180 137170 73210 138170
rect 73370 137170 76400 138170
rect 76560 137170 79590 138170
rect 79750 137170 82780 138170
rect 82940 137170 85970 138170
rect 86130 137170 89160 138170
rect 89320 137170 92350 138170
rect 92510 137170 95540 138170
rect 95700 137170 98730 138170
rect 98890 137170 101920 138170
rect 102080 137170 105110 138170
rect 105270 137170 108300 138170
rect 108460 137170 111490 138170
rect 111650 137170 114680 138170
rect 114840 137170 117870 138170
rect 118030 137170 121060 138170
rect 121220 137170 124250 138170
rect 124410 137170 127440 138170
rect 127600 137170 130630 138170
rect 130790 137170 133820 138170
rect 133980 137170 137010 138170
rect 9320 137010 9370 137170
rect 10570 137010 11570 137170
rect 13760 137010 14760 137170
rect 16950 137010 17950 137170
rect 20140 137010 21140 137170
rect 23330 137010 24330 137170
rect 26520 137010 27520 137170
rect 29710 137010 30710 137170
rect 32900 137010 33900 137170
rect 36090 137010 37090 137170
rect 39280 137010 40280 137170
rect 42470 137010 43470 137170
rect 45660 137010 46660 137170
rect 48850 137010 49850 137170
rect 52040 137010 53040 137170
rect 55230 137010 56230 137170
rect 58420 137010 59420 137170
rect 61610 137010 62610 137170
rect 64800 137010 65800 137170
rect 67990 137010 68990 137170
rect 71180 137010 72180 137170
rect 74370 137010 75370 137170
rect 77560 137010 78560 137170
rect 80750 137010 81750 137170
rect 83940 137010 84940 137170
rect 87130 137010 88130 137170
rect 90320 137010 91320 137170
rect 93510 137010 94510 137170
rect 96700 137010 97700 137170
rect 99890 137010 100890 137170
rect 103080 137010 104080 137170
rect 106270 137010 107270 137170
rect 109460 137010 110460 137170
rect 112650 137010 113650 137170
rect 115840 137010 116840 137170
rect 119030 137010 120030 137170
rect 122220 137010 123220 137170
rect 125410 137010 126410 137170
rect 128600 137010 129600 137170
rect 131790 137010 132790 137170
rect 134980 137010 135980 137170
rect 9320 135980 9410 137010
rect 9570 135980 12600 137010
rect 12760 135980 15790 137010
rect 15950 135980 18980 137010
rect 19140 135980 22170 137010
rect 22330 135980 25360 137010
rect 25520 135980 28550 137010
rect 28710 135980 31740 137010
rect 31900 135980 34930 137010
rect 35090 135980 38120 137010
rect 38280 135980 41310 137010
rect 41470 135980 44500 137010
rect 44660 135980 47690 137010
rect 47850 135980 50880 137010
rect 51040 135980 54070 137010
rect 54230 135980 57260 137010
rect 57420 135980 60450 137010
rect 60610 135980 63640 137010
rect 63800 135980 66830 137010
rect 66990 135980 70020 137010
rect 70180 135980 73210 137010
rect 73370 135980 76400 137010
rect 76560 135980 79590 137010
rect 79750 135980 82780 137010
rect 82940 135980 85970 137010
rect 86130 135980 89160 137010
rect 89320 135980 92350 137010
rect 92510 135980 95540 137010
rect 95700 135980 98730 137010
rect 98890 135980 101920 137010
rect 102080 135980 105110 137010
rect 105270 135980 108300 137010
rect 108460 135980 111490 137010
rect 111650 135980 114680 137010
rect 114840 135980 117870 137010
rect 118030 135980 121060 137010
rect 121220 135980 124250 137010
rect 124410 135980 127440 137010
rect 127600 135980 130630 137010
rect 130790 135980 133820 137010
rect 133980 135980 137010 137010
rect 9320 134980 137170 135980
rect 9320 133980 9410 134980
rect 9570 133980 12600 134980
rect 12760 133980 15790 134980
rect 15950 133980 18980 134980
rect 19140 133980 22170 134980
rect 22330 133980 25360 134980
rect 25520 133980 28550 134980
rect 28710 133980 31740 134980
rect 31900 133980 34930 134980
rect 35090 133980 38120 134980
rect 38280 133980 41310 134980
rect 41470 133980 44500 134980
rect 44660 133980 47690 134980
rect 47850 133980 50880 134980
rect 51040 133980 54070 134980
rect 54230 133980 57260 134980
rect 57420 133980 60450 134980
rect 60610 133980 63640 134980
rect 63800 133980 66830 134980
rect 66990 133980 70020 134980
rect 70180 133980 73210 134980
rect 73370 133980 76400 134980
rect 76560 133980 79590 134980
rect 79750 133980 82780 134980
rect 82940 133980 85970 134980
rect 86130 133980 89160 134980
rect 89320 133980 92350 134980
rect 92510 133980 95540 134980
rect 95700 133980 98730 134980
rect 98890 133980 101920 134980
rect 102080 133980 105110 134980
rect 105270 133980 108300 134980
rect 108460 133980 111490 134980
rect 111650 133980 114680 134980
rect 114840 133980 117870 134980
rect 118030 133980 121060 134980
rect 121220 133980 124250 134980
rect 124410 133980 127440 134980
rect 127600 133980 130630 134980
rect 130790 133980 133820 134980
rect 133980 133980 137010 134980
rect 9320 133820 9370 133980
rect 10570 133820 11570 133980
rect 13760 133820 14760 133980
rect 16950 133820 17950 133980
rect 20140 133820 21140 133980
rect 23330 133820 24330 133980
rect 26520 133820 27520 133980
rect 29710 133820 30710 133980
rect 32900 133820 33900 133980
rect 36090 133820 37090 133980
rect 39280 133820 40280 133980
rect 42470 133820 43470 133980
rect 45660 133820 46660 133980
rect 48850 133820 49850 133980
rect 52040 133820 53040 133980
rect 55230 133820 56230 133980
rect 58420 133820 59420 133980
rect 61610 133820 62610 133980
rect 64800 133820 65800 133980
rect 67990 133820 68990 133980
rect 71180 133820 72180 133980
rect 74370 133820 75370 133980
rect 77560 133820 78560 133980
rect 80750 133820 81750 133980
rect 83940 133820 84940 133980
rect 87130 133820 88130 133980
rect 90320 133820 91320 133980
rect 93510 133820 94510 133980
rect 96700 133820 97700 133980
rect 99890 133820 100890 133980
rect 103080 133820 104080 133980
rect 106270 133820 107270 133980
rect 109460 133820 110460 133980
rect 112650 133820 113650 133980
rect 115840 133820 116840 133980
rect 119030 133820 120030 133980
rect 122220 133820 123220 133980
rect 125410 133820 126410 133980
rect 128600 133820 129600 133980
rect 131790 133820 132790 133980
rect 134980 133820 135980 133980
rect 9320 132790 9410 133820
rect 9570 132790 12600 133820
rect 12760 132790 15790 133820
rect 15950 132790 18980 133820
rect 19140 132790 22170 133820
rect 22330 132790 25360 133820
rect 25520 132790 28550 133820
rect 28710 132790 31740 133820
rect 31900 132790 34930 133820
rect 35090 132790 38120 133820
rect 38280 132790 41310 133820
rect 41470 132790 44500 133820
rect 44660 132790 47690 133820
rect 47850 132790 50880 133820
rect 51040 132790 54070 133820
rect 54230 132790 57260 133820
rect 57420 132790 60450 133820
rect 60610 132790 63640 133820
rect 63800 132790 66830 133820
rect 66990 132790 70020 133820
rect 70180 132790 73210 133820
rect 73370 132790 76400 133820
rect 76560 132790 79590 133820
rect 79750 132790 82780 133820
rect 82940 132790 85970 133820
rect 86130 132790 89160 133820
rect 89320 132790 92350 133820
rect 92510 132790 95540 133820
rect 95700 132790 98730 133820
rect 98890 132790 101920 133820
rect 102080 132790 105110 133820
rect 105270 132790 108300 133820
rect 108460 132790 111490 133820
rect 111650 132790 114680 133820
rect 114840 132790 117870 133820
rect 118030 132790 121060 133820
rect 121220 132790 124250 133820
rect 124410 132790 127440 133820
rect 127600 132790 130630 133820
rect 130790 132790 133820 133820
rect 133980 132790 137010 133820
rect 9320 131790 137170 132790
rect 9320 130790 9410 131790
rect 9570 130790 12600 131790
rect 12760 130790 15790 131790
rect 15950 130790 18980 131790
rect 19140 130790 22170 131790
rect 22330 130790 25360 131790
rect 25520 130790 28550 131790
rect 28710 130790 31740 131790
rect 31900 130790 34930 131790
rect 35090 130790 38120 131790
rect 38280 130790 41310 131790
rect 41470 130790 44500 131790
rect 44660 130790 47690 131790
rect 47850 130790 50880 131790
rect 51040 130790 54070 131790
rect 54230 130790 57260 131790
rect 57420 130790 60450 131790
rect 60610 130790 63640 131790
rect 63800 130790 66830 131790
rect 66990 130790 70020 131790
rect 70180 130790 73210 131790
rect 73370 130790 76400 131790
rect 76560 130790 79590 131790
rect 79750 130790 82780 131790
rect 82940 130790 85970 131790
rect 86130 130790 89160 131790
rect 89320 130790 92350 131790
rect 92510 130790 95540 131790
rect 95700 130790 98730 131790
rect 98890 130790 101920 131790
rect 102080 130790 105110 131790
rect 105270 130790 108300 131790
rect 108460 130790 111490 131790
rect 111650 130790 114680 131790
rect 114840 130790 117870 131790
rect 118030 130790 121060 131790
rect 121220 130790 124250 131790
rect 124410 130790 127440 131790
rect 127600 130790 130630 131790
rect 130790 130790 133820 131790
rect 133980 130790 137010 131790
rect 9320 130630 9370 130790
rect 10570 130630 11570 130790
rect 13760 130630 14760 130790
rect 16950 130630 17950 130790
rect 20140 130630 21140 130790
rect 23330 130630 24330 130790
rect 26520 130630 27520 130790
rect 29710 130630 30710 130790
rect 32900 130630 33900 130790
rect 36090 130630 37090 130790
rect 39280 130630 40280 130790
rect 42470 130630 43470 130790
rect 45660 130630 46660 130790
rect 48850 130630 49850 130790
rect 52040 130630 53040 130790
rect 55230 130630 56230 130790
rect 58420 130630 59420 130790
rect 61610 130630 62610 130790
rect 64800 130630 65800 130790
rect 67990 130630 68990 130790
rect 71180 130630 72180 130790
rect 74370 130630 75370 130790
rect 77560 130630 78560 130790
rect 80750 130630 81750 130790
rect 83940 130630 84940 130790
rect 87130 130630 88130 130790
rect 90320 130630 91320 130790
rect 93510 130630 94510 130790
rect 96700 130630 97700 130790
rect 99890 130630 100890 130790
rect 103080 130630 104080 130790
rect 106270 130630 107270 130790
rect 109460 130630 110460 130790
rect 112650 130630 113650 130790
rect 115840 130630 116840 130790
rect 119030 130630 120030 130790
rect 122220 130630 123220 130790
rect 125410 130630 126410 130790
rect 128600 130630 129600 130790
rect 131790 130630 132790 130790
rect 134980 130630 135980 130790
rect 9320 129600 9410 130630
rect 9570 129600 12600 130630
rect 12760 129600 15790 130630
rect 15950 129600 18980 130630
rect 19140 129600 22170 130630
rect 22330 129600 25360 130630
rect 25520 129600 28550 130630
rect 28710 129600 31740 130630
rect 31900 129600 34930 130630
rect 35090 129600 38120 130630
rect 38280 129600 41310 130630
rect 41470 129600 44500 130630
rect 44660 129600 47690 130630
rect 47850 129600 50880 130630
rect 51040 129600 54070 130630
rect 54230 129600 57260 130630
rect 57420 129600 60450 130630
rect 60610 129600 63640 130630
rect 63800 129600 66830 130630
rect 66990 129600 70020 130630
rect 70180 129600 73210 130630
rect 73370 129600 76400 130630
rect 76560 129600 79590 130630
rect 79750 129600 82780 130630
rect 82940 129600 85970 130630
rect 86130 129600 89160 130630
rect 89320 129600 92350 130630
rect 92510 129600 95540 130630
rect 95700 129600 98730 130630
rect 98890 129600 101920 130630
rect 102080 129600 105110 130630
rect 105270 129600 108300 130630
rect 108460 129600 111490 130630
rect 111650 129600 114680 130630
rect 114840 129600 117870 130630
rect 118030 129600 121060 130630
rect 121220 129600 124250 130630
rect 124410 129600 127440 130630
rect 127600 129600 130630 130630
rect 130790 129600 133820 130630
rect 133980 129600 137010 130630
rect 9320 128600 137170 129600
rect 9320 127600 9410 128600
rect 9570 127600 12600 128600
rect 12760 127600 15790 128600
rect 15950 127600 18980 128600
rect 19140 127600 22170 128600
rect 22330 127600 25360 128600
rect 25520 127600 28550 128600
rect 28710 127600 31740 128600
rect 31900 127600 34930 128600
rect 35090 127600 38120 128600
rect 38280 127600 41310 128600
rect 41470 127600 44500 128600
rect 44660 127600 47690 128600
rect 47850 127600 50880 128600
rect 51040 127600 54070 128600
rect 54230 127600 57260 128600
rect 57420 127600 60450 128600
rect 60610 127600 63640 128600
rect 63800 127600 66830 128600
rect 66990 127600 70020 128600
rect 70180 127600 73210 128600
rect 73370 127600 76400 128600
rect 76560 127600 79590 128600
rect 79750 127600 82780 128600
rect 82940 127600 85970 128600
rect 86130 127600 89160 128600
rect 89320 127600 92350 128600
rect 92510 127600 95540 128600
rect 95700 127600 98730 128600
rect 98890 127600 101920 128600
rect 102080 127600 105110 128600
rect 105270 127600 108300 128600
rect 108460 127600 111490 128600
rect 111650 127600 114680 128600
rect 114840 127600 117870 128600
rect 118030 127600 121060 128600
rect 121220 127600 124250 128600
rect 124410 127600 127440 128600
rect 127600 127600 130630 128600
rect 130790 127600 133820 128600
rect 133980 127600 137010 128600
rect 9320 127440 9370 127600
rect 10570 127440 11570 127600
rect 13760 127440 14760 127600
rect 16950 127440 17950 127600
rect 20140 127440 21140 127600
rect 23330 127440 24330 127600
rect 26520 127440 27520 127600
rect 29710 127440 30710 127600
rect 32900 127440 33900 127600
rect 36090 127440 37090 127600
rect 39280 127440 40280 127600
rect 42470 127440 43470 127600
rect 45660 127440 46660 127600
rect 48850 127440 49850 127600
rect 52040 127440 53040 127600
rect 55230 127440 56230 127600
rect 58420 127440 59420 127600
rect 61610 127440 62610 127600
rect 64800 127440 65800 127600
rect 67990 127440 68990 127600
rect 71180 127440 72180 127600
rect 74370 127440 75370 127600
rect 77560 127440 78560 127600
rect 80750 127440 81750 127600
rect 83940 127440 84940 127600
rect 87130 127440 88130 127600
rect 90320 127440 91320 127600
rect 93510 127440 94510 127600
rect 96700 127440 97700 127600
rect 99890 127440 100890 127600
rect 103080 127440 104080 127600
rect 106270 127440 107270 127600
rect 109460 127440 110460 127600
rect 112650 127440 113650 127600
rect 115840 127440 116840 127600
rect 119030 127440 120030 127600
rect 122220 127440 123220 127600
rect 125410 127440 126410 127600
rect 128600 127440 129600 127600
rect 131790 127440 132790 127600
rect 134980 127440 135980 127600
rect 9320 126410 9410 127440
rect 9570 126410 12600 127440
rect 12760 126410 15790 127440
rect 15950 126410 18980 127440
rect 19140 126410 22170 127440
rect 22330 126410 25360 127440
rect 25520 126410 28550 127440
rect 28710 126410 31740 127440
rect 31900 126410 34930 127440
rect 35090 126410 38120 127440
rect 38280 126410 41310 127440
rect 41470 126410 44500 127440
rect 44660 126410 47690 127440
rect 47850 126410 50880 127440
rect 51040 126410 54070 127440
rect 54230 126410 57260 127440
rect 57420 126410 60450 127440
rect 60610 126410 63640 127440
rect 63800 126410 66830 127440
rect 66990 126410 70020 127440
rect 70180 126410 73210 127440
rect 73370 126410 76400 127440
rect 76560 126410 79590 127440
rect 79750 126410 82780 127440
rect 82940 126410 85970 127440
rect 86130 126410 89160 127440
rect 89320 126410 92350 127440
rect 92510 126410 95540 127440
rect 95700 126410 98730 127440
rect 98890 126410 101920 127440
rect 102080 126410 105110 127440
rect 105270 126410 108300 127440
rect 108460 126410 111490 127440
rect 111650 126410 114680 127440
rect 114840 126410 117870 127440
rect 118030 126410 121060 127440
rect 121220 126410 124250 127440
rect 124410 126410 127440 127440
rect 127600 126410 130630 127440
rect 130790 126410 133820 127440
rect 133980 126410 137010 127440
rect 9320 125410 137170 126410
rect 9320 124410 9410 125410
rect 9570 124410 12600 125410
rect 12760 124410 15790 125410
rect 15950 124410 18980 125410
rect 19140 124410 22170 125410
rect 22330 124410 25360 125410
rect 25520 124410 28550 125410
rect 28710 124410 31740 125410
rect 31900 124410 34930 125410
rect 35090 124410 38120 125410
rect 38280 124410 41310 125410
rect 41470 124410 44500 125410
rect 44660 124410 47690 125410
rect 47850 124410 50880 125410
rect 51040 124410 54070 125410
rect 54230 124410 57260 125410
rect 57420 124410 60450 125410
rect 60610 124410 63640 125410
rect 63800 124410 66830 125410
rect 66990 124410 70020 125410
rect 70180 124410 73210 125410
rect 73370 124410 76400 125410
rect 76560 124410 79590 125410
rect 79750 124410 82780 125410
rect 82940 124410 85970 125410
rect 86130 124410 89160 125410
rect 89320 124410 92350 125410
rect 92510 124410 95540 125410
rect 95700 124410 98730 125410
rect 98890 124410 101920 125410
rect 102080 124410 105110 125410
rect 105270 124410 108300 125410
rect 108460 124410 111490 125410
rect 111650 124410 114680 125410
rect 114840 124410 117870 125410
rect 118030 124410 121060 125410
rect 121220 124410 124250 125410
rect 124410 124410 127440 125410
rect 127600 124410 130630 125410
rect 130790 124410 133820 125410
rect 133980 124410 137010 125410
rect 9320 124250 9370 124410
rect 10570 124250 11570 124410
rect 13760 124250 14760 124410
rect 16950 124250 17950 124410
rect 20140 124250 21140 124410
rect 23330 124250 24330 124410
rect 26520 124250 27520 124410
rect 29710 124250 30710 124410
rect 32900 124250 33900 124410
rect 36090 124250 37090 124410
rect 39280 124250 40280 124410
rect 42470 124250 43470 124410
rect 45660 124250 46660 124410
rect 48850 124250 49850 124410
rect 52040 124250 53040 124410
rect 55230 124250 56230 124410
rect 58420 124250 59420 124410
rect 61610 124250 62610 124410
rect 64800 124250 65800 124410
rect 67990 124250 68990 124410
rect 71180 124250 72180 124410
rect 74370 124250 75370 124410
rect 77560 124250 78560 124410
rect 80750 124250 81750 124410
rect 83940 124250 84940 124410
rect 87130 124250 88130 124410
rect 90320 124250 91320 124410
rect 93510 124250 94510 124410
rect 96700 124250 97700 124410
rect 99890 124250 100890 124410
rect 103080 124250 104080 124410
rect 106270 124250 107270 124410
rect 109460 124250 110460 124410
rect 112650 124250 113650 124410
rect 115840 124250 116840 124410
rect 119030 124250 120030 124410
rect 122220 124250 123220 124410
rect 125410 124250 126410 124410
rect 128600 124250 129600 124410
rect 131790 124250 132790 124410
rect 134980 124250 135980 124410
rect 9320 123220 9410 124250
rect 9570 123220 12600 124250
rect 12760 123220 15790 124250
rect 15950 123220 18980 124250
rect 19140 123220 22170 124250
rect 22330 123220 25360 124250
rect 25520 123220 28550 124250
rect 28710 123220 31740 124250
rect 31900 123220 34930 124250
rect 35090 123220 38120 124250
rect 38280 123220 41310 124250
rect 41470 123220 44500 124250
rect 44660 123220 47690 124250
rect 47850 123220 50880 124250
rect 51040 123220 54070 124250
rect 54230 123220 57260 124250
rect 57420 123220 60450 124250
rect 60610 123220 63640 124250
rect 63800 123220 66830 124250
rect 66990 123220 70020 124250
rect 70180 123220 73210 124250
rect 73370 123220 76400 124250
rect 76560 123220 79590 124250
rect 79750 123220 82780 124250
rect 82940 123220 85970 124250
rect 86130 123220 89160 124250
rect 89320 123220 92350 124250
rect 92510 123220 95540 124250
rect 95700 123220 98730 124250
rect 98890 123220 101920 124250
rect 102080 123220 105110 124250
rect 105270 123220 108300 124250
rect 108460 123220 111490 124250
rect 111650 123220 114680 124250
rect 114840 123220 117870 124250
rect 118030 123220 121060 124250
rect 121220 123220 124250 124250
rect 124410 123220 127440 124250
rect 127600 123220 130630 124250
rect 130790 123220 133820 124250
rect 133980 123220 137010 124250
rect 9320 122220 137170 123220
rect 9320 121310 9410 122220
rect 0 121260 9410 121310
rect 0 121220 3030 121260
rect 3190 121220 6220 121260
rect 6380 121220 9410 121260
rect 9570 121220 12600 122220
rect 12760 121220 15790 122220
rect 15950 121220 18980 122220
rect 19140 121220 22170 122220
rect 22330 121220 25360 122220
rect 25520 121220 28550 122220
rect 28710 121220 31740 122220
rect 31900 121220 34930 122220
rect 35090 121220 38120 122220
rect 38280 121220 41310 122220
rect 41470 121220 44500 122220
rect 44660 121220 47690 122220
rect 47850 121220 50880 122220
rect 51040 121220 54070 122220
rect 54230 121220 57260 122220
rect 57420 121220 60450 122220
rect 60610 121220 63640 122220
rect 63800 121220 66830 122220
rect 66990 121220 70020 122220
rect 70180 121220 73210 122220
rect 73370 121220 76400 122220
rect 76560 121220 79590 122220
rect 79750 121220 82780 122220
rect 82940 121220 85970 122220
rect 86130 121220 89160 122220
rect 89320 121220 92350 122220
rect 92510 121220 95540 122220
rect 95700 121220 98730 122220
rect 98890 121220 101920 122220
rect 102080 121220 105110 122220
rect 105270 121220 108300 122220
rect 108460 121220 111490 122220
rect 111650 121220 114680 122220
rect 114840 121220 117870 122220
rect 118030 121220 121060 122220
rect 121220 121220 124250 122220
rect 124410 121220 127440 122220
rect 127600 121220 130630 122220
rect 130790 121220 133820 122220
rect 133980 121220 137010 122220
rect 1000 121060 2000 121220
rect 4190 121060 5190 121220
rect 7380 121060 8380 121220
rect 10570 121060 11570 121220
rect 13760 121060 14760 121220
rect 16950 121060 17950 121220
rect 20140 121060 21140 121220
rect 23330 121060 24330 121220
rect 26520 121060 27520 121220
rect 29710 121060 30710 121220
rect 32900 121060 33900 121220
rect 36090 121060 37090 121220
rect 39280 121060 40280 121220
rect 42470 121060 43470 121220
rect 45660 121060 46660 121220
rect 48850 121060 49850 121220
rect 52040 121060 53040 121220
rect 55230 121060 56230 121220
rect 58420 121060 59420 121220
rect 61610 121060 62610 121220
rect 64800 121060 65800 121220
rect 67990 121060 68990 121220
rect 71180 121060 72180 121220
rect 74370 121060 75370 121220
rect 77560 121060 78560 121220
rect 80750 121060 81750 121220
rect 83940 121060 84940 121220
rect 87130 121060 88130 121220
rect 90320 121060 91320 121220
rect 93510 121060 94510 121220
rect 96700 121060 97700 121220
rect 99890 121060 100890 121220
rect 103080 121060 104080 121220
rect 106270 121060 107270 121220
rect 109460 121060 110460 121220
rect 112650 121060 113650 121220
rect 115840 121060 116840 121220
rect 119030 121060 120030 121220
rect 122220 121060 123220 121220
rect 125410 121060 126410 121220
rect 128600 121060 129600 121220
rect 131790 121060 132790 121220
rect 134980 121060 135980 121220
rect 0 120030 3030 121060
rect 3190 120030 6220 121060
rect 6380 120030 9410 121060
rect 9570 120030 12600 121060
rect 12760 120030 15790 121060
rect 15950 120030 18980 121060
rect 19140 120030 22170 121060
rect 22330 120030 25360 121060
rect 25520 120030 28550 121060
rect 28710 120030 31740 121060
rect 31900 120030 34930 121060
rect 35090 120030 38120 121060
rect 38280 120030 41310 121060
rect 41470 120030 44500 121060
rect 44660 120030 47690 121060
rect 47850 120030 50880 121060
rect 51040 120030 54070 121060
rect 54230 120030 57260 121060
rect 57420 120030 60450 121060
rect 60610 120030 63640 121060
rect 63800 120030 66830 121060
rect 66990 120030 70020 121060
rect 70180 120030 73210 121060
rect 73370 120030 76400 121060
rect 76560 120030 79590 121060
rect 79750 120030 82780 121060
rect 82940 120030 85970 121060
rect 86130 120030 89160 121060
rect 89320 120030 92350 121060
rect 92510 120030 95540 121060
rect 95700 120030 98730 121060
rect 98890 120030 101920 121060
rect 102080 120030 105110 121060
rect 105270 120030 108300 121060
rect 108460 120030 111490 121060
rect 111650 120030 114680 121060
rect 114840 120030 117870 121060
rect 118030 120030 121060 121060
rect 121220 120030 124250 121060
rect 124410 120030 127440 121060
rect 127600 120030 130630 121060
rect 130790 120030 133820 121060
rect 133980 120030 137010 121060
rect 0 119030 137170 120030
rect 0 118030 3030 119030
rect 3190 118030 6220 119030
rect 6380 118030 9410 119030
rect 9570 118030 12600 119030
rect 12760 118030 15790 119030
rect 15950 118030 18980 119030
rect 19140 118030 22170 119030
rect 22330 118030 25360 119030
rect 25520 118030 28550 119030
rect 28710 118030 31740 119030
rect 31900 118030 34930 119030
rect 35090 118030 38120 119030
rect 38280 118030 41310 119030
rect 41470 118030 44500 119030
rect 44660 118030 47690 119030
rect 47850 118030 50880 119030
rect 51040 118030 54070 119030
rect 54230 118030 57260 119030
rect 57420 118030 60450 119030
rect 60610 118030 63640 119030
rect 63800 118030 66830 119030
rect 66990 118030 70020 119030
rect 70180 118030 73210 119030
rect 73370 118030 76400 119030
rect 76560 118030 79590 119030
rect 79750 118030 82780 119030
rect 82940 118030 85970 119030
rect 86130 118030 89160 119030
rect 89320 118030 92350 119030
rect 92510 118030 95540 119030
rect 95700 118030 98730 119030
rect 98890 118030 101920 119030
rect 102080 118030 105110 119030
rect 105270 118030 108300 119030
rect 108460 118030 111490 119030
rect 111650 118030 114680 119030
rect 114840 118030 117870 119030
rect 118030 118030 121060 119030
rect 121220 118030 124250 119030
rect 124410 118030 127440 119030
rect 127600 118030 130630 119030
rect 130790 118030 133820 119030
rect 133980 118030 137010 119030
rect 1000 117870 2000 118030
rect 4190 117870 5190 118030
rect 7380 117870 8380 118030
rect 10570 117870 11570 118030
rect 13760 117870 14760 118030
rect 16950 117870 17950 118030
rect 20140 117870 21140 118030
rect 23330 117870 24330 118030
rect 26520 117870 27520 118030
rect 29710 117870 30710 118030
rect 32900 117870 33900 118030
rect 36090 117870 37090 118030
rect 39280 117870 40280 118030
rect 42470 117870 43470 118030
rect 45660 117870 46660 118030
rect 48850 117870 49850 118030
rect 52040 117870 53040 118030
rect 55230 117870 56230 118030
rect 58420 117870 59420 118030
rect 61610 117870 62610 118030
rect 64800 117870 65800 118030
rect 67990 117870 68990 118030
rect 71180 117870 72180 118030
rect 74370 117870 75370 118030
rect 77560 117870 78560 118030
rect 80750 117870 81750 118030
rect 83940 117870 84940 118030
rect 87130 117870 88130 118030
rect 90320 117870 91320 118030
rect 93510 117870 94510 118030
rect 96700 117870 97700 118030
rect 99890 117870 100890 118030
rect 103080 117870 104080 118030
rect 106270 117870 107270 118030
rect 109460 117870 110460 118030
rect 112650 117870 113650 118030
rect 115840 117870 116840 118030
rect 119030 117870 120030 118030
rect 122220 117870 123220 118030
rect 125410 117870 126410 118030
rect 128600 117870 129600 118030
rect 131790 117870 132790 118030
rect 134980 117870 135980 118030
rect 0 116840 3030 117870
rect 3190 116840 6220 117870
rect 6380 116840 9410 117870
rect 9570 116840 12600 117870
rect 12760 116840 15790 117870
rect 15950 116840 18980 117870
rect 19140 116840 22170 117870
rect 22330 116840 25360 117870
rect 25520 116840 28550 117870
rect 28710 116840 31740 117870
rect 31900 116840 34930 117870
rect 35090 116840 38120 117870
rect 38280 116840 41310 117870
rect 41470 116840 44500 117870
rect 44660 116840 47690 117870
rect 47850 116840 50880 117870
rect 51040 116840 54070 117870
rect 54230 116840 57260 117870
rect 57420 116840 60450 117870
rect 60610 116840 63640 117870
rect 63800 116840 66830 117870
rect 66990 116840 70020 117870
rect 70180 116840 73210 117870
rect 73370 116840 76400 117870
rect 76560 116840 79590 117870
rect 79750 116840 82780 117870
rect 82940 116840 85970 117870
rect 86130 116840 89160 117870
rect 89320 116840 92350 117870
rect 92510 116840 95540 117870
rect 95700 116840 98730 117870
rect 98890 116840 101920 117870
rect 102080 116840 105110 117870
rect 105270 116840 108300 117870
rect 108460 116840 111490 117870
rect 111650 116840 114680 117870
rect 114840 116840 117870 117870
rect 118030 116840 121060 117870
rect 121220 116840 124250 117870
rect 124410 116840 127440 117870
rect 127600 116840 130630 117870
rect 130790 116840 133820 117870
rect 133980 116840 137010 117870
rect 0 115840 137170 116840
rect 0 114840 3030 115840
rect 3190 114840 6220 115840
rect 6380 114840 9410 115840
rect 9570 114840 12600 115840
rect 12760 114840 15790 115840
rect 15950 114840 18980 115840
rect 19140 114840 22170 115840
rect 22330 114840 25360 115840
rect 25520 114840 28550 115840
rect 28710 114840 31740 115840
rect 31900 114840 34930 115840
rect 35090 114840 38120 115840
rect 38280 114840 41310 115840
rect 41470 114840 44500 115840
rect 44660 114840 47690 115840
rect 47850 114840 50880 115840
rect 51040 114840 54070 115840
rect 54230 114840 57260 115840
rect 57420 114840 60450 115840
rect 60610 114840 63640 115840
rect 63800 114840 66830 115840
rect 66990 114840 70020 115840
rect 70180 114840 73210 115840
rect 73370 114840 76400 115840
rect 76560 114840 79590 115840
rect 79750 114840 82780 115840
rect 82940 114840 85970 115840
rect 86130 114840 89160 115840
rect 89320 114840 92350 115840
rect 92510 114840 95540 115840
rect 95700 114840 98730 115840
rect 98890 114840 101920 115840
rect 102080 114840 105110 115840
rect 105270 114840 108300 115840
rect 108460 114840 111490 115840
rect 111650 114840 114680 115840
rect 114840 114840 117870 115840
rect 118030 114840 121060 115840
rect 121220 114840 124250 115840
rect 124410 114840 127440 115840
rect 127600 114840 130630 115840
rect 130790 114840 133820 115840
rect 133980 114840 137010 115840
rect 1000 114680 2000 114840
rect 4190 114680 5190 114840
rect 7380 114680 8380 114840
rect 10570 114680 11570 114840
rect 13760 114680 14760 114840
rect 16950 114680 17950 114840
rect 20140 114680 21140 114840
rect 23330 114680 24330 114840
rect 26520 114680 27520 114840
rect 29710 114680 30710 114840
rect 32900 114680 33900 114840
rect 36090 114680 37090 114840
rect 39280 114680 40280 114840
rect 42470 114680 43470 114840
rect 45660 114680 46660 114840
rect 48850 114680 49850 114840
rect 52040 114680 53040 114840
rect 55230 114680 56230 114840
rect 58420 114680 59420 114840
rect 61610 114680 62610 114840
rect 64800 114680 65800 114840
rect 67990 114680 68990 114840
rect 71180 114680 72180 114840
rect 74370 114680 75370 114840
rect 77560 114680 78560 114840
rect 80750 114680 81750 114840
rect 83940 114680 84940 114840
rect 87130 114680 88130 114840
rect 90320 114680 91320 114840
rect 93510 114680 94510 114840
rect 96700 114680 97700 114840
rect 99890 114680 100890 114840
rect 103080 114680 104080 114840
rect 106270 114680 107270 114840
rect 109460 114680 110460 114840
rect 112650 114680 113650 114840
rect 115840 114680 116840 114840
rect 119030 114680 120030 114840
rect 122220 114680 123220 114840
rect 125410 114680 126410 114840
rect 128600 114680 129600 114840
rect 131790 114680 132790 114840
rect 134980 114680 135980 114840
rect 0 113650 3030 114680
rect 3190 113650 6220 114680
rect 6380 113650 9410 114680
rect 9570 113650 12600 114680
rect 12760 113650 15790 114680
rect 15950 113650 18980 114680
rect 19140 113650 22170 114680
rect 22330 113650 25360 114680
rect 25520 113650 28550 114680
rect 28710 113650 31740 114680
rect 31900 113650 34930 114680
rect 35090 113650 38120 114680
rect 38280 113650 41310 114680
rect 41470 113650 44500 114680
rect 44660 113650 47690 114680
rect 47850 113650 50880 114680
rect 51040 113650 54070 114680
rect 54230 113650 57260 114680
rect 57420 113650 60450 114680
rect 60610 113650 63640 114680
rect 63800 113650 66830 114680
rect 66990 113650 70020 114680
rect 70180 113650 73210 114680
rect 73370 113650 76400 114680
rect 76560 113650 79590 114680
rect 79750 113650 82780 114680
rect 82940 113650 85970 114680
rect 86130 113650 89160 114680
rect 89320 113650 92350 114680
rect 92510 113650 95540 114680
rect 95700 113650 98730 114680
rect 98890 113650 101920 114680
rect 102080 113650 105110 114680
rect 105270 113650 108300 114680
rect 108460 113650 111490 114680
rect 111650 113650 114680 114680
rect 114840 113650 117870 114680
rect 118030 113650 121060 114680
rect 121220 113650 124250 114680
rect 124410 113650 127440 114680
rect 127600 113650 130630 114680
rect 130790 113650 133820 114680
rect 133980 113650 137010 114680
rect 0 112650 137170 113650
rect 0 111650 3030 112650
rect 3190 111650 6220 112650
rect 6380 111650 9410 112650
rect 9570 111650 12600 112650
rect 12760 111650 15790 112650
rect 15950 111650 18980 112650
rect 19140 111650 22170 112650
rect 22330 111650 25360 112650
rect 25520 111650 28550 112650
rect 28710 111650 31740 112650
rect 31900 111650 34930 112650
rect 35090 111650 38120 112650
rect 38280 111650 41310 112650
rect 41470 111650 44500 112650
rect 44660 111650 47690 112650
rect 47850 111650 50880 112650
rect 51040 111650 54070 112650
rect 54230 111650 57260 112650
rect 57420 111650 60450 112650
rect 60610 111650 63640 112650
rect 63800 111650 66830 112650
rect 66990 111650 70020 112650
rect 70180 111650 73210 112650
rect 73370 111650 76400 112650
rect 76560 111650 79590 112650
rect 79750 111650 82780 112650
rect 82940 111650 85970 112650
rect 86130 111650 89160 112650
rect 89320 111650 92350 112650
rect 92510 111650 95540 112650
rect 95700 111650 98730 112650
rect 98890 111650 101920 112650
rect 102080 111650 105110 112650
rect 105270 111650 108300 112650
rect 108460 111650 111490 112650
rect 111650 111650 114680 112650
rect 114840 111650 117870 112650
rect 118030 111650 121060 112650
rect 121220 111650 124250 112650
rect 124410 111650 127440 112650
rect 127600 111650 130630 112650
rect 130790 111650 133820 112650
rect 133980 111650 137010 112650
rect 1000 111490 2000 111650
rect 4190 111490 5190 111650
rect 7380 111490 8380 111650
rect 10570 111490 11570 111650
rect 13760 111490 14760 111650
rect 16950 111490 17950 111650
rect 20140 111490 21140 111650
rect 23330 111490 24330 111650
rect 26520 111490 27520 111650
rect 29710 111490 30710 111650
rect 32900 111490 33900 111650
rect 36090 111490 37090 111650
rect 39280 111490 40280 111650
rect 42470 111490 43470 111650
rect 45660 111490 46660 111650
rect 48850 111490 49850 111650
rect 52040 111490 53040 111650
rect 55230 111490 56230 111650
rect 58420 111490 59420 111650
rect 61610 111490 62610 111650
rect 64800 111490 65800 111650
rect 67990 111490 68990 111650
rect 71180 111490 72180 111650
rect 74370 111490 75370 111650
rect 77560 111490 78560 111650
rect 80750 111490 81750 111650
rect 83940 111490 84940 111650
rect 87130 111490 88130 111650
rect 90320 111490 91320 111650
rect 93510 111490 94510 111650
rect 96700 111490 97700 111650
rect 99890 111490 100890 111650
rect 103080 111490 104080 111650
rect 106270 111490 107270 111650
rect 109460 111490 110460 111650
rect 112650 111490 113650 111650
rect 115840 111490 116840 111650
rect 119030 111490 120030 111650
rect 122220 111490 123220 111650
rect 125410 111490 126410 111650
rect 128600 111490 129600 111650
rect 131790 111490 132790 111650
rect 134980 111490 135980 111650
rect 0 110460 3030 111490
rect 3190 110460 6220 111490
rect 6380 110460 9410 111490
rect 9570 110460 12600 111490
rect 12760 110460 15790 111490
rect 15950 110460 18980 111490
rect 19140 110460 22170 111490
rect 22330 110460 25360 111490
rect 25520 110460 28550 111490
rect 28710 110460 31740 111490
rect 31900 110460 34930 111490
rect 35090 110460 38120 111490
rect 38280 110460 41310 111490
rect 41470 110460 44500 111490
rect 44660 110460 47690 111490
rect 47850 110460 50880 111490
rect 51040 110460 54070 111490
rect 54230 110460 57260 111490
rect 57420 110460 60450 111490
rect 60610 110460 63640 111490
rect 63800 110460 66830 111490
rect 66990 110460 70020 111490
rect 70180 110460 73210 111490
rect 73370 110460 76400 111490
rect 76560 110460 79590 111490
rect 79750 110460 82780 111490
rect 82940 110460 85970 111490
rect 86130 110460 89160 111490
rect 89320 110460 92350 111490
rect 92510 110460 95540 111490
rect 95700 110460 98730 111490
rect 98890 110460 101920 111490
rect 102080 110460 105110 111490
rect 105270 110460 108300 111490
rect 108460 110460 111490 111490
rect 111650 110460 114680 111490
rect 114840 110460 117870 111490
rect 118030 110460 121060 111490
rect 121220 110460 124250 111490
rect 124410 110460 127440 111490
rect 127600 110460 130630 111490
rect 130790 110460 133820 111490
rect 133980 110460 137010 111490
rect 0 109460 137170 110460
rect 0 108460 3030 109460
rect 3190 108460 6220 109460
rect 6380 108460 9410 109460
rect 9570 108460 12600 109460
rect 12760 108460 15790 109460
rect 15950 108460 18980 109460
rect 19140 108460 22170 109460
rect 22330 108460 25360 109460
rect 25520 108460 28550 109460
rect 28710 108460 31740 109460
rect 31900 108460 34930 109460
rect 35090 108460 38120 109460
rect 38280 108460 41310 109460
rect 41470 108460 44500 109460
rect 44660 108460 47690 109460
rect 47850 108460 50880 109460
rect 51040 108460 54070 109460
rect 54230 108460 57260 109460
rect 57420 108460 60450 109460
rect 60610 108460 63640 109460
rect 63800 108460 66830 109460
rect 66990 108460 70020 109460
rect 70180 108460 73210 109460
rect 73370 108460 76400 109460
rect 76560 108460 79590 109460
rect 79750 108460 82780 109460
rect 82940 108460 85970 109460
rect 86130 108460 89160 109460
rect 89320 108460 92350 109460
rect 92510 108460 95540 109460
rect 95700 108460 98730 109460
rect 98890 108460 101920 109460
rect 102080 108460 105110 109460
rect 105270 108460 108300 109460
rect 108460 108460 111490 109460
rect 111650 108460 114680 109460
rect 114840 108460 117870 109460
rect 118030 108460 121060 109460
rect 121220 108460 124250 109460
rect 124410 108460 127440 109460
rect 127600 108460 130630 109460
rect 130790 108460 133820 109460
rect 133980 108460 137010 109460
rect 1000 108300 2000 108460
rect 4190 108300 5190 108460
rect 7380 108300 8380 108460
rect 10570 108300 11570 108460
rect 13760 108300 14760 108460
rect 16950 108300 17950 108460
rect 20140 108300 21140 108460
rect 23330 108300 24330 108460
rect 26520 108300 27520 108460
rect 29710 108300 30710 108460
rect 32900 108300 33900 108460
rect 36090 108300 37090 108460
rect 39280 108300 40280 108460
rect 42470 108300 43470 108460
rect 45660 108300 46660 108460
rect 48850 108300 49850 108460
rect 52040 108300 53040 108460
rect 55230 108300 56230 108460
rect 58420 108300 59420 108460
rect 61610 108300 62610 108460
rect 64800 108300 65800 108460
rect 67990 108300 68990 108460
rect 71180 108300 72180 108460
rect 74370 108300 75370 108460
rect 77560 108300 78560 108460
rect 80750 108300 81750 108460
rect 83940 108300 84940 108460
rect 87130 108300 88130 108460
rect 90320 108300 91320 108460
rect 93510 108300 94510 108460
rect 96700 108300 97700 108460
rect 99890 108300 100890 108460
rect 103080 108300 104080 108460
rect 106270 108300 107270 108460
rect 109460 108300 110460 108460
rect 112650 108300 113650 108460
rect 115840 108300 116840 108460
rect 119030 108300 120030 108460
rect 122220 108300 123220 108460
rect 125410 108300 126410 108460
rect 128600 108300 129600 108460
rect 131790 108300 132790 108460
rect 134980 108300 135980 108460
rect 0 107270 3030 108300
rect 3190 107270 6220 108300
rect 6380 107270 9410 108300
rect 9570 107270 12600 108300
rect 12760 107270 15790 108300
rect 15950 107270 18980 108300
rect 19140 107270 22170 108300
rect 22330 107270 25360 108300
rect 25520 107270 28550 108300
rect 28710 107270 31740 108300
rect 31900 107270 34930 108300
rect 35090 107270 38120 108300
rect 38280 107270 41310 108300
rect 41470 107270 44500 108300
rect 44660 107270 47690 108300
rect 47850 107270 50880 108300
rect 51040 107270 54070 108300
rect 54230 107270 57260 108300
rect 57420 107270 60450 108300
rect 60610 107270 63640 108300
rect 63800 107270 66830 108300
rect 66990 107270 70020 108300
rect 70180 107270 73210 108300
rect 73370 107270 76400 108300
rect 76560 107270 79590 108300
rect 79750 107270 82780 108300
rect 82940 107270 85970 108300
rect 86130 107270 89160 108300
rect 89320 107270 92350 108300
rect 92510 107270 95540 108300
rect 95700 107270 98730 108300
rect 98890 107270 101920 108300
rect 102080 107270 105110 108300
rect 105270 107270 108300 108300
rect 108460 107270 111490 108300
rect 111650 107270 114680 108300
rect 114840 107270 117870 108300
rect 118030 107270 121060 108300
rect 121220 107270 124250 108300
rect 124410 107270 127440 108300
rect 127600 107270 130630 108300
rect 130790 107270 133820 108300
rect 133980 107270 137010 108300
rect 0 106270 137170 107270
rect 0 105270 3030 106270
rect 3190 105270 6220 106270
rect 6380 105270 9410 106270
rect 9570 105270 12600 106270
rect 12760 105270 15790 106270
rect 15950 105270 18980 106270
rect 19140 105270 22170 106270
rect 22330 105270 25360 106270
rect 25520 105270 28550 106270
rect 28710 105270 31740 106270
rect 31900 105270 34930 106270
rect 35090 105270 38120 106270
rect 38280 105270 41310 106270
rect 41470 105270 44500 106270
rect 44660 105270 47690 106270
rect 47850 105270 50880 106270
rect 51040 105270 54070 106270
rect 54230 105270 57260 106270
rect 57420 105270 60450 106270
rect 60610 105270 63640 106270
rect 63800 105270 66830 106270
rect 66990 105270 70020 106270
rect 70180 105270 73210 106270
rect 73370 105270 76400 106270
rect 76560 105270 79590 106270
rect 79750 105270 82780 106270
rect 82940 105270 85970 106270
rect 86130 105270 89160 106270
rect 89320 105270 92350 106270
rect 92510 105270 95540 106270
rect 95700 105270 98730 106270
rect 98890 105270 101920 106270
rect 102080 105270 105110 106270
rect 105270 105270 108300 106270
rect 108460 105270 111490 106270
rect 111650 105270 114680 106270
rect 114840 105270 117870 106270
rect 118030 105270 121060 106270
rect 121220 105270 124250 106270
rect 124410 105270 127440 106270
rect 127600 105270 130630 106270
rect 130790 105270 133820 106270
rect 133980 105270 137010 106270
rect 1000 105110 2000 105270
rect 4190 105110 5190 105270
rect 7380 105110 8380 105270
rect 10570 105110 11570 105270
rect 13760 105110 14760 105270
rect 16950 105110 17950 105270
rect 20140 105110 21140 105270
rect 23330 105110 24330 105270
rect 26520 105110 27520 105270
rect 29710 105110 30710 105270
rect 32900 105110 33900 105270
rect 36090 105110 37090 105270
rect 39280 105110 40280 105270
rect 42470 105110 43470 105270
rect 45660 105110 46660 105270
rect 48850 105110 49850 105270
rect 52040 105110 53040 105270
rect 55230 105110 56230 105270
rect 58420 105110 59420 105270
rect 61610 105110 62610 105270
rect 64800 105110 65800 105270
rect 67990 105110 68990 105270
rect 71180 105110 72180 105270
rect 74370 105110 75370 105270
rect 77560 105110 78560 105270
rect 80750 105110 81750 105270
rect 83940 105110 84940 105270
rect 87130 105110 88130 105270
rect 90320 105110 91320 105270
rect 93510 105110 94510 105270
rect 96700 105110 97700 105270
rect 99890 105110 100890 105270
rect 103080 105110 104080 105270
rect 106270 105110 107270 105270
rect 109460 105110 110460 105270
rect 112650 105110 113650 105270
rect 115840 105110 116840 105270
rect 119030 105110 120030 105270
rect 122220 105110 123220 105270
rect 125410 105110 126410 105270
rect 128600 105110 129600 105270
rect 131790 105110 132790 105270
rect 134980 105110 135980 105270
rect 0 104080 3030 105110
rect 3190 104080 6220 105110
rect 6380 104080 9410 105110
rect 9570 104080 12600 105110
rect 12760 104080 15790 105110
rect 15950 104080 18980 105110
rect 19140 104080 22170 105110
rect 22330 104080 25360 105110
rect 25520 104080 28550 105110
rect 28710 104080 31740 105110
rect 31900 104080 34930 105110
rect 35090 104080 38120 105110
rect 38280 104080 41310 105110
rect 41470 104080 44500 105110
rect 44660 104080 47690 105110
rect 47850 104080 50880 105110
rect 51040 104080 54070 105110
rect 54230 104080 57260 105110
rect 57420 104080 60450 105110
rect 60610 104080 63640 105110
rect 63800 104080 66830 105110
rect 66990 104080 70020 105110
rect 70180 104080 73210 105110
rect 73370 104080 76400 105110
rect 76560 104080 79590 105110
rect 79750 104080 82780 105110
rect 82940 104080 85970 105110
rect 86130 104080 89160 105110
rect 89320 104080 92350 105110
rect 92510 104080 95540 105110
rect 95700 104080 98730 105110
rect 98890 104080 101920 105110
rect 102080 104080 105110 105110
rect 105270 104080 108300 105110
rect 108460 104080 111490 105110
rect 111650 104080 114680 105110
rect 114840 104080 117870 105110
rect 118030 104080 121060 105110
rect 121220 104080 124250 105110
rect 124410 104080 127440 105110
rect 127600 104080 130630 105110
rect 130790 104080 133820 105110
rect 133980 104080 137010 105110
rect 0 103080 137170 104080
rect 0 102080 3030 103080
rect 3190 102080 6220 103080
rect 6380 102080 9410 103080
rect 9570 102080 12600 103080
rect 12760 102080 15790 103080
rect 15950 102080 18980 103080
rect 19140 102080 22170 103080
rect 22330 102080 25360 103080
rect 25520 102080 28550 103080
rect 28710 102080 31740 103080
rect 31900 102080 34930 103080
rect 35090 102080 38120 103080
rect 38280 102080 41310 103080
rect 41470 102080 44500 103080
rect 44660 102080 47690 103080
rect 47850 102080 50880 103080
rect 51040 102080 54070 103080
rect 54230 102080 57260 103080
rect 57420 102080 60450 103080
rect 60610 102080 63640 103080
rect 63800 102080 66830 103080
rect 66990 102080 70020 103080
rect 70180 102080 73210 103080
rect 73370 102080 76400 103080
rect 76560 102080 79590 103080
rect 79750 102080 82780 103080
rect 82940 102080 85970 103080
rect 86130 102080 89160 103080
rect 89320 102080 92350 103080
rect 92510 102080 95540 103080
rect 95700 102080 98730 103080
rect 98890 102080 101920 103080
rect 102080 102080 105110 103080
rect 105270 102080 108300 103080
rect 108460 102080 111490 103080
rect 111650 102080 114680 103080
rect 114840 102080 117870 103080
rect 118030 102080 121060 103080
rect 121220 102080 124250 103080
rect 124410 102080 127440 103080
rect 127600 102080 130630 103080
rect 130790 102080 133820 103080
rect 133980 102080 137010 103080
rect 1000 101920 2000 102080
rect 4190 101920 5190 102080
rect 7380 101920 8380 102080
rect 10570 101920 11570 102080
rect 13760 101920 14760 102080
rect 16950 101920 17950 102080
rect 20140 101920 21140 102080
rect 23330 101920 24330 102080
rect 26520 101920 27520 102080
rect 29710 101920 30710 102080
rect 32900 101920 33900 102080
rect 36090 101920 37090 102080
rect 39280 101920 40280 102080
rect 42470 101920 43470 102080
rect 45660 101920 46660 102080
rect 48850 101920 49850 102080
rect 52040 101920 53040 102080
rect 55230 101920 56230 102080
rect 58420 101920 59420 102080
rect 61610 101920 62610 102080
rect 64800 101920 65800 102080
rect 67990 101920 68990 102080
rect 71180 101920 72180 102080
rect 74370 101920 75370 102080
rect 77560 101920 78560 102080
rect 80750 101920 81750 102080
rect 83940 101920 84940 102080
rect 87130 101920 88130 102080
rect 90320 101920 91320 102080
rect 93510 101920 94510 102080
rect 96700 101920 97700 102080
rect 99890 101920 100890 102080
rect 103080 101920 104080 102080
rect 106270 101920 107270 102080
rect 109460 101920 110460 102080
rect 112650 101920 113650 102080
rect 115840 101920 116840 102080
rect 119030 101920 120030 102080
rect 122220 101920 123220 102080
rect 125410 101920 126410 102080
rect 128600 101920 129600 102080
rect 131790 101920 132790 102080
rect 134980 101920 135980 102080
rect 0 100890 3030 101920
rect 3190 100890 6220 101920
rect 6380 100890 9410 101920
rect 9570 100890 12600 101920
rect 12760 100890 15790 101920
rect 15950 100890 18980 101920
rect 19140 100890 22170 101920
rect 22330 100890 25360 101920
rect 25520 100890 28550 101920
rect 28710 100890 31740 101920
rect 31900 100890 34930 101920
rect 35090 100890 38120 101920
rect 38280 100890 41310 101920
rect 41470 100890 44500 101920
rect 44660 100890 47690 101920
rect 47850 100890 50880 101920
rect 51040 100890 54070 101920
rect 54230 100890 57260 101920
rect 57420 100890 60450 101920
rect 60610 100890 63640 101920
rect 63800 100890 66830 101920
rect 66990 100890 70020 101920
rect 70180 100890 73210 101920
rect 73370 100890 76400 101920
rect 76560 100890 79590 101920
rect 79750 100890 82780 101920
rect 82940 100890 85970 101920
rect 86130 100890 89160 101920
rect 89320 100890 92350 101920
rect 92510 100890 95540 101920
rect 95700 100890 98730 101920
rect 98890 100890 101920 101920
rect 102080 100890 105110 101920
rect 105270 100890 108300 101920
rect 108460 100890 111490 101920
rect 111650 100890 114680 101920
rect 114840 100890 117870 101920
rect 118030 100890 121060 101920
rect 121220 100890 124250 101920
rect 124410 100890 127440 101920
rect 127600 100890 130630 101920
rect 130790 100890 133820 101920
rect 133980 100890 137010 101920
rect 0 99890 137170 100890
rect 0 98890 3030 99890
rect 3190 98890 6220 99890
rect 6380 98890 9410 99890
rect 9570 98890 12600 99890
rect 12760 98890 15790 99890
rect 15950 98890 18980 99890
rect 19140 98890 22170 99890
rect 22330 98890 25360 99890
rect 25520 98890 28550 99890
rect 28710 98890 31740 99890
rect 31900 98890 34930 99890
rect 35090 98890 38120 99890
rect 38280 98890 41310 99890
rect 41470 98890 44500 99890
rect 44660 98890 47690 99890
rect 47850 98890 50880 99890
rect 51040 98890 54070 99890
rect 54230 98890 57260 99890
rect 57420 98890 60450 99890
rect 60610 98890 63640 99890
rect 63800 98890 66830 99890
rect 66990 98890 70020 99890
rect 70180 98890 73210 99890
rect 73370 98890 76400 99890
rect 76560 98890 79590 99890
rect 79750 98890 82780 99890
rect 82940 98890 85970 99890
rect 86130 98890 89160 99890
rect 89320 98890 92350 99890
rect 92510 98890 95540 99890
rect 95700 98890 98730 99890
rect 98890 98890 101920 99890
rect 102080 98890 105110 99890
rect 105270 98890 108300 99890
rect 108460 98890 111490 99890
rect 111650 98890 114680 99890
rect 114840 98890 117870 99890
rect 118030 98890 121060 99890
rect 121220 98890 124250 99890
rect 124410 98890 127440 99890
rect 127600 98890 130630 99890
rect 130790 98890 133820 99890
rect 133980 98890 137010 99890
rect 1000 98889 2000 98890
rect 4190 98889 5190 98890
rect 7380 98889 8380 98890
rect 10570 98730 11570 98890
rect 13760 98730 14760 98890
rect 16950 98730 17950 98890
rect 20140 98730 21140 98890
rect 23330 98730 24330 98890
rect 26520 98730 27520 98890
rect 29710 98730 30710 98890
rect 32900 98730 33900 98890
rect 36090 98730 37090 98890
rect 39280 98730 40280 98890
rect 42470 98730 43470 98890
rect 45660 98730 46660 98890
rect 48850 98730 49850 98890
rect 52040 98730 53040 98890
rect 55230 98730 56230 98890
rect 58420 98730 59420 98890
rect 61610 98730 62610 98890
rect 64800 98730 65800 98890
rect 67990 98730 68990 98890
rect 71180 98730 72180 98890
rect 74370 98730 75370 98890
rect 77560 98730 78560 98890
rect 80750 98730 81750 98890
rect 83940 98730 84940 98890
rect 87130 98730 88130 98890
rect 90320 98730 91320 98890
rect 93510 98730 94510 98890
rect 96700 98730 97700 98890
rect 99890 98730 100890 98890
rect 103080 98730 104080 98890
rect 106270 98730 107270 98890
rect 109460 98730 110460 98890
rect 112650 98730 113650 98890
rect 115840 98730 116840 98890
rect 119030 98730 120030 98890
rect 122220 98730 123220 98890
rect 125410 98730 126410 98890
rect 128600 98730 129600 98890
rect 131790 98730 132790 98890
rect 134980 98730 135980 98890
rect 0 98639 9370 98689
rect 0 79839 50 98639
rect 9320 79839 9370 98639
rect 9570 97700 12600 98730
rect 12760 97700 15790 98730
rect 15950 97700 18980 98730
rect 19140 97700 22170 98730
rect 22330 97700 25360 98730
rect 25520 97700 28550 98730
rect 28710 97700 31740 98730
rect 31900 97700 34930 98730
rect 35090 97700 38120 98730
rect 38280 97700 41310 98730
rect 41470 97700 44500 98730
rect 44660 97700 47690 98730
rect 47850 97700 50880 98730
rect 51040 97700 54070 98730
rect 54230 97700 57260 98730
rect 57420 97700 60450 98730
rect 60610 97700 63640 98730
rect 63800 97700 66830 98730
rect 66990 97700 70020 98730
rect 70180 97700 73210 98730
rect 73370 97700 76400 98730
rect 76560 97700 79590 98730
rect 79750 97700 82780 98730
rect 82940 97700 85970 98730
rect 86130 97700 89160 98730
rect 89320 97700 92350 98730
rect 92510 97700 95540 98730
rect 95700 97700 98730 98730
rect 98890 97700 101920 98730
rect 102080 97700 105110 98730
rect 105270 97700 108300 98730
rect 108460 97700 111490 98730
rect 111650 97700 114680 98730
rect 114840 97700 117870 98730
rect 118030 97700 121060 98730
rect 121220 97700 124250 98730
rect 124410 97700 127440 98730
rect 127600 97700 130630 98730
rect 130790 97700 133820 98730
rect 133980 97700 137010 98730
rect 9570 96700 137170 97700
rect 9570 95700 12600 96700
rect 12760 95700 15790 96700
rect 15950 95700 18980 96700
rect 19140 95700 22170 96700
rect 22330 95700 25360 96700
rect 25520 95700 28550 96700
rect 28710 95700 31740 96700
rect 31900 95700 34930 96700
rect 35090 95700 38120 96700
rect 38280 95700 41310 96700
rect 41470 95700 44500 96700
rect 44660 95700 47690 96700
rect 47850 95700 50880 96700
rect 51040 95700 54070 96700
rect 54230 95700 57260 96700
rect 57420 95700 60450 96700
rect 60610 95700 63640 96700
rect 63800 95700 66830 96700
rect 66990 95700 70020 96700
rect 70180 95700 73210 96700
rect 73370 95700 76400 96700
rect 76560 95700 79590 96700
rect 79750 95700 82780 96700
rect 82940 95700 85970 96700
rect 86130 95700 89160 96700
rect 89320 95700 92350 96700
rect 92510 95700 95540 96700
rect 95700 95700 98730 96700
rect 98890 95700 101920 96700
rect 102080 95700 105110 96700
rect 105270 95700 108300 96700
rect 108460 95700 111490 96700
rect 111650 95700 114680 96700
rect 114840 95700 117870 96700
rect 118030 95700 121060 96700
rect 121220 95700 124250 96700
rect 124410 95700 127440 96700
rect 127600 95700 130630 96700
rect 130790 95700 133820 96700
rect 133980 95700 137010 96700
rect 10570 95540 11570 95700
rect 13760 95540 14760 95700
rect 16950 95540 17950 95700
rect 20140 95540 21140 95700
rect 23330 95540 24330 95700
rect 26520 95540 27520 95700
rect 29710 95540 30710 95700
rect 32900 95540 33900 95700
rect 36090 95540 37090 95700
rect 39280 95540 40280 95700
rect 42470 95540 43470 95700
rect 45660 95540 46660 95700
rect 48850 95540 49850 95700
rect 52040 95540 53040 95700
rect 55230 95540 56230 95700
rect 58420 95540 59420 95700
rect 61610 95540 62610 95700
rect 64800 95540 65800 95700
rect 67990 95540 68990 95700
rect 71180 95540 72180 95700
rect 74370 95540 75370 95700
rect 77560 95540 78560 95700
rect 80750 95540 81750 95700
rect 83940 95540 84940 95700
rect 87130 95540 88130 95700
rect 90320 95540 91320 95700
rect 93510 95540 94510 95700
rect 96700 95540 97700 95700
rect 99890 95540 100890 95700
rect 103080 95540 104080 95700
rect 106270 95540 107270 95700
rect 109460 95540 110460 95700
rect 112650 95540 113650 95700
rect 115840 95540 116840 95700
rect 119030 95540 120030 95700
rect 122220 95540 123220 95700
rect 125410 95540 126410 95700
rect 128600 95540 129600 95700
rect 131790 95540 132790 95700
rect 134980 95540 135980 95700
rect 9570 94510 12600 95540
rect 12760 94510 15790 95540
rect 15950 94510 18980 95540
rect 19140 94510 22170 95540
rect 22330 94510 25360 95540
rect 25520 94510 28550 95540
rect 28710 94510 31740 95540
rect 31900 94510 34930 95540
rect 35090 94510 38120 95540
rect 38280 94510 41310 95540
rect 41470 94510 44500 95540
rect 44660 94510 47690 95540
rect 47850 94510 50880 95540
rect 51040 94510 54070 95540
rect 54230 94510 57260 95540
rect 57420 94510 60450 95540
rect 60610 94510 63640 95540
rect 63800 94510 66830 95540
rect 66990 94510 70020 95540
rect 70180 94510 73210 95540
rect 73370 94510 76400 95540
rect 76560 94510 79590 95540
rect 79750 94510 82780 95540
rect 82940 94510 85970 95540
rect 86130 94510 89160 95540
rect 89320 94510 92350 95540
rect 92510 94510 95540 95540
rect 95700 94510 98730 95540
rect 98890 94510 101920 95540
rect 102080 94510 105110 95540
rect 105270 94510 108300 95540
rect 108460 94510 111490 95540
rect 111650 94510 114680 95540
rect 114840 94510 117870 95540
rect 118030 94510 121060 95540
rect 121220 94510 124250 95540
rect 124410 94510 127440 95540
rect 127600 94510 130630 95540
rect 130790 94510 133820 95540
rect 133980 94510 137010 95540
rect 9570 93510 137170 94510
rect 9570 92510 12600 93510
rect 12760 92510 15790 93510
rect 15950 92510 18980 93510
rect 19140 92510 22170 93510
rect 22330 92510 25360 93510
rect 25520 92510 28550 93510
rect 28710 92510 31740 93510
rect 31900 92510 34930 93510
rect 35090 92510 38120 93510
rect 38280 92510 41310 93510
rect 41470 92510 44500 93510
rect 44660 92510 47690 93510
rect 47850 92510 50880 93510
rect 51040 92510 54070 93510
rect 54230 92510 57260 93510
rect 57420 92510 60450 93510
rect 60610 92510 63640 93510
rect 63800 92510 66830 93510
rect 66990 92510 70020 93510
rect 70180 92510 73210 93510
rect 73370 92510 76400 93510
rect 76560 92510 79590 93510
rect 79750 92510 82780 93510
rect 82940 92510 85970 93510
rect 86130 92510 89160 93510
rect 89320 92510 92350 93510
rect 92510 92510 95540 93510
rect 95700 92510 98730 93510
rect 98890 92510 101920 93510
rect 102080 92510 105110 93510
rect 105270 92510 108300 93510
rect 108460 92510 111490 93510
rect 111650 92510 114680 93510
rect 114840 92510 117870 93510
rect 118030 92510 121060 93510
rect 121220 92510 124250 93510
rect 124410 92510 127440 93510
rect 127600 92510 130630 93510
rect 130790 92510 133820 93510
rect 133980 92510 137010 93510
rect 10570 92350 11570 92510
rect 13760 92350 14760 92510
rect 16950 92350 17950 92510
rect 20140 92350 21140 92510
rect 23330 92350 24330 92510
rect 26520 92350 27520 92510
rect 29710 92350 30710 92510
rect 32900 92350 33900 92510
rect 36090 92350 37090 92510
rect 39280 92350 40280 92510
rect 42470 92350 43470 92510
rect 45660 92350 46660 92510
rect 48850 92350 49850 92510
rect 52040 92350 53040 92510
rect 55230 92350 56230 92510
rect 58420 92350 59420 92510
rect 61610 92350 62610 92510
rect 64800 92350 65800 92510
rect 67990 92350 68990 92510
rect 71180 92350 72180 92510
rect 74370 92350 75370 92510
rect 77560 92350 78560 92510
rect 80750 92350 81750 92510
rect 83940 92350 84940 92510
rect 87130 92350 88130 92510
rect 90320 92350 91320 92510
rect 93510 92350 94510 92510
rect 96700 92350 97700 92510
rect 99890 92350 100890 92510
rect 103080 92350 104080 92510
rect 106270 92350 107270 92510
rect 109460 92350 110460 92510
rect 112650 92350 113650 92510
rect 115840 92350 116840 92510
rect 119030 92350 120030 92510
rect 122220 92350 123220 92510
rect 125410 92350 126410 92510
rect 128600 92350 129600 92510
rect 131790 92350 132790 92510
rect 134980 92350 135980 92510
rect 9570 91320 12600 92350
rect 12760 91320 15790 92350
rect 15950 91320 18980 92350
rect 19140 91320 22170 92350
rect 22330 91320 25360 92350
rect 25520 91320 28550 92350
rect 28710 91320 31740 92350
rect 31900 91320 34930 92350
rect 35090 91320 38120 92350
rect 38280 91320 41310 92350
rect 41470 91320 44500 92350
rect 44660 91320 47690 92350
rect 47850 91320 50880 92350
rect 51040 91320 54070 92350
rect 54230 91320 57260 92350
rect 57420 91320 60450 92350
rect 60610 91320 63640 92350
rect 63800 91320 66830 92350
rect 66990 91320 70020 92350
rect 70180 91320 73210 92350
rect 73370 91320 76400 92350
rect 76560 91320 79590 92350
rect 79750 91320 82780 92350
rect 82940 91320 85970 92350
rect 86130 91320 89160 92350
rect 89320 91320 92350 92350
rect 92510 91320 95540 92350
rect 95700 91320 98730 92350
rect 98890 91320 101920 92350
rect 102080 91320 105110 92350
rect 105270 91320 108300 92350
rect 108460 91320 111490 92350
rect 111650 91320 114680 92350
rect 114840 91320 117870 92350
rect 118030 91320 121060 92350
rect 121220 91320 124250 92350
rect 124410 91320 127440 92350
rect 127600 91320 130630 92350
rect 130790 91320 133820 92350
rect 133980 91320 137010 92350
rect 9570 90320 137170 91320
rect 9570 89320 12600 90320
rect 12760 89320 15790 90320
rect 15950 89320 18980 90320
rect 19140 89320 22170 90320
rect 22330 89320 25360 90320
rect 25520 89320 28550 90320
rect 28710 89320 31740 90320
rect 31900 89320 34930 90320
rect 35090 89320 38120 90320
rect 38280 89320 41310 90320
rect 41470 89320 44500 90320
rect 44660 89320 47690 90320
rect 47850 89320 50880 90320
rect 51040 89320 54070 90320
rect 54230 89320 57260 90320
rect 57420 89320 60450 90320
rect 60610 89320 63640 90320
rect 63800 89320 66830 90320
rect 66990 89320 70020 90320
rect 70180 89320 73210 90320
rect 73370 89320 76400 90320
rect 76560 89320 79590 90320
rect 79750 89320 82780 90320
rect 82940 89320 85970 90320
rect 86130 89320 89160 90320
rect 89320 89320 92350 90320
rect 92510 89320 95540 90320
rect 95700 89320 98730 90320
rect 98890 89320 101920 90320
rect 102080 89320 105110 90320
rect 105270 89320 108300 90320
rect 108460 89320 111490 90320
rect 111650 89320 114680 90320
rect 114840 89320 117870 90320
rect 118030 89320 121060 90320
rect 121220 89320 124250 90320
rect 124410 89320 127440 90320
rect 127600 89320 130630 90320
rect 130790 89320 133820 90320
rect 133980 89320 137010 90320
rect 10570 89160 11570 89320
rect 13760 89160 14760 89320
rect 16950 89160 17950 89320
rect 20140 89160 21140 89320
rect 23330 89160 24330 89320
rect 26520 89160 27520 89320
rect 29710 89160 30710 89320
rect 32900 89160 33900 89320
rect 36090 89160 37090 89320
rect 39280 89160 40280 89320
rect 42470 89160 43470 89320
rect 45660 89160 46660 89320
rect 48850 89160 49850 89320
rect 52040 89160 53040 89320
rect 55230 89160 56230 89320
rect 58420 89160 59420 89320
rect 61610 89160 62610 89320
rect 64800 89160 65800 89320
rect 67990 89160 68990 89320
rect 71180 89160 72180 89320
rect 74370 89160 75370 89320
rect 77560 89160 78560 89320
rect 80750 89160 81750 89320
rect 83940 89160 84940 89320
rect 87130 89160 88130 89320
rect 90320 89160 91320 89320
rect 93510 89160 94510 89320
rect 96700 89160 97700 89320
rect 99890 89160 100890 89320
rect 103080 89160 104080 89320
rect 106270 89160 107270 89320
rect 109460 89160 110460 89320
rect 112650 89160 113650 89320
rect 115840 89160 116840 89320
rect 119030 89160 120030 89320
rect 122220 89160 123220 89320
rect 125410 89160 126410 89320
rect 128600 89160 129600 89320
rect 131790 89160 132790 89320
rect 134980 89160 135980 89320
rect 9570 88130 12600 89160
rect 12760 88130 15790 89160
rect 15950 88130 18980 89160
rect 19140 88130 22170 89160
rect 22330 88130 25360 89160
rect 25520 88130 28550 89160
rect 28710 88130 31740 89160
rect 31900 88130 34930 89160
rect 35090 88130 38120 89160
rect 38280 88130 41310 89160
rect 41470 88130 44500 89160
rect 44660 88130 47690 89160
rect 47850 88130 50880 89160
rect 51040 88130 54070 89160
rect 54230 88130 57260 89160
rect 57420 88130 60450 89160
rect 60610 88130 63640 89160
rect 63800 88130 66830 89160
rect 66990 88130 70020 89160
rect 70180 88130 73210 89160
rect 73370 88130 76400 89160
rect 76560 88130 79590 89160
rect 79750 88130 82780 89160
rect 82940 88130 85970 89160
rect 86130 88130 89160 89160
rect 89320 88130 92350 89160
rect 92510 88130 95540 89160
rect 95700 88130 98730 89160
rect 98890 88130 101920 89160
rect 102080 88130 105110 89160
rect 105270 88130 108300 89160
rect 108460 88130 111490 89160
rect 111650 88130 114680 89160
rect 114840 88130 117870 89160
rect 118030 88130 121060 89160
rect 121220 88130 124250 89160
rect 124410 88130 127440 89160
rect 127600 88130 130630 89160
rect 130790 88130 133820 89160
rect 133980 88130 137010 89160
rect 9570 87130 137170 88130
rect 9570 86130 12600 87130
rect 12760 86130 15790 87130
rect 15950 86130 18980 87130
rect 19140 86130 22170 87130
rect 22330 86130 25360 87130
rect 25520 86130 28550 87130
rect 28710 86130 31740 87130
rect 31900 86130 34930 87130
rect 35090 86130 38120 87130
rect 38280 86130 41310 87130
rect 41470 86130 44500 87130
rect 44660 86130 47690 87130
rect 47850 86130 50880 87130
rect 51040 86130 54070 87130
rect 54230 86130 57260 87130
rect 57420 86130 60450 87130
rect 60610 86130 63640 87130
rect 63800 86130 66830 87130
rect 66990 86130 70020 87130
rect 70180 86130 73210 87130
rect 73370 86130 76400 87130
rect 76560 86130 79590 87130
rect 79750 86130 82780 87130
rect 82940 86130 85970 87130
rect 86130 86130 89160 87130
rect 89320 86130 92350 87130
rect 92510 86130 95540 87130
rect 95700 86130 98730 87130
rect 98890 86130 101920 87130
rect 102080 86130 105110 87130
rect 105270 86130 108300 87130
rect 108460 86130 111490 87130
rect 111650 86130 114680 87130
rect 114840 86130 117870 87130
rect 118030 86130 121060 87130
rect 121220 86130 124250 87130
rect 124410 86130 127440 87130
rect 127600 86130 130630 87130
rect 130790 86130 133820 87130
rect 133980 86130 137010 87130
rect 10570 85970 11570 86130
rect 13760 85970 14760 86130
rect 16950 85970 17950 86130
rect 20140 85970 21140 86130
rect 23330 85970 24330 86130
rect 26520 85970 27520 86130
rect 29710 85970 30710 86130
rect 32900 85970 33900 86130
rect 36090 85970 37090 86130
rect 39280 85970 40280 86130
rect 42470 85970 43470 86130
rect 45660 85970 46660 86130
rect 48850 85970 49850 86130
rect 52040 85970 53040 86130
rect 55230 85970 56230 86130
rect 58420 85970 59420 86130
rect 61610 85970 62610 86130
rect 64800 85970 65800 86130
rect 67990 85970 68990 86130
rect 71180 85970 72180 86130
rect 74370 85970 75370 86130
rect 77560 85970 78560 86130
rect 80750 85970 81750 86130
rect 83940 85970 84940 86130
rect 87130 85970 88130 86130
rect 90320 85970 91320 86130
rect 93510 85970 94510 86130
rect 96700 85970 97700 86130
rect 99890 85970 100890 86130
rect 103080 85970 104080 86130
rect 106270 85970 107270 86130
rect 109460 85970 110460 86130
rect 112650 85970 113650 86130
rect 115840 85970 116840 86130
rect 119030 85970 120030 86130
rect 122220 85970 123220 86130
rect 125410 85970 126410 86130
rect 128600 85970 129600 86130
rect 131790 85970 132790 86130
rect 134980 85970 135980 86130
rect 9570 84940 12600 85970
rect 12760 84940 15790 85970
rect 15950 84940 18980 85970
rect 19140 84940 22170 85970
rect 22330 84940 25360 85970
rect 25520 84940 28550 85970
rect 28710 84940 31740 85970
rect 31900 84940 34930 85970
rect 35090 84940 38120 85970
rect 38280 84940 41310 85970
rect 41470 84940 44500 85970
rect 44660 84940 47690 85970
rect 47850 84940 50880 85970
rect 51040 84940 54070 85970
rect 54230 84940 57260 85970
rect 57420 84940 60450 85970
rect 60610 84940 63640 85970
rect 63800 84940 66830 85970
rect 66990 84940 70020 85970
rect 70180 84940 73210 85970
rect 73370 84940 76400 85970
rect 76560 84940 79590 85970
rect 79750 84940 82780 85970
rect 82940 84940 85970 85970
rect 86130 84940 89160 85970
rect 89320 84940 92350 85970
rect 92510 84940 95540 85970
rect 95700 84940 98730 85970
rect 98890 84940 101920 85970
rect 102080 84940 105110 85970
rect 105270 84940 108300 85970
rect 108460 84940 111490 85970
rect 111650 84940 114680 85970
rect 114840 84940 117870 85970
rect 118030 84940 121060 85970
rect 121220 84940 124250 85970
rect 124410 84940 127440 85970
rect 127600 84940 130630 85970
rect 130790 84940 133820 85970
rect 133980 84940 137010 85970
rect 9570 83940 137170 84940
rect 9570 82940 12600 83940
rect 12760 82940 15790 83940
rect 15950 82940 18980 83940
rect 19140 82940 22170 83940
rect 22330 82940 25360 83940
rect 25520 82940 28550 83940
rect 28710 82940 31740 83940
rect 31900 82940 34930 83940
rect 35090 82940 38120 83940
rect 38280 82940 41310 83940
rect 41470 82940 44500 83940
rect 44660 82940 47690 83940
rect 47850 82940 50880 83940
rect 51040 82940 54070 83940
rect 54230 82940 57260 83940
rect 57420 82940 60450 83940
rect 60610 82940 63640 83940
rect 63800 82940 66830 83940
rect 66990 82940 70020 83940
rect 70180 82940 73210 83940
rect 73370 82940 76400 83940
rect 76560 82940 79590 83940
rect 79750 82940 82780 83940
rect 82940 82940 85970 83940
rect 86130 82940 89160 83940
rect 89320 82940 92350 83940
rect 92510 82940 95540 83940
rect 95700 82940 98730 83940
rect 98890 82940 101920 83940
rect 102080 82940 105110 83940
rect 105270 82940 108300 83940
rect 108460 82940 111490 83940
rect 111650 82940 114680 83940
rect 114840 82940 117870 83940
rect 118030 82940 121060 83940
rect 121220 82940 124250 83940
rect 124410 82940 127440 83940
rect 127600 82940 130630 83940
rect 130790 82940 133820 83940
rect 133980 82940 137010 83940
rect 10570 82780 11570 82940
rect 13760 82780 14760 82940
rect 16950 82780 17950 82940
rect 20140 82780 21140 82940
rect 23330 82780 24330 82940
rect 26520 82780 27520 82940
rect 29710 82780 30710 82940
rect 32900 82780 33900 82940
rect 36090 82780 37090 82940
rect 39280 82780 40280 82940
rect 42470 82780 43470 82940
rect 45660 82780 46660 82940
rect 48850 82780 49850 82940
rect 52040 82780 53040 82940
rect 55230 82780 56230 82940
rect 58420 82780 59420 82940
rect 61610 82780 62610 82940
rect 64800 82780 65800 82940
rect 67990 82780 68990 82940
rect 71180 82780 72180 82940
rect 74370 82780 75370 82940
rect 77560 82780 78560 82940
rect 80750 82780 81750 82940
rect 83940 82780 84940 82940
rect 87130 82780 88130 82940
rect 90320 82780 91320 82940
rect 93510 82780 94510 82940
rect 96700 82780 97700 82940
rect 99890 82780 100890 82940
rect 103080 82780 104080 82940
rect 106270 82780 107270 82940
rect 109460 82780 110460 82940
rect 112650 82780 113650 82940
rect 115840 82780 116840 82940
rect 119030 82780 120030 82940
rect 122220 82780 123220 82940
rect 125410 82780 126410 82940
rect 128600 82780 129600 82940
rect 131790 82780 132790 82940
rect 134980 82780 135980 82940
rect 0 79789 9370 79839
rect 9570 81750 12600 82780
rect 12760 81750 15790 82780
rect 15950 81750 18980 82780
rect 19140 81750 22170 82780
rect 22330 81750 25360 82780
rect 25520 81750 28550 82780
rect 28710 81750 31740 82780
rect 31900 81750 34930 82780
rect 35090 81750 38120 82780
rect 38280 81750 41310 82780
rect 41470 81750 44500 82780
rect 44660 81750 47690 82780
rect 47850 81750 50880 82780
rect 51040 81750 54070 82780
rect 54230 81750 57260 82780
rect 57420 81750 60450 82780
rect 60610 81750 63640 82780
rect 63800 81750 66830 82780
rect 66990 81750 70020 82780
rect 70180 81750 73210 82780
rect 73370 81750 76400 82780
rect 76560 81750 79590 82780
rect 79750 81750 82780 82780
rect 82940 81750 85970 82780
rect 86130 81750 89160 82780
rect 89320 81750 92350 82780
rect 92510 81750 95540 82780
rect 95700 81750 98730 82780
rect 98890 81750 101920 82780
rect 102080 81750 105110 82780
rect 105270 81750 108300 82780
rect 108460 81750 111490 82780
rect 111650 81750 114680 82780
rect 114840 81750 117870 82780
rect 118030 81750 121060 82780
rect 121220 81750 124250 82780
rect 124410 81750 127440 82780
rect 127600 81750 130630 82780
rect 130790 81750 133820 82780
rect 133980 81750 137010 82780
rect 9570 80750 137170 81750
rect 9570 79750 12600 80750
rect 12760 79750 15790 80750
rect 15950 79750 18980 80750
rect 19140 79750 22170 80750
rect 22330 79750 25360 80750
rect 25520 79750 28550 80750
rect 28710 79750 31740 80750
rect 31900 79750 34930 80750
rect 35090 79750 38120 80750
rect 38280 79750 41310 80750
rect 41470 79750 44500 80750
rect 44660 79750 47690 80750
rect 47850 79750 50880 80750
rect 51040 79750 54070 80750
rect 54230 79750 57260 80750
rect 57420 79750 60450 80750
rect 60610 79750 63640 80750
rect 63800 79750 66830 80750
rect 66990 79750 70020 80750
rect 70180 79750 73210 80750
rect 73370 79750 76400 80750
rect 76560 79750 79590 80750
rect 79750 79750 82780 80750
rect 82940 79750 85970 80750
rect 86130 79750 89160 80750
rect 89320 79750 92350 80750
rect 92510 79750 95540 80750
rect 95700 79750 98730 80750
rect 98890 79750 101920 80750
rect 102080 79750 105110 80750
rect 105270 79750 108300 80750
rect 108460 79750 111490 80750
rect 111650 79750 114680 80750
rect 114840 79750 117870 80750
rect 118030 79750 121060 80750
rect 121220 79750 124250 80750
rect 124410 79750 127440 80750
rect 127600 79750 130630 80750
rect 130790 79750 133820 80750
rect 133980 79750 137010 80750
rect 10570 79590 11570 79750
rect 13760 79590 14760 79750
rect 16950 79590 17950 79750
rect 20140 79590 21140 79750
rect 23330 79590 24330 79750
rect 26520 79590 27520 79750
rect 29710 79590 30710 79750
rect 32900 79590 33900 79750
rect 36090 79590 37090 79750
rect 39280 79590 40280 79750
rect 42470 79590 43470 79750
rect 45660 79590 46660 79750
rect 48850 79590 49850 79750
rect 52040 79590 53040 79750
rect 55230 79590 56230 79750
rect 58420 79590 59420 79750
rect 61610 79590 62610 79750
rect 64800 79590 65800 79750
rect 67990 79590 68990 79750
rect 71180 79590 72180 79750
rect 74370 79590 75370 79750
rect 77560 79590 78560 79750
rect 80750 79590 81750 79750
rect 83940 79590 84940 79750
rect 87130 79590 88130 79750
rect 90320 79590 91320 79750
rect 93510 79590 94510 79750
rect 96700 79590 97700 79750
rect 99890 79590 100890 79750
rect 103080 79590 104080 79750
rect 106270 79590 107270 79750
rect 109460 79590 110460 79750
rect 112650 79590 113650 79750
rect 115840 79590 116840 79750
rect 119030 79590 120030 79750
rect 122220 79590 123220 79750
rect 125410 79590 126410 79750
rect 128600 79590 129600 79750
rect 131790 79590 132790 79750
rect 134980 79590 135980 79750
rect 0 78560 3030 79589
rect 3190 78560 6220 79589
rect 6380 78560 9410 79589
rect 9570 78560 12600 79590
rect 12760 78560 15790 79590
rect 15950 78560 18980 79590
rect 19140 78560 22170 79590
rect 22330 78560 25360 79590
rect 25520 78560 28550 79590
rect 28710 78560 31740 79590
rect 31900 78560 34930 79590
rect 35090 78560 38120 79590
rect 38280 78560 41310 79590
rect 41470 78560 44500 79590
rect 44660 78560 47690 79590
rect 47850 78560 50880 79590
rect 51040 78560 54070 79590
rect 54230 78560 57260 79590
rect 57420 78560 60450 79590
rect 60610 78560 63640 79590
rect 63800 78560 66830 79590
rect 66990 78560 70020 79590
rect 70180 78560 73210 79590
rect 73370 78560 76400 79590
rect 76560 78560 79590 79590
rect 79750 78560 82780 79590
rect 82940 78560 85970 79590
rect 86130 78560 89160 79590
rect 89320 78560 92350 79590
rect 92510 78560 95540 79590
rect 95700 78560 98730 79590
rect 98890 78560 101920 79590
rect 102080 78560 105110 79590
rect 105270 78560 108300 79590
rect 108460 78560 111490 79590
rect 111650 78560 114680 79590
rect 114840 78560 117870 79590
rect 118030 78560 121060 79590
rect 121220 78560 124250 79590
rect 124410 78560 127440 79590
rect 127600 78560 130630 79590
rect 130790 78560 133820 79590
rect 133980 78560 137010 79590
rect 0 77560 137170 78560
rect 0 76560 3030 77560
rect 3190 76560 6220 77560
rect 6380 76560 9410 77560
rect 9570 76560 12600 77560
rect 12760 76560 15790 77560
rect 15950 76560 18980 77560
rect 19140 76560 22170 77560
rect 22330 76560 25360 77560
rect 25520 76560 28550 77560
rect 28710 76560 31740 77560
rect 31900 76560 34930 77560
rect 35090 76560 38120 77560
rect 38280 76560 41310 77560
rect 41470 76560 44500 77560
rect 44660 76560 47690 77560
rect 47850 76560 50880 77560
rect 51040 76560 54070 77560
rect 54230 76560 57260 77560
rect 57420 76560 60450 77560
rect 60610 76560 63640 77560
rect 63800 76560 66830 77560
rect 66990 76560 70020 77560
rect 70180 76560 73210 77560
rect 73370 76560 76400 77560
rect 76560 76560 79590 77560
rect 79750 76560 82780 77560
rect 82940 76560 85970 77560
rect 86130 76560 89160 77560
rect 89320 76560 92350 77560
rect 92510 76560 95540 77560
rect 95700 76560 98730 77560
rect 98890 76560 101920 77560
rect 102080 76560 105110 77560
rect 105270 76560 108300 77560
rect 108460 76560 111490 77560
rect 111650 76560 114680 77560
rect 114840 76560 117870 77560
rect 118030 76560 121060 77560
rect 121220 76560 124250 77560
rect 124410 76560 127440 77560
rect 127600 76560 130630 77560
rect 130790 76560 133820 77560
rect 133980 76560 137010 77560
rect 1000 76400 2000 76560
rect 4190 76400 5190 76560
rect 7380 76400 8380 76560
rect 10570 76400 11570 76560
rect 13760 76400 14760 76560
rect 16950 76400 17950 76560
rect 20140 76400 21140 76560
rect 23330 76400 24330 76560
rect 26520 76400 27520 76560
rect 29710 76400 30710 76560
rect 32900 76400 33900 76560
rect 36090 76400 37090 76560
rect 39280 76400 40280 76560
rect 42470 76400 43470 76560
rect 45660 76400 46660 76560
rect 48850 76400 49850 76560
rect 52040 76400 53040 76560
rect 55230 76400 56230 76560
rect 58420 76400 59420 76560
rect 61610 76400 62610 76560
rect 64800 76400 65800 76560
rect 67990 76400 68990 76560
rect 71180 76400 72180 76560
rect 74370 76400 75370 76560
rect 77560 76400 78560 76560
rect 80750 76400 81750 76560
rect 83940 76400 84940 76560
rect 87130 76400 88130 76560
rect 90320 76400 91320 76560
rect 93510 76400 94510 76560
rect 96700 76400 97700 76560
rect 99890 76400 100890 76560
rect 103080 76400 104080 76560
rect 106270 76400 107270 76560
rect 109460 76400 110460 76560
rect 112650 76400 113650 76560
rect 115840 76400 116840 76560
rect 119030 76400 120030 76560
rect 122220 76400 123220 76560
rect 125410 76400 126410 76560
rect 128600 76400 129600 76560
rect 131790 76400 132790 76560
rect 134980 76400 135980 76560
rect 0 75370 3030 76400
rect 3190 75370 6220 76400
rect 6380 75370 9410 76400
rect 9570 75370 12600 76400
rect 12760 75370 15790 76400
rect 15950 75370 18980 76400
rect 19140 75370 22170 76400
rect 22330 75370 25360 76400
rect 25520 75370 28550 76400
rect 28710 75370 31740 76400
rect 31900 75370 34930 76400
rect 35090 75370 38120 76400
rect 38280 75370 41310 76400
rect 41470 75370 44500 76400
rect 44660 75370 47690 76400
rect 47850 75370 50880 76400
rect 51040 75370 54070 76400
rect 54230 75370 57260 76400
rect 57420 75370 60450 76400
rect 60610 75370 63640 76400
rect 63800 75370 66830 76400
rect 66990 75370 70020 76400
rect 70180 75370 73210 76400
rect 73370 75370 76400 76400
rect 76560 75370 79590 76400
rect 79750 75370 82780 76400
rect 82940 75370 85970 76400
rect 86130 75370 89160 76400
rect 89320 75370 92350 76400
rect 92510 75370 95540 76400
rect 95700 75370 98730 76400
rect 98890 75370 101920 76400
rect 102080 75370 105110 76400
rect 105270 75370 108300 76400
rect 108460 75370 111490 76400
rect 111650 75370 114680 76400
rect 114840 75370 117870 76400
rect 118030 75370 121060 76400
rect 121220 75370 124250 76400
rect 124410 75370 127440 76400
rect 127600 75370 130630 76400
rect 130790 75370 133820 76400
rect 133980 75370 137010 76400
rect 0 74370 137170 75370
rect 0 73370 3030 74370
rect 3190 73370 6220 74370
rect 6380 73370 9410 74370
rect 9570 73370 12600 74370
rect 12760 73370 15790 74370
rect 15950 73370 18980 74370
rect 19140 73370 22170 74370
rect 22330 73370 25360 74370
rect 25520 73370 28550 74370
rect 28710 73370 31740 74370
rect 31900 73370 34930 74370
rect 35090 73370 38120 74370
rect 38280 73370 41310 74370
rect 41470 73370 44500 74370
rect 44660 73370 47690 74370
rect 47850 73370 50880 74370
rect 51040 73370 54070 74370
rect 54230 73370 57260 74370
rect 57420 73370 60450 74370
rect 60610 73370 63640 74370
rect 63800 73370 66830 74370
rect 66990 73370 70020 74370
rect 70180 73370 73210 74370
rect 73370 73370 76400 74370
rect 76560 73370 79590 74370
rect 79750 73370 82780 74370
rect 82940 73370 85970 74370
rect 86130 73370 89160 74370
rect 89320 73370 92350 74370
rect 92510 73370 95540 74370
rect 95700 73370 98730 74370
rect 98890 73370 101920 74370
rect 102080 73370 105110 74370
rect 105270 73370 108300 74370
rect 108460 73370 111490 74370
rect 111650 73370 114680 74370
rect 114840 73370 117870 74370
rect 118030 73370 121060 74370
rect 121220 73370 124250 74370
rect 124410 73370 127440 74370
rect 127600 73370 130630 74370
rect 130790 73370 133820 74370
rect 133980 73370 137010 74370
rect 1000 73210 2000 73370
rect 4190 73210 5190 73370
rect 7380 73210 8380 73370
rect 10570 73210 11570 73370
rect 13760 73210 14760 73370
rect 16950 73210 17950 73370
rect 20140 73210 21140 73370
rect 23330 73210 24330 73370
rect 26520 73210 27520 73370
rect 29710 73210 30710 73370
rect 32900 73210 33900 73370
rect 36090 73210 37090 73370
rect 39280 73210 40280 73370
rect 42470 73210 43470 73370
rect 45660 73210 46660 73370
rect 48850 73210 49850 73370
rect 52040 73210 53040 73370
rect 55230 73210 56230 73370
rect 58420 73210 59420 73370
rect 61610 73210 62610 73370
rect 64800 73210 65800 73370
rect 67990 73210 68990 73370
rect 71180 73210 72180 73370
rect 74370 73210 75370 73370
rect 77560 73210 78560 73370
rect 80750 73210 81750 73370
rect 83940 73210 84940 73370
rect 87130 73210 88130 73370
rect 90320 73210 91320 73370
rect 93510 73210 94510 73370
rect 96700 73210 97700 73370
rect 99890 73210 100890 73370
rect 103080 73210 104080 73370
rect 106270 73210 107270 73370
rect 109460 73210 110460 73370
rect 112650 73210 113650 73370
rect 115840 73210 116840 73370
rect 119030 73210 120030 73370
rect 122220 73210 123220 73370
rect 125410 73210 126410 73370
rect 128600 73210 129600 73370
rect 131790 73210 132790 73370
rect 134980 73210 135980 73370
rect 0 72180 3030 73210
rect 3190 72180 6220 73210
rect 6380 72180 9410 73210
rect 9570 72180 12600 73210
rect 12760 72180 15790 73210
rect 15950 72180 18980 73210
rect 19140 72180 22170 73210
rect 22330 72180 25360 73210
rect 25520 72180 28550 73210
rect 28710 72180 31740 73210
rect 31900 72180 34930 73210
rect 35090 72180 38120 73210
rect 38280 72180 41310 73210
rect 41470 72180 44500 73210
rect 44660 72180 47690 73210
rect 47850 72180 50880 73210
rect 51040 72180 54070 73210
rect 54230 72180 57260 73210
rect 57420 72180 60450 73210
rect 60610 72180 63640 73210
rect 63800 72180 66830 73210
rect 66990 72180 70020 73210
rect 70180 72180 73210 73210
rect 73370 72180 76400 73210
rect 76560 72180 79590 73210
rect 79750 72180 82780 73210
rect 82940 72180 85970 73210
rect 86130 72180 89160 73210
rect 89320 72180 92350 73210
rect 92510 72180 95540 73210
rect 95700 72180 98730 73210
rect 98890 72180 101920 73210
rect 102080 72180 105110 73210
rect 105270 72180 108300 73210
rect 108460 72180 111490 73210
rect 111650 72180 114680 73210
rect 114840 72180 117870 73210
rect 118030 72180 121060 73210
rect 121220 72180 124250 73210
rect 124410 72180 127440 73210
rect 127600 72180 130630 73210
rect 130790 72180 133820 73210
rect 133980 72180 137010 73210
rect 0 71180 137170 72180
rect 0 70180 3030 71180
rect 3190 70180 6220 71180
rect 6380 70180 9410 71180
rect 9570 70180 12600 71180
rect 12760 70180 15790 71180
rect 15950 70180 18980 71180
rect 19140 70180 22170 71180
rect 22330 70180 25360 71180
rect 25520 70180 28550 71180
rect 28710 70180 31740 71180
rect 31900 70180 34930 71180
rect 35090 70180 38120 71180
rect 38280 70180 41310 71180
rect 41470 70180 44500 71180
rect 44660 70180 47690 71180
rect 47850 70180 50880 71180
rect 51040 70180 54070 71180
rect 54230 70180 57260 71180
rect 57420 70180 60450 71180
rect 60610 70180 63640 71180
rect 63800 70180 66830 71180
rect 66990 70180 70020 71180
rect 70180 70180 73210 71180
rect 73370 70180 76400 71180
rect 76560 70180 79590 71180
rect 79750 70180 82780 71180
rect 82940 70180 85970 71180
rect 86130 70180 89160 71180
rect 89320 70180 92350 71180
rect 92510 70180 95540 71180
rect 95700 70180 98730 71180
rect 98890 70180 101920 71180
rect 102080 70180 105110 71180
rect 105270 70180 108300 71180
rect 108460 70180 111490 71180
rect 111650 70180 114680 71180
rect 114840 70180 117870 71180
rect 118030 70180 121060 71180
rect 121220 70180 124250 71180
rect 124410 70180 127440 71180
rect 127600 70180 130630 71180
rect 130790 70180 133820 71180
rect 133980 70180 137010 71180
rect 1000 70020 2000 70180
rect 4190 70020 5190 70180
rect 7380 70020 8380 70180
rect 10570 70020 11570 70180
rect 13760 70020 14760 70180
rect 16950 70020 17950 70180
rect 20140 70020 21140 70180
rect 23330 70020 24330 70180
rect 26520 70020 27520 70180
rect 29710 70020 30710 70180
rect 32900 70020 33900 70180
rect 36090 70020 37090 70180
rect 39280 70020 40280 70180
rect 42470 70020 43470 70180
rect 45660 70020 46660 70180
rect 48850 70020 49850 70180
rect 52040 70020 53040 70180
rect 55230 70020 56230 70180
rect 58420 70020 59420 70180
rect 61610 70020 62610 70180
rect 64800 70020 65800 70180
rect 67990 70020 68990 70180
rect 71180 70020 72180 70180
rect 74370 70020 75370 70180
rect 77560 70020 78560 70180
rect 80750 70020 81750 70180
rect 83940 70020 84940 70180
rect 87130 70020 88130 70180
rect 90320 70020 91320 70180
rect 93510 70020 94510 70180
rect 96700 70020 97700 70180
rect 99890 70020 100890 70180
rect 103080 70020 104080 70180
rect 106270 70020 107270 70180
rect 109460 70020 110460 70180
rect 112650 70020 113650 70180
rect 115840 70020 116840 70180
rect 119030 70020 120030 70180
rect 122220 70020 123220 70180
rect 125410 70020 126410 70180
rect 128600 70020 129600 70180
rect 131790 70020 132790 70180
rect 134980 70020 135980 70180
rect 0 68990 3030 70020
rect 3190 68990 6220 70020
rect 6380 68990 9410 70020
rect 9570 68990 12600 70020
rect 12760 68990 15790 70020
rect 15950 68990 18980 70020
rect 19140 68990 22170 70020
rect 22330 68990 25360 70020
rect 25520 68990 28550 70020
rect 28710 68990 31740 70020
rect 31900 68990 34930 70020
rect 35090 68990 38120 70020
rect 38280 68990 41310 70020
rect 41470 68990 44500 70020
rect 44660 68990 47690 70020
rect 47850 68990 50880 70020
rect 51040 68990 54070 70020
rect 54230 68990 57260 70020
rect 57420 68990 60450 70020
rect 60610 68990 63640 70020
rect 63800 68990 66830 70020
rect 66990 68990 70020 70020
rect 70180 68990 73210 70020
rect 73370 68990 76400 70020
rect 76560 68990 79590 70020
rect 79750 68990 82780 70020
rect 82940 68990 85970 70020
rect 86130 68990 89160 70020
rect 89320 68990 92350 70020
rect 92510 68990 95540 70020
rect 95700 68990 98730 70020
rect 98890 68990 101920 70020
rect 102080 68990 105110 70020
rect 105270 68990 108300 70020
rect 108460 68990 111490 70020
rect 111650 68990 114680 70020
rect 114840 68990 117870 70020
rect 118030 68990 121060 70020
rect 121220 68990 124250 70020
rect 124410 68990 127440 70020
rect 127600 68990 130630 70020
rect 130790 68990 133820 70020
rect 133980 68990 137010 70020
rect 0 67990 137170 68990
rect 0 66990 3030 67990
rect 3190 66990 6220 67990
rect 6380 66990 9410 67990
rect 9570 66990 12600 67990
rect 12760 66990 15790 67990
rect 15950 66990 18980 67990
rect 19140 66990 22170 67990
rect 22330 66990 25360 67990
rect 25520 66990 28550 67990
rect 28710 66990 31740 67990
rect 31900 66990 34930 67990
rect 35090 66990 38120 67990
rect 38280 66990 41310 67990
rect 41470 66990 44500 67990
rect 44660 66990 47690 67990
rect 47850 66990 50880 67990
rect 51040 66990 54070 67990
rect 54230 66990 57260 67990
rect 57420 66990 60450 67990
rect 60610 66990 63640 67990
rect 63800 66990 66830 67990
rect 66990 66990 70020 67990
rect 70180 66990 73210 67990
rect 73370 66990 76400 67990
rect 76560 66990 79590 67990
rect 79750 66990 82780 67990
rect 82940 66990 85970 67990
rect 86130 66990 89160 67990
rect 89320 66990 92350 67990
rect 92510 66990 95540 67990
rect 95700 66990 98730 67990
rect 98890 66990 101920 67990
rect 102080 66990 105110 67990
rect 105270 66990 108300 67990
rect 108460 66990 111490 67990
rect 111650 66990 114680 67990
rect 114840 66990 117870 67990
rect 118030 66990 121060 67990
rect 121220 66990 124250 67990
rect 124410 66990 127440 67990
rect 127600 66990 130630 67990
rect 130790 66990 133820 67990
rect 133980 66990 137010 67990
rect 1000 66830 2000 66990
rect 4190 66830 5190 66990
rect 7380 66830 8380 66990
rect 10570 66830 11570 66990
rect 13760 66830 14760 66990
rect 16950 66830 17950 66990
rect 20140 66830 21140 66990
rect 23330 66830 24330 66990
rect 26520 66830 27520 66990
rect 29710 66830 30710 66990
rect 32900 66830 33900 66990
rect 36090 66830 37090 66990
rect 39280 66830 40280 66990
rect 42470 66830 43470 66990
rect 45660 66830 46660 66990
rect 48850 66830 49850 66990
rect 52040 66830 53040 66990
rect 55230 66830 56230 66990
rect 58420 66830 59420 66990
rect 61610 66830 62610 66990
rect 64800 66830 65800 66990
rect 67990 66830 68990 66990
rect 71180 66830 72180 66990
rect 74370 66830 75370 66990
rect 77560 66830 78560 66990
rect 80750 66830 81750 66990
rect 83940 66830 84940 66990
rect 87130 66830 88130 66990
rect 90320 66830 91320 66990
rect 93510 66830 94510 66990
rect 96700 66830 97700 66990
rect 99890 66830 100890 66990
rect 103080 66830 104080 66990
rect 106270 66830 107270 66990
rect 109460 66830 110460 66990
rect 112650 66830 113650 66990
rect 115840 66830 116840 66990
rect 119030 66830 120030 66990
rect 122220 66830 123220 66990
rect 125410 66830 126410 66990
rect 128600 66830 129600 66990
rect 131790 66830 132790 66990
rect 134980 66830 135980 66990
rect 0 65800 3030 66830
rect 3190 65800 6220 66830
rect 6380 65800 9410 66830
rect 9570 65800 12600 66830
rect 12760 65800 15790 66830
rect 15950 65800 18980 66830
rect 19140 65800 22170 66830
rect 22330 65800 25360 66830
rect 25520 65800 28550 66830
rect 28710 65800 31740 66830
rect 31900 65800 34930 66830
rect 35090 65800 38120 66830
rect 38280 65800 41310 66830
rect 41470 65800 44500 66830
rect 44660 65800 47690 66830
rect 47850 65800 50880 66830
rect 51040 65800 54070 66830
rect 54230 65800 57260 66830
rect 57420 65800 60450 66830
rect 60610 65800 63640 66830
rect 63800 65800 66830 66830
rect 66990 65800 70020 66830
rect 70180 65800 73210 66830
rect 73370 65800 76400 66830
rect 76560 65800 79590 66830
rect 79750 65800 82780 66830
rect 82940 65800 85970 66830
rect 86130 65800 89160 66830
rect 89320 65800 92350 66830
rect 92510 65800 95540 66830
rect 95700 65800 98730 66830
rect 98890 65800 101920 66830
rect 102080 65800 105110 66830
rect 105270 65800 108300 66830
rect 108460 65800 111490 66830
rect 111650 65800 114680 66830
rect 114840 65800 117870 66830
rect 118030 65800 121060 66830
rect 121220 65800 124250 66830
rect 124410 65800 127440 66830
rect 127600 65800 130630 66830
rect 130790 65800 133820 66830
rect 133980 65800 137010 66830
rect 0 64800 137170 65800
rect 0 63800 3030 64800
rect 3190 63800 6220 64800
rect 6380 63800 9410 64800
rect 9570 63800 12600 64800
rect 12760 63800 15790 64800
rect 15950 63800 18980 64800
rect 19140 63800 22170 64800
rect 22330 63800 25360 64800
rect 25520 63800 28550 64800
rect 28710 63800 31740 64800
rect 31900 63800 34930 64800
rect 35090 63800 38120 64800
rect 38280 63800 41310 64800
rect 41470 63800 44500 64800
rect 44660 63800 47690 64800
rect 47850 63800 50880 64800
rect 51040 63800 54070 64800
rect 54230 63800 57260 64800
rect 57420 63800 60450 64800
rect 60610 63800 63640 64800
rect 63800 63800 66830 64800
rect 66990 63800 70020 64800
rect 70180 63800 73210 64800
rect 73370 63800 76400 64800
rect 76560 63800 79590 64800
rect 79750 63800 82780 64800
rect 82940 63800 85970 64800
rect 86130 63800 89160 64800
rect 89320 63800 92350 64800
rect 92510 63800 95540 64800
rect 95700 63800 98730 64800
rect 98890 63800 101920 64800
rect 102080 63800 105110 64800
rect 105270 63800 108300 64800
rect 108460 63800 111490 64800
rect 111650 63800 114680 64800
rect 114840 63800 117870 64800
rect 118030 63800 121060 64800
rect 121220 63800 124250 64800
rect 124410 63800 127440 64800
rect 127600 63800 130630 64800
rect 130790 63800 133820 64800
rect 133980 63800 137010 64800
rect 1000 63640 2000 63800
rect 4190 63640 5190 63800
rect 7380 63640 8380 63800
rect 10570 63640 11570 63800
rect 13760 63640 14760 63800
rect 16950 63640 17950 63800
rect 20140 63640 21140 63800
rect 23330 63640 24330 63800
rect 26520 63640 27520 63800
rect 29710 63640 30710 63800
rect 32900 63640 33900 63800
rect 36090 63640 37090 63800
rect 39280 63640 40280 63800
rect 42470 63640 43470 63800
rect 45660 63640 46660 63800
rect 48850 63640 49850 63800
rect 52040 63640 53040 63800
rect 55230 63640 56230 63800
rect 58420 63640 59420 63800
rect 61610 63640 62610 63800
rect 64800 63640 65800 63800
rect 67990 63640 68990 63800
rect 71180 63640 72180 63800
rect 74370 63640 75370 63800
rect 77560 63640 78560 63800
rect 80750 63640 81750 63800
rect 83940 63640 84940 63800
rect 87130 63640 88130 63800
rect 90320 63640 91320 63800
rect 93510 63640 94510 63800
rect 96700 63640 97700 63800
rect 99890 63640 100890 63800
rect 103080 63640 104080 63800
rect 106270 63640 107270 63800
rect 109460 63640 110460 63800
rect 112650 63640 113650 63800
rect 115840 63640 116840 63800
rect 119030 63640 120030 63800
rect 122220 63640 123220 63800
rect 125410 63640 126410 63800
rect 128600 63640 129600 63800
rect 131790 63640 132790 63800
rect 134980 63640 135980 63800
rect 0 62610 3030 63640
rect 3190 62610 6220 63640
rect 6380 62610 9410 63640
rect 9570 62610 12600 63640
rect 12760 62610 15790 63640
rect 15950 62610 18980 63640
rect 19140 62610 22170 63640
rect 22330 62610 25360 63640
rect 25520 62610 28550 63640
rect 28710 62610 31740 63640
rect 31900 62610 34930 63640
rect 35090 62610 38120 63640
rect 38280 62610 41310 63640
rect 41470 62610 44500 63640
rect 44660 62610 47690 63640
rect 47850 62610 50880 63640
rect 51040 62610 54070 63640
rect 54230 62610 57260 63640
rect 57420 62610 60450 63640
rect 60610 62610 63640 63640
rect 63800 62610 66830 63640
rect 66990 62610 70020 63640
rect 70180 62610 73210 63640
rect 73370 62610 76400 63640
rect 76560 62610 79590 63640
rect 79750 62610 82780 63640
rect 82940 62610 85970 63640
rect 86130 62610 89160 63640
rect 89320 62610 92350 63640
rect 92510 62610 95540 63640
rect 95700 62610 98730 63640
rect 98890 62610 101920 63640
rect 102080 62610 105110 63640
rect 105270 62610 108300 63640
rect 108460 62610 111490 63640
rect 111650 62610 114680 63640
rect 114840 62610 117870 63640
rect 118030 62610 121060 63640
rect 121220 62610 124250 63640
rect 124410 62610 127440 63640
rect 127600 62610 130630 63640
rect 130790 62610 133820 63640
rect 133980 62610 137010 63640
rect 0 61610 137170 62610
rect 0 60610 3030 61610
rect 3190 60610 6220 61610
rect 6380 60610 9410 61610
rect 9570 60610 12600 61610
rect 12760 60610 15790 61610
rect 15950 60610 18980 61610
rect 19140 60610 22170 61610
rect 22330 60610 25360 61610
rect 25520 60610 28550 61610
rect 28710 60610 31740 61610
rect 31900 60610 34930 61610
rect 35090 60610 38120 61610
rect 38280 60610 41310 61610
rect 41470 60610 44500 61610
rect 44660 60610 47690 61610
rect 47850 60610 50880 61610
rect 51040 60610 54070 61610
rect 54230 60610 57260 61610
rect 57420 60610 60450 61610
rect 60610 60610 63640 61610
rect 63800 60610 66830 61610
rect 66990 60610 70020 61610
rect 70180 60610 73210 61610
rect 73370 60610 76400 61610
rect 76560 60610 79590 61610
rect 79750 60610 82780 61610
rect 82940 60610 85970 61610
rect 86130 60610 89160 61610
rect 89320 60610 92350 61610
rect 92510 60610 95540 61610
rect 95700 60610 98730 61610
rect 98890 60610 101920 61610
rect 102080 60610 105110 61610
rect 105270 60610 108300 61610
rect 108460 60610 111490 61610
rect 111650 60610 114680 61610
rect 114840 60610 117870 61610
rect 118030 60610 121060 61610
rect 121220 60610 124250 61610
rect 124410 60610 127440 61610
rect 127600 60610 130630 61610
rect 130790 60610 133820 61610
rect 133980 60610 137010 61610
rect 1000 60450 2000 60610
rect 4190 60450 5190 60610
rect 7380 60450 8380 60610
rect 10570 60450 11570 60610
rect 13760 60450 14760 60610
rect 16950 60450 17950 60610
rect 20140 60450 21140 60610
rect 23330 60450 24330 60610
rect 26520 60450 27520 60610
rect 29710 60450 30710 60610
rect 32900 60450 33900 60610
rect 36090 60450 37090 60610
rect 39280 60450 40280 60610
rect 42470 60450 43470 60610
rect 45660 60450 46660 60610
rect 48850 60450 49850 60610
rect 52040 60450 53040 60610
rect 55230 60450 56230 60610
rect 58420 60450 59420 60610
rect 61610 60450 62610 60610
rect 64800 60450 65800 60610
rect 67990 60450 68990 60610
rect 71180 60450 72180 60610
rect 74370 60450 75370 60610
rect 77560 60450 78560 60610
rect 80750 60450 81750 60610
rect 83940 60450 84940 60610
rect 87130 60450 88130 60610
rect 90320 60450 91320 60610
rect 93510 60450 94510 60610
rect 96700 60450 97700 60610
rect 99890 60450 100890 60610
rect 103080 60450 104080 60610
rect 106270 60450 107270 60610
rect 109460 60450 110460 60610
rect 112650 60450 113650 60610
rect 115840 60450 116840 60610
rect 119030 60450 120030 60610
rect 122220 60450 123220 60610
rect 125410 60450 126410 60610
rect 128600 60450 129600 60610
rect 131790 60450 132790 60610
rect 134980 60450 135980 60610
rect 0 59420 3030 60450
rect 3190 59420 6220 60450
rect 6380 59420 9410 60450
rect 9570 59420 12600 60450
rect 12760 59420 15790 60450
rect 15950 59420 18980 60450
rect 19140 59420 22170 60450
rect 22330 59420 25360 60450
rect 25520 59420 28550 60450
rect 28710 59420 31740 60450
rect 31900 59420 34930 60450
rect 35090 59420 38120 60450
rect 38280 59420 41310 60450
rect 41470 59420 44500 60450
rect 44660 59420 47690 60450
rect 47850 59420 50880 60450
rect 51040 59420 54070 60450
rect 54230 59420 57260 60450
rect 57420 59420 60450 60450
rect 60610 59420 63640 60450
rect 63800 59420 66830 60450
rect 66990 59420 70020 60450
rect 70180 59420 73210 60450
rect 73370 59420 76400 60450
rect 76560 59420 79590 60450
rect 79750 59420 82780 60450
rect 82940 59420 85970 60450
rect 86130 59420 89160 60450
rect 89320 59420 92350 60450
rect 92510 59420 95540 60450
rect 95700 59420 98730 60450
rect 98890 59420 101920 60450
rect 102080 59420 105110 60450
rect 105270 59420 108300 60450
rect 108460 59420 111490 60450
rect 111650 59420 114680 60450
rect 114840 59420 117870 60450
rect 118030 59420 121060 60450
rect 121220 59420 124250 60450
rect 124410 59420 127440 60450
rect 127600 59420 130630 60450
rect 130790 59420 133820 60450
rect 133980 59420 137010 60450
rect 0 58420 137170 59420
rect 0 57420 3030 58420
rect 3190 57420 6220 58420
rect 6380 57420 9410 58420
rect 9570 57420 12600 58420
rect 12760 57420 15790 58420
rect 15950 57420 18980 58420
rect 19140 57420 22170 58420
rect 22330 57420 25360 58420
rect 25520 57420 28550 58420
rect 28710 57420 31740 58420
rect 31900 57420 34930 58420
rect 35090 57420 38120 58420
rect 38280 57420 41310 58420
rect 41470 57420 44500 58420
rect 44660 57420 47690 58420
rect 47850 57420 50880 58420
rect 51040 57420 54070 58420
rect 54230 57420 57260 58420
rect 57420 57420 60450 58420
rect 60610 57420 63640 58420
rect 63800 57420 66830 58420
rect 66990 57420 70020 58420
rect 70180 57420 73210 58420
rect 73370 57420 76400 58420
rect 76560 57420 79590 58420
rect 79750 57420 82780 58420
rect 82940 57420 85970 58420
rect 86130 57420 89160 58420
rect 89320 57420 92350 58420
rect 92510 57420 95540 58420
rect 95700 57420 98730 58420
rect 98890 57420 101920 58420
rect 102080 57420 105110 58420
rect 105270 57420 108300 58420
rect 108460 57420 111490 58420
rect 111650 57420 114680 58420
rect 114840 57420 117870 58420
rect 118030 57420 121060 58420
rect 121220 57420 124250 58420
rect 124410 57420 127440 58420
rect 127600 57420 130630 58420
rect 130790 57420 133820 58420
rect 133980 57420 137010 58420
rect 1000 57260 2000 57420
rect 4190 57260 5190 57420
rect 7380 57260 8380 57420
rect 10570 57260 11570 57420
rect 13760 57260 14760 57420
rect 16950 57260 17950 57420
rect 20140 57260 21140 57420
rect 23330 57260 24330 57420
rect 26520 57260 27520 57420
rect 29710 57260 30710 57420
rect 32900 57260 33900 57420
rect 36090 57260 37090 57420
rect 39280 57260 40280 57420
rect 42470 57260 43470 57420
rect 45660 57260 46660 57420
rect 48850 57260 49850 57420
rect 52040 57260 53040 57420
rect 55230 57260 56230 57420
rect 58420 57260 59420 57420
rect 61610 57260 62610 57420
rect 64800 57260 65800 57420
rect 67990 57260 68990 57420
rect 71180 57260 72180 57420
rect 74370 57260 75370 57420
rect 77560 57260 78560 57420
rect 80750 57260 81750 57420
rect 83940 57260 84940 57420
rect 87130 57260 88130 57420
rect 90320 57260 91320 57420
rect 93510 57260 94510 57420
rect 96700 57260 97700 57420
rect 99890 57260 100890 57420
rect 103080 57260 104080 57420
rect 106270 57260 107270 57420
rect 109460 57260 110460 57420
rect 112650 57260 113650 57420
rect 115840 57260 116840 57420
rect 119030 57260 120030 57420
rect 122220 57260 123220 57420
rect 125410 57260 126410 57420
rect 128600 57260 129600 57420
rect 131790 57260 132790 57420
rect 134980 57260 135980 57420
rect 0 56230 3030 57260
rect 3190 56230 6220 57260
rect 6380 56230 9410 57260
rect 9570 56230 12600 57260
rect 12760 56230 15790 57260
rect 15950 56230 18980 57260
rect 19140 56230 22170 57260
rect 22330 56230 25360 57260
rect 25520 56230 28550 57260
rect 28710 56230 31740 57260
rect 31900 56230 34930 57260
rect 35090 56230 38120 57260
rect 38280 56230 41310 57260
rect 41470 56230 44500 57260
rect 44660 56230 47690 57260
rect 47850 56230 50880 57260
rect 51040 56230 54070 57260
rect 54230 56230 57260 57260
rect 57420 56230 60450 57260
rect 60610 56230 63640 57260
rect 63800 56230 66830 57260
rect 66990 56230 70020 57260
rect 70180 56230 73210 57260
rect 73370 56230 76400 57260
rect 76560 56230 79590 57260
rect 79750 56230 82780 57260
rect 82940 56230 85970 57260
rect 86130 56230 89160 57260
rect 89320 56230 92350 57260
rect 92510 56230 95540 57260
rect 95700 56230 98730 57260
rect 98890 56230 101920 57260
rect 102080 56230 105110 57260
rect 105270 56230 108300 57260
rect 108460 56230 111490 57260
rect 111650 56230 114680 57260
rect 114840 56230 117870 57260
rect 118030 56230 121060 57260
rect 121220 56230 124250 57260
rect 124410 56230 127440 57260
rect 127600 56230 130630 57260
rect 130790 56230 133820 57260
rect 133980 56230 137010 57260
rect 0 55230 137170 56230
rect 0 54230 3030 55230
rect 3190 54230 6220 55230
rect 6380 54230 9410 55230
rect 9570 54230 12600 55230
rect 12760 54230 15790 55230
rect 15950 54230 18980 55230
rect 19140 54230 22170 55230
rect 22330 54230 25360 55230
rect 25520 54230 28550 55230
rect 28710 54230 31740 55230
rect 31900 54230 34930 55230
rect 35090 54230 38120 55230
rect 38280 54230 41310 55230
rect 41470 54230 44500 55230
rect 44660 54230 47690 55230
rect 47850 54230 50880 55230
rect 51040 54230 54070 55230
rect 54230 54230 57260 55230
rect 57420 54230 60450 55230
rect 60610 54230 63640 55230
rect 63800 54230 66830 55230
rect 66990 54230 70020 55230
rect 70180 54230 73210 55230
rect 73370 54230 76400 55230
rect 76560 54230 79590 55230
rect 79750 54230 82780 55230
rect 82940 54230 85970 55230
rect 86130 54230 89160 55230
rect 89320 54230 92350 55230
rect 92510 54230 95540 55230
rect 95700 54230 98730 55230
rect 98890 54230 101920 55230
rect 102080 54230 105110 55230
rect 105270 54230 108300 55230
rect 108460 54230 111490 55230
rect 111650 54230 114680 55230
rect 114840 54230 117870 55230
rect 118030 54230 121060 55230
rect 121220 54230 124250 55230
rect 124410 54230 127440 55230
rect 127600 54230 130630 55230
rect 130790 54230 133820 55230
rect 133980 54230 137010 55230
rect 1000 54070 2000 54230
rect 4190 54070 5190 54230
rect 7380 54070 8380 54230
rect 10570 54070 11570 54230
rect 13760 54070 14760 54230
rect 16950 54070 17950 54230
rect 20140 54070 21140 54230
rect 23330 54070 24330 54230
rect 26520 54070 27520 54230
rect 29710 54070 30710 54230
rect 32900 54070 33900 54230
rect 36090 54070 37090 54230
rect 39280 54070 40280 54230
rect 42470 54070 43470 54230
rect 45660 54070 46660 54230
rect 48850 54070 49850 54230
rect 52040 54070 53040 54230
rect 55230 54070 56230 54230
rect 58420 54070 59420 54230
rect 61610 54070 62610 54230
rect 64800 54070 65800 54230
rect 67990 54070 68990 54230
rect 71180 54070 72180 54230
rect 74370 54070 75370 54230
rect 77560 54070 78560 54230
rect 80750 54070 81750 54230
rect 83940 54070 84940 54230
rect 87130 54070 88130 54230
rect 90320 54070 91320 54230
rect 93510 54070 94510 54230
rect 96700 54070 97700 54230
rect 99890 54070 100890 54230
rect 103080 54070 104080 54230
rect 106270 54070 107270 54230
rect 109460 54070 110460 54230
rect 112650 54070 113650 54230
rect 115840 54070 116840 54230
rect 119030 54070 120030 54230
rect 122220 54070 123220 54230
rect 125410 54070 126410 54230
rect 128600 54070 129600 54230
rect 131790 54070 132790 54230
rect 134980 54070 135980 54230
rect 0 53040 3030 54070
rect 3190 53040 6220 54070
rect 6380 53040 9410 54070
rect 9570 53040 12600 54070
rect 12760 53040 15790 54070
rect 15950 53040 18980 54070
rect 19140 53040 22170 54070
rect 22330 53040 25360 54070
rect 25520 53040 28550 54070
rect 28710 53040 31740 54070
rect 31900 53040 34930 54070
rect 35090 53040 38120 54070
rect 38280 53040 41310 54070
rect 41470 53040 44500 54070
rect 44660 53040 47690 54070
rect 47850 53040 50880 54070
rect 51040 53040 54070 54070
rect 54230 53040 57260 54070
rect 57420 53040 60450 54070
rect 60610 53040 63640 54070
rect 63800 53040 66830 54070
rect 66990 53040 70020 54070
rect 70180 53040 73210 54070
rect 73370 53040 76400 54070
rect 76560 53040 79590 54070
rect 79750 53040 82780 54070
rect 82940 53040 85970 54070
rect 86130 53040 89160 54070
rect 89320 53040 92350 54070
rect 92510 53040 95540 54070
rect 95700 53040 98730 54070
rect 98890 53040 101920 54070
rect 102080 53040 105110 54070
rect 105270 53040 108300 54070
rect 108460 53040 111490 54070
rect 111650 53040 114680 54070
rect 114840 53040 117870 54070
rect 118030 53040 121060 54070
rect 121220 53040 124250 54070
rect 124410 53040 127440 54070
rect 127600 53040 130630 54070
rect 130790 53040 133820 54070
rect 133980 53040 137010 54070
rect 0 52040 137170 53040
rect 0 51040 3030 52040
rect 3190 51040 6220 52040
rect 6380 51040 9410 52040
rect 9570 51040 12600 52040
rect 12760 51040 15790 52040
rect 15950 51040 18980 52040
rect 19140 51040 22170 52040
rect 22330 51040 25360 52040
rect 25520 51040 28550 52040
rect 28710 51040 31740 52040
rect 31900 51040 34930 52040
rect 35090 51040 38120 52040
rect 38280 51040 41310 52040
rect 41470 51040 44500 52040
rect 44660 51040 47690 52040
rect 47850 51040 50880 52040
rect 51040 51040 54070 52040
rect 54230 51040 57260 52040
rect 57420 51040 60450 52040
rect 60610 51040 63640 52040
rect 63800 51040 66830 52040
rect 66990 51040 70020 52040
rect 70180 51040 73210 52040
rect 73370 51040 76400 52040
rect 76560 51040 79590 52040
rect 79750 51040 82780 52040
rect 82940 51040 85970 52040
rect 86130 51040 89160 52040
rect 89320 51040 92350 52040
rect 92510 51040 95540 52040
rect 95700 51040 98730 52040
rect 98890 51040 101920 52040
rect 102080 51040 105110 52040
rect 105270 51040 108300 52040
rect 108460 51040 111490 52040
rect 111650 51040 114680 52040
rect 114840 51040 117870 52040
rect 118030 51040 121060 52040
rect 121220 51040 124250 52040
rect 124410 51040 127440 52040
rect 127600 51040 130630 52040
rect 130790 51040 133820 52040
rect 133980 51040 137010 52040
rect 1000 50880 2000 51040
rect 4190 50880 5190 51040
rect 7380 50880 8380 51040
rect 10570 50880 11570 51040
rect 13760 50880 14760 51040
rect 16950 50880 17950 51040
rect 20140 50880 21140 51040
rect 23330 50880 24330 51040
rect 26520 50880 27520 51040
rect 29710 50880 30710 51040
rect 32900 50880 33900 51040
rect 36090 50880 37090 51040
rect 39280 50880 40280 51040
rect 42470 50880 43470 51040
rect 45660 50880 46660 51040
rect 48850 50880 49850 51040
rect 52040 50880 53040 51040
rect 55230 50880 56230 51040
rect 58420 50880 59420 51040
rect 61610 50880 62610 51040
rect 64800 50880 65800 51040
rect 67990 50880 68990 51040
rect 71180 50880 72180 51040
rect 74370 50880 75370 51040
rect 77560 50880 78560 51040
rect 80750 50880 81750 51040
rect 83940 50880 84940 51040
rect 87130 50880 88130 51040
rect 90320 50880 91320 51040
rect 93510 50880 94510 51040
rect 96700 50880 97700 51040
rect 99890 50880 100890 51040
rect 103080 50880 104080 51040
rect 106270 50880 107270 51040
rect 109460 50880 110460 51040
rect 112650 50880 113650 51040
rect 115840 50880 116840 51040
rect 119030 50880 120030 51040
rect 122220 50880 123220 51040
rect 125410 50880 126410 51040
rect 128600 50880 129600 51040
rect 131790 50880 132790 51040
rect 134980 50880 135980 51040
rect 0 49850 3030 50880
rect 3190 49850 6220 50880
rect 6380 49850 9410 50880
rect 9570 49850 12600 50880
rect 12760 49850 15790 50880
rect 15950 49850 18980 50880
rect 19140 49850 22170 50880
rect 22330 49850 25360 50880
rect 25520 49850 28550 50880
rect 28710 49850 31740 50880
rect 31900 49850 34930 50880
rect 35090 49850 38120 50880
rect 38280 49850 41310 50880
rect 41470 49850 44500 50880
rect 44660 49850 47690 50880
rect 47850 49850 50880 50880
rect 51040 49850 54070 50880
rect 54230 49850 57260 50880
rect 57420 49850 60450 50880
rect 60610 49850 63640 50880
rect 63800 49850 66830 50880
rect 66990 49850 70020 50880
rect 70180 49850 73210 50880
rect 73370 49850 76400 50880
rect 76560 49850 79590 50880
rect 79750 49850 82780 50880
rect 82940 49850 85970 50880
rect 86130 49850 89160 50880
rect 89320 49850 92350 50880
rect 92510 49850 95540 50880
rect 95700 49850 98730 50880
rect 98890 49850 101920 50880
rect 102080 49850 105110 50880
rect 105270 49850 108300 50880
rect 108460 49850 111490 50880
rect 111650 49850 114680 50880
rect 114840 49850 117870 50880
rect 118030 49850 121060 50880
rect 121220 49850 124250 50880
rect 124410 49850 127440 50880
rect 127600 49850 130630 50880
rect 130790 49850 133820 50880
rect 133980 49850 137010 50880
rect 0 48850 137170 49850
rect 0 47850 3030 48850
rect 3190 47850 6220 48850
rect 6380 47850 9410 48850
rect 9570 47850 12600 48850
rect 12760 47850 15790 48850
rect 15950 47850 18980 48850
rect 19140 47850 22170 48850
rect 22330 47850 25360 48850
rect 25520 47850 28550 48850
rect 28710 47850 31740 48850
rect 31900 47850 34930 48850
rect 35090 47850 38120 48850
rect 38280 47850 41310 48850
rect 41470 47850 44500 48850
rect 44660 47850 47690 48850
rect 47850 47850 50880 48850
rect 51040 47850 54070 48850
rect 54230 47850 57260 48850
rect 57420 47850 60450 48850
rect 60610 47850 63640 48850
rect 63800 47850 66830 48850
rect 66990 47850 70020 48850
rect 70180 47850 73210 48850
rect 73370 47850 76400 48850
rect 76560 47850 79590 48850
rect 79750 47850 82780 48850
rect 82940 47850 85970 48850
rect 86130 47850 89160 48850
rect 89320 47850 92350 48850
rect 92510 47850 95540 48850
rect 95700 47850 98730 48850
rect 98890 47850 101920 48850
rect 102080 47850 105110 48850
rect 105270 47850 108300 48850
rect 108460 47850 111490 48850
rect 111650 47850 114680 48850
rect 114840 47850 117870 48850
rect 118030 47850 121060 48850
rect 121220 47850 124250 48850
rect 124410 47850 127440 48850
rect 127600 47850 130630 48850
rect 130790 47850 133820 48850
rect 133980 47850 137010 48850
rect 1000 47690 2000 47850
rect 4190 47690 5190 47850
rect 7380 47690 8380 47850
rect 10570 47690 11570 47850
rect 13760 47690 14760 47850
rect 16950 47690 17950 47850
rect 20140 47690 21140 47850
rect 23330 47690 24330 47850
rect 26520 47690 27520 47850
rect 29710 47690 30710 47850
rect 32900 47690 33900 47850
rect 36090 47690 37090 47850
rect 39280 47690 40280 47850
rect 42470 47690 43470 47850
rect 45660 47690 46660 47850
rect 48850 47690 49850 47850
rect 52040 47690 53040 47850
rect 55230 47690 56230 47850
rect 58420 47690 59420 47850
rect 61610 47690 62610 47850
rect 64800 47690 65800 47850
rect 67990 47690 68990 47850
rect 71180 47690 72180 47850
rect 74370 47690 75370 47850
rect 77560 47690 78560 47850
rect 80750 47690 81750 47850
rect 83940 47690 84940 47850
rect 87130 47690 88130 47850
rect 90320 47690 91320 47850
rect 93510 47690 94510 47850
rect 96700 47690 97700 47850
rect 99890 47690 100890 47850
rect 103080 47690 104080 47850
rect 106270 47690 107270 47850
rect 109460 47690 110460 47850
rect 112650 47690 113650 47850
rect 115840 47690 116840 47850
rect 119030 47690 120030 47850
rect 122220 47690 123220 47850
rect 125410 47690 126410 47850
rect 128600 47690 129600 47850
rect 131790 47690 132790 47850
rect 134980 47690 135980 47850
rect 0 46660 3030 47690
rect 3190 46660 6220 47690
rect 6380 46660 9410 47690
rect 9570 46660 12600 47690
rect 12760 46660 15790 47690
rect 15950 46660 18980 47690
rect 19140 46660 22170 47690
rect 22330 46660 25360 47690
rect 25520 46660 28550 47690
rect 28710 46660 31740 47690
rect 31900 46660 34930 47690
rect 35090 46660 38120 47690
rect 38280 46660 41310 47690
rect 41470 46660 44500 47690
rect 44660 46660 47690 47690
rect 47850 46660 50880 47690
rect 51040 46660 54070 47690
rect 54230 46660 57260 47690
rect 57420 46660 60450 47690
rect 60610 46660 63640 47690
rect 63800 46660 66830 47690
rect 66990 46660 70020 47690
rect 70180 46660 73210 47690
rect 73370 46660 76400 47690
rect 76560 46660 79590 47690
rect 79750 46660 82780 47690
rect 82940 46660 85970 47690
rect 86130 46660 89160 47690
rect 89320 46660 92350 47690
rect 92510 46660 95540 47690
rect 95700 46660 98730 47690
rect 98890 46660 101920 47690
rect 102080 46660 105110 47690
rect 105270 46660 108300 47690
rect 108460 46660 111490 47690
rect 111650 46660 114680 47690
rect 114840 46660 117870 47690
rect 118030 46660 121060 47690
rect 121220 46660 124250 47690
rect 124410 46660 127440 47690
rect 127600 46660 130630 47690
rect 130790 46660 133820 47690
rect 133980 46660 137010 47690
rect 0 45660 137170 46660
rect 0 44660 3030 45660
rect 3190 44660 6220 45660
rect 6380 44660 9410 45660
rect 9570 44660 12600 45660
rect 12760 44660 15790 45660
rect 15950 44660 18980 45660
rect 19140 44660 22170 45660
rect 22330 44660 25360 45660
rect 25520 44660 28550 45660
rect 28710 44660 31740 45660
rect 31900 44660 34930 45660
rect 35090 44660 38120 45660
rect 38280 44660 41310 45660
rect 41470 44660 44500 45660
rect 44660 44660 47690 45660
rect 47850 44660 50880 45660
rect 51040 44660 54070 45660
rect 54230 44660 57260 45660
rect 57420 44660 60450 45660
rect 60610 44660 63640 45660
rect 63800 44660 66830 45660
rect 66990 44660 70020 45660
rect 70180 44660 73210 45660
rect 73370 44660 76400 45660
rect 76560 44660 79590 45660
rect 79750 44660 82780 45660
rect 82940 44660 85970 45660
rect 86130 44660 89160 45660
rect 89320 44660 92350 45660
rect 92510 44660 95540 45660
rect 95700 44660 98730 45660
rect 98890 44660 101920 45660
rect 102080 44660 105110 45660
rect 105270 44660 108300 45660
rect 108460 44660 111490 45660
rect 111650 44660 114680 45660
rect 114840 44660 117870 45660
rect 118030 44660 121060 45660
rect 121220 44660 124250 45660
rect 124410 44660 127440 45660
rect 127600 44660 130630 45660
rect 130790 44660 133820 45660
rect 133980 44660 137010 45660
rect 1000 44500 2000 44660
rect 4190 44500 5190 44660
rect 7380 44500 8380 44660
rect 10570 44500 11570 44660
rect 13760 44500 14760 44660
rect 16950 44500 17950 44660
rect 20140 44500 21140 44660
rect 23330 44500 24330 44660
rect 26520 44500 27520 44660
rect 29710 44500 30710 44660
rect 32900 44500 33900 44660
rect 36090 44500 37090 44660
rect 39280 44500 40280 44660
rect 42470 44500 43470 44660
rect 45660 44500 46660 44660
rect 48850 44500 49850 44660
rect 52040 44500 53040 44660
rect 55230 44500 56230 44660
rect 58420 44500 59420 44660
rect 61610 44500 62610 44660
rect 64800 44500 65800 44660
rect 67990 44500 68990 44660
rect 71180 44500 72180 44660
rect 74370 44500 75370 44660
rect 77560 44500 78560 44660
rect 80750 44500 81750 44660
rect 83940 44500 84940 44660
rect 87130 44500 88130 44660
rect 90320 44500 91320 44660
rect 93510 44500 94510 44660
rect 96700 44500 97700 44660
rect 99890 44500 100890 44660
rect 103080 44500 104080 44660
rect 106270 44500 107270 44660
rect 109460 44500 110460 44660
rect 112650 44500 113650 44660
rect 115840 44500 116840 44660
rect 119030 44500 120030 44660
rect 122220 44500 123220 44660
rect 125410 44500 126410 44660
rect 128600 44500 129600 44660
rect 131790 44500 132790 44660
rect 134980 44500 135980 44660
rect 0 43470 3030 44500
rect 3190 43470 6220 44500
rect 6380 43470 9410 44500
rect 9570 43470 12600 44500
rect 12760 43470 15790 44500
rect 15950 43470 18980 44500
rect 19140 43470 22170 44500
rect 22330 43470 25360 44500
rect 25520 43470 28550 44500
rect 28710 43470 31740 44500
rect 31900 43470 34930 44500
rect 35090 43470 38120 44500
rect 38280 43470 41310 44500
rect 41470 43470 44500 44500
rect 44660 43470 47690 44500
rect 47850 43470 50880 44500
rect 51040 43470 54070 44500
rect 54230 43470 57260 44500
rect 57420 43470 60450 44500
rect 60610 43470 63640 44500
rect 63800 43470 66830 44500
rect 66990 43470 70020 44500
rect 70180 43470 73210 44500
rect 73370 43470 76400 44500
rect 76560 43470 79590 44500
rect 79750 43470 82780 44500
rect 82940 43470 85970 44500
rect 86130 43470 89160 44500
rect 89320 43470 92350 44500
rect 92510 43470 95540 44500
rect 95700 43470 98730 44500
rect 98890 43470 101920 44500
rect 102080 43470 105110 44500
rect 105270 43470 108300 44500
rect 108460 43470 111490 44500
rect 111650 43470 114680 44500
rect 114840 43470 117870 44500
rect 118030 43470 121060 44500
rect 121220 43470 124250 44500
rect 124410 43470 127440 44500
rect 127600 43470 130630 44500
rect 130790 43470 133820 44500
rect 133980 43470 137010 44500
rect 0 42470 137170 43470
rect 0 41470 3030 42470
rect 3190 41470 6220 42470
rect 6380 41470 9410 42470
rect 9570 41470 12600 42470
rect 12760 41470 15790 42470
rect 15950 41470 18980 42470
rect 19140 41470 22170 42470
rect 22330 41470 25360 42470
rect 25520 41470 28550 42470
rect 28710 41470 31740 42470
rect 31900 41470 34930 42470
rect 35090 41470 38120 42470
rect 38280 41470 41310 42470
rect 41470 41470 44500 42470
rect 44660 41470 47690 42470
rect 47850 41470 50880 42470
rect 51040 41470 54070 42470
rect 54230 41470 57260 42470
rect 57420 41470 60450 42470
rect 60610 41470 63640 42470
rect 63800 41470 66830 42470
rect 66990 41470 70020 42470
rect 70180 41470 73210 42470
rect 73370 41470 76400 42470
rect 76560 41470 79590 42470
rect 79750 41470 82780 42470
rect 82940 41470 85970 42470
rect 86130 41470 89160 42470
rect 89320 41470 92350 42470
rect 92510 41470 95540 42470
rect 95700 41470 98730 42470
rect 98890 41470 101920 42470
rect 102080 41470 105110 42470
rect 105270 41470 108300 42470
rect 108460 41470 111490 42470
rect 111650 41470 114680 42470
rect 114840 41470 117870 42470
rect 118030 41470 121060 42470
rect 121220 41470 124250 42470
rect 124410 41470 127440 42470
rect 127600 41470 130630 42470
rect 130790 41470 133820 42470
rect 133980 41470 137010 42470
rect 1000 41310 2000 41470
rect 4190 41310 5190 41470
rect 7380 41310 8380 41470
rect 10570 41310 11570 41470
rect 13760 41310 14760 41470
rect 16950 41310 17950 41470
rect 20140 41310 21140 41470
rect 23330 41310 24330 41470
rect 26520 41310 27520 41470
rect 29710 41310 30710 41470
rect 32900 41310 33900 41470
rect 36090 41310 37090 41470
rect 39280 41310 40280 41470
rect 42470 41310 43470 41470
rect 45660 41310 46660 41470
rect 48850 41310 49850 41470
rect 52040 41310 53040 41470
rect 55230 41310 56230 41470
rect 58420 41310 59420 41470
rect 61610 41310 62610 41470
rect 64800 41310 65800 41470
rect 67990 41310 68990 41470
rect 71180 41310 72180 41470
rect 74370 41310 75370 41470
rect 77560 41310 78560 41470
rect 80750 41310 81750 41470
rect 83940 41310 84940 41470
rect 87130 41310 88130 41470
rect 90320 41310 91320 41470
rect 93510 41310 94510 41470
rect 96700 41310 97700 41470
rect 99890 41310 100890 41470
rect 103080 41310 104080 41470
rect 106270 41310 107270 41470
rect 109460 41310 110460 41470
rect 112650 41310 113650 41470
rect 115840 41310 116840 41470
rect 119030 41310 120030 41470
rect 122220 41310 123220 41470
rect 125410 41310 126410 41470
rect 128600 41310 129600 41470
rect 131790 41310 132790 41470
rect 134980 41310 135980 41470
rect 0 40280 3030 41310
rect 3190 40280 6220 41310
rect 6380 40280 9410 41310
rect 9570 40280 12600 41310
rect 12760 40280 15790 41310
rect 15950 40280 18980 41310
rect 19140 40280 22170 41310
rect 22330 40280 25360 41310
rect 25520 40280 28550 41310
rect 28710 40280 31740 41310
rect 31900 40280 34930 41310
rect 35090 40280 38120 41310
rect 38280 40280 41310 41310
rect 41470 40280 44500 41310
rect 44660 40280 47690 41310
rect 47850 40280 50880 41310
rect 51040 40280 54070 41310
rect 54230 40280 57260 41310
rect 57420 40280 60450 41310
rect 60610 40280 63640 41310
rect 63800 40280 66830 41310
rect 66990 40280 70020 41310
rect 70180 40280 73210 41310
rect 73370 40280 76400 41310
rect 76560 40280 79590 41310
rect 79750 40280 82780 41310
rect 82940 40280 85970 41310
rect 86130 40280 89160 41310
rect 89320 40280 92350 41310
rect 92510 40280 95540 41310
rect 95700 40280 98730 41310
rect 98890 40280 101920 41310
rect 102080 40280 105110 41310
rect 105270 40280 108300 41310
rect 108460 40280 111490 41310
rect 111650 40280 114680 41310
rect 114840 40280 117870 41310
rect 118030 40280 121060 41310
rect 121220 40280 124250 41310
rect 124410 40280 127440 41310
rect 127600 40280 130630 41310
rect 130790 40280 133820 41310
rect 133980 40280 137010 41310
rect 0 39280 137170 40280
rect 0 38280 3030 39280
rect 3190 38280 6220 39280
rect 6380 38280 9410 39280
rect 9570 38280 12600 39280
rect 12760 38280 15790 39280
rect 15950 38280 18980 39280
rect 19140 38280 22170 39280
rect 22330 38280 25360 39280
rect 25520 38280 28550 39280
rect 28710 38280 31740 39280
rect 31900 38280 34930 39280
rect 35090 38280 38120 39280
rect 38280 38280 41310 39280
rect 41470 38280 44500 39280
rect 44660 38280 47690 39280
rect 47850 38280 50880 39280
rect 51040 38280 54070 39280
rect 54230 38280 57260 39280
rect 57420 38280 60450 39280
rect 60610 38280 63640 39280
rect 63800 38280 66830 39280
rect 66990 38280 70020 39280
rect 70180 38280 73210 39280
rect 73370 38280 76400 39280
rect 76560 38280 79590 39280
rect 79750 38280 82780 39280
rect 82940 38280 85970 39280
rect 86130 38280 89160 39280
rect 89320 38280 92350 39280
rect 92510 38280 95540 39280
rect 95700 38280 98730 39280
rect 98890 38280 101920 39280
rect 102080 38280 105110 39280
rect 105270 38280 108300 39280
rect 108460 38280 111490 39280
rect 111650 38280 114680 39280
rect 114840 38280 117870 39280
rect 118030 38280 121060 39280
rect 121220 38280 124250 39280
rect 124410 38280 127440 39280
rect 127600 38280 130630 39280
rect 130790 38280 133820 39280
rect 133980 38280 137010 39280
rect 1000 38120 2000 38280
rect 4190 38120 5190 38280
rect 7380 38120 8380 38280
rect 10570 38120 11570 38280
rect 13760 38120 14760 38280
rect 16950 38120 17950 38280
rect 20140 38120 21140 38280
rect 23330 38120 24330 38280
rect 26520 38120 27520 38280
rect 29710 38120 30710 38280
rect 32900 38120 33900 38280
rect 36090 38120 37090 38280
rect 39280 38120 40280 38280
rect 42470 38120 43470 38280
rect 45660 38120 46660 38280
rect 48850 38120 49850 38280
rect 52040 38120 53040 38280
rect 55230 38120 56230 38280
rect 58420 38120 59420 38280
rect 61610 38120 62610 38280
rect 64800 38120 65800 38280
rect 67990 38120 68990 38280
rect 71180 38120 72180 38280
rect 74370 38120 75370 38280
rect 77560 38120 78560 38280
rect 80750 38120 81750 38280
rect 83940 38120 84940 38280
rect 87130 38120 88130 38280
rect 90320 38120 91320 38280
rect 93510 38120 94510 38280
rect 96700 38120 97700 38280
rect 99890 38120 100890 38280
rect 103080 38120 104080 38280
rect 106270 38120 107270 38280
rect 109460 38120 110460 38280
rect 112650 38120 113650 38280
rect 115840 38120 116840 38280
rect 119030 38120 120030 38280
rect 122220 38120 123220 38280
rect 125410 38120 126410 38280
rect 128600 38120 129600 38280
rect 131790 38120 132790 38280
rect 134980 38120 135980 38280
rect 0 37090 3030 38120
rect 3190 37090 6220 38120
rect 6380 37090 9410 38120
rect 9570 37090 12600 38120
rect 12760 37090 15790 38120
rect 15950 37090 18980 38120
rect 19140 37090 22170 38120
rect 22330 37090 25360 38120
rect 25520 37090 28550 38120
rect 28710 37090 31740 38120
rect 31900 37090 34930 38120
rect 35090 37090 38120 38120
rect 38280 37090 41310 38120
rect 41470 37090 44500 38120
rect 44660 37090 47690 38120
rect 47850 37090 50880 38120
rect 51040 37090 54070 38120
rect 54230 37090 57260 38120
rect 57420 37090 60450 38120
rect 60610 37090 63640 38120
rect 63800 37090 66830 38120
rect 66990 37090 70020 38120
rect 70180 37090 73210 38120
rect 73370 37090 76400 38120
rect 76560 37090 79590 38120
rect 79750 37090 82780 38120
rect 82940 37090 85970 38120
rect 86130 37090 89160 38120
rect 89320 37090 92350 38120
rect 92510 37090 95540 38120
rect 95700 37090 98730 38120
rect 98890 37090 101920 38120
rect 102080 37090 105110 38120
rect 105270 37090 108300 38120
rect 108460 37090 111490 38120
rect 111650 37090 114680 38120
rect 114840 37090 117870 38120
rect 118030 37090 121060 38120
rect 121220 37090 124250 38120
rect 124410 37090 127440 38120
rect 127600 37090 130630 38120
rect 130790 37090 133820 38120
rect 133980 37090 137010 38120
rect 0 36090 137170 37090
rect 0 35090 3030 36090
rect 3190 35090 6220 36090
rect 6380 35090 9410 36090
rect 9570 35090 12600 36090
rect 12760 35090 15790 36090
rect 15950 35090 18980 36090
rect 19140 35090 22170 36090
rect 22330 35090 25360 36090
rect 25520 35090 28550 36090
rect 28710 35090 31740 36090
rect 31900 35090 34930 36090
rect 35090 35090 38120 36090
rect 38280 35090 41310 36090
rect 41470 35090 44500 36090
rect 44660 35090 47690 36090
rect 47850 35090 50880 36090
rect 51040 35090 54070 36090
rect 54230 35090 57260 36090
rect 57420 35090 60450 36090
rect 60610 35090 63640 36090
rect 63800 35090 66830 36090
rect 66990 35090 70020 36090
rect 70180 35090 73210 36090
rect 73370 35090 76400 36090
rect 76560 35090 79590 36090
rect 79750 35090 82780 36090
rect 82940 35090 85970 36090
rect 86130 35090 89160 36090
rect 89320 35090 92350 36090
rect 92510 35090 95540 36090
rect 95700 35090 98730 36090
rect 98890 35090 101920 36090
rect 102080 35090 105110 36090
rect 105270 35090 108300 36090
rect 108460 35090 111490 36090
rect 111650 35090 114680 36090
rect 114840 35090 117870 36090
rect 118030 35090 121060 36090
rect 121220 35090 124250 36090
rect 124410 35090 127440 36090
rect 127600 35090 130630 36090
rect 130790 35090 133820 36090
rect 133980 35090 137010 36090
rect 1000 34930 2000 35090
rect 4190 34930 5190 35090
rect 7380 34930 8380 35090
rect 10570 34930 11570 35090
rect 13760 34930 14760 35090
rect 16950 34930 17950 35090
rect 20140 34930 21140 35090
rect 23330 34930 24330 35090
rect 26520 34930 27520 35090
rect 29710 34930 30710 35090
rect 32900 34930 33900 35090
rect 36090 34930 37090 35090
rect 39280 34930 40280 35090
rect 42470 34930 43470 35090
rect 45660 34930 46660 35090
rect 48850 34930 49850 35090
rect 52040 34930 53040 35090
rect 55230 34930 56230 35090
rect 58420 34930 59420 35090
rect 61610 34930 62610 35090
rect 64800 34930 65800 35090
rect 67990 34930 68990 35090
rect 71180 34930 72180 35090
rect 74370 34930 75370 35090
rect 77560 34930 78560 35090
rect 80750 34930 81750 35090
rect 83940 34930 84940 35090
rect 87130 34930 88130 35090
rect 90320 34930 91320 35090
rect 93510 34930 94510 35090
rect 96700 34930 97700 35090
rect 99890 34930 100890 35090
rect 103080 34930 104080 35090
rect 106270 34930 107270 35090
rect 109460 34930 110460 35090
rect 112650 34930 113650 35090
rect 115840 34930 116840 35090
rect 119030 34930 120030 35090
rect 122220 34930 123220 35090
rect 125410 34930 126410 35090
rect 128600 34930 129600 35090
rect 131790 34930 132790 35090
rect 134980 34930 135980 35090
rect 0 33900 3030 34930
rect 3190 33900 6220 34930
rect 6380 33900 9410 34930
rect 9570 33900 12600 34930
rect 12760 33900 15790 34930
rect 15950 33900 18980 34930
rect 19140 33900 22170 34930
rect 22330 33900 25360 34930
rect 25520 33900 28550 34930
rect 28710 33900 31740 34930
rect 31900 33900 34930 34930
rect 35090 33900 38120 34930
rect 38280 33900 41310 34930
rect 41470 33900 44500 34930
rect 44660 33900 47690 34930
rect 47850 33900 50880 34930
rect 51040 33900 54070 34930
rect 54230 33900 57260 34930
rect 57420 33900 60450 34930
rect 60610 33900 63640 34930
rect 63800 33900 66830 34930
rect 66990 33900 70020 34930
rect 70180 33900 73210 34930
rect 73370 33900 76400 34930
rect 76560 33900 79590 34930
rect 79750 33900 82780 34930
rect 82940 33900 85970 34930
rect 86130 33900 89160 34930
rect 89320 33900 92350 34930
rect 92510 33900 95540 34930
rect 95700 33900 98730 34930
rect 98890 33900 101920 34930
rect 102080 33900 105110 34930
rect 105270 33900 108300 34930
rect 108460 33900 111490 34930
rect 111650 33900 114680 34930
rect 114840 33900 117870 34930
rect 118030 33900 121060 34930
rect 121220 33900 124250 34930
rect 124410 33900 127440 34930
rect 127600 33900 130630 34930
rect 130790 33900 133820 34930
rect 133980 33900 137010 34930
rect 0 32900 137170 33900
rect 0 31900 3030 32900
rect 3190 31900 6220 32900
rect 6380 31900 9410 32900
rect 9570 31900 12600 32900
rect 12760 31900 15790 32900
rect 15950 31900 18980 32900
rect 19140 31900 22170 32900
rect 22330 31900 25360 32900
rect 25520 31900 28550 32900
rect 28710 31900 31740 32900
rect 31900 31900 34930 32900
rect 35090 31900 38120 32900
rect 38280 31900 41310 32900
rect 41470 31900 44500 32900
rect 44660 31900 47690 32900
rect 47850 31900 50880 32900
rect 51040 31900 54070 32900
rect 54230 31900 57260 32900
rect 57420 31900 60450 32900
rect 60610 31900 63640 32900
rect 63800 31900 66830 32900
rect 66990 31900 70020 32900
rect 70180 31900 73210 32900
rect 73370 31900 76400 32900
rect 76560 31900 79590 32900
rect 79750 31900 82780 32900
rect 82940 31900 85970 32900
rect 86130 31900 89160 32900
rect 89320 31900 92350 32900
rect 92510 31900 95540 32900
rect 95700 31900 98730 32900
rect 98890 31900 101920 32900
rect 102080 31900 105110 32900
rect 105270 31900 108300 32900
rect 108460 31900 111490 32900
rect 111650 31900 114680 32900
rect 114840 31900 117870 32900
rect 118030 31900 121060 32900
rect 121220 31900 124250 32900
rect 124410 31900 127440 32900
rect 127600 31900 130630 32900
rect 130790 31900 133820 32900
rect 133980 31900 137010 32900
rect 1000 31740 2000 31900
rect 4190 31740 5190 31900
rect 7380 31740 8380 31900
rect 10570 31740 11570 31900
rect 13760 31740 14760 31900
rect 16950 31740 17950 31900
rect 20140 31740 21140 31900
rect 23330 31740 24330 31900
rect 26520 31740 27520 31900
rect 29710 31740 30710 31900
rect 32900 31740 33900 31900
rect 36090 31740 37090 31900
rect 39280 31740 40280 31900
rect 42470 31740 43470 31900
rect 45660 31740 46660 31900
rect 48850 31740 49850 31900
rect 52040 31740 53040 31900
rect 55230 31740 56230 31900
rect 58420 31740 59420 31900
rect 61610 31740 62610 31900
rect 64800 31740 65800 31900
rect 67990 31740 68990 31900
rect 71180 31740 72180 31900
rect 74370 31740 75370 31900
rect 77560 31740 78560 31900
rect 80750 31740 81750 31900
rect 83940 31740 84940 31900
rect 87130 31740 88130 31900
rect 90320 31740 91320 31900
rect 93510 31740 94510 31900
rect 96700 31740 97700 31900
rect 99890 31740 100890 31900
rect 103080 31740 104080 31900
rect 106270 31740 107270 31900
rect 109460 31740 110460 31900
rect 112650 31740 113650 31900
rect 115840 31740 116840 31900
rect 119030 31740 120030 31900
rect 122220 31740 123220 31900
rect 125410 31740 126410 31900
rect 128600 31740 129600 31900
rect 131790 31740 132790 31900
rect 134980 31740 135980 31900
rect 0 30710 3030 31740
rect 3190 30710 6220 31740
rect 6380 30710 9410 31740
rect 9570 30710 12600 31740
rect 12760 30710 15790 31740
rect 15950 30710 18980 31740
rect 19140 30710 22170 31740
rect 22330 30710 25360 31740
rect 25520 30710 28550 31740
rect 28710 30710 31740 31740
rect 31900 30710 34930 31740
rect 35090 30710 38120 31740
rect 38280 30710 41310 31740
rect 41470 30710 44500 31740
rect 44660 30710 47690 31740
rect 47850 30710 50880 31740
rect 51040 30710 54070 31740
rect 54230 30710 57260 31740
rect 57420 30710 60450 31740
rect 60610 30710 63640 31740
rect 63800 30710 66830 31740
rect 66990 30710 70020 31740
rect 70180 30710 73210 31740
rect 73370 30710 76400 31740
rect 76560 30710 79590 31740
rect 79750 30710 82780 31740
rect 82940 30710 85970 31740
rect 86130 30710 89160 31740
rect 89320 30710 92350 31740
rect 92510 30710 95540 31740
rect 95700 30710 98730 31740
rect 98890 30710 101920 31740
rect 102080 30710 105110 31740
rect 105270 30710 108300 31740
rect 108460 30710 111490 31740
rect 111650 30710 114680 31740
rect 114840 30710 117870 31740
rect 118030 30710 121060 31740
rect 121220 30710 124250 31740
rect 124410 30710 127440 31740
rect 127600 30710 130630 31740
rect 130790 30710 133820 31740
rect 133980 30710 137010 31740
rect 0 29710 137170 30710
rect 0 28710 3030 29710
rect 3190 28710 6220 29710
rect 6380 28710 9410 29710
rect 9570 28710 12600 29710
rect 12760 28710 15790 29710
rect 15950 28710 18980 29710
rect 19140 28710 22170 29710
rect 22330 28710 25360 29710
rect 25520 28710 28550 29710
rect 28710 28710 31740 29710
rect 31900 28710 34930 29710
rect 35090 28710 38120 29710
rect 38280 28710 41310 29710
rect 41470 28710 44500 29710
rect 44660 28710 47690 29710
rect 47850 28710 50880 29710
rect 51040 28710 54070 29710
rect 54230 28710 57260 29710
rect 57420 28710 60450 29710
rect 60610 28710 63640 29710
rect 63800 28710 66830 29710
rect 66990 28710 70020 29710
rect 70180 28710 73210 29710
rect 73370 28710 76400 29710
rect 76560 28710 79590 29710
rect 79750 28710 82780 29710
rect 82940 28710 85970 29710
rect 86130 28710 89160 29710
rect 89320 28710 92350 29710
rect 92510 28710 95540 29710
rect 95700 28710 98730 29710
rect 98890 28710 101920 29710
rect 102080 28710 105110 29710
rect 105270 28710 108300 29710
rect 108460 28710 111490 29710
rect 111650 28710 114680 29710
rect 114840 28710 117870 29710
rect 118030 28710 121060 29710
rect 121220 28710 124250 29710
rect 124410 28710 127440 29710
rect 127600 28710 130630 29710
rect 130790 28710 133820 29710
rect 133980 28710 137010 29710
rect 1000 28550 2000 28710
rect 4190 28550 5190 28710
rect 7380 28550 8380 28710
rect 10570 28550 11570 28710
rect 13760 28550 14760 28710
rect 16950 28550 17950 28710
rect 20140 28550 21140 28710
rect 23330 28550 24330 28710
rect 26520 28550 27520 28710
rect 29710 28550 30710 28710
rect 32900 28550 33900 28710
rect 36090 28550 37090 28710
rect 39280 28550 40280 28710
rect 42470 28550 43470 28710
rect 45660 28550 46660 28710
rect 48850 28550 49850 28710
rect 52040 28550 53040 28710
rect 55230 28550 56230 28710
rect 58420 28550 59420 28710
rect 61610 28550 62610 28710
rect 64800 28550 65800 28710
rect 67990 28550 68990 28710
rect 71180 28550 72180 28710
rect 74370 28550 75370 28710
rect 77560 28550 78560 28710
rect 80750 28550 81750 28710
rect 83940 28550 84940 28710
rect 87130 28550 88130 28710
rect 90320 28550 91320 28710
rect 93510 28550 94510 28710
rect 96700 28550 97700 28710
rect 99890 28550 100890 28710
rect 103080 28550 104080 28710
rect 106270 28550 107270 28710
rect 109460 28550 110460 28710
rect 112650 28550 113650 28710
rect 115840 28550 116840 28710
rect 119030 28550 120030 28710
rect 122220 28550 123220 28710
rect 125410 28550 126410 28710
rect 128600 28550 129600 28710
rect 131790 28550 132790 28710
rect 134980 28550 135980 28710
rect 0 27520 3030 28550
rect 3190 27520 6220 28550
rect 6380 27520 9410 28550
rect 9570 27520 12600 28550
rect 12760 27520 15790 28550
rect 15950 27520 18980 28550
rect 19140 27520 22170 28550
rect 22330 27520 25360 28550
rect 25520 27520 28550 28550
rect 28710 27520 31740 28550
rect 31900 27520 34930 28550
rect 35090 27520 38120 28550
rect 38280 27520 41310 28550
rect 41470 27520 44500 28550
rect 44660 27520 47690 28550
rect 47850 27520 50880 28550
rect 51040 27520 54070 28550
rect 54230 27520 57260 28550
rect 57420 27520 60450 28550
rect 60610 27520 63640 28550
rect 63800 27520 66830 28550
rect 66990 27520 70020 28550
rect 70180 27520 73210 28550
rect 73370 27520 76400 28550
rect 76560 27520 79590 28550
rect 79750 27520 82780 28550
rect 82940 27520 85970 28550
rect 86130 27520 89160 28550
rect 89320 27520 92350 28550
rect 92510 27520 95540 28550
rect 95700 27520 98730 28550
rect 98890 27520 101920 28550
rect 102080 27520 105110 28550
rect 105270 27520 108300 28550
rect 108460 27520 111490 28550
rect 111650 27520 114680 28550
rect 114840 27520 117870 28550
rect 118030 27520 121060 28550
rect 121220 27520 124250 28550
rect 124410 27520 127440 28550
rect 127600 27520 130630 28550
rect 130790 27520 133820 28550
rect 133980 27520 137010 28550
rect 0 26520 137170 27520
rect 0 25520 3030 26520
rect 3190 25520 6220 26520
rect 6380 25520 9410 26520
rect 9570 25520 12600 26520
rect 12760 25520 15790 26520
rect 15950 25520 18980 26520
rect 19140 25520 22170 26520
rect 22330 25520 25360 26520
rect 25520 25520 28550 26520
rect 28710 25520 31740 26520
rect 31900 25520 34930 26520
rect 35090 25520 38120 26520
rect 38280 25520 41310 26520
rect 41470 25520 44500 26520
rect 44660 25520 47690 26520
rect 47850 25520 50880 26520
rect 51040 25520 54070 26520
rect 54230 25520 57260 26520
rect 57420 25520 60450 26520
rect 60610 25520 63640 26520
rect 63800 25520 66830 26520
rect 66990 25520 70020 26520
rect 70180 25520 73210 26520
rect 73370 25520 76400 26520
rect 76560 25520 79590 26520
rect 79750 25520 82780 26520
rect 82940 25520 85970 26520
rect 86130 25520 89160 26520
rect 89320 25520 92350 26520
rect 92510 25520 95540 26520
rect 95700 25520 98730 26520
rect 98890 25520 101920 26520
rect 102080 25520 105110 26520
rect 105270 25520 108300 26520
rect 108460 25520 111490 26520
rect 111650 25520 114680 26520
rect 114840 25520 117870 26520
rect 118030 25520 121060 26520
rect 121220 25520 124250 26520
rect 124410 25520 127440 26520
rect 127600 25520 130630 26520
rect 130790 25520 133820 26520
rect 133980 25520 137010 26520
rect 1000 25360 2000 25520
rect 4190 25360 5190 25520
rect 7380 25360 8380 25520
rect 10570 25360 11570 25520
rect 13760 25360 14760 25520
rect 16950 25360 17950 25520
rect 20140 25360 21140 25520
rect 23330 25360 24330 25520
rect 26520 25360 27520 25520
rect 29710 25360 30710 25520
rect 32900 25360 33900 25520
rect 36090 25360 37090 25520
rect 39280 25360 40280 25520
rect 42470 25360 43470 25520
rect 45660 25360 46660 25520
rect 48850 25360 49850 25520
rect 52040 25360 53040 25520
rect 55230 25360 56230 25520
rect 58420 25360 59420 25520
rect 61610 25360 62610 25520
rect 64800 25360 65800 25520
rect 67990 25360 68990 25520
rect 71180 25360 72180 25520
rect 74370 25360 75370 25520
rect 77560 25360 78560 25520
rect 80750 25360 81750 25520
rect 83940 25360 84940 25520
rect 87130 25360 88130 25520
rect 90320 25360 91320 25520
rect 93510 25360 94510 25520
rect 96700 25360 97700 25520
rect 99890 25360 100890 25520
rect 103080 25360 104080 25520
rect 106270 25360 107270 25520
rect 109460 25360 110460 25520
rect 112650 25360 113650 25520
rect 115840 25360 116840 25520
rect 119030 25360 120030 25520
rect 122220 25360 123220 25520
rect 125410 25360 126410 25520
rect 128600 25360 129600 25520
rect 131790 25360 132790 25520
rect 134980 25360 135980 25520
rect 0 24330 3030 25360
rect 3190 24330 6220 25360
rect 6380 24330 9410 25360
rect 9570 24330 12600 25360
rect 12760 24330 15790 25360
rect 15950 24330 18980 25360
rect 19140 24330 22170 25360
rect 22330 24330 25360 25360
rect 25520 24330 28550 25360
rect 28710 24330 31740 25360
rect 31900 24330 34930 25360
rect 35090 24330 38120 25360
rect 38280 24330 41310 25360
rect 41470 24330 44500 25360
rect 44660 24330 47690 25360
rect 47850 24330 50880 25360
rect 51040 24330 54070 25360
rect 54230 24330 57260 25360
rect 57420 24330 60450 25360
rect 60610 24330 63640 25360
rect 63800 24330 66830 25360
rect 66990 24330 70020 25360
rect 70180 24330 73210 25360
rect 73370 24330 76400 25360
rect 76560 24330 79590 25360
rect 79750 24330 82780 25360
rect 82940 24330 85970 25360
rect 86130 24330 89160 25360
rect 89320 24330 92350 25360
rect 92510 24330 95540 25360
rect 95700 24330 98730 25360
rect 98890 24330 101920 25360
rect 102080 24330 105110 25360
rect 105270 24330 108300 25360
rect 108460 24330 111490 25360
rect 111650 24330 114680 25360
rect 114840 24330 117870 25360
rect 118030 24330 121060 25360
rect 121220 24330 124250 25360
rect 124410 24330 127440 25360
rect 127600 24330 130630 25360
rect 130790 24330 133820 25360
rect 133980 24330 137010 25360
rect 0 23330 137170 24330
rect 0 22330 3030 23330
rect 3190 22330 6220 23330
rect 6380 22330 9410 23330
rect 9570 22330 12600 23330
rect 12760 22330 15790 23330
rect 15950 22330 18980 23330
rect 19140 22330 22170 23330
rect 22330 22330 25360 23330
rect 25520 22330 28550 23330
rect 28710 22330 31740 23330
rect 31900 22330 34930 23330
rect 35090 22330 38120 23330
rect 38280 22330 41310 23330
rect 41470 22330 44500 23330
rect 44660 22330 47690 23330
rect 47850 22330 50880 23330
rect 51040 22330 54070 23330
rect 54230 22330 57260 23330
rect 57420 22330 60450 23330
rect 60610 22330 63640 23330
rect 63800 22330 66830 23330
rect 66990 22330 70020 23330
rect 70180 22330 73210 23330
rect 73370 22330 76400 23330
rect 76560 22330 79590 23330
rect 79750 22330 82780 23330
rect 82940 22330 85970 23330
rect 86130 22330 89160 23330
rect 89320 22330 92350 23330
rect 92510 22330 95540 23330
rect 95700 22330 98730 23330
rect 98890 22330 101920 23330
rect 102080 22330 105110 23330
rect 105270 22330 108300 23330
rect 108460 22330 111490 23330
rect 111650 22330 114680 23330
rect 114840 22330 117870 23330
rect 118030 22330 121060 23330
rect 121220 22330 124250 23330
rect 124410 22330 127440 23330
rect 127600 22330 130630 23330
rect 130790 22330 133820 23330
rect 133980 22330 137010 23330
rect 1000 22170 2000 22330
rect 4190 22170 5190 22330
rect 7380 22170 8380 22330
rect 10570 22170 11570 22330
rect 13760 22170 14760 22330
rect 16950 22170 17950 22330
rect 20140 22170 21140 22330
rect 23330 22170 24330 22330
rect 26520 22170 27520 22330
rect 29710 22170 30710 22330
rect 32900 22170 33900 22330
rect 36090 22170 37090 22330
rect 39280 22170 40280 22330
rect 42470 22170 43470 22330
rect 45660 22170 46660 22330
rect 48850 22170 49850 22330
rect 52040 22170 53040 22330
rect 55230 22170 56230 22330
rect 58420 22170 59420 22330
rect 61610 22170 62610 22330
rect 64800 22170 65800 22330
rect 67990 22170 68990 22330
rect 71180 22170 72180 22330
rect 74370 22170 75370 22330
rect 77560 22170 78560 22330
rect 80750 22170 81750 22330
rect 83940 22170 84940 22330
rect 87130 22170 88130 22330
rect 90320 22170 91320 22330
rect 93510 22170 94510 22330
rect 96700 22170 97700 22330
rect 99890 22170 100890 22330
rect 103080 22170 104080 22330
rect 106270 22170 107270 22330
rect 109460 22170 110460 22330
rect 112650 22170 113650 22330
rect 115840 22170 116840 22330
rect 119030 22170 120030 22330
rect 122220 22170 123220 22330
rect 125410 22170 126410 22330
rect 128600 22170 129600 22330
rect 131790 22170 132790 22330
rect 134980 22170 135980 22330
rect 0 21140 3030 22170
rect 3190 21140 6220 22170
rect 6380 21140 9410 22170
rect 9570 21140 12600 22170
rect 12760 21140 15790 22170
rect 15950 21140 18980 22170
rect 19140 21140 22170 22170
rect 22330 21140 25360 22170
rect 25520 21140 28550 22170
rect 28710 21140 31740 22170
rect 31900 21140 34930 22170
rect 35090 21140 38120 22170
rect 38280 21140 41310 22170
rect 41470 21140 44500 22170
rect 44660 21140 47690 22170
rect 47850 21140 50880 22170
rect 51040 21140 54070 22170
rect 54230 21140 57260 22170
rect 57420 21140 60450 22170
rect 60610 21140 63640 22170
rect 63800 21140 66830 22170
rect 66990 21140 70020 22170
rect 70180 21140 73210 22170
rect 73370 21140 76400 22170
rect 76560 21140 79590 22170
rect 79750 21140 82780 22170
rect 82940 21140 85970 22170
rect 86130 21140 89160 22170
rect 89320 21140 92350 22170
rect 92510 21140 95540 22170
rect 95700 21140 98730 22170
rect 98890 21140 101920 22170
rect 102080 21140 105110 22170
rect 105270 21140 108300 22170
rect 108460 21140 111490 22170
rect 111650 21140 114680 22170
rect 114840 21140 117870 22170
rect 118030 21140 121060 22170
rect 121220 21140 124250 22170
rect 124410 21140 127440 22170
rect 127600 21140 130630 22170
rect 130790 21140 133820 22170
rect 133980 21140 137010 22170
rect 0 20140 137170 21140
rect 0 19140 3030 20140
rect 3190 19140 6220 20140
rect 6380 19140 9410 20140
rect 9570 19140 12600 20140
rect 12760 19140 15790 20140
rect 15950 19140 18980 20140
rect 19140 19140 22170 20140
rect 22330 19140 25360 20140
rect 25520 19140 28550 20140
rect 28710 19140 31740 20140
rect 31900 19140 34930 20140
rect 35090 19140 38120 20140
rect 38280 19140 41310 20140
rect 41470 19140 44500 20140
rect 44660 19140 47690 20140
rect 47850 19140 50880 20140
rect 51040 19140 54070 20140
rect 54230 19140 57260 20140
rect 57420 19140 60450 20140
rect 60610 19140 63640 20140
rect 63800 19140 66830 20140
rect 66990 19140 70020 20140
rect 70180 19140 73210 20140
rect 73370 19140 76400 20140
rect 76560 19140 79590 20140
rect 79750 19140 82780 20140
rect 82940 19140 85970 20140
rect 86130 19140 89160 20140
rect 89320 19140 92350 20140
rect 92510 19140 95540 20140
rect 95700 19140 98730 20140
rect 98890 19140 101920 20140
rect 102080 19140 105110 20140
rect 105270 19140 108300 20140
rect 108460 19140 111490 20140
rect 111650 19140 114680 20140
rect 114840 19140 117870 20140
rect 118030 19140 121060 20140
rect 121220 19140 124250 20140
rect 124410 19140 127440 20140
rect 127600 19140 130630 20140
rect 130790 19140 133820 20140
rect 133980 19140 137010 20140
rect 1000 18980 2000 19140
rect 4190 18980 5190 19140
rect 7380 18980 8380 19140
rect 10570 18980 11570 19140
rect 13760 18980 14760 19140
rect 16950 18980 17950 19140
rect 20140 18980 21140 19140
rect 23330 18980 24330 19140
rect 26520 18980 27520 19140
rect 29710 18980 30710 19140
rect 32900 18980 33900 19140
rect 36090 18980 37090 19140
rect 39280 18980 40280 19140
rect 42470 18980 43470 19140
rect 45660 18980 46660 19140
rect 48850 18980 49850 19140
rect 52040 18980 53040 19140
rect 55230 18980 56230 19140
rect 58420 18980 59420 19140
rect 61610 18980 62610 19140
rect 64800 18980 65800 19140
rect 67990 18980 68990 19140
rect 71180 18980 72180 19140
rect 74370 18980 75370 19140
rect 77560 18980 78560 19140
rect 80750 18980 81750 19140
rect 83940 18980 84940 19140
rect 87130 18980 88130 19140
rect 90320 18980 91320 19140
rect 93510 18980 94510 19140
rect 96700 18980 97700 19140
rect 99890 18980 100890 19140
rect 103080 18980 104080 19140
rect 106270 18980 107270 19140
rect 109460 18980 110460 19140
rect 112650 18980 113650 19140
rect 115840 18980 116840 19140
rect 119030 18980 120030 19140
rect 122220 18980 123220 19140
rect 125410 18980 126410 19140
rect 128600 18980 129600 19140
rect 131790 18980 132790 19140
rect 134980 18980 135980 19140
rect 0 17950 3030 18980
rect 3190 17950 6220 18980
rect 6380 17950 9410 18980
rect 9570 17950 12600 18980
rect 12760 17950 15790 18980
rect 15950 17950 18980 18980
rect 19140 17950 22170 18980
rect 22330 17950 25360 18980
rect 25520 17950 28550 18980
rect 28710 17950 31740 18980
rect 31900 17950 34930 18980
rect 35090 17950 38120 18980
rect 38280 17950 41310 18980
rect 41470 17950 44500 18980
rect 44660 17950 47690 18980
rect 47850 17950 50880 18980
rect 51040 17950 54070 18980
rect 54230 17950 57260 18980
rect 57420 17950 60450 18980
rect 60610 17950 63640 18980
rect 63800 17950 66830 18980
rect 66990 17950 70020 18980
rect 70180 17950 73210 18980
rect 73370 17950 76400 18980
rect 76560 17950 79590 18980
rect 79750 17950 82780 18980
rect 82940 17950 85970 18980
rect 86130 17950 89160 18980
rect 89320 17950 92350 18980
rect 92510 17950 95540 18980
rect 95700 17950 98730 18980
rect 98890 17950 101920 18980
rect 102080 17950 105110 18980
rect 105270 17950 108300 18980
rect 108460 17950 111490 18980
rect 111650 17950 114680 18980
rect 114840 17950 117870 18980
rect 118030 17950 121060 18980
rect 121220 17950 124250 18980
rect 124410 17950 127440 18980
rect 127600 17950 130630 18980
rect 130790 17950 133820 18980
rect 133980 17950 137010 18980
rect 0 16950 137170 17950
rect 0 15950 3030 16950
rect 3190 15950 6220 16950
rect 6380 15950 9410 16950
rect 9570 15950 12600 16950
rect 12760 15950 15790 16950
rect 15950 15950 18980 16950
rect 19140 15950 22170 16950
rect 22330 15950 25360 16950
rect 25520 15950 28550 16950
rect 28710 15950 31740 16950
rect 31900 15950 34930 16950
rect 35090 15950 38120 16950
rect 38280 15950 41310 16950
rect 41470 15950 44500 16950
rect 44660 15950 47690 16950
rect 47850 15950 50880 16950
rect 51040 15950 54070 16950
rect 54230 15950 57260 16950
rect 57420 15950 60450 16950
rect 60610 15950 63640 16950
rect 63800 15950 66830 16950
rect 66990 15950 70020 16950
rect 70180 15950 73210 16950
rect 73370 15950 76400 16950
rect 76560 15950 79590 16950
rect 79750 15950 82780 16950
rect 82940 15950 85970 16950
rect 86130 15950 89160 16950
rect 89320 15950 92350 16950
rect 92510 15950 95540 16950
rect 95700 15950 98730 16950
rect 98890 15950 101920 16950
rect 102080 15950 105110 16950
rect 105270 15950 108300 16950
rect 108460 15950 111490 16950
rect 111650 15950 114680 16950
rect 114840 15950 117870 16950
rect 118030 15950 121060 16950
rect 121220 15950 124250 16950
rect 124410 15950 127440 16950
rect 127600 15950 130630 16950
rect 130790 15950 133820 16950
rect 133980 15950 137010 16950
rect 1000 15790 2000 15950
rect 4190 15790 5190 15950
rect 7380 15790 8380 15950
rect 10570 15790 11570 15950
rect 13760 15790 14760 15950
rect 16950 15790 17950 15950
rect 20140 15790 21140 15950
rect 23330 15790 24330 15950
rect 26520 15790 27520 15950
rect 29710 15790 30710 15950
rect 32900 15790 33900 15950
rect 36090 15790 37090 15950
rect 39280 15790 40280 15950
rect 42470 15790 43470 15950
rect 45660 15790 46660 15950
rect 48850 15790 49850 15950
rect 52040 15790 53040 15950
rect 55230 15790 56230 15950
rect 58420 15790 59420 15950
rect 61610 15790 62610 15950
rect 64800 15790 65800 15950
rect 67990 15790 68990 15950
rect 71180 15790 72180 15950
rect 74370 15790 75370 15950
rect 77560 15790 78560 15950
rect 80750 15790 81750 15950
rect 83940 15790 84940 15950
rect 87130 15790 88130 15950
rect 90320 15790 91320 15950
rect 93510 15790 94510 15950
rect 96700 15790 97700 15950
rect 99890 15790 100890 15950
rect 103080 15790 104080 15950
rect 106270 15790 107270 15950
rect 109460 15790 110460 15950
rect 112650 15790 113650 15950
rect 115840 15790 116840 15950
rect 119030 15790 120030 15950
rect 122220 15790 123220 15950
rect 125410 15790 126410 15950
rect 128600 15790 129600 15950
rect 131790 15790 132790 15950
rect 134980 15790 135980 15950
rect 0 14760 3030 15790
rect 3190 14760 6220 15790
rect 6380 14760 9410 15790
rect 9570 14760 12600 15790
rect 12760 14760 15790 15790
rect 15950 14760 18980 15790
rect 19140 14760 22170 15790
rect 22330 14760 25360 15790
rect 25520 14760 28550 15790
rect 28710 14760 31740 15790
rect 31900 14760 34930 15790
rect 35090 14760 38120 15790
rect 38280 14760 41310 15790
rect 41470 14760 44500 15790
rect 44660 14760 47690 15790
rect 47850 14760 50880 15790
rect 51040 14760 54070 15790
rect 54230 14760 57260 15790
rect 57420 14760 60450 15790
rect 60610 14760 63640 15790
rect 63800 14760 66830 15790
rect 66990 14760 70020 15790
rect 70180 14760 73210 15790
rect 73370 14760 76400 15790
rect 76560 14760 79590 15790
rect 79750 14760 82780 15790
rect 82940 14760 85970 15790
rect 86130 14760 89160 15790
rect 89320 14760 92350 15790
rect 92510 14760 95540 15790
rect 95700 14760 98730 15790
rect 98890 14760 101920 15790
rect 102080 14760 105110 15790
rect 105270 14760 108300 15790
rect 108460 14760 111490 15790
rect 111650 14760 114680 15790
rect 114840 14760 117870 15790
rect 118030 14760 121060 15790
rect 121220 14760 124250 15790
rect 124410 14760 127440 15790
rect 127600 14760 130630 15790
rect 130790 14760 133820 15790
rect 133980 14760 137010 15790
rect 0 13760 137170 14760
rect 0 12760 3030 13760
rect 3190 12760 6220 13760
rect 6380 12760 9410 13760
rect 9570 12760 12600 13760
rect 12760 12760 15790 13760
rect 15950 12760 18980 13760
rect 19140 12760 22170 13760
rect 22330 12760 25360 13760
rect 25520 12760 28550 13760
rect 28710 12760 31740 13760
rect 31900 12760 34930 13760
rect 35090 12760 38120 13760
rect 38280 12760 41310 13760
rect 41470 12760 44500 13760
rect 44660 12760 47690 13760
rect 47850 12760 50880 13760
rect 51040 12760 54070 13760
rect 54230 12760 57260 13760
rect 57420 12760 60450 13760
rect 60610 12760 63640 13760
rect 63800 12760 66830 13760
rect 66990 12760 70020 13760
rect 70180 12760 73210 13760
rect 73370 12760 76400 13760
rect 76560 12760 79590 13760
rect 79750 12760 82780 13760
rect 82940 12760 85970 13760
rect 86130 12760 89160 13760
rect 89320 12760 92350 13760
rect 92510 12760 95540 13760
rect 95700 12760 98730 13760
rect 98890 12760 101920 13760
rect 102080 12760 105110 13760
rect 105270 12760 108300 13760
rect 108460 12760 111490 13760
rect 111650 12760 114680 13760
rect 114840 12760 117870 13760
rect 118030 12760 121060 13760
rect 121220 12760 124250 13760
rect 124410 12760 127440 13760
rect 127600 12760 130630 13760
rect 130790 12760 133820 13760
rect 133980 12760 137010 13760
rect 1000 12600 2000 12760
rect 4190 12600 5190 12760
rect 7380 12600 8380 12760
rect 10570 12600 11570 12760
rect 13760 12600 14760 12760
rect 16950 12600 17950 12760
rect 20140 12600 21140 12760
rect 23330 12600 24330 12760
rect 26520 12600 27520 12760
rect 29710 12600 30710 12760
rect 32900 12600 33900 12760
rect 36090 12600 37090 12760
rect 39280 12600 40280 12760
rect 42470 12600 43470 12760
rect 45660 12600 46660 12760
rect 48850 12600 49850 12760
rect 52040 12600 53040 12760
rect 55230 12600 56230 12760
rect 58420 12600 59420 12760
rect 61610 12600 62610 12760
rect 64800 12600 65800 12760
rect 67990 12600 68990 12760
rect 71180 12600 72180 12760
rect 74370 12600 75370 12760
rect 77560 12600 78560 12760
rect 80750 12600 81750 12760
rect 83940 12600 84940 12760
rect 87130 12600 88130 12760
rect 90320 12600 91320 12760
rect 93510 12600 94510 12760
rect 96700 12600 97700 12760
rect 99890 12600 100890 12760
rect 103080 12600 104080 12760
rect 106270 12600 107270 12760
rect 109460 12600 110460 12760
rect 112650 12600 113650 12760
rect 115840 12600 116840 12760
rect 119030 12600 120030 12760
rect 122220 12600 123220 12760
rect 125410 12600 126410 12760
rect 128600 12600 129600 12760
rect 131790 12600 132790 12760
rect 134980 12600 135980 12760
rect 0 11570 3030 12600
rect 3190 11570 6220 12600
rect 6380 11570 9410 12600
rect 9570 11570 12600 12600
rect 12760 11570 15790 12600
rect 15950 11570 18980 12600
rect 19140 11570 22170 12600
rect 22330 11570 25360 12600
rect 25520 11570 28550 12600
rect 28710 11570 31740 12600
rect 31900 11570 34930 12600
rect 35090 11570 38120 12600
rect 38280 11570 41310 12600
rect 41470 11570 44500 12600
rect 44660 11570 47690 12600
rect 47850 11570 50880 12600
rect 51040 11570 54070 12600
rect 54230 11570 57260 12600
rect 57420 11570 60450 12600
rect 60610 11570 63640 12600
rect 63800 11570 66830 12600
rect 66990 11570 70020 12600
rect 70180 11570 73210 12600
rect 73370 11570 76400 12600
rect 76560 11570 79590 12600
rect 79750 11570 82780 12600
rect 82940 11570 85970 12600
rect 86130 11570 89160 12600
rect 89320 11570 92350 12600
rect 92510 11570 95540 12600
rect 95700 11570 98730 12600
rect 98890 11570 101920 12600
rect 102080 11570 105110 12600
rect 105270 11570 108300 12600
rect 108460 11570 111490 12600
rect 111650 11570 114680 12600
rect 114840 11570 117870 12600
rect 118030 11570 121060 12600
rect 121220 11570 124250 12600
rect 124410 11570 127440 12600
rect 127600 11570 130630 12600
rect 130790 11570 133820 12600
rect 133980 11570 137010 12600
rect 0 10570 137170 11570
rect 0 9570 3030 10570
rect 3190 9570 6220 10570
rect 6380 9570 9410 10570
rect 9570 9570 12600 10570
rect 12760 9570 15790 10570
rect 15950 9570 18980 10570
rect 19140 9570 22170 10570
rect 22330 9570 25360 10570
rect 25520 9570 28550 10570
rect 28710 9570 31740 10570
rect 31900 9570 34930 10570
rect 35090 9570 38120 10570
rect 38280 9570 41310 10570
rect 41470 9570 44500 10570
rect 44660 9570 47690 10570
rect 47850 9570 50880 10570
rect 51040 9570 54070 10570
rect 54230 9570 57260 10570
rect 57420 9570 60450 10570
rect 60610 9570 63640 10570
rect 63800 9570 66830 10570
rect 66990 9570 70020 10570
rect 70180 9570 73210 10570
rect 73370 9570 76400 10570
rect 76560 9570 79590 10570
rect 79750 9570 82780 10570
rect 82940 9570 85970 10570
rect 86130 9570 89160 10570
rect 89320 9570 92350 10570
rect 92510 9570 95540 10570
rect 95700 9570 98730 10570
rect 98890 9570 101920 10570
rect 102080 9570 105110 10570
rect 105270 9570 108300 10570
rect 108460 9570 111490 10570
rect 111650 9570 114680 10570
rect 114840 9570 117870 10570
rect 118030 9570 121060 10570
rect 121220 9570 124250 10570
rect 124410 9570 127440 10570
rect 127600 9570 130630 10570
rect 130790 9570 133820 10570
rect 133980 9570 137010 10570
rect 1000 9410 2000 9570
rect 4190 9410 5190 9570
rect 7380 9410 8380 9570
rect 10570 9410 11570 9570
rect 13760 9410 14760 9570
rect 16950 9410 17950 9570
rect 20140 9410 21140 9570
rect 23330 9410 24330 9570
rect 26520 9410 27520 9570
rect 29710 9410 30710 9570
rect 32900 9410 33900 9570
rect 36090 9410 37090 9570
rect 39280 9410 40280 9570
rect 42470 9410 43470 9570
rect 45660 9410 46660 9570
rect 48850 9410 49850 9570
rect 52040 9410 53040 9570
rect 55230 9410 56230 9570
rect 58420 9410 59420 9570
rect 61610 9410 62610 9570
rect 64800 9410 65800 9570
rect 67990 9410 68990 9570
rect 71180 9410 72180 9570
rect 74370 9410 75370 9570
rect 77560 9410 78560 9570
rect 80750 9410 81750 9570
rect 83940 9410 84940 9570
rect 87130 9410 88130 9570
rect 90320 9410 91320 9570
rect 93510 9410 94510 9570
rect 96700 9410 97700 9570
rect 99890 9410 100890 9570
rect 103080 9410 104080 9570
rect 106270 9410 107270 9570
rect 109460 9410 110460 9570
rect 112650 9410 113650 9570
rect 115840 9410 116840 9570
rect 119030 9410 120030 9570
rect 122220 9410 123220 9570
rect 125410 9410 126410 9570
rect 128600 9410 129600 9570
rect 131790 9410 132790 9570
rect 134980 9410 135980 9570
rect 0 8380 3030 9410
rect 3190 8380 6220 9410
rect 6380 8380 9410 9410
rect 9570 8380 12600 9410
rect 12760 8380 15790 9410
rect 15950 8380 18980 9410
rect 19140 8380 22170 9410
rect 22330 8380 25360 9410
rect 25520 8380 28550 9410
rect 28710 8380 31740 9410
rect 31900 8380 34930 9410
rect 35090 8380 38120 9410
rect 38280 8380 41310 9410
rect 41470 8380 44500 9410
rect 44660 8380 47690 9410
rect 47850 8380 50880 9410
rect 51040 8380 54070 9410
rect 54230 8380 57260 9410
rect 57420 8380 60450 9410
rect 60610 8380 63640 9410
rect 63800 8380 66830 9410
rect 66990 8380 70020 9410
rect 70180 8380 73210 9410
rect 73370 8380 76400 9410
rect 76560 8380 79590 9410
rect 79750 8380 82780 9410
rect 82940 8380 85970 9410
rect 86130 8380 89160 9410
rect 89320 8380 92350 9410
rect 92510 8380 95540 9410
rect 95700 8380 98730 9410
rect 98890 8380 101920 9410
rect 102080 8380 105110 9410
rect 105270 8380 108300 9410
rect 108460 8380 111490 9410
rect 111650 8380 114680 9410
rect 114840 8380 117870 9410
rect 118030 8380 121060 9410
rect 121220 8380 124250 9410
rect 124410 8380 127440 9410
rect 127600 8380 130630 9410
rect 130790 8380 133820 9410
rect 133980 8380 137010 9410
rect 0 7380 137170 8380
rect 0 6380 3030 7380
rect 3190 6380 6220 7380
rect 6380 6380 9410 7380
rect 9570 6380 12600 7380
rect 12760 6380 15790 7380
rect 15950 6380 18980 7380
rect 19140 6380 22170 7380
rect 22330 6380 25360 7380
rect 25520 6380 28550 7380
rect 28710 6380 31740 7380
rect 31900 6380 34930 7380
rect 35090 6380 38120 7380
rect 38280 6380 41310 7380
rect 41470 6380 44500 7380
rect 44660 6380 47690 7380
rect 47850 6380 50880 7380
rect 51040 6380 54070 7380
rect 54230 6380 57260 7380
rect 57420 6380 60450 7380
rect 60610 6380 63640 7380
rect 63800 6380 66830 7380
rect 66990 6380 70020 7380
rect 70180 6380 73210 7380
rect 73370 6380 76400 7380
rect 76560 6380 79590 7380
rect 79750 6380 82780 7380
rect 82940 6380 85970 7380
rect 86130 6380 89160 7380
rect 89320 6380 92350 7380
rect 92510 6380 95540 7380
rect 95700 6380 98730 7380
rect 98890 6380 101920 7380
rect 102080 6380 105110 7380
rect 105270 6380 108300 7380
rect 108460 6380 111490 7380
rect 111650 6380 114680 7380
rect 114840 6380 117870 7380
rect 118030 6380 121060 7380
rect 121220 6380 124250 7380
rect 124410 6380 127440 7380
rect 127600 6380 130630 7380
rect 130790 6380 133820 7380
rect 133980 6380 137010 7380
rect 1000 6220 2000 6380
rect 4190 6220 5190 6380
rect 7380 6220 8380 6380
rect 10570 6220 11570 6380
rect 13760 6220 14760 6380
rect 16950 6220 17950 6380
rect 20140 6220 21140 6380
rect 23330 6220 24330 6380
rect 26520 6220 27520 6380
rect 29710 6220 30710 6380
rect 32900 6220 33900 6380
rect 36090 6220 37090 6380
rect 39280 6220 40280 6380
rect 42470 6220 43470 6380
rect 45660 6220 46660 6380
rect 48850 6220 49850 6380
rect 52040 6220 53040 6380
rect 55230 6220 56230 6380
rect 58420 6220 59420 6380
rect 61610 6220 62610 6380
rect 64800 6220 65800 6380
rect 67990 6220 68990 6380
rect 71180 6220 72180 6380
rect 74370 6220 75370 6380
rect 77560 6220 78560 6380
rect 80750 6220 81750 6380
rect 83940 6220 84940 6380
rect 87130 6220 88130 6380
rect 90320 6220 91320 6380
rect 93510 6220 94510 6380
rect 96700 6220 97700 6380
rect 99890 6220 100890 6380
rect 103080 6220 104080 6380
rect 106270 6220 107270 6380
rect 109460 6220 110460 6380
rect 112650 6220 113650 6380
rect 115840 6220 116840 6380
rect 119030 6220 120030 6380
rect 122220 6220 123220 6380
rect 125410 6220 126410 6380
rect 128600 6220 129600 6380
rect 131790 6220 132790 6380
rect 134980 6220 135980 6380
rect 0 5190 3030 6220
rect 3190 5190 6220 6220
rect 6380 5190 9410 6220
rect 9570 5190 12600 6220
rect 12760 5190 15790 6220
rect 15950 5190 18980 6220
rect 19140 5190 22170 6220
rect 22330 5190 25360 6220
rect 25520 5190 28550 6220
rect 28710 5190 31740 6220
rect 31900 5190 34930 6220
rect 35090 5190 38120 6220
rect 38280 5190 41310 6220
rect 41470 5190 44500 6220
rect 44660 5190 47690 6220
rect 47850 5190 50880 6220
rect 51040 5190 54070 6220
rect 54230 5190 57260 6220
rect 57420 5190 60450 6220
rect 60610 5190 63640 6220
rect 63800 5190 66830 6220
rect 66990 5190 70020 6220
rect 70180 5190 73210 6220
rect 73370 5190 76400 6220
rect 76560 5190 79590 6220
rect 79750 5190 82780 6220
rect 82940 5190 85970 6220
rect 86130 5190 89160 6220
rect 89320 5190 92350 6220
rect 92510 5190 95540 6220
rect 95700 5190 98730 6220
rect 98890 5190 101920 6220
rect 102080 5190 105110 6220
rect 105270 5190 108300 6220
rect 108460 5190 111490 6220
rect 111650 5190 114680 6220
rect 114840 5190 117870 6220
rect 118030 5190 121060 6220
rect 121220 5190 124250 6220
rect 124410 5190 127440 6220
rect 127600 5190 130630 6220
rect 130790 5190 133820 6220
rect 133980 5190 137010 6220
rect 0 4190 137170 5190
rect 0 3190 3030 4190
rect 3190 3190 6220 4190
rect 6380 3190 9410 4190
rect 9570 3190 12600 4190
rect 12760 3190 15790 4190
rect 15950 3190 18980 4190
rect 19140 3190 22170 4190
rect 22330 3190 25360 4190
rect 25520 3190 28550 4190
rect 28710 3190 31740 4190
rect 31900 3190 34930 4190
rect 35090 3190 38120 4190
rect 38280 3190 41310 4190
rect 41470 3190 44500 4190
rect 44660 3190 47690 4190
rect 47850 3190 50880 4190
rect 51040 3190 54070 4190
rect 54230 3190 57260 4190
rect 57420 3190 60450 4190
rect 60610 3190 63640 4190
rect 63800 3190 66830 4190
rect 66990 3190 70020 4190
rect 70180 3190 73210 4190
rect 73370 3190 76400 4190
rect 76560 3190 79590 4190
rect 79750 3190 82780 4190
rect 82940 3190 85970 4190
rect 86130 3190 89160 4190
rect 89320 3190 92350 4190
rect 92510 3190 95540 4190
rect 95700 3190 98730 4190
rect 98890 3190 101920 4190
rect 102080 3190 105110 4190
rect 105270 3190 108300 4190
rect 108460 3190 111490 4190
rect 111650 3190 114680 4190
rect 114840 3190 117870 4190
rect 118030 3190 121060 4190
rect 121220 3190 124250 4190
rect 124410 3190 127440 4190
rect 127600 3190 130630 4190
rect 130790 3190 133820 4190
rect 133980 3190 137010 4190
rect 1000 3030 2000 3190
rect 4190 3030 5190 3190
rect 7380 3030 8380 3190
rect 10570 3030 11570 3190
rect 13760 3030 14760 3190
rect 16950 3030 17950 3190
rect 20140 3030 21140 3190
rect 23330 3030 24330 3190
rect 26520 3030 27520 3190
rect 29710 3030 30710 3190
rect 32900 3030 33900 3190
rect 36090 3030 37090 3190
rect 39280 3030 40280 3190
rect 42470 3030 43470 3190
rect 45660 3030 46660 3190
rect 48850 3030 49850 3190
rect 52040 3030 53040 3190
rect 55230 3030 56230 3190
rect 58420 3030 59420 3190
rect 61610 3030 62610 3190
rect 64800 3030 65800 3190
rect 67990 3030 68990 3190
rect 71180 3030 72180 3190
rect 74370 3030 75370 3190
rect 77560 3030 78560 3190
rect 80750 3030 81750 3190
rect 83940 3030 84940 3190
rect 87130 3030 88130 3190
rect 90320 3030 91320 3190
rect 93510 3030 94510 3190
rect 96700 3030 97700 3190
rect 99890 3030 100890 3190
rect 103080 3030 104080 3190
rect 106270 3030 107270 3190
rect 109460 3030 110460 3190
rect 112650 3030 113650 3190
rect 115840 3030 116840 3190
rect 119030 3030 120030 3190
rect 122220 3030 123220 3190
rect 125410 3030 126410 3190
rect 128600 3030 129600 3190
rect 131790 3030 132790 3190
rect 134980 3030 135980 3190
rect 0 2000 3030 3030
rect 3190 2000 6220 3030
rect 6380 2000 9410 3030
rect 9570 2000 12600 3030
rect 12760 2000 15790 3030
rect 15950 2000 18980 3030
rect 19140 2000 22170 3030
rect 22330 2000 25360 3030
rect 25520 2000 28550 3030
rect 28710 2000 31740 3030
rect 31900 2000 34930 3030
rect 35090 2000 38120 3030
rect 38280 2000 41310 3030
rect 41470 2000 44500 3030
rect 44660 2000 47690 3030
rect 47850 2000 50880 3030
rect 51040 2000 54070 3030
rect 54230 2000 57260 3030
rect 57420 2000 60450 3030
rect 60610 2000 63640 3030
rect 63800 2000 66830 3030
rect 66990 2000 70020 3030
rect 70180 2000 73210 3030
rect 73370 2000 76400 3030
rect 76560 2000 79590 3030
rect 79750 2000 82780 3030
rect 82940 2000 85970 3030
rect 86130 2000 89160 3030
rect 89320 2000 92350 3030
rect 92510 2000 95540 3030
rect 95700 2000 98730 3030
rect 98890 2000 101920 3030
rect 102080 2000 105110 3030
rect 105270 2000 108300 3030
rect 108460 2000 111490 3030
rect 111650 2000 114680 3030
rect 114840 2000 117870 3030
rect 118030 2000 121060 3030
rect 121220 2000 124250 3030
rect 124410 2000 127440 3030
rect 127600 2000 130630 3030
rect 130790 2000 133820 3030
rect 133980 2000 137010 3030
rect 0 1000 137170 2000
rect 0 0 3030 1000
rect 3190 0 6220 1000
rect 6380 0 9410 1000
rect 9570 0 12600 1000
rect 12760 0 15790 1000
rect 15950 0 18980 1000
rect 19140 0 22170 1000
rect 22330 0 25360 1000
rect 25520 0 28550 1000
rect 28710 0 31740 1000
rect 31900 0 34930 1000
rect 35090 0 38120 1000
rect 38280 0 41310 1000
rect 41470 0 44500 1000
rect 44660 0 47690 1000
rect 47850 0 50880 1000
rect 51040 0 54070 1000
rect 54230 0 57260 1000
rect 57420 0 60450 1000
rect 60610 0 63640 1000
rect 63800 0 66830 1000
rect 66990 0 70020 1000
rect 70180 0 73210 1000
rect 73370 0 76400 1000
rect 76560 0 79590 1000
rect 79750 0 82780 1000
rect 82940 0 85970 1000
rect 86130 0 89160 1000
rect 89320 0 92350 1000
rect 92510 0 95540 1000
rect 95700 0 98730 1000
rect 98890 0 101920 1000
rect 102080 0 105110 1000
rect 105270 0 108300 1000
rect 108460 0 111490 1000
rect 111650 0 114680 1000
rect 114840 0 117870 1000
rect 118030 0 121060 1000
rect 121220 0 124250 1000
rect 124410 0 127440 1000
rect 127600 0 130630 1000
rect 130790 0 133820 1000
rect 133980 0 137010 1000
<< via3 >>
rect 1020 166020 68970 166980
rect 71200 166020 135960 166980
rect 50 121310 9320 140110
rect 50 79839 9320 98639
<< mimcap >>
rect 15 165697 3015 165705
rect 15 162713 23 165697
rect 3007 162713 3015 165697
rect 15 162705 3015 162713
rect 3205 165697 6205 165705
rect 3205 162713 3213 165697
rect 6197 162713 6205 165697
rect 3205 162705 6205 162713
rect 6395 165697 9395 165705
rect 6395 162713 6403 165697
rect 9387 162713 9395 165697
rect 6395 162705 9395 162713
rect 9585 165697 12585 165705
rect 9585 162713 9593 165697
rect 12577 162713 12585 165697
rect 9585 162705 12585 162713
rect 12775 165697 15775 165705
rect 12775 162713 12783 165697
rect 15767 162713 15775 165697
rect 12775 162705 15775 162713
rect 15965 165697 18965 165705
rect 15965 162713 15973 165697
rect 18957 162713 18965 165697
rect 15965 162705 18965 162713
rect 19155 165697 22155 165705
rect 19155 162713 19163 165697
rect 22147 162713 22155 165697
rect 19155 162705 22155 162713
rect 22345 165697 25345 165705
rect 22345 162713 22353 165697
rect 25337 162713 25345 165697
rect 22345 162705 25345 162713
rect 25535 165697 28535 165705
rect 25535 162713 25543 165697
rect 28527 162713 28535 165697
rect 25535 162705 28535 162713
rect 28725 165697 31725 165705
rect 28725 162713 28733 165697
rect 31717 162713 31725 165697
rect 28725 162705 31725 162713
rect 31915 165697 34915 165705
rect 31915 162713 31923 165697
rect 34907 162713 34915 165697
rect 31915 162705 34915 162713
rect 35105 165697 38105 165705
rect 35105 162713 35113 165697
rect 38097 162713 38105 165697
rect 35105 162705 38105 162713
rect 38295 165697 41295 165705
rect 38295 162713 38303 165697
rect 41287 162713 41295 165697
rect 38295 162705 41295 162713
rect 41485 165697 44485 165705
rect 41485 162713 41493 165697
rect 44477 162713 44485 165697
rect 41485 162705 44485 162713
rect 44675 165697 47675 165705
rect 44675 162713 44683 165697
rect 47667 162713 47675 165697
rect 44675 162705 47675 162713
rect 47865 165697 50865 165705
rect 47865 162713 47873 165697
rect 50857 162713 50865 165697
rect 47865 162705 50865 162713
rect 51055 165697 54055 165705
rect 51055 162713 51063 165697
rect 54047 162713 54055 165697
rect 51055 162705 54055 162713
rect 54245 165697 57245 165705
rect 54245 162713 54253 165697
rect 57237 162713 57245 165697
rect 54245 162705 57245 162713
rect 57435 165697 60435 165705
rect 57435 162713 57443 165697
rect 60427 162713 60435 165697
rect 57435 162705 60435 162713
rect 60625 165697 63625 165705
rect 60625 162713 60633 165697
rect 63617 162713 63625 165697
rect 60625 162705 63625 162713
rect 63815 165697 66815 165705
rect 63815 162713 63823 165697
rect 66807 162713 66815 165697
rect 63815 162705 66815 162713
rect 67005 165697 70005 165705
rect 67005 162713 67013 165697
rect 69997 162713 70005 165697
rect 67005 162705 70005 162713
rect 70195 165697 73195 165705
rect 70195 162713 70203 165697
rect 73187 162713 73195 165697
rect 70195 162705 73195 162713
rect 73385 165697 76385 165705
rect 73385 162713 73393 165697
rect 76377 162713 76385 165697
rect 73385 162705 76385 162713
rect 76575 165697 79575 165705
rect 76575 162713 76583 165697
rect 79567 162713 79575 165697
rect 76575 162705 79575 162713
rect 79765 165697 82765 165705
rect 79765 162713 79773 165697
rect 82757 162713 82765 165697
rect 79765 162705 82765 162713
rect 82955 165697 85955 165705
rect 82955 162713 82963 165697
rect 85947 162713 85955 165697
rect 82955 162705 85955 162713
rect 86145 165697 89145 165705
rect 86145 162713 86153 165697
rect 89137 162713 89145 165697
rect 86145 162705 89145 162713
rect 89335 165697 92335 165705
rect 89335 162713 89343 165697
rect 92327 162713 92335 165697
rect 89335 162705 92335 162713
rect 92525 165697 95525 165705
rect 92525 162713 92533 165697
rect 95517 162713 95525 165697
rect 92525 162705 95525 162713
rect 95715 165697 98715 165705
rect 95715 162713 95723 165697
rect 98707 162713 98715 165697
rect 95715 162705 98715 162713
rect 98905 165697 101905 165705
rect 98905 162713 98913 165697
rect 101897 162713 101905 165697
rect 98905 162705 101905 162713
rect 102095 165697 105095 165705
rect 102095 162713 102103 165697
rect 105087 162713 105095 165697
rect 102095 162705 105095 162713
rect 105285 165697 108285 165705
rect 105285 162713 105293 165697
rect 108277 162713 108285 165697
rect 105285 162705 108285 162713
rect 108475 165697 111475 165705
rect 108475 162713 108483 165697
rect 111467 162713 111475 165697
rect 108475 162705 111475 162713
rect 111665 165697 114665 165705
rect 111665 162713 111673 165697
rect 114657 162713 114665 165697
rect 111665 162705 114665 162713
rect 114855 165697 117855 165705
rect 114855 162713 114863 165697
rect 117847 162713 117855 165697
rect 114855 162705 117855 162713
rect 118045 165697 121045 165705
rect 118045 162713 118053 165697
rect 121037 162713 121045 165697
rect 118045 162705 121045 162713
rect 121235 165697 124235 165705
rect 121235 162713 121243 165697
rect 124227 162713 124235 165697
rect 121235 162705 124235 162713
rect 124425 165697 127425 165705
rect 124425 162713 124433 165697
rect 127417 162713 127425 165697
rect 124425 162705 127425 162713
rect 127615 165697 130615 165705
rect 127615 162713 127623 165697
rect 130607 162713 130615 165697
rect 127615 162705 130615 162713
rect 130805 165697 133805 165705
rect 130805 162713 130813 165697
rect 133797 162713 133805 165697
rect 130805 162705 133805 162713
rect 133995 165697 136995 165705
rect 133995 162713 134003 165697
rect 136987 162713 136995 165697
rect 133995 162705 136995 162713
rect 15 162507 3015 162515
rect 15 159523 23 162507
rect 3007 159523 3015 162507
rect 15 159515 3015 159523
rect 3205 162507 6205 162515
rect 3205 159523 3213 162507
rect 6197 159523 6205 162507
rect 3205 159515 6205 159523
rect 6395 162507 9395 162515
rect 6395 159523 6403 162507
rect 9387 159523 9395 162507
rect 6395 159515 9395 159523
rect 9585 162507 12585 162515
rect 9585 159523 9593 162507
rect 12577 159523 12585 162507
rect 9585 159515 12585 159523
rect 12775 162507 15775 162515
rect 12775 159523 12783 162507
rect 15767 159523 15775 162507
rect 12775 159515 15775 159523
rect 15965 162507 18965 162515
rect 15965 159523 15973 162507
rect 18957 159523 18965 162507
rect 15965 159515 18965 159523
rect 19155 162507 22155 162515
rect 19155 159523 19163 162507
rect 22147 159523 22155 162507
rect 19155 159515 22155 159523
rect 22345 162507 25345 162515
rect 22345 159523 22353 162507
rect 25337 159523 25345 162507
rect 22345 159515 25345 159523
rect 25535 162507 28535 162515
rect 25535 159523 25543 162507
rect 28527 159523 28535 162507
rect 25535 159515 28535 159523
rect 28725 162507 31725 162515
rect 28725 159523 28733 162507
rect 31717 159523 31725 162507
rect 28725 159515 31725 159523
rect 31915 162507 34915 162515
rect 31915 159523 31923 162507
rect 34907 159523 34915 162507
rect 31915 159515 34915 159523
rect 35105 162507 38105 162515
rect 35105 159523 35113 162507
rect 38097 159523 38105 162507
rect 35105 159515 38105 159523
rect 38295 162507 41295 162515
rect 38295 159523 38303 162507
rect 41287 159523 41295 162507
rect 38295 159515 41295 159523
rect 41485 162507 44485 162515
rect 41485 159523 41493 162507
rect 44477 159523 44485 162507
rect 41485 159515 44485 159523
rect 44675 162507 47675 162515
rect 44675 159523 44683 162507
rect 47667 159523 47675 162507
rect 44675 159515 47675 159523
rect 47865 162507 50865 162515
rect 47865 159523 47873 162507
rect 50857 159523 50865 162507
rect 47865 159515 50865 159523
rect 51055 162507 54055 162515
rect 51055 159523 51063 162507
rect 54047 159523 54055 162507
rect 51055 159515 54055 159523
rect 54245 162507 57245 162515
rect 54245 159523 54253 162507
rect 57237 159523 57245 162507
rect 54245 159515 57245 159523
rect 57435 162507 60435 162515
rect 57435 159523 57443 162507
rect 60427 159523 60435 162507
rect 57435 159515 60435 159523
rect 60625 162507 63625 162515
rect 60625 159523 60633 162507
rect 63617 159523 63625 162507
rect 60625 159515 63625 159523
rect 63815 162507 66815 162515
rect 63815 159523 63823 162507
rect 66807 159523 66815 162507
rect 63815 159515 66815 159523
rect 67005 162507 70005 162515
rect 67005 159523 67013 162507
rect 69997 159523 70005 162507
rect 67005 159515 70005 159523
rect 70195 162507 73195 162515
rect 70195 159523 70203 162507
rect 73187 159523 73195 162507
rect 70195 159515 73195 159523
rect 73385 162507 76385 162515
rect 73385 159523 73393 162507
rect 76377 159523 76385 162507
rect 73385 159515 76385 159523
rect 76575 162507 79575 162515
rect 76575 159523 76583 162507
rect 79567 159523 79575 162507
rect 76575 159515 79575 159523
rect 79765 162507 82765 162515
rect 79765 159523 79773 162507
rect 82757 159523 82765 162507
rect 79765 159515 82765 159523
rect 82955 162507 85955 162515
rect 82955 159523 82963 162507
rect 85947 159523 85955 162507
rect 82955 159515 85955 159523
rect 86145 162507 89145 162515
rect 86145 159523 86153 162507
rect 89137 159523 89145 162507
rect 86145 159515 89145 159523
rect 89335 162507 92335 162515
rect 89335 159523 89343 162507
rect 92327 159523 92335 162507
rect 89335 159515 92335 159523
rect 92525 162507 95525 162515
rect 92525 159523 92533 162507
rect 95517 159523 95525 162507
rect 92525 159515 95525 159523
rect 95715 162507 98715 162515
rect 95715 159523 95723 162507
rect 98707 159523 98715 162507
rect 95715 159515 98715 159523
rect 98905 162507 101905 162515
rect 98905 159523 98913 162507
rect 101897 159523 101905 162507
rect 98905 159515 101905 159523
rect 102095 162507 105095 162515
rect 102095 159523 102103 162507
rect 105087 159523 105095 162507
rect 102095 159515 105095 159523
rect 105285 162507 108285 162515
rect 105285 159523 105293 162507
rect 108277 159523 108285 162507
rect 105285 159515 108285 159523
rect 108475 162507 111475 162515
rect 108475 159523 108483 162507
rect 111467 159523 111475 162507
rect 108475 159515 111475 159523
rect 111665 162507 114665 162515
rect 111665 159523 111673 162507
rect 114657 159523 114665 162507
rect 111665 159515 114665 159523
rect 114855 162507 117855 162515
rect 114855 159523 114863 162507
rect 117847 159523 117855 162507
rect 114855 159515 117855 159523
rect 118045 162507 121045 162515
rect 118045 159523 118053 162507
rect 121037 159523 121045 162507
rect 118045 159515 121045 159523
rect 121235 162507 124235 162515
rect 121235 159523 121243 162507
rect 124227 159523 124235 162507
rect 121235 159515 124235 159523
rect 124425 162507 127425 162515
rect 124425 159523 124433 162507
rect 127417 159523 127425 162507
rect 124425 159515 127425 159523
rect 127615 162507 130615 162515
rect 127615 159523 127623 162507
rect 130607 159523 130615 162507
rect 127615 159515 130615 159523
rect 130805 162507 133805 162515
rect 130805 159523 130813 162507
rect 133797 159523 133805 162507
rect 130805 159515 133805 159523
rect 133995 162507 136995 162515
rect 133995 159523 134003 162507
rect 136987 159523 136995 162507
rect 133995 159515 136995 159523
rect 15 159317 3015 159325
rect 15 156333 23 159317
rect 3007 156333 3015 159317
rect 15 156325 3015 156333
rect 3205 159317 6205 159325
rect 3205 156333 3213 159317
rect 6197 156333 6205 159317
rect 3205 156325 6205 156333
rect 6395 159317 9395 159325
rect 6395 156333 6403 159317
rect 9387 156333 9395 159317
rect 6395 156325 9395 156333
rect 9585 159317 12585 159325
rect 9585 156333 9593 159317
rect 12577 156333 12585 159317
rect 9585 156325 12585 156333
rect 12775 159317 15775 159325
rect 12775 156333 12783 159317
rect 15767 156333 15775 159317
rect 12775 156325 15775 156333
rect 15965 159317 18965 159325
rect 15965 156333 15973 159317
rect 18957 156333 18965 159317
rect 15965 156325 18965 156333
rect 19155 159317 22155 159325
rect 19155 156333 19163 159317
rect 22147 156333 22155 159317
rect 19155 156325 22155 156333
rect 22345 159317 25345 159325
rect 22345 156333 22353 159317
rect 25337 156333 25345 159317
rect 22345 156325 25345 156333
rect 25535 159317 28535 159325
rect 25535 156333 25543 159317
rect 28527 156333 28535 159317
rect 25535 156325 28535 156333
rect 28725 159317 31725 159325
rect 28725 156333 28733 159317
rect 31717 156333 31725 159317
rect 28725 156325 31725 156333
rect 31915 159317 34915 159325
rect 31915 156333 31923 159317
rect 34907 156333 34915 159317
rect 31915 156325 34915 156333
rect 35105 159317 38105 159325
rect 35105 156333 35113 159317
rect 38097 156333 38105 159317
rect 35105 156325 38105 156333
rect 38295 159317 41295 159325
rect 38295 156333 38303 159317
rect 41287 156333 41295 159317
rect 38295 156325 41295 156333
rect 41485 159317 44485 159325
rect 41485 156333 41493 159317
rect 44477 156333 44485 159317
rect 41485 156325 44485 156333
rect 44675 159317 47675 159325
rect 44675 156333 44683 159317
rect 47667 156333 47675 159317
rect 44675 156325 47675 156333
rect 47865 159317 50865 159325
rect 47865 156333 47873 159317
rect 50857 156333 50865 159317
rect 47865 156325 50865 156333
rect 51055 159317 54055 159325
rect 51055 156333 51063 159317
rect 54047 156333 54055 159317
rect 51055 156325 54055 156333
rect 54245 159317 57245 159325
rect 54245 156333 54253 159317
rect 57237 156333 57245 159317
rect 54245 156325 57245 156333
rect 57435 159317 60435 159325
rect 57435 156333 57443 159317
rect 60427 156333 60435 159317
rect 57435 156325 60435 156333
rect 60625 159317 63625 159325
rect 60625 156333 60633 159317
rect 63617 156333 63625 159317
rect 60625 156325 63625 156333
rect 63815 159317 66815 159325
rect 63815 156333 63823 159317
rect 66807 156333 66815 159317
rect 63815 156325 66815 156333
rect 67005 159317 70005 159325
rect 67005 156333 67013 159317
rect 69997 156333 70005 159317
rect 67005 156325 70005 156333
rect 70195 159317 73195 159325
rect 70195 156333 70203 159317
rect 73187 156333 73195 159317
rect 70195 156325 73195 156333
rect 73385 159317 76385 159325
rect 73385 156333 73393 159317
rect 76377 156333 76385 159317
rect 73385 156325 76385 156333
rect 76575 159317 79575 159325
rect 76575 156333 76583 159317
rect 79567 156333 79575 159317
rect 76575 156325 79575 156333
rect 79765 159317 82765 159325
rect 79765 156333 79773 159317
rect 82757 156333 82765 159317
rect 79765 156325 82765 156333
rect 82955 159317 85955 159325
rect 82955 156333 82963 159317
rect 85947 156333 85955 159317
rect 82955 156325 85955 156333
rect 86145 159317 89145 159325
rect 86145 156333 86153 159317
rect 89137 156333 89145 159317
rect 86145 156325 89145 156333
rect 89335 159317 92335 159325
rect 89335 156333 89343 159317
rect 92327 156333 92335 159317
rect 89335 156325 92335 156333
rect 92525 159317 95525 159325
rect 92525 156333 92533 159317
rect 95517 156333 95525 159317
rect 92525 156325 95525 156333
rect 95715 159317 98715 159325
rect 95715 156333 95723 159317
rect 98707 156333 98715 159317
rect 95715 156325 98715 156333
rect 98905 159317 101905 159325
rect 98905 156333 98913 159317
rect 101897 156333 101905 159317
rect 98905 156325 101905 156333
rect 102095 159317 105095 159325
rect 102095 156333 102103 159317
rect 105087 156333 105095 159317
rect 102095 156325 105095 156333
rect 105285 159317 108285 159325
rect 105285 156333 105293 159317
rect 108277 156333 108285 159317
rect 105285 156325 108285 156333
rect 108475 159317 111475 159325
rect 108475 156333 108483 159317
rect 111467 156333 111475 159317
rect 108475 156325 111475 156333
rect 111665 159317 114665 159325
rect 111665 156333 111673 159317
rect 114657 156333 114665 159317
rect 111665 156325 114665 156333
rect 114855 159317 117855 159325
rect 114855 156333 114863 159317
rect 117847 156333 117855 159317
rect 114855 156325 117855 156333
rect 118045 159317 121045 159325
rect 118045 156333 118053 159317
rect 121037 156333 121045 159317
rect 118045 156325 121045 156333
rect 121235 159317 124235 159325
rect 121235 156333 121243 159317
rect 124227 156333 124235 159317
rect 121235 156325 124235 156333
rect 124425 159317 127425 159325
rect 124425 156333 124433 159317
rect 127417 156333 127425 159317
rect 124425 156325 127425 156333
rect 127615 159317 130615 159325
rect 127615 156333 127623 159317
rect 130607 156333 130615 159317
rect 127615 156325 130615 156333
rect 130805 159317 133805 159325
rect 130805 156333 130813 159317
rect 133797 156333 133805 159317
rect 130805 156325 133805 156333
rect 133995 159317 136995 159325
rect 133995 156333 134003 159317
rect 136987 156333 136995 159317
rect 133995 156325 136995 156333
rect 15 156127 3015 156135
rect 15 153143 23 156127
rect 3007 153143 3015 156127
rect 15 153135 3015 153143
rect 3205 156127 6205 156135
rect 3205 153143 3213 156127
rect 6197 153143 6205 156127
rect 3205 153135 6205 153143
rect 6395 156127 9395 156135
rect 6395 153143 6403 156127
rect 9387 153143 9395 156127
rect 6395 153135 9395 153143
rect 9585 156127 12585 156135
rect 9585 153143 9593 156127
rect 12577 153143 12585 156127
rect 9585 153135 12585 153143
rect 12775 156127 15775 156135
rect 12775 153143 12783 156127
rect 15767 153143 15775 156127
rect 12775 153135 15775 153143
rect 15965 156127 18965 156135
rect 15965 153143 15973 156127
rect 18957 153143 18965 156127
rect 15965 153135 18965 153143
rect 19155 156127 22155 156135
rect 19155 153143 19163 156127
rect 22147 153143 22155 156127
rect 19155 153135 22155 153143
rect 22345 156127 25345 156135
rect 22345 153143 22353 156127
rect 25337 153143 25345 156127
rect 22345 153135 25345 153143
rect 25535 156127 28535 156135
rect 25535 153143 25543 156127
rect 28527 153143 28535 156127
rect 25535 153135 28535 153143
rect 28725 156127 31725 156135
rect 28725 153143 28733 156127
rect 31717 153143 31725 156127
rect 28725 153135 31725 153143
rect 31915 156127 34915 156135
rect 31915 153143 31923 156127
rect 34907 153143 34915 156127
rect 31915 153135 34915 153143
rect 35105 156127 38105 156135
rect 35105 153143 35113 156127
rect 38097 153143 38105 156127
rect 35105 153135 38105 153143
rect 38295 156127 41295 156135
rect 38295 153143 38303 156127
rect 41287 153143 41295 156127
rect 38295 153135 41295 153143
rect 41485 156127 44485 156135
rect 41485 153143 41493 156127
rect 44477 153143 44485 156127
rect 41485 153135 44485 153143
rect 44675 156127 47675 156135
rect 44675 153143 44683 156127
rect 47667 153143 47675 156127
rect 44675 153135 47675 153143
rect 47865 156127 50865 156135
rect 47865 153143 47873 156127
rect 50857 153143 50865 156127
rect 47865 153135 50865 153143
rect 51055 156127 54055 156135
rect 51055 153143 51063 156127
rect 54047 153143 54055 156127
rect 51055 153135 54055 153143
rect 54245 156127 57245 156135
rect 54245 153143 54253 156127
rect 57237 153143 57245 156127
rect 54245 153135 57245 153143
rect 57435 156127 60435 156135
rect 57435 153143 57443 156127
rect 60427 153143 60435 156127
rect 57435 153135 60435 153143
rect 60625 156127 63625 156135
rect 60625 153143 60633 156127
rect 63617 153143 63625 156127
rect 60625 153135 63625 153143
rect 63815 156127 66815 156135
rect 63815 153143 63823 156127
rect 66807 153143 66815 156127
rect 63815 153135 66815 153143
rect 67005 156127 70005 156135
rect 67005 153143 67013 156127
rect 69997 153143 70005 156127
rect 67005 153135 70005 153143
rect 70195 156127 73195 156135
rect 70195 153143 70203 156127
rect 73187 153143 73195 156127
rect 70195 153135 73195 153143
rect 73385 156127 76385 156135
rect 73385 153143 73393 156127
rect 76377 153143 76385 156127
rect 73385 153135 76385 153143
rect 76575 156127 79575 156135
rect 76575 153143 76583 156127
rect 79567 153143 79575 156127
rect 76575 153135 79575 153143
rect 79765 156127 82765 156135
rect 79765 153143 79773 156127
rect 82757 153143 82765 156127
rect 79765 153135 82765 153143
rect 82955 156127 85955 156135
rect 82955 153143 82963 156127
rect 85947 153143 85955 156127
rect 82955 153135 85955 153143
rect 86145 156127 89145 156135
rect 86145 153143 86153 156127
rect 89137 153143 89145 156127
rect 86145 153135 89145 153143
rect 89335 156127 92335 156135
rect 89335 153143 89343 156127
rect 92327 153143 92335 156127
rect 89335 153135 92335 153143
rect 92525 156127 95525 156135
rect 92525 153143 92533 156127
rect 95517 153143 95525 156127
rect 92525 153135 95525 153143
rect 95715 156127 98715 156135
rect 95715 153143 95723 156127
rect 98707 153143 98715 156127
rect 95715 153135 98715 153143
rect 98905 156127 101905 156135
rect 98905 153143 98913 156127
rect 101897 153143 101905 156127
rect 98905 153135 101905 153143
rect 102095 156127 105095 156135
rect 102095 153143 102103 156127
rect 105087 153143 105095 156127
rect 102095 153135 105095 153143
rect 105285 156127 108285 156135
rect 105285 153143 105293 156127
rect 108277 153143 108285 156127
rect 105285 153135 108285 153143
rect 108475 156127 111475 156135
rect 108475 153143 108483 156127
rect 111467 153143 111475 156127
rect 108475 153135 111475 153143
rect 111665 156127 114665 156135
rect 111665 153143 111673 156127
rect 114657 153143 114665 156127
rect 111665 153135 114665 153143
rect 114855 156127 117855 156135
rect 114855 153143 114863 156127
rect 117847 153143 117855 156127
rect 114855 153135 117855 153143
rect 118045 156127 121045 156135
rect 118045 153143 118053 156127
rect 121037 153143 121045 156127
rect 118045 153135 121045 153143
rect 121235 156127 124235 156135
rect 121235 153143 121243 156127
rect 124227 153143 124235 156127
rect 121235 153135 124235 153143
rect 124425 156127 127425 156135
rect 124425 153143 124433 156127
rect 127417 153143 127425 156127
rect 124425 153135 127425 153143
rect 127615 156127 130615 156135
rect 127615 153143 127623 156127
rect 130607 153143 130615 156127
rect 127615 153135 130615 153143
rect 130805 156127 133805 156135
rect 130805 153143 130813 156127
rect 133797 153143 133805 156127
rect 130805 153135 133805 153143
rect 133995 156127 136995 156135
rect 133995 153143 134003 156127
rect 136987 153143 136995 156127
rect 133995 153135 136995 153143
rect 15 152937 3015 152945
rect 15 149953 23 152937
rect 3007 149953 3015 152937
rect 15 149945 3015 149953
rect 3205 152937 6205 152945
rect 3205 149953 3213 152937
rect 6197 149953 6205 152937
rect 3205 149945 6205 149953
rect 6395 152937 9395 152945
rect 6395 149953 6403 152937
rect 9387 149953 9395 152937
rect 6395 149945 9395 149953
rect 9585 152937 12585 152945
rect 9585 149953 9593 152937
rect 12577 149953 12585 152937
rect 9585 149945 12585 149953
rect 12775 152937 15775 152945
rect 12775 149953 12783 152937
rect 15767 149953 15775 152937
rect 12775 149945 15775 149953
rect 15965 152937 18965 152945
rect 15965 149953 15973 152937
rect 18957 149953 18965 152937
rect 15965 149945 18965 149953
rect 19155 152937 22155 152945
rect 19155 149953 19163 152937
rect 22147 149953 22155 152937
rect 19155 149945 22155 149953
rect 22345 152937 25345 152945
rect 22345 149953 22353 152937
rect 25337 149953 25345 152937
rect 22345 149945 25345 149953
rect 25535 152937 28535 152945
rect 25535 149953 25543 152937
rect 28527 149953 28535 152937
rect 25535 149945 28535 149953
rect 28725 152937 31725 152945
rect 28725 149953 28733 152937
rect 31717 149953 31725 152937
rect 28725 149945 31725 149953
rect 31915 152937 34915 152945
rect 31915 149953 31923 152937
rect 34907 149953 34915 152937
rect 31915 149945 34915 149953
rect 35105 152937 38105 152945
rect 35105 149953 35113 152937
rect 38097 149953 38105 152937
rect 35105 149945 38105 149953
rect 38295 152937 41295 152945
rect 38295 149953 38303 152937
rect 41287 149953 41295 152937
rect 38295 149945 41295 149953
rect 41485 152937 44485 152945
rect 41485 149953 41493 152937
rect 44477 149953 44485 152937
rect 41485 149945 44485 149953
rect 44675 152937 47675 152945
rect 44675 149953 44683 152937
rect 47667 149953 47675 152937
rect 44675 149945 47675 149953
rect 47865 152937 50865 152945
rect 47865 149953 47873 152937
rect 50857 149953 50865 152937
rect 47865 149945 50865 149953
rect 51055 152937 54055 152945
rect 51055 149953 51063 152937
rect 54047 149953 54055 152937
rect 51055 149945 54055 149953
rect 54245 152937 57245 152945
rect 54245 149953 54253 152937
rect 57237 149953 57245 152937
rect 54245 149945 57245 149953
rect 57435 152937 60435 152945
rect 57435 149953 57443 152937
rect 60427 149953 60435 152937
rect 57435 149945 60435 149953
rect 60625 152937 63625 152945
rect 60625 149953 60633 152937
rect 63617 149953 63625 152937
rect 60625 149945 63625 149953
rect 63815 152937 66815 152945
rect 63815 149953 63823 152937
rect 66807 149953 66815 152937
rect 63815 149945 66815 149953
rect 67005 152937 70005 152945
rect 67005 149953 67013 152937
rect 69997 149953 70005 152937
rect 67005 149945 70005 149953
rect 70195 152937 73195 152945
rect 70195 149953 70203 152937
rect 73187 149953 73195 152937
rect 70195 149945 73195 149953
rect 73385 152937 76385 152945
rect 73385 149953 73393 152937
rect 76377 149953 76385 152937
rect 73385 149945 76385 149953
rect 76575 152937 79575 152945
rect 76575 149953 76583 152937
rect 79567 149953 79575 152937
rect 76575 149945 79575 149953
rect 79765 152937 82765 152945
rect 79765 149953 79773 152937
rect 82757 149953 82765 152937
rect 79765 149945 82765 149953
rect 82955 152937 85955 152945
rect 82955 149953 82963 152937
rect 85947 149953 85955 152937
rect 82955 149945 85955 149953
rect 86145 152937 89145 152945
rect 86145 149953 86153 152937
rect 89137 149953 89145 152937
rect 86145 149945 89145 149953
rect 89335 152937 92335 152945
rect 89335 149953 89343 152937
rect 92327 149953 92335 152937
rect 89335 149945 92335 149953
rect 92525 152937 95525 152945
rect 92525 149953 92533 152937
rect 95517 149953 95525 152937
rect 92525 149945 95525 149953
rect 95715 152937 98715 152945
rect 95715 149953 95723 152937
rect 98707 149953 98715 152937
rect 95715 149945 98715 149953
rect 98905 152937 101905 152945
rect 98905 149953 98913 152937
rect 101897 149953 101905 152937
rect 98905 149945 101905 149953
rect 102095 152937 105095 152945
rect 102095 149953 102103 152937
rect 105087 149953 105095 152937
rect 102095 149945 105095 149953
rect 105285 152937 108285 152945
rect 105285 149953 105293 152937
rect 108277 149953 108285 152937
rect 105285 149945 108285 149953
rect 108475 152937 111475 152945
rect 108475 149953 108483 152937
rect 111467 149953 111475 152937
rect 108475 149945 111475 149953
rect 111665 152937 114665 152945
rect 111665 149953 111673 152937
rect 114657 149953 114665 152937
rect 111665 149945 114665 149953
rect 114855 152937 117855 152945
rect 114855 149953 114863 152937
rect 117847 149953 117855 152937
rect 114855 149945 117855 149953
rect 118045 152937 121045 152945
rect 118045 149953 118053 152937
rect 121037 149953 121045 152937
rect 118045 149945 121045 149953
rect 121235 152937 124235 152945
rect 121235 149953 121243 152937
rect 124227 149953 124235 152937
rect 121235 149945 124235 149953
rect 124425 152937 127425 152945
rect 124425 149953 124433 152937
rect 127417 149953 127425 152937
rect 124425 149945 127425 149953
rect 127615 152937 130615 152945
rect 127615 149953 127623 152937
rect 130607 149953 130615 152937
rect 127615 149945 130615 149953
rect 130805 152937 133805 152945
rect 130805 149953 130813 152937
rect 133797 149953 133805 152937
rect 130805 149945 133805 149953
rect 133995 152937 136995 152945
rect 133995 149953 134003 152937
rect 136987 149953 136995 152937
rect 133995 149945 136995 149953
rect 15 149747 3015 149755
rect 15 146763 23 149747
rect 3007 146763 3015 149747
rect 15 146755 3015 146763
rect 3205 149747 6205 149755
rect 3205 146763 3213 149747
rect 6197 146763 6205 149747
rect 3205 146755 6205 146763
rect 6395 149747 9395 149755
rect 6395 146763 6403 149747
rect 9387 146763 9395 149747
rect 6395 146755 9395 146763
rect 9585 149747 12585 149755
rect 9585 146763 9593 149747
rect 12577 146763 12585 149747
rect 9585 146755 12585 146763
rect 12775 149747 15775 149755
rect 12775 146763 12783 149747
rect 15767 146763 15775 149747
rect 12775 146755 15775 146763
rect 15965 149747 18965 149755
rect 15965 146763 15973 149747
rect 18957 146763 18965 149747
rect 15965 146755 18965 146763
rect 19155 149747 22155 149755
rect 19155 146763 19163 149747
rect 22147 146763 22155 149747
rect 19155 146755 22155 146763
rect 22345 149747 25345 149755
rect 22345 146763 22353 149747
rect 25337 146763 25345 149747
rect 22345 146755 25345 146763
rect 25535 149747 28535 149755
rect 25535 146763 25543 149747
rect 28527 146763 28535 149747
rect 25535 146755 28535 146763
rect 28725 149747 31725 149755
rect 28725 146763 28733 149747
rect 31717 146763 31725 149747
rect 28725 146755 31725 146763
rect 31915 149747 34915 149755
rect 31915 146763 31923 149747
rect 34907 146763 34915 149747
rect 31915 146755 34915 146763
rect 35105 149747 38105 149755
rect 35105 146763 35113 149747
rect 38097 146763 38105 149747
rect 35105 146755 38105 146763
rect 38295 149747 41295 149755
rect 38295 146763 38303 149747
rect 41287 146763 41295 149747
rect 38295 146755 41295 146763
rect 41485 149747 44485 149755
rect 41485 146763 41493 149747
rect 44477 146763 44485 149747
rect 41485 146755 44485 146763
rect 44675 149747 47675 149755
rect 44675 146763 44683 149747
rect 47667 146763 47675 149747
rect 44675 146755 47675 146763
rect 47865 149747 50865 149755
rect 47865 146763 47873 149747
rect 50857 146763 50865 149747
rect 47865 146755 50865 146763
rect 51055 149747 54055 149755
rect 51055 146763 51063 149747
rect 54047 146763 54055 149747
rect 51055 146755 54055 146763
rect 54245 149747 57245 149755
rect 54245 146763 54253 149747
rect 57237 146763 57245 149747
rect 54245 146755 57245 146763
rect 57435 149747 60435 149755
rect 57435 146763 57443 149747
rect 60427 146763 60435 149747
rect 57435 146755 60435 146763
rect 60625 149747 63625 149755
rect 60625 146763 60633 149747
rect 63617 146763 63625 149747
rect 60625 146755 63625 146763
rect 63815 149747 66815 149755
rect 63815 146763 63823 149747
rect 66807 146763 66815 149747
rect 63815 146755 66815 146763
rect 67005 149747 70005 149755
rect 67005 146763 67013 149747
rect 69997 146763 70005 149747
rect 67005 146755 70005 146763
rect 70195 149747 73195 149755
rect 70195 146763 70203 149747
rect 73187 146763 73195 149747
rect 70195 146755 73195 146763
rect 73385 149747 76385 149755
rect 73385 146763 73393 149747
rect 76377 146763 76385 149747
rect 73385 146755 76385 146763
rect 76575 149747 79575 149755
rect 76575 146763 76583 149747
rect 79567 146763 79575 149747
rect 76575 146755 79575 146763
rect 79765 149747 82765 149755
rect 79765 146763 79773 149747
rect 82757 146763 82765 149747
rect 79765 146755 82765 146763
rect 82955 149747 85955 149755
rect 82955 146763 82963 149747
rect 85947 146763 85955 149747
rect 82955 146755 85955 146763
rect 86145 149747 89145 149755
rect 86145 146763 86153 149747
rect 89137 146763 89145 149747
rect 86145 146755 89145 146763
rect 89335 149747 92335 149755
rect 89335 146763 89343 149747
rect 92327 146763 92335 149747
rect 89335 146755 92335 146763
rect 92525 149747 95525 149755
rect 92525 146763 92533 149747
rect 95517 146763 95525 149747
rect 92525 146755 95525 146763
rect 95715 149747 98715 149755
rect 95715 146763 95723 149747
rect 98707 146763 98715 149747
rect 95715 146755 98715 146763
rect 98905 149747 101905 149755
rect 98905 146763 98913 149747
rect 101897 146763 101905 149747
rect 98905 146755 101905 146763
rect 102095 149747 105095 149755
rect 102095 146763 102103 149747
rect 105087 146763 105095 149747
rect 102095 146755 105095 146763
rect 105285 149747 108285 149755
rect 105285 146763 105293 149747
rect 108277 146763 108285 149747
rect 105285 146755 108285 146763
rect 108475 149747 111475 149755
rect 108475 146763 108483 149747
rect 111467 146763 111475 149747
rect 108475 146755 111475 146763
rect 111665 149747 114665 149755
rect 111665 146763 111673 149747
rect 114657 146763 114665 149747
rect 111665 146755 114665 146763
rect 114855 149747 117855 149755
rect 114855 146763 114863 149747
rect 117847 146763 117855 149747
rect 114855 146755 117855 146763
rect 118045 149747 121045 149755
rect 118045 146763 118053 149747
rect 121037 146763 121045 149747
rect 118045 146755 121045 146763
rect 121235 149747 124235 149755
rect 121235 146763 121243 149747
rect 124227 146763 124235 149747
rect 121235 146755 124235 146763
rect 124425 149747 127425 149755
rect 124425 146763 124433 149747
rect 127417 146763 127425 149747
rect 124425 146755 127425 146763
rect 127615 149747 130615 149755
rect 127615 146763 127623 149747
rect 130607 146763 130615 149747
rect 127615 146755 130615 146763
rect 130805 149747 133805 149755
rect 130805 146763 130813 149747
rect 133797 146763 133805 149747
rect 130805 146755 133805 146763
rect 133995 149747 136995 149755
rect 133995 146763 134003 149747
rect 136987 146763 136995 149747
rect 133995 146755 136995 146763
rect 15 146557 3015 146565
rect 15 143573 23 146557
rect 3007 143573 3015 146557
rect 15 143565 3015 143573
rect 3205 146557 6205 146565
rect 3205 143573 3213 146557
rect 6197 143573 6205 146557
rect 3205 143565 6205 143573
rect 6395 146557 9395 146565
rect 6395 143573 6403 146557
rect 9387 143573 9395 146557
rect 6395 143565 9395 143573
rect 9585 146557 12585 146565
rect 9585 143573 9593 146557
rect 12577 143573 12585 146557
rect 9585 143565 12585 143573
rect 12775 146557 15775 146565
rect 12775 143573 12783 146557
rect 15767 143573 15775 146557
rect 12775 143565 15775 143573
rect 15965 146557 18965 146565
rect 15965 143573 15973 146557
rect 18957 143573 18965 146557
rect 15965 143565 18965 143573
rect 19155 146557 22155 146565
rect 19155 143573 19163 146557
rect 22147 143573 22155 146557
rect 19155 143565 22155 143573
rect 22345 146557 25345 146565
rect 22345 143573 22353 146557
rect 25337 143573 25345 146557
rect 22345 143565 25345 143573
rect 25535 146557 28535 146565
rect 25535 143573 25543 146557
rect 28527 143573 28535 146557
rect 25535 143565 28535 143573
rect 28725 146557 31725 146565
rect 28725 143573 28733 146557
rect 31717 143573 31725 146557
rect 28725 143565 31725 143573
rect 31915 146557 34915 146565
rect 31915 143573 31923 146557
rect 34907 143573 34915 146557
rect 31915 143565 34915 143573
rect 35105 146557 38105 146565
rect 35105 143573 35113 146557
rect 38097 143573 38105 146557
rect 35105 143565 38105 143573
rect 38295 146557 41295 146565
rect 38295 143573 38303 146557
rect 41287 143573 41295 146557
rect 38295 143565 41295 143573
rect 41485 146557 44485 146565
rect 41485 143573 41493 146557
rect 44477 143573 44485 146557
rect 41485 143565 44485 143573
rect 44675 146557 47675 146565
rect 44675 143573 44683 146557
rect 47667 143573 47675 146557
rect 44675 143565 47675 143573
rect 47865 146557 50865 146565
rect 47865 143573 47873 146557
rect 50857 143573 50865 146557
rect 47865 143565 50865 143573
rect 51055 146557 54055 146565
rect 51055 143573 51063 146557
rect 54047 143573 54055 146557
rect 51055 143565 54055 143573
rect 54245 146557 57245 146565
rect 54245 143573 54253 146557
rect 57237 143573 57245 146557
rect 54245 143565 57245 143573
rect 57435 146557 60435 146565
rect 57435 143573 57443 146557
rect 60427 143573 60435 146557
rect 57435 143565 60435 143573
rect 60625 146557 63625 146565
rect 60625 143573 60633 146557
rect 63617 143573 63625 146557
rect 60625 143565 63625 143573
rect 63815 146557 66815 146565
rect 63815 143573 63823 146557
rect 66807 143573 66815 146557
rect 63815 143565 66815 143573
rect 67005 146557 70005 146565
rect 67005 143573 67013 146557
rect 69997 143573 70005 146557
rect 67005 143565 70005 143573
rect 70195 146557 73195 146565
rect 70195 143573 70203 146557
rect 73187 143573 73195 146557
rect 70195 143565 73195 143573
rect 73385 146557 76385 146565
rect 73385 143573 73393 146557
rect 76377 143573 76385 146557
rect 73385 143565 76385 143573
rect 76575 146557 79575 146565
rect 76575 143573 76583 146557
rect 79567 143573 79575 146557
rect 76575 143565 79575 143573
rect 79765 146557 82765 146565
rect 79765 143573 79773 146557
rect 82757 143573 82765 146557
rect 79765 143565 82765 143573
rect 82955 146557 85955 146565
rect 82955 143573 82963 146557
rect 85947 143573 85955 146557
rect 82955 143565 85955 143573
rect 86145 146557 89145 146565
rect 86145 143573 86153 146557
rect 89137 143573 89145 146557
rect 86145 143565 89145 143573
rect 89335 146557 92335 146565
rect 89335 143573 89343 146557
rect 92327 143573 92335 146557
rect 89335 143565 92335 143573
rect 92525 146557 95525 146565
rect 92525 143573 92533 146557
rect 95517 143573 95525 146557
rect 92525 143565 95525 143573
rect 95715 146557 98715 146565
rect 95715 143573 95723 146557
rect 98707 143573 98715 146557
rect 95715 143565 98715 143573
rect 98905 146557 101905 146565
rect 98905 143573 98913 146557
rect 101897 143573 101905 146557
rect 98905 143565 101905 143573
rect 102095 146557 105095 146565
rect 102095 143573 102103 146557
rect 105087 143573 105095 146557
rect 102095 143565 105095 143573
rect 105285 146557 108285 146565
rect 105285 143573 105293 146557
rect 108277 143573 108285 146557
rect 105285 143565 108285 143573
rect 108475 146557 111475 146565
rect 108475 143573 108483 146557
rect 111467 143573 111475 146557
rect 108475 143565 111475 143573
rect 111665 146557 114665 146565
rect 111665 143573 111673 146557
rect 114657 143573 114665 146557
rect 111665 143565 114665 143573
rect 114855 146557 117855 146565
rect 114855 143573 114863 146557
rect 117847 143573 117855 146557
rect 114855 143565 117855 143573
rect 118045 146557 121045 146565
rect 118045 143573 118053 146557
rect 121037 143573 121045 146557
rect 118045 143565 121045 143573
rect 121235 146557 124235 146565
rect 121235 143573 121243 146557
rect 124227 143573 124235 146557
rect 121235 143565 124235 143573
rect 124425 146557 127425 146565
rect 124425 143573 124433 146557
rect 127417 143573 127425 146557
rect 124425 143565 127425 143573
rect 127615 146557 130615 146565
rect 127615 143573 127623 146557
rect 130607 143573 130615 146557
rect 127615 143565 130615 143573
rect 130805 146557 133805 146565
rect 130805 143573 130813 146557
rect 133797 143573 133805 146557
rect 130805 143565 133805 143573
rect 133995 146557 136995 146565
rect 133995 143573 134003 146557
rect 136987 143573 136995 146557
rect 133995 143565 136995 143573
rect 15 143367 3015 143375
rect 15 140383 23 143367
rect 3007 140383 3015 143367
rect 15 140375 3015 140383
rect 3205 143367 6205 143375
rect 3205 140383 3213 143367
rect 6197 140383 6205 143367
rect 3205 140375 6205 140383
rect 6395 143367 9395 143375
rect 6395 140383 6403 143367
rect 9387 140383 9395 143367
rect 6395 140375 9395 140383
rect 9585 143367 12585 143375
rect 9585 140383 9593 143367
rect 12577 140383 12585 143367
rect 9585 140375 12585 140383
rect 12775 143367 15775 143375
rect 12775 140383 12783 143367
rect 15767 140383 15775 143367
rect 12775 140375 15775 140383
rect 15965 143367 18965 143375
rect 15965 140383 15973 143367
rect 18957 140383 18965 143367
rect 15965 140375 18965 140383
rect 19155 143367 22155 143375
rect 19155 140383 19163 143367
rect 22147 140383 22155 143367
rect 19155 140375 22155 140383
rect 22345 143367 25345 143375
rect 22345 140383 22353 143367
rect 25337 140383 25345 143367
rect 22345 140375 25345 140383
rect 25535 143367 28535 143375
rect 25535 140383 25543 143367
rect 28527 140383 28535 143367
rect 25535 140375 28535 140383
rect 28725 143367 31725 143375
rect 28725 140383 28733 143367
rect 31717 140383 31725 143367
rect 28725 140375 31725 140383
rect 31915 143367 34915 143375
rect 31915 140383 31923 143367
rect 34907 140383 34915 143367
rect 31915 140375 34915 140383
rect 35105 143367 38105 143375
rect 35105 140383 35113 143367
rect 38097 140383 38105 143367
rect 35105 140375 38105 140383
rect 38295 143367 41295 143375
rect 38295 140383 38303 143367
rect 41287 140383 41295 143367
rect 38295 140375 41295 140383
rect 41485 143367 44485 143375
rect 41485 140383 41493 143367
rect 44477 140383 44485 143367
rect 41485 140375 44485 140383
rect 44675 143367 47675 143375
rect 44675 140383 44683 143367
rect 47667 140383 47675 143367
rect 44675 140375 47675 140383
rect 47865 143367 50865 143375
rect 47865 140383 47873 143367
rect 50857 140383 50865 143367
rect 47865 140375 50865 140383
rect 51055 143367 54055 143375
rect 51055 140383 51063 143367
rect 54047 140383 54055 143367
rect 51055 140375 54055 140383
rect 54245 143367 57245 143375
rect 54245 140383 54253 143367
rect 57237 140383 57245 143367
rect 54245 140375 57245 140383
rect 57435 143367 60435 143375
rect 57435 140383 57443 143367
rect 60427 140383 60435 143367
rect 57435 140375 60435 140383
rect 60625 143367 63625 143375
rect 60625 140383 60633 143367
rect 63617 140383 63625 143367
rect 60625 140375 63625 140383
rect 63815 143367 66815 143375
rect 63815 140383 63823 143367
rect 66807 140383 66815 143367
rect 63815 140375 66815 140383
rect 67005 143367 70005 143375
rect 67005 140383 67013 143367
rect 69997 140383 70005 143367
rect 67005 140375 70005 140383
rect 70195 143367 73195 143375
rect 70195 140383 70203 143367
rect 73187 140383 73195 143367
rect 70195 140375 73195 140383
rect 73385 143367 76385 143375
rect 73385 140383 73393 143367
rect 76377 140383 76385 143367
rect 73385 140375 76385 140383
rect 76575 143367 79575 143375
rect 76575 140383 76583 143367
rect 79567 140383 79575 143367
rect 76575 140375 79575 140383
rect 79765 143367 82765 143375
rect 79765 140383 79773 143367
rect 82757 140383 82765 143367
rect 79765 140375 82765 140383
rect 82955 143367 85955 143375
rect 82955 140383 82963 143367
rect 85947 140383 85955 143367
rect 82955 140375 85955 140383
rect 86145 143367 89145 143375
rect 86145 140383 86153 143367
rect 89137 140383 89145 143367
rect 86145 140375 89145 140383
rect 89335 143367 92335 143375
rect 89335 140383 89343 143367
rect 92327 140383 92335 143367
rect 89335 140375 92335 140383
rect 92525 143367 95525 143375
rect 92525 140383 92533 143367
rect 95517 140383 95525 143367
rect 92525 140375 95525 140383
rect 95715 143367 98715 143375
rect 95715 140383 95723 143367
rect 98707 140383 98715 143367
rect 95715 140375 98715 140383
rect 98905 143367 101905 143375
rect 98905 140383 98913 143367
rect 101897 140383 101905 143367
rect 98905 140375 101905 140383
rect 102095 143367 105095 143375
rect 102095 140383 102103 143367
rect 105087 140383 105095 143367
rect 102095 140375 105095 140383
rect 105285 143367 108285 143375
rect 105285 140383 105293 143367
rect 108277 140383 108285 143367
rect 105285 140375 108285 140383
rect 108475 143367 111475 143375
rect 108475 140383 108483 143367
rect 111467 140383 111475 143367
rect 108475 140375 111475 140383
rect 111665 143367 114665 143375
rect 111665 140383 111673 143367
rect 114657 140383 114665 143367
rect 111665 140375 114665 140383
rect 114855 143367 117855 143375
rect 114855 140383 114863 143367
rect 117847 140383 117855 143367
rect 114855 140375 117855 140383
rect 118045 143367 121045 143375
rect 118045 140383 118053 143367
rect 121037 140383 121045 143367
rect 118045 140375 121045 140383
rect 121235 143367 124235 143375
rect 121235 140383 121243 143367
rect 124227 140383 124235 143367
rect 121235 140375 124235 140383
rect 124425 143367 127425 143375
rect 124425 140383 124433 143367
rect 127417 140383 127425 143367
rect 124425 140375 127425 140383
rect 127615 143367 130615 143375
rect 127615 140383 127623 143367
rect 130607 140383 130615 143367
rect 127615 140375 130615 140383
rect 130805 143367 133805 143375
rect 130805 140383 130813 143367
rect 133797 140383 133805 143367
rect 130805 140375 133805 140383
rect 133995 143367 136995 143375
rect 133995 140383 134003 143367
rect 136987 140383 136995 143367
rect 133995 140375 136995 140383
rect 9585 140177 12585 140185
rect 9585 137193 9593 140177
rect 12577 137193 12585 140177
rect 9585 137185 12585 137193
rect 12775 140177 15775 140185
rect 12775 137193 12783 140177
rect 15767 137193 15775 140177
rect 12775 137185 15775 137193
rect 15965 140177 18965 140185
rect 15965 137193 15973 140177
rect 18957 137193 18965 140177
rect 15965 137185 18965 137193
rect 19155 140177 22155 140185
rect 19155 137193 19163 140177
rect 22147 137193 22155 140177
rect 19155 137185 22155 137193
rect 22345 140177 25345 140185
rect 22345 137193 22353 140177
rect 25337 137193 25345 140177
rect 22345 137185 25345 137193
rect 25535 140177 28535 140185
rect 25535 137193 25543 140177
rect 28527 137193 28535 140177
rect 25535 137185 28535 137193
rect 28725 140177 31725 140185
rect 28725 137193 28733 140177
rect 31717 137193 31725 140177
rect 28725 137185 31725 137193
rect 31915 140177 34915 140185
rect 31915 137193 31923 140177
rect 34907 137193 34915 140177
rect 31915 137185 34915 137193
rect 35105 140177 38105 140185
rect 35105 137193 35113 140177
rect 38097 137193 38105 140177
rect 35105 137185 38105 137193
rect 38295 140177 41295 140185
rect 38295 137193 38303 140177
rect 41287 137193 41295 140177
rect 38295 137185 41295 137193
rect 41485 140177 44485 140185
rect 41485 137193 41493 140177
rect 44477 137193 44485 140177
rect 41485 137185 44485 137193
rect 44675 140177 47675 140185
rect 44675 137193 44683 140177
rect 47667 137193 47675 140177
rect 44675 137185 47675 137193
rect 47865 140177 50865 140185
rect 47865 137193 47873 140177
rect 50857 137193 50865 140177
rect 47865 137185 50865 137193
rect 51055 140177 54055 140185
rect 51055 137193 51063 140177
rect 54047 137193 54055 140177
rect 51055 137185 54055 137193
rect 54245 140177 57245 140185
rect 54245 137193 54253 140177
rect 57237 137193 57245 140177
rect 54245 137185 57245 137193
rect 57435 140177 60435 140185
rect 57435 137193 57443 140177
rect 60427 137193 60435 140177
rect 57435 137185 60435 137193
rect 60625 140177 63625 140185
rect 60625 137193 60633 140177
rect 63617 137193 63625 140177
rect 60625 137185 63625 137193
rect 63815 140177 66815 140185
rect 63815 137193 63823 140177
rect 66807 137193 66815 140177
rect 63815 137185 66815 137193
rect 67005 140177 70005 140185
rect 67005 137193 67013 140177
rect 69997 137193 70005 140177
rect 67005 137185 70005 137193
rect 70195 140177 73195 140185
rect 70195 137193 70203 140177
rect 73187 137193 73195 140177
rect 70195 137185 73195 137193
rect 73385 140177 76385 140185
rect 73385 137193 73393 140177
rect 76377 137193 76385 140177
rect 73385 137185 76385 137193
rect 76575 140177 79575 140185
rect 76575 137193 76583 140177
rect 79567 137193 79575 140177
rect 76575 137185 79575 137193
rect 79765 140177 82765 140185
rect 79765 137193 79773 140177
rect 82757 137193 82765 140177
rect 79765 137185 82765 137193
rect 82955 140177 85955 140185
rect 82955 137193 82963 140177
rect 85947 137193 85955 140177
rect 82955 137185 85955 137193
rect 86145 140177 89145 140185
rect 86145 137193 86153 140177
rect 89137 137193 89145 140177
rect 86145 137185 89145 137193
rect 89335 140177 92335 140185
rect 89335 137193 89343 140177
rect 92327 137193 92335 140177
rect 89335 137185 92335 137193
rect 92525 140177 95525 140185
rect 92525 137193 92533 140177
rect 95517 137193 95525 140177
rect 92525 137185 95525 137193
rect 95715 140177 98715 140185
rect 95715 137193 95723 140177
rect 98707 137193 98715 140177
rect 95715 137185 98715 137193
rect 98905 140177 101905 140185
rect 98905 137193 98913 140177
rect 101897 137193 101905 140177
rect 98905 137185 101905 137193
rect 102095 140177 105095 140185
rect 102095 137193 102103 140177
rect 105087 137193 105095 140177
rect 102095 137185 105095 137193
rect 105285 140177 108285 140185
rect 105285 137193 105293 140177
rect 108277 137193 108285 140177
rect 105285 137185 108285 137193
rect 108475 140177 111475 140185
rect 108475 137193 108483 140177
rect 111467 137193 111475 140177
rect 108475 137185 111475 137193
rect 111665 140177 114665 140185
rect 111665 137193 111673 140177
rect 114657 137193 114665 140177
rect 111665 137185 114665 137193
rect 114855 140177 117855 140185
rect 114855 137193 114863 140177
rect 117847 137193 117855 140177
rect 114855 137185 117855 137193
rect 118045 140177 121045 140185
rect 118045 137193 118053 140177
rect 121037 137193 121045 140177
rect 118045 137185 121045 137193
rect 121235 140177 124235 140185
rect 121235 137193 121243 140177
rect 124227 137193 124235 140177
rect 121235 137185 124235 137193
rect 124425 140177 127425 140185
rect 124425 137193 124433 140177
rect 127417 137193 127425 140177
rect 124425 137185 127425 137193
rect 127615 140177 130615 140185
rect 127615 137193 127623 140177
rect 130607 137193 130615 140177
rect 127615 137185 130615 137193
rect 130805 140177 133805 140185
rect 130805 137193 130813 140177
rect 133797 137193 133805 140177
rect 130805 137185 133805 137193
rect 133995 140177 136995 140185
rect 133995 137193 134003 140177
rect 136987 137193 136995 140177
rect 133995 137185 136995 137193
rect 9585 136987 12585 136995
rect 9585 134003 9593 136987
rect 12577 134003 12585 136987
rect 9585 133995 12585 134003
rect 12775 136987 15775 136995
rect 12775 134003 12783 136987
rect 15767 134003 15775 136987
rect 12775 133995 15775 134003
rect 15965 136987 18965 136995
rect 15965 134003 15973 136987
rect 18957 134003 18965 136987
rect 15965 133995 18965 134003
rect 19155 136987 22155 136995
rect 19155 134003 19163 136987
rect 22147 134003 22155 136987
rect 19155 133995 22155 134003
rect 22345 136987 25345 136995
rect 22345 134003 22353 136987
rect 25337 134003 25345 136987
rect 22345 133995 25345 134003
rect 25535 136987 28535 136995
rect 25535 134003 25543 136987
rect 28527 134003 28535 136987
rect 25535 133995 28535 134003
rect 28725 136987 31725 136995
rect 28725 134003 28733 136987
rect 31717 134003 31725 136987
rect 28725 133995 31725 134003
rect 31915 136987 34915 136995
rect 31915 134003 31923 136987
rect 34907 134003 34915 136987
rect 31915 133995 34915 134003
rect 35105 136987 38105 136995
rect 35105 134003 35113 136987
rect 38097 134003 38105 136987
rect 35105 133995 38105 134003
rect 38295 136987 41295 136995
rect 38295 134003 38303 136987
rect 41287 134003 41295 136987
rect 38295 133995 41295 134003
rect 41485 136987 44485 136995
rect 41485 134003 41493 136987
rect 44477 134003 44485 136987
rect 41485 133995 44485 134003
rect 44675 136987 47675 136995
rect 44675 134003 44683 136987
rect 47667 134003 47675 136987
rect 44675 133995 47675 134003
rect 47865 136987 50865 136995
rect 47865 134003 47873 136987
rect 50857 134003 50865 136987
rect 47865 133995 50865 134003
rect 51055 136987 54055 136995
rect 51055 134003 51063 136987
rect 54047 134003 54055 136987
rect 51055 133995 54055 134003
rect 54245 136987 57245 136995
rect 54245 134003 54253 136987
rect 57237 134003 57245 136987
rect 54245 133995 57245 134003
rect 57435 136987 60435 136995
rect 57435 134003 57443 136987
rect 60427 134003 60435 136987
rect 57435 133995 60435 134003
rect 60625 136987 63625 136995
rect 60625 134003 60633 136987
rect 63617 134003 63625 136987
rect 60625 133995 63625 134003
rect 63815 136987 66815 136995
rect 63815 134003 63823 136987
rect 66807 134003 66815 136987
rect 63815 133995 66815 134003
rect 67005 136987 70005 136995
rect 67005 134003 67013 136987
rect 69997 134003 70005 136987
rect 67005 133995 70005 134003
rect 70195 136987 73195 136995
rect 70195 134003 70203 136987
rect 73187 134003 73195 136987
rect 70195 133995 73195 134003
rect 73385 136987 76385 136995
rect 73385 134003 73393 136987
rect 76377 134003 76385 136987
rect 73385 133995 76385 134003
rect 76575 136987 79575 136995
rect 76575 134003 76583 136987
rect 79567 134003 79575 136987
rect 76575 133995 79575 134003
rect 79765 136987 82765 136995
rect 79765 134003 79773 136987
rect 82757 134003 82765 136987
rect 79765 133995 82765 134003
rect 82955 136987 85955 136995
rect 82955 134003 82963 136987
rect 85947 134003 85955 136987
rect 82955 133995 85955 134003
rect 86145 136987 89145 136995
rect 86145 134003 86153 136987
rect 89137 134003 89145 136987
rect 86145 133995 89145 134003
rect 89335 136987 92335 136995
rect 89335 134003 89343 136987
rect 92327 134003 92335 136987
rect 89335 133995 92335 134003
rect 92525 136987 95525 136995
rect 92525 134003 92533 136987
rect 95517 134003 95525 136987
rect 92525 133995 95525 134003
rect 95715 136987 98715 136995
rect 95715 134003 95723 136987
rect 98707 134003 98715 136987
rect 95715 133995 98715 134003
rect 98905 136987 101905 136995
rect 98905 134003 98913 136987
rect 101897 134003 101905 136987
rect 98905 133995 101905 134003
rect 102095 136987 105095 136995
rect 102095 134003 102103 136987
rect 105087 134003 105095 136987
rect 102095 133995 105095 134003
rect 105285 136987 108285 136995
rect 105285 134003 105293 136987
rect 108277 134003 108285 136987
rect 105285 133995 108285 134003
rect 108475 136987 111475 136995
rect 108475 134003 108483 136987
rect 111467 134003 111475 136987
rect 108475 133995 111475 134003
rect 111665 136987 114665 136995
rect 111665 134003 111673 136987
rect 114657 134003 114665 136987
rect 111665 133995 114665 134003
rect 114855 136987 117855 136995
rect 114855 134003 114863 136987
rect 117847 134003 117855 136987
rect 114855 133995 117855 134003
rect 118045 136987 121045 136995
rect 118045 134003 118053 136987
rect 121037 134003 121045 136987
rect 118045 133995 121045 134003
rect 121235 136987 124235 136995
rect 121235 134003 121243 136987
rect 124227 134003 124235 136987
rect 121235 133995 124235 134003
rect 124425 136987 127425 136995
rect 124425 134003 124433 136987
rect 127417 134003 127425 136987
rect 124425 133995 127425 134003
rect 127615 136987 130615 136995
rect 127615 134003 127623 136987
rect 130607 134003 130615 136987
rect 127615 133995 130615 134003
rect 130805 136987 133805 136995
rect 130805 134003 130813 136987
rect 133797 134003 133805 136987
rect 130805 133995 133805 134003
rect 133995 136987 136995 136995
rect 133995 134003 134003 136987
rect 136987 134003 136995 136987
rect 133995 133995 136995 134003
rect 9585 133797 12585 133805
rect 9585 130813 9593 133797
rect 12577 130813 12585 133797
rect 9585 130805 12585 130813
rect 12775 133797 15775 133805
rect 12775 130813 12783 133797
rect 15767 130813 15775 133797
rect 12775 130805 15775 130813
rect 15965 133797 18965 133805
rect 15965 130813 15973 133797
rect 18957 130813 18965 133797
rect 15965 130805 18965 130813
rect 19155 133797 22155 133805
rect 19155 130813 19163 133797
rect 22147 130813 22155 133797
rect 19155 130805 22155 130813
rect 22345 133797 25345 133805
rect 22345 130813 22353 133797
rect 25337 130813 25345 133797
rect 22345 130805 25345 130813
rect 25535 133797 28535 133805
rect 25535 130813 25543 133797
rect 28527 130813 28535 133797
rect 25535 130805 28535 130813
rect 28725 133797 31725 133805
rect 28725 130813 28733 133797
rect 31717 130813 31725 133797
rect 28725 130805 31725 130813
rect 31915 133797 34915 133805
rect 31915 130813 31923 133797
rect 34907 130813 34915 133797
rect 31915 130805 34915 130813
rect 35105 133797 38105 133805
rect 35105 130813 35113 133797
rect 38097 130813 38105 133797
rect 35105 130805 38105 130813
rect 38295 133797 41295 133805
rect 38295 130813 38303 133797
rect 41287 130813 41295 133797
rect 38295 130805 41295 130813
rect 41485 133797 44485 133805
rect 41485 130813 41493 133797
rect 44477 130813 44485 133797
rect 41485 130805 44485 130813
rect 44675 133797 47675 133805
rect 44675 130813 44683 133797
rect 47667 130813 47675 133797
rect 44675 130805 47675 130813
rect 47865 133797 50865 133805
rect 47865 130813 47873 133797
rect 50857 130813 50865 133797
rect 47865 130805 50865 130813
rect 51055 133797 54055 133805
rect 51055 130813 51063 133797
rect 54047 130813 54055 133797
rect 51055 130805 54055 130813
rect 54245 133797 57245 133805
rect 54245 130813 54253 133797
rect 57237 130813 57245 133797
rect 54245 130805 57245 130813
rect 57435 133797 60435 133805
rect 57435 130813 57443 133797
rect 60427 130813 60435 133797
rect 57435 130805 60435 130813
rect 60625 133797 63625 133805
rect 60625 130813 60633 133797
rect 63617 130813 63625 133797
rect 60625 130805 63625 130813
rect 63815 133797 66815 133805
rect 63815 130813 63823 133797
rect 66807 130813 66815 133797
rect 63815 130805 66815 130813
rect 67005 133797 70005 133805
rect 67005 130813 67013 133797
rect 69997 130813 70005 133797
rect 67005 130805 70005 130813
rect 70195 133797 73195 133805
rect 70195 130813 70203 133797
rect 73187 130813 73195 133797
rect 70195 130805 73195 130813
rect 73385 133797 76385 133805
rect 73385 130813 73393 133797
rect 76377 130813 76385 133797
rect 73385 130805 76385 130813
rect 76575 133797 79575 133805
rect 76575 130813 76583 133797
rect 79567 130813 79575 133797
rect 76575 130805 79575 130813
rect 79765 133797 82765 133805
rect 79765 130813 79773 133797
rect 82757 130813 82765 133797
rect 79765 130805 82765 130813
rect 82955 133797 85955 133805
rect 82955 130813 82963 133797
rect 85947 130813 85955 133797
rect 82955 130805 85955 130813
rect 86145 133797 89145 133805
rect 86145 130813 86153 133797
rect 89137 130813 89145 133797
rect 86145 130805 89145 130813
rect 89335 133797 92335 133805
rect 89335 130813 89343 133797
rect 92327 130813 92335 133797
rect 89335 130805 92335 130813
rect 92525 133797 95525 133805
rect 92525 130813 92533 133797
rect 95517 130813 95525 133797
rect 92525 130805 95525 130813
rect 95715 133797 98715 133805
rect 95715 130813 95723 133797
rect 98707 130813 98715 133797
rect 95715 130805 98715 130813
rect 98905 133797 101905 133805
rect 98905 130813 98913 133797
rect 101897 130813 101905 133797
rect 98905 130805 101905 130813
rect 102095 133797 105095 133805
rect 102095 130813 102103 133797
rect 105087 130813 105095 133797
rect 102095 130805 105095 130813
rect 105285 133797 108285 133805
rect 105285 130813 105293 133797
rect 108277 130813 108285 133797
rect 105285 130805 108285 130813
rect 108475 133797 111475 133805
rect 108475 130813 108483 133797
rect 111467 130813 111475 133797
rect 108475 130805 111475 130813
rect 111665 133797 114665 133805
rect 111665 130813 111673 133797
rect 114657 130813 114665 133797
rect 111665 130805 114665 130813
rect 114855 133797 117855 133805
rect 114855 130813 114863 133797
rect 117847 130813 117855 133797
rect 114855 130805 117855 130813
rect 118045 133797 121045 133805
rect 118045 130813 118053 133797
rect 121037 130813 121045 133797
rect 118045 130805 121045 130813
rect 121235 133797 124235 133805
rect 121235 130813 121243 133797
rect 124227 130813 124235 133797
rect 121235 130805 124235 130813
rect 124425 133797 127425 133805
rect 124425 130813 124433 133797
rect 127417 130813 127425 133797
rect 124425 130805 127425 130813
rect 127615 133797 130615 133805
rect 127615 130813 127623 133797
rect 130607 130813 130615 133797
rect 127615 130805 130615 130813
rect 130805 133797 133805 133805
rect 130805 130813 130813 133797
rect 133797 130813 133805 133797
rect 130805 130805 133805 130813
rect 133995 133797 136995 133805
rect 133995 130813 134003 133797
rect 136987 130813 136995 133797
rect 133995 130805 136995 130813
rect 9585 130607 12585 130615
rect 9585 127623 9593 130607
rect 12577 127623 12585 130607
rect 9585 127615 12585 127623
rect 12775 130607 15775 130615
rect 12775 127623 12783 130607
rect 15767 127623 15775 130607
rect 12775 127615 15775 127623
rect 15965 130607 18965 130615
rect 15965 127623 15973 130607
rect 18957 127623 18965 130607
rect 15965 127615 18965 127623
rect 19155 130607 22155 130615
rect 19155 127623 19163 130607
rect 22147 127623 22155 130607
rect 19155 127615 22155 127623
rect 22345 130607 25345 130615
rect 22345 127623 22353 130607
rect 25337 127623 25345 130607
rect 22345 127615 25345 127623
rect 25535 130607 28535 130615
rect 25535 127623 25543 130607
rect 28527 127623 28535 130607
rect 25535 127615 28535 127623
rect 28725 130607 31725 130615
rect 28725 127623 28733 130607
rect 31717 127623 31725 130607
rect 28725 127615 31725 127623
rect 31915 130607 34915 130615
rect 31915 127623 31923 130607
rect 34907 127623 34915 130607
rect 31915 127615 34915 127623
rect 35105 130607 38105 130615
rect 35105 127623 35113 130607
rect 38097 127623 38105 130607
rect 35105 127615 38105 127623
rect 38295 130607 41295 130615
rect 38295 127623 38303 130607
rect 41287 127623 41295 130607
rect 38295 127615 41295 127623
rect 41485 130607 44485 130615
rect 41485 127623 41493 130607
rect 44477 127623 44485 130607
rect 41485 127615 44485 127623
rect 44675 130607 47675 130615
rect 44675 127623 44683 130607
rect 47667 127623 47675 130607
rect 44675 127615 47675 127623
rect 47865 130607 50865 130615
rect 47865 127623 47873 130607
rect 50857 127623 50865 130607
rect 47865 127615 50865 127623
rect 51055 130607 54055 130615
rect 51055 127623 51063 130607
rect 54047 127623 54055 130607
rect 51055 127615 54055 127623
rect 54245 130607 57245 130615
rect 54245 127623 54253 130607
rect 57237 127623 57245 130607
rect 54245 127615 57245 127623
rect 57435 130607 60435 130615
rect 57435 127623 57443 130607
rect 60427 127623 60435 130607
rect 57435 127615 60435 127623
rect 60625 130607 63625 130615
rect 60625 127623 60633 130607
rect 63617 127623 63625 130607
rect 60625 127615 63625 127623
rect 63815 130607 66815 130615
rect 63815 127623 63823 130607
rect 66807 127623 66815 130607
rect 63815 127615 66815 127623
rect 67005 130607 70005 130615
rect 67005 127623 67013 130607
rect 69997 127623 70005 130607
rect 67005 127615 70005 127623
rect 70195 130607 73195 130615
rect 70195 127623 70203 130607
rect 73187 127623 73195 130607
rect 70195 127615 73195 127623
rect 73385 130607 76385 130615
rect 73385 127623 73393 130607
rect 76377 127623 76385 130607
rect 73385 127615 76385 127623
rect 76575 130607 79575 130615
rect 76575 127623 76583 130607
rect 79567 127623 79575 130607
rect 76575 127615 79575 127623
rect 79765 130607 82765 130615
rect 79765 127623 79773 130607
rect 82757 127623 82765 130607
rect 79765 127615 82765 127623
rect 82955 130607 85955 130615
rect 82955 127623 82963 130607
rect 85947 127623 85955 130607
rect 82955 127615 85955 127623
rect 86145 130607 89145 130615
rect 86145 127623 86153 130607
rect 89137 127623 89145 130607
rect 86145 127615 89145 127623
rect 89335 130607 92335 130615
rect 89335 127623 89343 130607
rect 92327 127623 92335 130607
rect 89335 127615 92335 127623
rect 92525 130607 95525 130615
rect 92525 127623 92533 130607
rect 95517 127623 95525 130607
rect 92525 127615 95525 127623
rect 95715 130607 98715 130615
rect 95715 127623 95723 130607
rect 98707 127623 98715 130607
rect 95715 127615 98715 127623
rect 98905 130607 101905 130615
rect 98905 127623 98913 130607
rect 101897 127623 101905 130607
rect 98905 127615 101905 127623
rect 102095 130607 105095 130615
rect 102095 127623 102103 130607
rect 105087 127623 105095 130607
rect 102095 127615 105095 127623
rect 105285 130607 108285 130615
rect 105285 127623 105293 130607
rect 108277 127623 108285 130607
rect 105285 127615 108285 127623
rect 108475 130607 111475 130615
rect 108475 127623 108483 130607
rect 111467 127623 111475 130607
rect 108475 127615 111475 127623
rect 111665 130607 114665 130615
rect 111665 127623 111673 130607
rect 114657 127623 114665 130607
rect 111665 127615 114665 127623
rect 114855 130607 117855 130615
rect 114855 127623 114863 130607
rect 117847 127623 117855 130607
rect 114855 127615 117855 127623
rect 118045 130607 121045 130615
rect 118045 127623 118053 130607
rect 121037 127623 121045 130607
rect 118045 127615 121045 127623
rect 121235 130607 124235 130615
rect 121235 127623 121243 130607
rect 124227 127623 124235 130607
rect 121235 127615 124235 127623
rect 124425 130607 127425 130615
rect 124425 127623 124433 130607
rect 127417 127623 127425 130607
rect 124425 127615 127425 127623
rect 127615 130607 130615 130615
rect 127615 127623 127623 130607
rect 130607 127623 130615 130607
rect 127615 127615 130615 127623
rect 130805 130607 133805 130615
rect 130805 127623 130813 130607
rect 133797 127623 133805 130607
rect 130805 127615 133805 127623
rect 133995 130607 136995 130615
rect 133995 127623 134003 130607
rect 136987 127623 136995 130607
rect 133995 127615 136995 127623
rect 9585 127417 12585 127425
rect 9585 124433 9593 127417
rect 12577 124433 12585 127417
rect 9585 124425 12585 124433
rect 12775 127417 15775 127425
rect 12775 124433 12783 127417
rect 15767 124433 15775 127417
rect 12775 124425 15775 124433
rect 15965 127417 18965 127425
rect 15965 124433 15973 127417
rect 18957 124433 18965 127417
rect 15965 124425 18965 124433
rect 19155 127417 22155 127425
rect 19155 124433 19163 127417
rect 22147 124433 22155 127417
rect 19155 124425 22155 124433
rect 22345 127417 25345 127425
rect 22345 124433 22353 127417
rect 25337 124433 25345 127417
rect 22345 124425 25345 124433
rect 25535 127417 28535 127425
rect 25535 124433 25543 127417
rect 28527 124433 28535 127417
rect 25535 124425 28535 124433
rect 28725 127417 31725 127425
rect 28725 124433 28733 127417
rect 31717 124433 31725 127417
rect 28725 124425 31725 124433
rect 31915 127417 34915 127425
rect 31915 124433 31923 127417
rect 34907 124433 34915 127417
rect 31915 124425 34915 124433
rect 35105 127417 38105 127425
rect 35105 124433 35113 127417
rect 38097 124433 38105 127417
rect 35105 124425 38105 124433
rect 38295 127417 41295 127425
rect 38295 124433 38303 127417
rect 41287 124433 41295 127417
rect 38295 124425 41295 124433
rect 41485 127417 44485 127425
rect 41485 124433 41493 127417
rect 44477 124433 44485 127417
rect 41485 124425 44485 124433
rect 44675 127417 47675 127425
rect 44675 124433 44683 127417
rect 47667 124433 47675 127417
rect 44675 124425 47675 124433
rect 47865 127417 50865 127425
rect 47865 124433 47873 127417
rect 50857 124433 50865 127417
rect 47865 124425 50865 124433
rect 51055 127417 54055 127425
rect 51055 124433 51063 127417
rect 54047 124433 54055 127417
rect 51055 124425 54055 124433
rect 54245 127417 57245 127425
rect 54245 124433 54253 127417
rect 57237 124433 57245 127417
rect 54245 124425 57245 124433
rect 57435 127417 60435 127425
rect 57435 124433 57443 127417
rect 60427 124433 60435 127417
rect 57435 124425 60435 124433
rect 60625 127417 63625 127425
rect 60625 124433 60633 127417
rect 63617 124433 63625 127417
rect 60625 124425 63625 124433
rect 63815 127417 66815 127425
rect 63815 124433 63823 127417
rect 66807 124433 66815 127417
rect 63815 124425 66815 124433
rect 67005 127417 70005 127425
rect 67005 124433 67013 127417
rect 69997 124433 70005 127417
rect 67005 124425 70005 124433
rect 70195 127417 73195 127425
rect 70195 124433 70203 127417
rect 73187 124433 73195 127417
rect 70195 124425 73195 124433
rect 73385 127417 76385 127425
rect 73385 124433 73393 127417
rect 76377 124433 76385 127417
rect 73385 124425 76385 124433
rect 76575 127417 79575 127425
rect 76575 124433 76583 127417
rect 79567 124433 79575 127417
rect 76575 124425 79575 124433
rect 79765 127417 82765 127425
rect 79765 124433 79773 127417
rect 82757 124433 82765 127417
rect 79765 124425 82765 124433
rect 82955 127417 85955 127425
rect 82955 124433 82963 127417
rect 85947 124433 85955 127417
rect 82955 124425 85955 124433
rect 86145 127417 89145 127425
rect 86145 124433 86153 127417
rect 89137 124433 89145 127417
rect 86145 124425 89145 124433
rect 89335 127417 92335 127425
rect 89335 124433 89343 127417
rect 92327 124433 92335 127417
rect 89335 124425 92335 124433
rect 92525 127417 95525 127425
rect 92525 124433 92533 127417
rect 95517 124433 95525 127417
rect 92525 124425 95525 124433
rect 95715 127417 98715 127425
rect 95715 124433 95723 127417
rect 98707 124433 98715 127417
rect 95715 124425 98715 124433
rect 98905 127417 101905 127425
rect 98905 124433 98913 127417
rect 101897 124433 101905 127417
rect 98905 124425 101905 124433
rect 102095 127417 105095 127425
rect 102095 124433 102103 127417
rect 105087 124433 105095 127417
rect 102095 124425 105095 124433
rect 105285 127417 108285 127425
rect 105285 124433 105293 127417
rect 108277 124433 108285 127417
rect 105285 124425 108285 124433
rect 108475 127417 111475 127425
rect 108475 124433 108483 127417
rect 111467 124433 111475 127417
rect 108475 124425 111475 124433
rect 111665 127417 114665 127425
rect 111665 124433 111673 127417
rect 114657 124433 114665 127417
rect 111665 124425 114665 124433
rect 114855 127417 117855 127425
rect 114855 124433 114863 127417
rect 117847 124433 117855 127417
rect 114855 124425 117855 124433
rect 118045 127417 121045 127425
rect 118045 124433 118053 127417
rect 121037 124433 121045 127417
rect 118045 124425 121045 124433
rect 121235 127417 124235 127425
rect 121235 124433 121243 127417
rect 124227 124433 124235 127417
rect 121235 124425 124235 124433
rect 124425 127417 127425 127425
rect 124425 124433 124433 127417
rect 127417 124433 127425 127417
rect 124425 124425 127425 124433
rect 127615 127417 130615 127425
rect 127615 124433 127623 127417
rect 130607 124433 130615 127417
rect 127615 124425 130615 124433
rect 130805 127417 133805 127425
rect 130805 124433 130813 127417
rect 133797 124433 133805 127417
rect 130805 124425 133805 124433
rect 133995 127417 136995 127425
rect 133995 124433 134003 127417
rect 136987 124433 136995 127417
rect 133995 124425 136995 124433
rect 9585 124227 12585 124235
rect 9585 121243 9593 124227
rect 12577 121243 12585 124227
rect 9585 121235 12585 121243
rect 12775 124227 15775 124235
rect 12775 121243 12783 124227
rect 15767 121243 15775 124227
rect 12775 121235 15775 121243
rect 15965 124227 18965 124235
rect 15965 121243 15973 124227
rect 18957 121243 18965 124227
rect 15965 121235 18965 121243
rect 19155 124227 22155 124235
rect 19155 121243 19163 124227
rect 22147 121243 22155 124227
rect 19155 121235 22155 121243
rect 22345 124227 25345 124235
rect 22345 121243 22353 124227
rect 25337 121243 25345 124227
rect 22345 121235 25345 121243
rect 25535 124227 28535 124235
rect 25535 121243 25543 124227
rect 28527 121243 28535 124227
rect 25535 121235 28535 121243
rect 28725 124227 31725 124235
rect 28725 121243 28733 124227
rect 31717 121243 31725 124227
rect 28725 121235 31725 121243
rect 31915 124227 34915 124235
rect 31915 121243 31923 124227
rect 34907 121243 34915 124227
rect 31915 121235 34915 121243
rect 35105 124227 38105 124235
rect 35105 121243 35113 124227
rect 38097 121243 38105 124227
rect 35105 121235 38105 121243
rect 38295 124227 41295 124235
rect 38295 121243 38303 124227
rect 41287 121243 41295 124227
rect 38295 121235 41295 121243
rect 41485 124227 44485 124235
rect 41485 121243 41493 124227
rect 44477 121243 44485 124227
rect 41485 121235 44485 121243
rect 44675 124227 47675 124235
rect 44675 121243 44683 124227
rect 47667 121243 47675 124227
rect 44675 121235 47675 121243
rect 47865 124227 50865 124235
rect 47865 121243 47873 124227
rect 50857 121243 50865 124227
rect 47865 121235 50865 121243
rect 51055 124227 54055 124235
rect 51055 121243 51063 124227
rect 54047 121243 54055 124227
rect 51055 121235 54055 121243
rect 54245 124227 57245 124235
rect 54245 121243 54253 124227
rect 57237 121243 57245 124227
rect 54245 121235 57245 121243
rect 57435 124227 60435 124235
rect 57435 121243 57443 124227
rect 60427 121243 60435 124227
rect 57435 121235 60435 121243
rect 60625 124227 63625 124235
rect 60625 121243 60633 124227
rect 63617 121243 63625 124227
rect 60625 121235 63625 121243
rect 63815 124227 66815 124235
rect 63815 121243 63823 124227
rect 66807 121243 66815 124227
rect 63815 121235 66815 121243
rect 67005 124227 70005 124235
rect 67005 121243 67013 124227
rect 69997 121243 70005 124227
rect 67005 121235 70005 121243
rect 70195 124227 73195 124235
rect 70195 121243 70203 124227
rect 73187 121243 73195 124227
rect 70195 121235 73195 121243
rect 73385 124227 76385 124235
rect 73385 121243 73393 124227
rect 76377 121243 76385 124227
rect 73385 121235 76385 121243
rect 76575 124227 79575 124235
rect 76575 121243 76583 124227
rect 79567 121243 79575 124227
rect 76575 121235 79575 121243
rect 79765 124227 82765 124235
rect 79765 121243 79773 124227
rect 82757 121243 82765 124227
rect 79765 121235 82765 121243
rect 82955 124227 85955 124235
rect 82955 121243 82963 124227
rect 85947 121243 85955 124227
rect 82955 121235 85955 121243
rect 86145 124227 89145 124235
rect 86145 121243 86153 124227
rect 89137 121243 89145 124227
rect 86145 121235 89145 121243
rect 89335 124227 92335 124235
rect 89335 121243 89343 124227
rect 92327 121243 92335 124227
rect 89335 121235 92335 121243
rect 92525 124227 95525 124235
rect 92525 121243 92533 124227
rect 95517 121243 95525 124227
rect 92525 121235 95525 121243
rect 95715 124227 98715 124235
rect 95715 121243 95723 124227
rect 98707 121243 98715 124227
rect 95715 121235 98715 121243
rect 98905 124227 101905 124235
rect 98905 121243 98913 124227
rect 101897 121243 101905 124227
rect 98905 121235 101905 121243
rect 102095 124227 105095 124235
rect 102095 121243 102103 124227
rect 105087 121243 105095 124227
rect 102095 121235 105095 121243
rect 105285 124227 108285 124235
rect 105285 121243 105293 124227
rect 108277 121243 108285 124227
rect 105285 121235 108285 121243
rect 108475 124227 111475 124235
rect 108475 121243 108483 124227
rect 111467 121243 111475 124227
rect 108475 121235 111475 121243
rect 111665 124227 114665 124235
rect 111665 121243 111673 124227
rect 114657 121243 114665 124227
rect 111665 121235 114665 121243
rect 114855 124227 117855 124235
rect 114855 121243 114863 124227
rect 117847 121243 117855 124227
rect 114855 121235 117855 121243
rect 118045 124227 121045 124235
rect 118045 121243 118053 124227
rect 121037 121243 121045 124227
rect 118045 121235 121045 121243
rect 121235 124227 124235 124235
rect 121235 121243 121243 124227
rect 124227 121243 124235 124227
rect 121235 121235 124235 121243
rect 124425 124227 127425 124235
rect 124425 121243 124433 124227
rect 127417 121243 127425 124227
rect 124425 121235 127425 121243
rect 127615 124227 130615 124235
rect 127615 121243 127623 124227
rect 130607 121243 130615 124227
rect 127615 121235 130615 121243
rect 130805 124227 133805 124235
rect 130805 121243 130813 124227
rect 133797 121243 133805 124227
rect 130805 121235 133805 121243
rect 133995 124227 136995 124235
rect 133995 121243 134003 124227
rect 136987 121243 136995 124227
rect 133995 121235 136995 121243
rect 15 121037 3015 121045
rect 15 118053 23 121037
rect 3007 118053 3015 121037
rect 15 118045 3015 118053
rect 3205 121037 6205 121045
rect 3205 118053 3213 121037
rect 6197 118053 6205 121037
rect 3205 118045 6205 118053
rect 6395 121037 9395 121045
rect 6395 118053 6403 121037
rect 9387 118053 9395 121037
rect 6395 118045 9395 118053
rect 9585 121037 12585 121045
rect 9585 118053 9593 121037
rect 12577 118053 12585 121037
rect 9585 118045 12585 118053
rect 12775 121037 15775 121045
rect 12775 118053 12783 121037
rect 15767 118053 15775 121037
rect 12775 118045 15775 118053
rect 15965 121037 18965 121045
rect 15965 118053 15973 121037
rect 18957 118053 18965 121037
rect 15965 118045 18965 118053
rect 19155 121037 22155 121045
rect 19155 118053 19163 121037
rect 22147 118053 22155 121037
rect 19155 118045 22155 118053
rect 22345 121037 25345 121045
rect 22345 118053 22353 121037
rect 25337 118053 25345 121037
rect 22345 118045 25345 118053
rect 25535 121037 28535 121045
rect 25535 118053 25543 121037
rect 28527 118053 28535 121037
rect 25535 118045 28535 118053
rect 28725 121037 31725 121045
rect 28725 118053 28733 121037
rect 31717 118053 31725 121037
rect 28725 118045 31725 118053
rect 31915 121037 34915 121045
rect 31915 118053 31923 121037
rect 34907 118053 34915 121037
rect 31915 118045 34915 118053
rect 35105 121037 38105 121045
rect 35105 118053 35113 121037
rect 38097 118053 38105 121037
rect 35105 118045 38105 118053
rect 38295 121037 41295 121045
rect 38295 118053 38303 121037
rect 41287 118053 41295 121037
rect 38295 118045 41295 118053
rect 41485 121037 44485 121045
rect 41485 118053 41493 121037
rect 44477 118053 44485 121037
rect 41485 118045 44485 118053
rect 44675 121037 47675 121045
rect 44675 118053 44683 121037
rect 47667 118053 47675 121037
rect 44675 118045 47675 118053
rect 47865 121037 50865 121045
rect 47865 118053 47873 121037
rect 50857 118053 50865 121037
rect 47865 118045 50865 118053
rect 51055 121037 54055 121045
rect 51055 118053 51063 121037
rect 54047 118053 54055 121037
rect 51055 118045 54055 118053
rect 54245 121037 57245 121045
rect 54245 118053 54253 121037
rect 57237 118053 57245 121037
rect 54245 118045 57245 118053
rect 57435 121037 60435 121045
rect 57435 118053 57443 121037
rect 60427 118053 60435 121037
rect 57435 118045 60435 118053
rect 60625 121037 63625 121045
rect 60625 118053 60633 121037
rect 63617 118053 63625 121037
rect 60625 118045 63625 118053
rect 63815 121037 66815 121045
rect 63815 118053 63823 121037
rect 66807 118053 66815 121037
rect 63815 118045 66815 118053
rect 67005 121037 70005 121045
rect 67005 118053 67013 121037
rect 69997 118053 70005 121037
rect 67005 118045 70005 118053
rect 70195 121037 73195 121045
rect 70195 118053 70203 121037
rect 73187 118053 73195 121037
rect 70195 118045 73195 118053
rect 73385 121037 76385 121045
rect 73385 118053 73393 121037
rect 76377 118053 76385 121037
rect 73385 118045 76385 118053
rect 76575 121037 79575 121045
rect 76575 118053 76583 121037
rect 79567 118053 79575 121037
rect 76575 118045 79575 118053
rect 79765 121037 82765 121045
rect 79765 118053 79773 121037
rect 82757 118053 82765 121037
rect 79765 118045 82765 118053
rect 82955 121037 85955 121045
rect 82955 118053 82963 121037
rect 85947 118053 85955 121037
rect 82955 118045 85955 118053
rect 86145 121037 89145 121045
rect 86145 118053 86153 121037
rect 89137 118053 89145 121037
rect 86145 118045 89145 118053
rect 89335 121037 92335 121045
rect 89335 118053 89343 121037
rect 92327 118053 92335 121037
rect 89335 118045 92335 118053
rect 92525 121037 95525 121045
rect 92525 118053 92533 121037
rect 95517 118053 95525 121037
rect 92525 118045 95525 118053
rect 95715 121037 98715 121045
rect 95715 118053 95723 121037
rect 98707 118053 98715 121037
rect 95715 118045 98715 118053
rect 98905 121037 101905 121045
rect 98905 118053 98913 121037
rect 101897 118053 101905 121037
rect 98905 118045 101905 118053
rect 102095 121037 105095 121045
rect 102095 118053 102103 121037
rect 105087 118053 105095 121037
rect 102095 118045 105095 118053
rect 105285 121037 108285 121045
rect 105285 118053 105293 121037
rect 108277 118053 108285 121037
rect 105285 118045 108285 118053
rect 108475 121037 111475 121045
rect 108475 118053 108483 121037
rect 111467 118053 111475 121037
rect 108475 118045 111475 118053
rect 111665 121037 114665 121045
rect 111665 118053 111673 121037
rect 114657 118053 114665 121037
rect 111665 118045 114665 118053
rect 114855 121037 117855 121045
rect 114855 118053 114863 121037
rect 117847 118053 117855 121037
rect 114855 118045 117855 118053
rect 118045 121037 121045 121045
rect 118045 118053 118053 121037
rect 121037 118053 121045 121037
rect 118045 118045 121045 118053
rect 121235 121037 124235 121045
rect 121235 118053 121243 121037
rect 124227 118053 124235 121037
rect 121235 118045 124235 118053
rect 124425 121037 127425 121045
rect 124425 118053 124433 121037
rect 127417 118053 127425 121037
rect 124425 118045 127425 118053
rect 127615 121037 130615 121045
rect 127615 118053 127623 121037
rect 130607 118053 130615 121037
rect 127615 118045 130615 118053
rect 130805 121037 133805 121045
rect 130805 118053 130813 121037
rect 133797 118053 133805 121037
rect 130805 118045 133805 118053
rect 133995 121037 136995 121045
rect 133995 118053 134003 121037
rect 136987 118053 136995 121037
rect 133995 118045 136995 118053
rect 15 117847 3015 117855
rect 15 114863 23 117847
rect 3007 114863 3015 117847
rect 15 114855 3015 114863
rect 3205 117847 6205 117855
rect 3205 114863 3213 117847
rect 6197 114863 6205 117847
rect 3205 114855 6205 114863
rect 6395 117847 9395 117855
rect 6395 114863 6403 117847
rect 9387 114863 9395 117847
rect 6395 114855 9395 114863
rect 9585 117847 12585 117855
rect 9585 114863 9593 117847
rect 12577 114863 12585 117847
rect 9585 114855 12585 114863
rect 12775 117847 15775 117855
rect 12775 114863 12783 117847
rect 15767 114863 15775 117847
rect 12775 114855 15775 114863
rect 15965 117847 18965 117855
rect 15965 114863 15973 117847
rect 18957 114863 18965 117847
rect 15965 114855 18965 114863
rect 19155 117847 22155 117855
rect 19155 114863 19163 117847
rect 22147 114863 22155 117847
rect 19155 114855 22155 114863
rect 22345 117847 25345 117855
rect 22345 114863 22353 117847
rect 25337 114863 25345 117847
rect 22345 114855 25345 114863
rect 25535 117847 28535 117855
rect 25535 114863 25543 117847
rect 28527 114863 28535 117847
rect 25535 114855 28535 114863
rect 28725 117847 31725 117855
rect 28725 114863 28733 117847
rect 31717 114863 31725 117847
rect 28725 114855 31725 114863
rect 31915 117847 34915 117855
rect 31915 114863 31923 117847
rect 34907 114863 34915 117847
rect 31915 114855 34915 114863
rect 35105 117847 38105 117855
rect 35105 114863 35113 117847
rect 38097 114863 38105 117847
rect 35105 114855 38105 114863
rect 38295 117847 41295 117855
rect 38295 114863 38303 117847
rect 41287 114863 41295 117847
rect 38295 114855 41295 114863
rect 41485 117847 44485 117855
rect 41485 114863 41493 117847
rect 44477 114863 44485 117847
rect 41485 114855 44485 114863
rect 44675 117847 47675 117855
rect 44675 114863 44683 117847
rect 47667 114863 47675 117847
rect 44675 114855 47675 114863
rect 47865 117847 50865 117855
rect 47865 114863 47873 117847
rect 50857 114863 50865 117847
rect 47865 114855 50865 114863
rect 51055 117847 54055 117855
rect 51055 114863 51063 117847
rect 54047 114863 54055 117847
rect 51055 114855 54055 114863
rect 54245 117847 57245 117855
rect 54245 114863 54253 117847
rect 57237 114863 57245 117847
rect 54245 114855 57245 114863
rect 57435 117847 60435 117855
rect 57435 114863 57443 117847
rect 60427 114863 60435 117847
rect 57435 114855 60435 114863
rect 60625 117847 63625 117855
rect 60625 114863 60633 117847
rect 63617 114863 63625 117847
rect 60625 114855 63625 114863
rect 63815 117847 66815 117855
rect 63815 114863 63823 117847
rect 66807 114863 66815 117847
rect 63815 114855 66815 114863
rect 67005 117847 70005 117855
rect 67005 114863 67013 117847
rect 69997 114863 70005 117847
rect 67005 114855 70005 114863
rect 70195 117847 73195 117855
rect 70195 114863 70203 117847
rect 73187 114863 73195 117847
rect 70195 114855 73195 114863
rect 73385 117847 76385 117855
rect 73385 114863 73393 117847
rect 76377 114863 76385 117847
rect 73385 114855 76385 114863
rect 76575 117847 79575 117855
rect 76575 114863 76583 117847
rect 79567 114863 79575 117847
rect 76575 114855 79575 114863
rect 79765 117847 82765 117855
rect 79765 114863 79773 117847
rect 82757 114863 82765 117847
rect 79765 114855 82765 114863
rect 82955 117847 85955 117855
rect 82955 114863 82963 117847
rect 85947 114863 85955 117847
rect 82955 114855 85955 114863
rect 86145 117847 89145 117855
rect 86145 114863 86153 117847
rect 89137 114863 89145 117847
rect 86145 114855 89145 114863
rect 89335 117847 92335 117855
rect 89335 114863 89343 117847
rect 92327 114863 92335 117847
rect 89335 114855 92335 114863
rect 92525 117847 95525 117855
rect 92525 114863 92533 117847
rect 95517 114863 95525 117847
rect 92525 114855 95525 114863
rect 95715 117847 98715 117855
rect 95715 114863 95723 117847
rect 98707 114863 98715 117847
rect 95715 114855 98715 114863
rect 98905 117847 101905 117855
rect 98905 114863 98913 117847
rect 101897 114863 101905 117847
rect 98905 114855 101905 114863
rect 102095 117847 105095 117855
rect 102095 114863 102103 117847
rect 105087 114863 105095 117847
rect 102095 114855 105095 114863
rect 105285 117847 108285 117855
rect 105285 114863 105293 117847
rect 108277 114863 108285 117847
rect 105285 114855 108285 114863
rect 108475 117847 111475 117855
rect 108475 114863 108483 117847
rect 111467 114863 111475 117847
rect 108475 114855 111475 114863
rect 111665 117847 114665 117855
rect 111665 114863 111673 117847
rect 114657 114863 114665 117847
rect 111665 114855 114665 114863
rect 114855 117847 117855 117855
rect 114855 114863 114863 117847
rect 117847 114863 117855 117847
rect 114855 114855 117855 114863
rect 118045 117847 121045 117855
rect 118045 114863 118053 117847
rect 121037 114863 121045 117847
rect 118045 114855 121045 114863
rect 121235 117847 124235 117855
rect 121235 114863 121243 117847
rect 124227 114863 124235 117847
rect 121235 114855 124235 114863
rect 124425 117847 127425 117855
rect 124425 114863 124433 117847
rect 127417 114863 127425 117847
rect 124425 114855 127425 114863
rect 127615 117847 130615 117855
rect 127615 114863 127623 117847
rect 130607 114863 130615 117847
rect 127615 114855 130615 114863
rect 130805 117847 133805 117855
rect 130805 114863 130813 117847
rect 133797 114863 133805 117847
rect 130805 114855 133805 114863
rect 133995 117847 136995 117855
rect 133995 114863 134003 117847
rect 136987 114863 136995 117847
rect 133995 114855 136995 114863
rect 15 114657 3015 114665
rect 15 111673 23 114657
rect 3007 111673 3015 114657
rect 15 111665 3015 111673
rect 3205 114657 6205 114665
rect 3205 111673 3213 114657
rect 6197 111673 6205 114657
rect 3205 111665 6205 111673
rect 6395 114657 9395 114665
rect 6395 111673 6403 114657
rect 9387 111673 9395 114657
rect 6395 111665 9395 111673
rect 9585 114657 12585 114665
rect 9585 111673 9593 114657
rect 12577 111673 12585 114657
rect 9585 111665 12585 111673
rect 12775 114657 15775 114665
rect 12775 111673 12783 114657
rect 15767 111673 15775 114657
rect 12775 111665 15775 111673
rect 15965 114657 18965 114665
rect 15965 111673 15973 114657
rect 18957 111673 18965 114657
rect 15965 111665 18965 111673
rect 19155 114657 22155 114665
rect 19155 111673 19163 114657
rect 22147 111673 22155 114657
rect 19155 111665 22155 111673
rect 22345 114657 25345 114665
rect 22345 111673 22353 114657
rect 25337 111673 25345 114657
rect 22345 111665 25345 111673
rect 25535 114657 28535 114665
rect 25535 111673 25543 114657
rect 28527 111673 28535 114657
rect 25535 111665 28535 111673
rect 28725 114657 31725 114665
rect 28725 111673 28733 114657
rect 31717 111673 31725 114657
rect 28725 111665 31725 111673
rect 31915 114657 34915 114665
rect 31915 111673 31923 114657
rect 34907 111673 34915 114657
rect 31915 111665 34915 111673
rect 35105 114657 38105 114665
rect 35105 111673 35113 114657
rect 38097 111673 38105 114657
rect 35105 111665 38105 111673
rect 38295 114657 41295 114665
rect 38295 111673 38303 114657
rect 41287 111673 41295 114657
rect 38295 111665 41295 111673
rect 41485 114657 44485 114665
rect 41485 111673 41493 114657
rect 44477 111673 44485 114657
rect 41485 111665 44485 111673
rect 44675 114657 47675 114665
rect 44675 111673 44683 114657
rect 47667 111673 47675 114657
rect 44675 111665 47675 111673
rect 47865 114657 50865 114665
rect 47865 111673 47873 114657
rect 50857 111673 50865 114657
rect 47865 111665 50865 111673
rect 51055 114657 54055 114665
rect 51055 111673 51063 114657
rect 54047 111673 54055 114657
rect 51055 111665 54055 111673
rect 54245 114657 57245 114665
rect 54245 111673 54253 114657
rect 57237 111673 57245 114657
rect 54245 111665 57245 111673
rect 57435 114657 60435 114665
rect 57435 111673 57443 114657
rect 60427 111673 60435 114657
rect 57435 111665 60435 111673
rect 60625 114657 63625 114665
rect 60625 111673 60633 114657
rect 63617 111673 63625 114657
rect 60625 111665 63625 111673
rect 63815 114657 66815 114665
rect 63815 111673 63823 114657
rect 66807 111673 66815 114657
rect 63815 111665 66815 111673
rect 67005 114657 70005 114665
rect 67005 111673 67013 114657
rect 69997 111673 70005 114657
rect 67005 111665 70005 111673
rect 70195 114657 73195 114665
rect 70195 111673 70203 114657
rect 73187 111673 73195 114657
rect 70195 111665 73195 111673
rect 73385 114657 76385 114665
rect 73385 111673 73393 114657
rect 76377 111673 76385 114657
rect 73385 111665 76385 111673
rect 76575 114657 79575 114665
rect 76575 111673 76583 114657
rect 79567 111673 79575 114657
rect 76575 111665 79575 111673
rect 79765 114657 82765 114665
rect 79765 111673 79773 114657
rect 82757 111673 82765 114657
rect 79765 111665 82765 111673
rect 82955 114657 85955 114665
rect 82955 111673 82963 114657
rect 85947 111673 85955 114657
rect 82955 111665 85955 111673
rect 86145 114657 89145 114665
rect 86145 111673 86153 114657
rect 89137 111673 89145 114657
rect 86145 111665 89145 111673
rect 89335 114657 92335 114665
rect 89335 111673 89343 114657
rect 92327 111673 92335 114657
rect 89335 111665 92335 111673
rect 92525 114657 95525 114665
rect 92525 111673 92533 114657
rect 95517 111673 95525 114657
rect 92525 111665 95525 111673
rect 95715 114657 98715 114665
rect 95715 111673 95723 114657
rect 98707 111673 98715 114657
rect 95715 111665 98715 111673
rect 98905 114657 101905 114665
rect 98905 111673 98913 114657
rect 101897 111673 101905 114657
rect 98905 111665 101905 111673
rect 102095 114657 105095 114665
rect 102095 111673 102103 114657
rect 105087 111673 105095 114657
rect 102095 111665 105095 111673
rect 105285 114657 108285 114665
rect 105285 111673 105293 114657
rect 108277 111673 108285 114657
rect 105285 111665 108285 111673
rect 108475 114657 111475 114665
rect 108475 111673 108483 114657
rect 111467 111673 111475 114657
rect 108475 111665 111475 111673
rect 111665 114657 114665 114665
rect 111665 111673 111673 114657
rect 114657 111673 114665 114657
rect 111665 111665 114665 111673
rect 114855 114657 117855 114665
rect 114855 111673 114863 114657
rect 117847 111673 117855 114657
rect 114855 111665 117855 111673
rect 118045 114657 121045 114665
rect 118045 111673 118053 114657
rect 121037 111673 121045 114657
rect 118045 111665 121045 111673
rect 121235 114657 124235 114665
rect 121235 111673 121243 114657
rect 124227 111673 124235 114657
rect 121235 111665 124235 111673
rect 124425 114657 127425 114665
rect 124425 111673 124433 114657
rect 127417 111673 127425 114657
rect 124425 111665 127425 111673
rect 127615 114657 130615 114665
rect 127615 111673 127623 114657
rect 130607 111673 130615 114657
rect 127615 111665 130615 111673
rect 130805 114657 133805 114665
rect 130805 111673 130813 114657
rect 133797 111673 133805 114657
rect 130805 111665 133805 111673
rect 133995 114657 136995 114665
rect 133995 111673 134003 114657
rect 136987 111673 136995 114657
rect 133995 111665 136995 111673
rect 15 111467 3015 111475
rect 15 108483 23 111467
rect 3007 108483 3015 111467
rect 15 108475 3015 108483
rect 3205 111467 6205 111475
rect 3205 108483 3213 111467
rect 6197 108483 6205 111467
rect 3205 108475 6205 108483
rect 6395 111467 9395 111475
rect 6395 108483 6403 111467
rect 9387 108483 9395 111467
rect 6395 108475 9395 108483
rect 9585 111467 12585 111475
rect 9585 108483 9593 111467
rect 12577 108483 12585 111467
rect 9585 108475 12585 108483
rect 12775 111467 15775 111475
rect 12775 108483 12783 111467
rect 15767 108483 15775 111467
rect 12775 108475 15775 108483
rect 15965 111467 18965 111475
rect 15965 108483 15973 111467
rect 18957 108483 18965 111467
rect 15965 108475 18965 108483
rect 19155 111467 22155 111475
rect 19155 108483 19163 111467
rect 22147 108483 22155 111467
rect 19155 108475 22155 108483
rect 22345 111467 25345 111475
rect 22345 108483 22353 111467
rect 25337 108483 25345 111467
rect 22345 108475 25345 108483
rect 25535 111467 28535 111475
rect 25535 108483 25543 111467
rect 28527 108483 28535 111467
rect 25535 108475 28535 108483
rect 28725 111467 31725 111475
rect 28725 108483 28733 111467
rect 31717 108483 31725 111467
rect 28725 108475 31725 108483
rect 31915 111467 34915 111475
rect 31915 108483 31923 111467
rect 34907 108483 34915 111467
rect 31915 108475 34915 108483
rect 35105 111467 38105 111475
rect 35105 108483 35113 111467
rect 38097 108483 38105 111467
rect 35105 108475 38105 108483
rect 38295 111467 41295 111475
rect 38295 108483 38303 111467
rect 41287 108483 41295 111467
rect 38295 108475 41295 108483
rect 41485 111467 44485 111475
rect 41485 108483 41493 111467
rect 44477 108483 44485 111467
rect 41485 108475 44485 108483
rect 44675 111467 47675 111475
rect 44675 108483 44683 111467
rect 47667 108483 47675 111467
rect 44675 108475 47675 108483
rect 47865 111467 50865 111475
rect 47865 108483 47873 111467
rect 50857 108483 50865 111467
rect 47865 108475 50865 108483
rect 51055 111467 54055 111475
rect 51055 108483 51063 111467
rect 54047 108483 54055 111467
rect 51055 108475 54055 108483
rect 54245 111467 57245 111475
rect 54245 108483 54253 111467
rect 57237 108483 57245 111467
rect 54245 108475 57245 108483
rect 57435 111467 60435 111475
rect 57435 108483 57443 111467
rect 60427 108483 60435 111467
rect 57435 108475 60435 108483
rect 60625 111467 63625 111475
rect 60625 108483 60633 111467
rect 63617 108483 63625 111467
rect 60625 108475 63625 108483
rect 63815 111467 66815 111475
rect 63815 108483 63823 111467
rect 66807 108483 66815 111467
rect 63815 108475 66815 108483
rect 67005 111467 70005 111475
rect 67005 108483 67013 111467
rect 69997 108483 70005 111467
rect 67005 108475 70005 108483
rect 70195 111467 73195 111475
rect 70195 108483 70203 111467
rect 73187 108483 73195 111467
rect 70195 108475 73195 108483
rect 73385 111467 76385 111475
rect 73385 108483 73393 111467
rect 76377 108483 76385 111467
rect 73385 108475 76385 108483
rect 76575 111467 79575 111475
rect 76575 108483 76583 111467
rect 79567 108483 79575 111467
rect 76575 108475 79575 108483
rect 79765 111467 82765 111475
rect 79765 108483 79773 111467
rect 82757 108483 82765 111467
rect 79765 108475 82765 108483
rect 82955 111467 85955 111475
rect 82955 108483 82963 111467
rect 85947 108483 85955 111467
rect 82955 108475 85955 108483
rect 86145 111467 89145 111475
rect 86145 108483 86153 111467
rect 89137 108483 89145 111467
rect 86145 108475 89145 108483
rect 89335 111467 92335 111475
rect 89335 108483 89343 111467
rect 92327 108483 92335 111467
rect 89335 108475 92335 108483
rect 92525 111467 95525 111475
rect 92525 108483 92533 111467
rect 95517 108483 95525 111467
rect 92525 108475 95525 108483
rect 95715 111467 98715 111475
rect 95715 108483 95723 111467
rect 98707 108483 98715 111467
rect 95715 108475 98715 108483
rect 98905 111467 101905 111475
rect 98905 108483 98913 111467
rect 101897 108483 101905 111467
rect 98905 108475 101905 108483
rect 102095 111467 105095 111475
rect 102095 108483 102103 111467
rect 105087 108483 105095 111467
rect 102095 108475 105095 108483
rect 105285 111467 108285 111475
rect 105285 108483 105293 111467
rect 108277 108483 108285 111467
rect 105285 108475 108285 108483
rect 108475 111467 111475 111475
rect 108475 108483 108483 111467
rect 111467 108483 111475 111467
rect 108475 108475 111475 108483
rect 111665 111467 114665 111475
rect 111665 108483 111673 111467
rect 114657 108483 114665 111467
rect 111665 108475 114665 108483
rect 114855 111467 117855 111475
rect 114855 108483 114863 111467
rect 117847 108483 117855 111467
rect 114855 108475 117855 108483
rect 118045 111467 121045 111475
rect 118045 108483 118053 111467
rect 121037 108483 121045 111467
rect 118045 108475 121045 108483
rect 121235 111467 124235 111475
rect 121235 108483 121243 111467
rect 124227 108483 124235 111467
rect 121235 108475 124235 108483
rect 124425 111467 127425 111475
rect 124425 108483 124433 111467
rect 127417 108483 127425 111467
rect 124425 108475 127425 108483
rect 127615 111467 130615 111475
rect 127615 108483 127623 111467
rect 130607 108483 130615 111467
rect 127615 108475 130615 108483
rect 130805 111467 133805 111475
rect 130805 108483 130813 111467
rect 133797 108483 133805 111467
rect 130805 108475 133805 108483
rect 133995 111467 136995 111475
rect 133995 108483 134003 111467
rect 136987 108483 136995 111467
rect 133995 108475 136995 108483
rect 15 108277 3015 108285
rect 15 105293 23 108277
rect 3007 105293 3015 108277
rect 15 105285 3015 105293
rect 3205 108277 6205 108285
rect 3205 105293 3213 108277
rect 6197 105293 6205 108277
rect 3205 105285 6205 105293
rect 6395 108277 9395 108285
rect 6395 105293 6403 108277
rect 9387 105293 9395 108277
rect 6395 105285 9395 105293
rect 9585 108277 12585 108285
rect 9585 105293 9593 108277
rect 12577 105293 12585 108277
rect 9585 105285 12585 105293
rect 12775 108277 15775 108285
rect 12775 105293 12783 108277
rect 15767 105293 15775 108277
rect 12775 105285 15775 105293
rect 15965 108277 18965 108285
rect 15965 105293 15973 108277
rect 18957 105293 18965 108277
rect 15965 105285 18965 105293
rect 19155 108277 22155 108285
rect 19155 105293 19163 108277
rect 22147 105293 22155 108277
rect 19155 105285 22155 105293
rect 22345 108277 25345 108285
rect 22345 105293 22353 108277
rect 25337 105293 25345 108277
rect 22345 105285 25345 105293
rect 25535 108277 28535 108285
rect 25535 105293 25543 108277
rect 28527 105293 28535 108277
rect 25535 105285 28535 105293
rect 28725 108277 31725 108285
rect 28725 105293 28733 108277
rect 31717 105293 31725 108277
rect 28725 105285 31725 105293
rect 31915 108277 34915 108285
rect 31915 105293 31923 108277
rect 34907 105293 34915 108277
rect 31915 105285 34915 105293
rect 35105 108277 38105 108285
rect 35105 105293 35113 108277
rect 38097 105293 38105 108277
rect 35105 105285 38105 105293
rect 38295 108277 41295 108285
rect 38295 105293 38303 108277
rect 41287 105293 41295 108277
rect 38295 105285 41295 105293
rect 41485 108277 44485 108285
rect 41485 105293 41493 108277
rect 44477 105293 44485 108277
rect 41485 105285 44485 105293
rect 44675 108277 47675 108285
rect 44675 105293 44683 108277
rect 47667 105293 47675 108277
rect 44675 105285 47675 105293
rect 47865 108277 50865 108285
rect 47865 105293 47873 108277
rect 50857 105293 50865 108277
rect 47865 105285 50865 105293
rect 51055 108277 54055 108285
rect 51055 105293 51063 108277
rect 54047 105293 54055 108277
rect 51055 105285 54055 105293
rect 54245 108277 57245 108285
rect 54245 105293 54253 108277
rect 57237 105293 57245 108277
rect 54245 105285 57245 105293
rect 57435 108277 60435 108285
rect 57435 105293 57443 108277
rect 60427 105293 60435 108277
rect 57435 105285 60435 105293
rect 60625 108277 63625 108285
rect 60625 105293 60633 108277
rect 63617 105293 63625 108277
rect 60625 105285 63625 105293
rect 63815 108277 66815 108285
rect 63815 105293 63823 108277
rect 66807 105293 66815 108277
rect 63815 105285 66815 105293
rect 67005 108277 70005 108285
rect 67005 105293 67013 108277
rect 69997 105293 70005 108277
rect 67005 105285 70005 105293
rect 70195 108277 73195 108285
rect 70195 105293 70203 108277
rect 73187 105293 73195 108277
rect 70195 105285 73195 105293
rect 73385 108277 76385 108285
rect 73385 105293 73393 108277
rect 76377 105293 76385 108277
rect 73385 105285 76385 105293
rect 76575 108277 79575 108285
rect 76575 105293 76583 108277
rect 79567 105293 79575 108277
rect 76575 105285 79575 105293
rect 79765 108277 82765 108285
rect 79765 105293 79773 108277
rect 82757 105293 82765 108277
rect 79765 105285 82765 105293
rect 82955 108277 85955 108285
rect 82955 105293 82963 108277
rect 85947 105293 85955 108277
rect 82955 105285 85955 105293
rect 86145 108277 89145 108285
rect 86145 105293 86153 108277
rect 89137 105293 89145 108277
rect 86145 105285 89145 105293
rect 89335 108277 92335 108285
rect 89335 105293 89343 108277
rect 92327 105293 92335 108277
rect 89335 105285 92335 105293
rect 92525 108277 95525 108285
rect 92525 105293 92533 108277
rect 95517 105293 95525 108277
rect 92525 105285 95525 105293
rect 95715 108277 98715 108285
rect 95715 105293 95723 108277
rect 98707 105293 98715 108277
rect 95715 105285 98715 105293
rect 98905 108277 101905 108285
rect 98905 105293 98913 108277
rect 101897 105293 101905 108277
rect 98905 105285 101905 105293
rect 102095 108277 105095 108285
rect 102095 105293 102103 108277
rect 105087 105293 105095 108277
rect 102095 105285 105095 105293
rect 105285 108277 108285 108285
rect 105285 105293 105293 108277
rect 108277 105293 108285 108277
rect 105285 105285 108285 105293
rect 108475 108277 111475 108285
rect 108475 105293 108483 108277
rect 111467 105293 111475 108277
rect 108475 105285 111475 105293
rect 111665 108277 114665 108285
rect 111665 105293 111673 108277
rect 114657 105293 114665 108277
rect 111665 105285 114665 105293
rect 114855 108277 117855 108285
rect 114855 105293 114863 108277
rect 117847 105293 117855 108277
rect 114855 105285 117855 105293
rect 118045 108277 121045 108285
rect 118045 105293 118053 108277
rect 121037 105293 121045 108277
rect 118045 105285 121045 105293
rect 121235 108277 124235 108285
rect 121235 105293 121243 108277
rect 124227 105293 124235 108277
rect 121235 105285 124235 105293
rect 124425 108277 127425 108285
rect 124425 105293 124433 108277
rect 127417 105293 127425 108277
rect 124425 105285 127425 105293
rect 127615 108277 130615 108285
rect 127615 105293 127623 108277
rect 130607 105293 130615 108277
rect 127615 105285 130615 105293
rect 130805 108277 133805 108285
rect 130805 105293 130813 108277
rect 133797 105293 133805 108277
rect 130805 105285 133805 105293
rect 133995 108277 136995 108285
rect 133995 105293 134003 108277
rect 136987 105293 136995 108277
rect 133995 105285 136995 105293
rect 15 105087 3015 105095
rect 15 102103 23 105087
rect 3007 102103 3015 105087
rect 15 102095 3015 102103
rect 3205 105087 6205 105095
rect 3205 102103 3213 105087
rect 6197 102103 6205 105087
rect 3205 102095 6205 102103
rect 6395 105087 9395 105095
rect 6395 102103 6403 105087
rect 9387 102103 9395 105087
rect 6395 102095 9395 102103
rect 9585 105087 12585 105095
rect 9585 102103 9593 105087
rect 12577 102103 12585 105087
rect 9585 102095 12585 102103
rect 12775 105087 15775 105095
rect 12775 102103 12783 105087
rect 15767 102103 15775 105087
rect 12775 102095 15775 102103
rect 15965 105087 18965 105095
rect 15965 102103 15973 105087
rect 18957 102103 18965 105087
rect 15965 102095 18965 102103
rect 19155 105087 22155 105095
rect 19155 102103 19163 105087
rect 22147 102103 22155 105087
rect 19155 102095 22155 102103
rect 22345 105087 25345 105095
rect 22345 102103 22353 105087
rect 25337 102103 25345 105087
rect 22345 102095 25345 102103
rect 25535 105087 28535 105095
rect 25535 102103 25543 105087
rect 28527 102103 28535 105087
rect 25535 102095 28535 102103
rect 28725 105087 31725 105095
rect 28725 102103 28733 105087
rect 31717 102103 31725 105087
rect 28725 102095 31725 102103
rect 31915 105087 34915 105095
rect 31915 102103 31923 105087
rect 34907 102103 34915 105087
rect 31915 102095 34915 102103
rect 35105 105087 38105 105095
rect 35105 102103 35113 105087
rect 38097 102103 38105 105087
rect 35105 102095 38105 102103
rect 38295 105087 41295 105095
rect 38295 102103 38303 105087
rect 41287 102103 41295 105087
rect 38295 102095 41295 102103
rect 41485 105087 44485 105095
rect 41485 102103 41493 105087
rect 44477 102103 44485 105087
rect 41485 102095 44485 102103
rect 44675 105087 47675 105095
rect 44675 102103 44683 105087
rect 47667 102103 47675 105087
rect 44675 102095 47675 102103
rect 47865 105087 50865 105095
rect 47865 102103 47873 105087
rect 50857 102103 50865 105087
rect 47865 102095 50865 102103
rect 51055 105087 54055 105095
rect 51055 102103 51063 105087
rect 54047 102103 54055 105087
rect 51055 102095 54055 102103
rect 54245 105087 57245 105095
rect 54245 102103 54253 105087
rect 57237 102103 57245 105087
rect 54245 102095 57245 102103
rect 57435 105087 60435 105095
rect 57435 102103 57443 105087
rect 60427 102103 60435 105087
rect 57435 102095 60435 102103
rect 60625 105087 63625 105095
rect 60625 102103 60633 105087
rect 63617 102103 63625 105087
rect 60625 102095 63625 102103
rect 63815 105087 66815 105095
rect 63815 102103 63823 105087
rect 66807 102103 66815 105087
rect 63815 102095 66815 102103
rect 67005 105087 70005 105095
rect 67005 102103 67013 105087
rect 69997 102103 70005 105087
rect 67005 102095 70005 102103
rect 70195 105087 73195 105095
rect 70195 102103 70203 105087
rect 73187 102103 73195 105087
rect 70195 102095 73195 102103
rect 73385 105087 76385 105095
rect 73385 102103 73393 105087
rect 76377 102103 76385 105087
rect 73385 102095 76385 102103
rect 76575 105087 79575 105095
rect 76575 102103 76583 105087
rect 79567 102103 79575 105087
rect 76575 102095 79575 102103
rect 79765 105087 82765 105095
rect 79765 102103 79773 105087
rect 82757 102103 82765 105087
rect 79765 102095 82765 102103
rect 82955 105087 85955 105095
rect 82955 102103 82963 105087
rect 85947 102103 85955 105087
rect 82955 102095 85955 102103
rect 86145 105087 89145 105095
rect 86145 102103 86153 105087
rect 89137 102103 89145 105087
rect 86145 102095 89145 102103
rect 89335 105087 92335 105095
rect 89335 102103 89343 105087
rect 92327 102103 92335 105087
rect 89335 102095 92335 102103
rect 92525 105087 95525 105095
rect 92525 102103 92533 105087
rect 95517 102103 95525 105087
rect 92525 102095 95525 102103
rect 95715 105087 98715 105095
rect 95715 102103 95723 105087
rect 98707 102103 98715 105087
rect 95715 102095 98715 102103
rect 98905 105087 101905 105095
rect 98905 102103 98913 105087
rect 101897 102103 101905 105087
rect 98905 102095 101905 102103
rect 102095 105087 105095 105095
rect 102095 102103 102103 105087
rect 105087 102103 105095 105087
rect 102095 102095 105095 102103
rect 105285 105087 108285 105095
rect 105285 102103 105293 105087
rect 108277 102103 108285 105087
rect 105285 102095 108285 102103
rect 108475 105087 111475 105095
rect 108475 102103 108483 105087
rect 111467 102103 111475 105087
rect 108475 102095 111475 102103
rect 111665 105087 114665 105095
rect 111665 102103 111673 105087
rect 114657 102103 114665 105087
rect 111665 102095 114665 102103
rect 114855 105087 117855 105095
rect 114855 102103 114863 105087
rect 117847 102103 117855 105087
rect 114855 102095 117855 102103
rect 118045 105087 121045 105095
rect 118045 102103 118053 105087
rect 121037 102103 121045 105087
rect 118045 102095 121045 102103
rect 121235 105087 124235 105095
rect 121235 102103 121243 105087
rect 124227 102103 124235 105087
rect 121235 102095 124235 102103
rect 124425 105087 127425 105095
rect 124425 102103 124433 105087
rect 127417 102103 127425 105087
rect 124425 102095 127425 102103
rect 127615 105087 130615 105095
rect 127615 102103 127623 105087
rect 130607 102103 130615 105087
rect 127615 102095 130615 102103
rect 130805 105087 133805 105095
rect 130805 102103 130813 105087
rect 133797 102103 133805 105087
rect 130805 102095 133805 102103
rect 133995 105087 136995 105095
rect 133995 102103 134003 105087
rect 136987 102103 136995 105087
rect 133995 102095 136995 102103
rect 15 101897 3015 101905
rect 15 98913 23 101897
rect 3007 98913 3015 101897
rect 15 98905 3015 98913
rect 3205 101897 6205 101905
rect 3205 98913 3213 101897
rect 6197 98913 6205 101897
rect 3205 98905 6205 98913
rect 6395 101897 9395 101905
rect 6395 98913 6403 101897
rect 9387 98913 9395 101897
rect 6395 98905 9395 98913
rect 9585 101897 12585 101905
rect 9585 98913 9593 101897
rect 12577 98913 12585 101897
rect 9585 98905 12585 98913
rect 12775 101897 15775 101905
rect 12775 98913 12783 101897
rect 15767 98913 15775 101897
rect 12775 98905 15775 98913
rect 15965 101897 18965 101905
rect 15965 98913 15973 101897
rect 18957 98913 18965 101897
rect 15965 98905 18965 98913
rect 19155 101897 22155 101905
rect 19155 98913 19163 101897
rect 22147 98913 22155 101897
rect 19155 98905 22155 98913
rect 22345 101897 25345 101905
rect 22345 98913 22353 101897
rect 25337 98913 25345 101897
rect 22345 98905 25345 98913
rect 25535 101897 28535 101905
rect 25535 98913 25543 101897
rect 28527 98913 28535 101897
rect 25535 98905 28535 98913
rect 28725 101897 31725 101905
rect 28725 98913 28733 101897
rect 31717 98913 31725 101897
rect 28725 98905 31725 98913
rect 31915 101897 34915 101905
rect 31915 98913 31923 101897
rect 34907 98913 34915 101897
rect 31915 98905 34915 98913
rect 35105 101897 38105 101905
rect 35105 98913 35113 101897
rect 38097 98913 38105 101897
rect 35105 98905 38105 98913
rect 38295 101897 41295 101905
rect 38295 98913 38303 101897
rect 41287 98913 41295 101897
rect 38295 98905 41295 98913
rect 41485 101897 44485 101905
rect 41485 98913 41493 101897
rect 44477 98913 44485 101897
rect 41485 98905 44485 98913
rect 44675 101897 47675 101905
rect 44675 98913 44683 101897
rect 47667 98913 47675 101897
rect 44675 98905 47675 98913
rect 47865 101897 50865 101905
rect 47865 98913 47873 101897
rect 50857 98913 50865 101897
rect 47865 98905 50865 98913
rect 51055 101897 54055 101905
rect 51055 98913 51063 101897
rect 54047 98913 54055 101897
rect 51055 98905 54055 98913
rect 54245 101897 57245 101905
rect 54245 98913 54253 101897
rect 57237 98913 57245 101897
rect 54245 98905 57245 98913
rect 57435 101897 60435 101905
rect 57435 98913 57443 101897
rect 60427 98913 60435 101897
rect 57435 98905 60435 98913
rect 60625 101897 63625 101905
rect 60625 98913 60633 101897
rect 63617 98913 63625 101897
rect 60625 98905 63625 98913
rect 63815 101897 66815 101905
rect 63815 98913 63823 101897
rect 66807 98913 66815 101897
rect 63815 98905 66815 98913
rect 67005 101897 70005 101905
rect 67005 98913 67013 101897
rect 69997 98913 70005 101897
rect 67005 98905 70005 98913
rect 70195 101897 73195 101905
rect 70195 98913 70203 101897
rect 73187 98913 73195 101897
rect 70195 98905 73195 98913
rect 73385 101897 76385 101905
rect 73385 98913 73393 101897
rect 76377 98913 76385 101897
rect 73385 98905 76385 98913
rect 76575 101897 79575 101905
rect 76575 98913 76583 101897
rect 79567 98913 79575 101897
rect 76575 98905 79575 98913
rect 79765 101897 82765 101905
rect 79765 98913 79773 101897
rect 82757 98913 82765 101897
rect 79765 98905 82765 98913
rect 82955 101897 85955 101905
rect 82955 98913 82963 101897
rect 85947 98913 85955 101897
rect 82955 98905 85955 98913
rect 86145 101897 89145 101905
rect 86145 98913 86153 101897
rect 89137 98913 89145 101897
rect 86145 98905 89145 98913
rect 89335 101897 92335 101905
rect 89335 98913 89343 101897
rect 92327 98913 92335 101897
rect 89335 98905 92335 98913
rect 92525 101897 95525 101905
rect 92525 98913 92533 101897
rect 95517 98913 95525 101897
rect 92525 98905 95525 98913
rect 95715 101897 98715 101905
rect 95715 98913 95723 101897
rect 98707 98913 98715 101897
rect 95715 98905 98715 98913
rect 98905 101897 101905 101905
rect 98905 98913 98913 101897
rect 101897 98913 101905 101897
rect 98905 98905 101905 98913
rect 102095 101897 105095 101905
rect 102095 98913 102103 101897
rect 105087 98913 105095 101897
rect 102095 98905 105095 98913
rect 105285 101897 108285 101905
rect 105285 98913 105293 101897
rect 108277 98913 108285 101897
rect 105285 98905 108285 98913
rect 108475 101897 111475 101905
rect 108475 98913 108483 101897
rect 111467 98913 111475 101897
rect 108475 98905 111475 98913
rect 111665 101897 114665 101905
rect 111665 98913 111673 101897
rect 114657 98913 114665 101897
rect 111665 98905 114665 98913
rect 114855 101897 117855 101905
rect 114855 98913 114863 101897
rect 117847 98913 117855 101897
rect 114855 98905 117855 98913
rect 118045 101897 121045 101905
rect 118045 98913 118053 101897
rect 121037 98913 121045 101897
rect 118045 98905 121045 98913
rect 121235 101897 124235 101905
rect 121235 98913 121243 101897
rect 124227 98913 124235 101897
rect 121235 98905 124235 98913
rect 124425 101897 127425 101905
rect 124425 98913 124433 101897
rect 127417 98913 127425 101897
rect 124425 98905 127425 98913
rect 127615 101897 130615 101905
rect 127615 98913 127623 101897
rect 130607 98913 130615 101897
rect 127615 98905 130615 98913
rect 130805 101897 133805 101905
rect 130805 98913 130813 101897
rect 133797 98913 133805 101897
rect 130805 98905 133805 98913
rect 133995 101897 136995 101905
rect 133995 98913 134003 101897
rect 136987 98913 136995 101897
rect 133995 98905 136995 98913
rect 9585 98707 12585 98715
rect 9585 95723 9593 98707
rect 12577 95723 12585 98707
rect 9585 95715 12585 95723
rect 12775 98707 15775 98715
rect 12775 95723 12783 98707
rect 15767 95723 15775 98707
rect 12775 95715 15775 95723
rect 15965 98707 18965 98715
rect 15965 95723 15973 98707
rect 18957 95723 18965 98707
rect 15965 95715 18965 95723
rect 19155 98707 22155 98715
rect 19155 95723 19163 98707
rect 22147 95723 22155 98707
rect 19155 95715 22155 95723
rect 22345 98707 25345 98715
rect 22345 95723 22353 98707
rect 25337 95723 25345 98707
rect 22345 95715 25345 95723
rect 25535 98707 28535 98715
rect 25535 95723 25543 98707
rect 28527 95723 28535 98707
rect 25535 95715 28535 95723
rect 28725 98707 31725 98715
rect 28725 95723 28733 98707
rect 31717 95723 31725 98707
rect 28725 95715 31725 95723
rect 31915 98707 34915 98715
rect 31915 95723 31923 98707
rect 34907 95723 34915 98707
rect 31915 95715 34915 95723
rect 35105 98707 38105 98715
rect 35105 95723 35113 98707
rect 38097 95723 38105 98707
rect 35105 95715 38105 95723
rect 38295 98707 41295 98715
rect 38295 95723 38303 98707
rect 41287 95723 41295 98707
rect 38295 95715 41295 95723
rect 41485 98707 44485 98715
rect 41485 95723 41493 98707
rect 44477 95723 44485 98707
rect 41485 95715 44485 95723
rect 44675 98707 47675 98715
rect 44675 95723 44683 98707
rect 47667 95723 47675 98707
rect 44675 95715 47675 95723
rect 47865 98707 50865 98715
rect 47865 95723 47873 98707
rect 50857 95723 50865 98707
rect 47865 95715 50865 95723
rect 51055 98707 54055 98715
rect 51055 95723 51063 98707
rect 54047 95723 54055 98707
rect 51055 95715 54055 95723
rect 54245 98707 57245 98715
rect 54245 95723 54253 98707
rect 57237 95723 57245 98707
rect 54245 95715 57245 95723
rect 57435 98707 60435 98715
rect 57435 95723 57443 98707
rect 60427 95723 60435 98707
rect 57435 95715 60435 95723
rect 60625 98707 63625 98715
rect 60625 95723 60633 98707
rect 63617 95723 63625 98707
rect 60625 95715 63625 95723
rect 63815 98707 66815 98715
rect 63815 95723 63823 98707
rect 66807 95723 66815 98707
rect 63815 95715 66815 95723
rect 67005 98707 70005 98715
rect 67005 95723 67013 98707
rect 69997 95723 70005 98707
rect 67005 95715 70005 95723
rect 70195 98707 73195 98715
rect 70195 95723 70203 98707
rect 73187 95723 73195 98707
rect 70195 95715 73195 95723
rect 73385 98707 76385 98715
rect 73385 95723 73393 98707
rect 76377 95723 76385 98707
rect 73385 95715 76385 95723
rect 76575 98707 79575 98715
rect 76575 95723 76583 98707
rect 79567 95723 79575 98707
rect 76575 95715 79575 95723
rect 79765 98707 82765 98715
rect 79765 95723 79773 98707
rect 82757 95723 82765 98707
rect 79765 95715 82765 95723
rect 82955 98707 85955 98715
rect 82955 95723 82963 98707
rect 85947 95723 85955 98707
rect 82955 95715 85955 95723
rect 86145 98707 89145 98715
rect 86145 95723 86153 98707
rect 89137 95723 89145 98707
rect 86145 95715 89145 95723
rect 89335 98707 92335 98715
rect 89335 95723 89343 98707
rect 92327 95723 92335 98707
rect 89335 95715 92335 95723
rect 92525 98707 95525 98715
rect 92525 95723 92533 98707
rect 95517 95723 95525 98707
rect 92525 95715 95525 95723
rect 95715 98707 98715 98715
rect 95715 95723 95723 98707
rect 98707 95723 98715 98707
rect 95715 95715 98715 95723
rect 98905 98707 101905 98715
rect 98905 95723 98913 98707
rect 101897 95723 101905 98707
rect 98905 95715 101905 95723
rect 102095 98707 105095 98715
rect 102095 95723 102103 98707
rect 105087 95723 105095 98707
rect 102095 95715 105095 95723
rect 105285 98707 108285 98715
rect 105285 95723 105293 98707
rect 108277 95723 108285 98707
rect 105285 95715 108285 95723
rect 108475 98707 111475 98715
rect 108475 95723 108483 98707
rect 111467 95723 111475 98707
rect 108475 95715 111475 95723
rect 111665 98707 114665 98715
rect 111665 95723 111673 98707
rect 114657 95723 114665 98707
rect 111665 95715 114665 95723
rect 114855 98707 117855 98715
rect 114855 95723 114863 98707
rect 117847 95723 117855 98707
rect 114855 95715 117855 95723
rect 118045 98707 121045 98715
rect 118045 95723 118053 98707
rect 121037 95723 121045 98707
rect 118045 95715 121045 95723
rect 121235 98707 124235 98715
rect 121235 95723 121243 98707
rect 124227 95723 124235 98707
rect 121235 95715 124235 95723
rect 124425 98707 127425 98715
rect 124425 95723 124433 98707
rect 127417 95723 127425 98707
rect 124425 95715 127425 95723
rect 127615 98707 130615 98715
rect 127615 95723 127623 98707
rect 130607 95723 130615 98707
rect 127615 95715 130615 95723
rect 130805 98707 133805 98715
rect 130805 95723 130813 98707
rect 133797 95723 133805 98707
rect 130805 95715 133805 95723
rect 133995 98707 136995 98715
rect 133995 95723 134003 98707
rect 136987 95723 136995 98707
rect 133995 95715 136995 95723
rect 9585 95517 12585 95525
rect 9585 92533 9593 95517
rect 12577 92533 12585 95517
rect 9585 92525 12585 92533
rect 12775 95517 15775 95525
rect 12775 92533 12783 95517
rect 15767 92533 15775 95517
rect 12775 92525 15775 92533
rect 15965 95517 18965 95525
rect 15965 92533 15973 95517
rect 18957 92533 18965 95517
rect 15965 92525 18965 92533
rect 19155 95517 22155 95525
rect 19155 92533 19163 95517
rect 22147 92533 22155 95517
rect 19155 92525 22155 92533
rect 22345 95517 25345 95525
rect 22345 92533 22353 95517
rect 25337 92533 25345 95517
rect 22345 92525 25345 92533
rect 25535 95517 28535 95525
rect 25535 92533 25543 95517
rect 28527 92533 28535 95517
rect 25535 92525 28535 92533
rect 28725 95517 31725 95525
rect 28725 92533 28733 95517
rect 31717 92533 31725 95517
rect 28725 92525 31725 92533
rect 31915 95517 34915 95525
rect 31915 92533 31923 95517
rect 34907 92533 34915 95517
rect 31915 92525 34915 92533
rect 35105 95517 38105 95525
rect 35105 92533 35113 95517
rect 38097 92533 38105 95517
rect 35105 92525 38105 92533
rect 38295 95517 41295 95525
rect 38295 92533 38303 95517
rect 41287 92533 41295 95517
rect 38295 92525 41295 92533
rect 41485 95517 44485 95525
rect 41485 92533 41493 95517
rect 44477 92533 44485 95517
rect 41485 92525 44485 92533
rect 44675 95517 47675 95525
rect 44675 92533 44683 95517
rect 47667 92533 47675 95517
rect 44675 92525 47675 92533
rect 47865 95517 50865 95525
rect 47865 92533 47873 95517
rect 50857 92533 50865 95517
rect 47865 92525 50865 92533
rect 51055 95517 54055 95525
rect 51055 92533 51063 95517
rect 54047 92533 54055 95517
rect 51055 92525 54055 92533
rect 54245 95517 57245 95525
rect 54245 92533 54253 95517
rect 57237 92533 57245 95517
rect 54245 92525 57245 92533
rect 57435 95517 60435 95525
rect 57435 92533 57443 95517
rect 60427 92533 60435 95517
rect 57435 92525 60435 92533
rect 60625 95517 63625 95525
rect 60625 92533 60633 95517
rect 63617 92533 63625 95517
rect 60625 92525 63625 92533
rect 63815 95517 66815 95525
rect 63815 92533 63823 95517
rect 66807 92533 66815 95517
rect 63815 92525 66815 92533
rect 67005 95517 70005 95525
rect 67005 92533 67013 95517
rect 69997 92533 70005 95517
rect 67005 92525 70005 92533
rect 70195 95517 73195 95525
rect 70195 92533 70203 95517
rect 73187 92533 73195 95517
rect 70195 92525 73195 92533
rect 73385 95517 76385 95525
rect 73385 92533 73393 95517
rect 76377 92533 76385 95517
rect 73385 92525 76385 92533
rect 76575 95517 79575 95525
rect 76575 92533 76583 95517
rect 79567 92533 79575 95517
rect 76575 92525 79575 92533
rect 79765 95517 82765 95525
rect 79765 92533 79773 95517
rect 82757 92533 82765 95517
rect 79765 92525 82765 92533
rect 82955 95517 85955 95525
rect 82955 92533 82963 95517
rect 85947 92533 85955 95517
rect 82955 92525 85955 92533
rect 86145 95517 89145 95525
rect 86145 92533 86153 95517
rect 89137 92533 89145 95517
rect 86145 92525 89145 92533
rect 89335 95517 92335 95525
rect 89335 92533 89343 95517
rect 92327 92533 92335 95517
rect 89335 92525 92335 92533
rect 92525 95517 95525 95525
rect 92525 92533 92533 95517
rect 95517 92533 95525 95517
rect 92525 92525 95525 92533
rect 95715 95517 98715 95525
rect 95715 92533 95723 95517
rect 98707 92533 98715 95517
rect 95715 92525 98715 92533
rect 98905 95517 101905 95525
rect 98905 92533 98913 95517
rect 101897 92533 101905 95517
rect 98905 92525 101905 92533
rect 102095 95517 105095 95525
rect 102095 92533 102103 95517
rect 105087 92533 105095 95517
rect 102095 92525 105095 92533
rect 105285 95517 108285 95525
rect 105285 92533 105293 95517
rect 108277 92533 108285 95517
rect 105285 92525 108285 92533
rect 108475 95517 111475 95525
rect 108475 92533 108483 95517
rect 111467 92533 111475 95517
rect 108475 92525 111475 92533
rect 111665 95517 114665 95525
rect 111665 92533 111673 95517
rect 114657 92533 114665 95517
rect 111665 92525 114665 92533
rect 114855 95517 117855 95525
rect 114855 92533 114863 95517
rect 117847 92533 117855 95517
rect 114855 92525 117855 92533
rect 118045 95517 121045 95525
rect 118045 92533 118053 95517
rect 121037 92533 121045 95517
rect 118045 92525 121045 92533
rect 121235 95517 124235 95525
rect 121235 92533 121243 95517
rect 124227 92533 124235 95517
rect 121235 92525 124235 92533
rect 124425 95517 127425 95525
rect 124425 92533 124433 95517
rect 127417 92533 127425 95517
rect 124425 92525 127425 92533
rect 127615 95517 130615 95525
rect 127615 92533 127623 95517
rect 130607 92533 130615 95517
rect 127615 92525 130615 92533
rect 130805 95517 133805 95525
rect 130805 92533 130813 95517
rect 133797 92533 133805 95517
rect 130805 92525 133805 92533
rect 133995 95517 136995 95525
rect 133995 92533 134003 95517
rect 136987 92533 136995 95517
rect 133995 92525 136995 92533
rect 9585 92327 12585 92335
rect 9585 89343 9593 92327
rect 12577 89343 12585 92327
rect 9585 89335 12585 89343
rect 12775 92327 15775 92335
rect 12775 89343 12783 92327
rect 15767 89343 15775 92327
rect 12775 89335 15775 89343
rect 15965 92327 18965 92335
rect 15965 89343 15973 92327
rect 18957 89343 18965 92327
rect 15965 89335 18965 89343
rect 19155 92327 22155 92335
rect 19155 89343 19163 92327
rect 22147 89343 22155 92327
rect 19155 89335 22155 89343
rect 22345 92327 25345 92335
rect 22345 89343 22353 92327
rect 25337 89343 25345 92327
rect 22345 89335 25345 89343
rect 25535 92327 28535 92335
rect 25535 89343 25543 92327
rect 28527 89343 28535 92327
rect 25535 89335 28535 89343
rect 28725 92327 31725 92335
rect 28725 89343 28733 92327
rect 31717 89343 31725 92327
rect 28725 89335 31725 89343
rect 31915 92327 34915 92335
rect 31915 89343 31923 92327
rect 34907 89343 34915 92327
rect 31915 89335 34915 89343
rect 35105 92327 38105 92335
rect 35105 89343 35113 92327
rect 38097 89343 38105 92327
rect 35105 89335 38105 89343
rect 38295 92327 41295 92335
rect 38295 89343 38303 92327
rect 41287 89343 41295 92327
rect 38295 89335 41295 89343
rect 41485 92327 44485 92335
rect 41485 89343 41493 92327
rect 44477 89343 44485 92327
rect 41485 89335 44485 89343
rect 44675 92327 47675 92335
rect 44675 89343 44683 92327
rect 47667 89343 47675 92327
rect 44675 89335 47675 89343
rect 47865 92327 50865 92335
rect 47865 89343 47873 92327
rect 50857 89343 50865 92327
rect 47865 89335 50865 89343
rect 51055 92327 54055 92335
rect 51055 89343 51063 92327
rect 54047 89343 54055 92327
rect 51055 89335 54055 89343
rect 54245 92327 57245 92335
rect 54245 89343 54253 92327
rect 57237 89343 57245 92327
rect 54245 89335 57245 89343
rect 57435 92327 60435 92335
rect 57435 89343 57443 92327
rect 60427 89343 60435 92327
rect 57435 89335 60435 89343
rect 60625 92327 63625 92335
rect 60625 89343 60633 92327
rect 63617 89343 63625 92327
rect 60625 89335 63625 89343
rect 63815 92327 66815 92335
rect 63815 89343 63823 92327
rect 66807 89343 66815 92327
rect 63815 89335 66815 89343
rect 67005 92327 70005 92335
rect 67005 89343 67013 92327
rect 69997 89343 70005 92327
rect 67005 89335 70005 89343
rect 70195 92327 73195 92335
rect 70195 89343 70203 92327
rect 73187 89343 73195 92327
rect 70195 89335 73195 89343
rect 73385 92327 76385 92335
rect 73385 89343 73393 92327
rect 76377 89343 76385 92327
rect 73385 89335 76385 89343
rect 76575 92327 79575 92335
rect 76575 89343 76583 92327
rect 79567 89343 79575 92327
rect 76575 89335 79575 89343
rect 79765 92327 82765 92335
rect 79765 89343 79773 92327
rect 82757 89343 82765 92327
rect 79765 89335 82765 89343
rect 82955 92327 85955 92335
rect 82955 89343 82963 92327
rect 85947 89343 85955 92327
rect 82955 89335 85955 89343
rect 86145 92327 89145 92335
rect 86145 89343 86153 92327
rect 89137 89343 89145 92327
rect 86145 89335 89145 89343
rect 89335 92327 92335 92335
rect 89335 89343 89343 92327
rect 92327 89343 92335 92327
rect 89335 89335 92335 89343
rect 92525 92327 95525 92335
rect 92525 89343 92533 92327
rect 95517 89343 95525 92327
rect 92525 89335 95525 89343
rect 95715 92327 98715 92335
rect 95715 89343 95723 92327
rect 98707 89343 98715 92327
rect 95715 89335 98715 89343
rect 98905 92327 101905 92335
rect 98905 89343 98913 92327
rect 101897 89343 101905 92327
rect 98905 89335 101905 89343
rect 102095 92327 105095 92335
rect 102095 89343 102103 92327
rect 105087 89343 105095 92327
rect 102095 89335 105095 89343
rect 105285 92327 108285 92335
rect 105285 89343 105293 92327
rect 108277 89343 108285 92327
rect 105285 89335 108285 89343
rect 108475 92327 111475 92335
rect 108475 89343 108483 92327
rect 111467 89343 111475 92327
rect 108475 89335 111475 89343
rect 111665 92327 114665 92335
rect 111665 89343 111673 92327
rect 114657 89343 114665 92327
rect 111665 89335 114665 89343
rect 114855 92327 117855 92335
rect 114855 89343 114863 92327
rect 117847 89343 117855 92327
rect 114855 89335 117855 89343
rect 118045 92327 121045 92335
rect 118045 89343 118053 92327
rect 121037 89343 121045 92327
rect 118045 89335 121045 89343
rect 121235 92327 124235 92335
rect 121235 89343 121243 92327
rect 124227 89343 124235 92327
rect 121235 89335 124235 89343
rect 124425 92327 127425 92335
rect 124425 89343 124433 92327
rect 127417 89343 127425 92327
rect 124425 89335 127425 89343
rect 127615 92327 130615 92335
rect 127615 89343 127623 92327
rect 130607 89343 130615 92327
rect 127615 89335 130615 89343
rect 130805 92327 133805 92335
rect 130805 89343 130813 92327
rect 133797 89343 133805 92327
rect 130805 89335 133805 89343
rect 133995 92327 136995 92335
rect 133995 89343 134003 92327
rect 136987 89343 136995 92327
rect 133995 89335 136995 89343
rect 9585 89137 12585 89145
rect 9585 86153 9593 89137
rect 12577 86153 12585 89137
rect 9585 86145 12585 86153
rect 12775 89137 15775 89145
rect 12775 86153 12783 89137
rect 15767 86153 15775 89137
rect 12775 86145 15775 86153
rect 15965 89137 18965 89145
rect 15965 86153 15973 89137
rect 18957 86153 18965 89137
rect 15965 86145 18965 86153
rect 19155 89137 22155 89145
rect 19155 86153 19163 89137
rect 22147 86153 22155 89137
rect 19155 86145 22155 86153
rect 22345 89137 25345 89145
rect 22345 86153 22353 89137
rect 25337 86153 25345 89137
rect 22345 86145 25345 86153
rect 25535 89137 28535 89145
rect 25535 86153 25543 89137
rect 28527 86153 28535 89137
rect 25535 86145 28535 86153
rect 28725 89137 31725 89145
rect 28725 86153 28733 89137
rect 31717 86153 31725 89137
rect 28725 86145 31725 86153
rect 31915 89137 34915 89145
rect 31915 86153 31923 89137
rect 34907 86153 34915 89137
rect 31915 86145 34915 86153
rect 35105 89137 38105 89145
rect 35105 86153 35113 89137
rect 38097 86153 38105 89137
rect 35105 86145 38105 86153
rect 38295 89137 41295 89145
rect 38295 86153 38303 89137
rect 41287 86153 41295 89137
rect 38295 86145 41295 86153
rect 41485 89137 44485 89145
rect 41485 86153 41493 89137
rect 44477 86153 44485 89137
rect 41485 86145 44485 86153
rect 44675 89137 47675 89145
rect 44675 86153 44683 89137
rect 47667 86153 47675 89137
rect 44675 86145 47675 86153
rect 47865 89137 50865 89145
rect 47865 86153 47873 89137
rect 50857 86153 50865 89137
rect 47865 86145 50865 86153
rect 51055 89137 54055 89145
rect 51055 86153 51063 89137
rect 54047 86153 54055 89137
rect 51055 86145 54055 86153
rect 54245 89137 57245 89145
rect 54245 86153 54253 89137
rect 57237 86153 57245 89137
rect 54245 86145 57245 86153
rect 57435 89137 60435 89145
rect 57435 86153 57443 89137
rect 60427 86153 60435 89137
rect 57435 86145 60435 86153
rect 60625 89137 63625 89145
rect 60625 86153 60633 89137
rect 63617 86153 63625 89137
rect 60625 86145 63625 86153
rect 63815 89137 66815 89145
rect 63815 86153 63823 89137
rect 66807 86153 66815 89137
rect 63815 86145 66815 86153
rect 67005 89137 70005 89145
rect 67005 86153 67013 89137
rect 69997 86153 70005 89137
rect 67005 86145 70005 86153
rect 70195 89137 73195 89145
rect 70195 86153 70203 89137
rect 73187 86153 73195 89137
rect 70195 86145 73195 86153
rect 73385 89137 76385 89145
rect 73385 86153 73393 89137
rect 76377 86153 76385 89137
rect 73385 86145 76385 86153
rect 76575 89137 79575 89145
rect 76575 86153 76583 89137
rect 79567 86153 79575 89137
rect 76575 86145 79575 86153
rect 79765 89137 82765 89145
rect 79765 86153 79773 89137
rect 82757 86153 82765 89137
rect 79765 86145 82765 86153
rect 82955 89137 85955 89145
rect 82955 86153 82963 89137
rect 85947 86153 85955 89137
rect 82955 86145 85955 86153
rect 86145 89137 89145 89145
rect 86145 86153 86153 89137
rect 89137 86153 89145 89137
rect 86145 86145 89145 86153
rect 89335 89137 92335 89145
rect 89335 86153 89343 89137
rect 92327 86153 92335 89137
rect 89335 86145 92335 86153
rect 92525 89137 95525 89145
rect 92525 86153 92533 89137
rect 95517 86153 95525 89137
rect 92525 86145 95525 86153
rect 95715 89137 98715 89145
rect 95715 86153 95723 89137
rect 98707 86153 98715 89137
rect 95715 86145 98715 86153
rect 98905 89137 101905 89145
rect 98905 86153 98913 89137
rect 101897 86153 101905 89137
rect 98905 86145 101905 86153
rect 102095 89137 105095 89145
rect 102095 86153 102103 89137
rect 105087 86153 105095 89137
rect 102095 86145 105095 86153
rect 105285 89137 108285 89145
rect 105285 86153 105293 89137
rect 108277 86153 108285 89137
rect 105285 86145 108285 86153
rect 108475 89137 111475 89145
rect 108475 86153 108483 89137
rect 111467 86153 111475 89137
rect 108475 86145 111475 86153
rect 111665 89137 114665 89145
rect 111665 86153 111673 89137
rect 114657 86153 114665 89137
rect 111665 86145 114665 86153
rect 114855 89137 117855 89145
rect 114855 86153 114863 89137
rect 117847 86153 117855 89137
rect 114855 86145 117855 86153
rect 118045 89137 121045 89145
rect 118045 86153 118053 89137
rect 121037 86153 121045 89137
rect 118045 86145 121045 86153
rect 121235 89137 124235 89145
rect 121235 86153 121243 89137
rect 124227 86153 124235 89137
rect 121235 86145 124235 86153
rect 124425 89137 127425 89145
rect 124425 86153 124433 89137
rect 127417 86153 127425 89137
rect 124425 86145 127425 86153
rect 127615 89137 130615 89145
rect 127615 86153 127623 89137
rect 130607 86153 130615 89137
rect 127615 86145 130615 86153
rect 130805 89137 133805 89145
rect 130805 86153 130813 89137
rect 133797 86153 133805 89137
rect 130805 86145 133805 86153
rect 133995 89137 136995 89145
rect 133995 86153 134003 89137
rect 136987 86153 136995 89137
rect 133995 86145 136995 86153
rect 9585 85947 12585 85955
rect 9585 82963 9593 85947
rect 12577 82963 12585 85947
rect 9585 82955 12585 82963
rect 12775 85947 15775 85955
rect 12775 82963 12783 85947
rect 15767 82963 15775 85947
rect 12775 82955 15775 82963
rect 15965 85947 18965 85955
rect 15965 82963 15973 85947
rect 18957 82963 18965 85947
rect 15965 82955 18965 82963
rect 19155 85947 22155 85955
rect 19155 82963 19163 85947
rect 22147 82963 22155 85947
rect 19155 82955 22155 82963
rect 22345 85947 25345 85955
rect 22345 82963 22353 85947
rect 25337 82963 25345 85947
rect 22345 82955 25345 82963
rect 25535 85947 28535 85955
rect 25535 82963 25543 85947
rect 28527 82963 28535 85947
rect 25535 82955 28535 82963
rect 28725 85947 31725 85955
rect 28725 82963 28733 85947
rect 31717 82963 31725 85947
rect 28725 82955 31725 82963
rect 31915 85947 34915 85955
rect 31915 82963 31923 85947
rect 34907 82963 34915 85947
rect 31915 82955 34915 82963
rect 35105 85947 38105 85955
rect 35105 82963 35113 85947
rect 38097 82963 38105 85947
rect 35105 82955 38105 82963
rect 38295 85947 41295 85955
rect 38295 82963 38303 85947
rect 41287 82963 41295 85947
rect 38295 82955 41295 82963
rect 41485 85947 44485 85955
rect 41485 82963 41493 85947
rect 44477 82963 44485 85947
rect 41485 82955 44485 82963
rect 44675 85947 47675 85955
rect 44675 82963 44683 85947
rect 47667 82963 47675 85947
rect 44675 82955 47675 82963
rect 47865 85947 50865 85955
rect 47865 82963 47873 85947
rect 50857 82963 50865 85947
rect 47865 82955 50865 82963
rect 51055 85947 54055 85955
rect 51055 82963 51063 85947
rect 54047 82963 54055 85947
rect 51055 82955 54055 82963
rect 54245 85947 57245 85955
rect 54245 82963 54253 85947
rect 57237 82963 57245 85947
rect 54245 82955 57245 82963
rect 57435 85947 60435 85955
rect 57435 82963 57443 85947
rect 60427 82963 60435 85947
rect 57435 82955 60435 82963
rect 60625 85947 63625 85955
rect 60625 82963 60633 85947
rect 63617 82963 63625 85947
rect 60625 82955 63625 82963
rect 63815 85947 66815 85955
rect 63815 82963 63823 85947
rect 66807 82963 66815 85947
rect 63815 82955 66815 82963
rect 67005 85947 70005 85955
rect 67005 82963 67013 85947
rect 69997 82963 70005 85947
rect 67005 82955 70005 82963
rect 70195 85947 73195 85955
rect 70195 82963 70203 85947
rect 73187 82963 73195 85947
rect 70195 82955 73195 82963
rect 73385 85947 76385 85955
rect 73385 82963 73393 85947
rect 76377 82963 76385 85947
rect 73385 82955 76385 82963
rect 76575 85947 79575 85955
rect 76575 82963 76583 85947
rect 79567 82963 79575 85947
rect 76575 82955 79575 82963
rect 79765 85947 82765 85955
rect 79765 82963 79773 85947
rect 82757 82963 82765 85947
rect 79765 82955 82765 82963
rect 82955 85947 85955 85955
rect 82955 82963 82963 85947
rect 85947 82963 85955 85947
rect 82955 82955 85955 82963
rect 86145 85947 89145 85955
rect 86145 82963 86153 85947
rect 89137 82963 89145 85947
rect 86145 82955 89145 82963
rect 89335 85947 92335 85955
rect 89335 82963 89343 85947
rect 92327 82963 92335 85947
rect 89335 82955 92335 82963
rect 92525 85947 95525 85955
rect 92525 82963 92533 85947
rect 95517 82963 95525 85947
rect 92525 82955 95525 82963
rect 95715 85947 98715 85955
rect 95715 82963 95723 85947
rect 98707 82963 98715 85947
rect 95715 82955 98715 82963
rect 98905 85947 101905 85955
rect 98905 82963 98913 85947
rect 101897 82963 101905 85947
rect 98905 82955 101905 82963
rect 102095 85947 105095 85955
rect 102095 82963 102103 85947
rect 105087 82963 105095 85947
rect 102095 82955 105095 82963
rect 105285 85947 108285 85955
rect 105285 82963 105293 85947
rect 108277 82963 108285 85947
rect 105285 82955 108285 82963
rect 108475 85947 111475 85955
rect 108475 82963 108483 85947
rect 111467 82963 111475 85947
rect 108475 82955 111475 82963
rect 111665 85947 114665 85955
rect 111665 82963 111673 85947
rect 114657 82963 114665 85947
rect 111665 82955 114665 82963
rect 114855 85947 117855 85955
rect 114855 82963 114863 85947
rect 117847 82963 117855 85947
rect 114855 82955 117855 82963
rect 118045 85947 121045 85955
rect 118045 82963 118053 85947
rect 121037 82963 121045 85947
rect 118045 82955 121045 82963
rect 121235 85947 124235 85955
rect 121235 82963 121243 85947
rect 124227 82963 124235 85947
rect 121235 82955 124235 82963
rect 124425 85947 127425 85955
rect 124425 82963 124433 85947
rect 127417 82963 127425 85947
rect 124425 82955 127425 82963
rect 127615 85947 130615 85955
rect 127615 82963 127623 85947
rect 130607 82963 130615 85947
rect 127615 82955 130615 82963
rect 130805 85947 133805 85955
rect 130805 82963 130813 85947
rect 133797 82963 133805 85947
rect 130805 82955 133805 82963
rect 133995 85947 136995 85955
rect 133995 82963 134003 85947
rect 136987 82963 136995 85947
rect 133995 82955 136995 82963
rect 9585 82757 12585 82765
rect 9585 79773 9593 82757
rect 12577 79773 12585 82757
rect 9585 79765 12585 79773
rect 12775 82757 15775 82765
rect 12775 79773 12783 82757
rect 15767 79773 15775 82757
rect 12775 79765 15775 79773
rect 15965 82757 18965 82765
rect 15965 79773 15973 82757
rect 18957 79773 18965 82757
rect 15965 79765 18965 79773
rect 19155 82757 22155 82765
rect 19155 79773 19163 82757
rect 22147 79773 22155 82757
rect 19155 79765 22155 79773
rect 22345 82757 25345 82765
rect 22345 79773 22353 82757
rect 25337 79773 25345 82757
rect 22345 79765 25345 79773
rect 25535 82757 28535 82765
rect 25535 79773 25543 82757
rect 28527 79773 28535 82757
rect 25535 79765 28535 79773
rect 28725 82757 31725 82765
rect 28725 79773 28733 82757
rect 31717 79773 31725 82757
rect 28725 79765 31725 79773
rect 31915 82757 34915 82765
rect 31915 79773 31923 82757
rect 34907 79773 34915 82757
rect 31915 79765 34915 79773
rect 35105 82757 38105 82765
rect 35105 79773 35113 82757
rect 38097 79773 38105 82757
rect 35105 79765 38105 79773
rect 38295 82757 41295 82765
rect 38295 79773 38303 82757
rect 41287 79773 41295 82757
rect 38295 79765 41295 79773
rect 41485 82757 44485 82765
rect 41485 79773 41493 82757
rect 44477 79773 44485 82757
rect 41485 79765 44485 79773
rect 44675 82757 47675 82765
rect 44675 79773 44683 82757
rect 47667 79773 47675 82757
rect 44675 79765 47675 79773
rect 47865 82757 50865 82765
rect 47865 79773 47873 82757
rect 50857 79773 50865 82757
rect 47865 79765 50865 79773
rect 51055 82757 54055 82765
rect 51055 79773 51063 82757
rect 54047 79773 54055 82757
rect 51055 79765 54055 79773
rect 54245 82757 57245 82765
rect 54245 79773 54253 82757
rect 57237 79773 57245 82757
rect 54245 79765 57245 79773
rect 57435 82757 60435 82765
rect 57435 79773 57443 82757
rect 60427 79773 60435 82757
rect 57435 79765 60435 79773
rect 60625 82757 63625 82765
rect 60625 79773 60633 82757
rect 63617 79773 63625 82757
rect 60625 79765 63625 79773
rect 63815 82757 66815 82765
rect 63815 79773 63823 82757
rect 66807 79773 66815 82757
rect 63815 79765 66815 79773
rect 67005 82757 70005 82765
rect 67005 79773 67013 82757
rect 69997 79773 70005 82757
rect 67005 79765 70005 79773
rect 70195 82757 73195 82765
rect 70195 79773 70203 82757
rect 73187 79773 73195 82757
rect 70195 79765 73195 79773
rect 73385 82757 76385 82765
rect 73385 79773 73393 82757
rect 76377 79773 76385 82757
rect 73385 79765 76385 79773
rect 76575 82757 79575 82765
rect 76575 79773 76583 82757
rect 79567 79773 79575 82757
rect 76575 79765 79575 79773
rect 79765 82757 82765 82765
rect 79765 79773 79773 82757
rect 82757 79773 82765 82757
rect 79765 79765 82765 79773
rect 82955 82757 85955 82765
rect 82955 79773 82963 82757
rect 85947 79773 85955 82757
rect 82955 79765 85955 79773
rect 86145 82757 89145 82765
rect 86145 79773 86153 82757
rect 89137 79773 89145 82757
rect 86145 79765 89145 79773
rect 89335 82757 92335 82765
rect 89335 79773 89343 82757
rect 92327 79773 92335 82757
rect 89335 79765 92335 79773
rect 92525 82757 95525 82765
rect 92525 79773 92533 82757
rect 95517 79773 95525 82757
rect 92525 79765 95525 79773
rect 95715 82757 98715 82765
rect 95715 79773 95723 82757
rect 98707 79773 98715 82757
rect 95715 79765 98715 79773
rect 98905 82757 101905 82765
rect 98905 79773 98913 82757
rect 101897 79773 101905 82757
rect 98905 79765 101905 79773
rect 102095 82757 105095 82765
rect 102095 79773 102103 82757
rect 105087 79773 105095 82757
rect 102095 79765 105095 79773
rect 105285 82757 108285 82765
rect 105285 79773 105293 82757
rect 108277 79773 108285 82757
rect 105285 79765 108285 79773
rect 108475 82757 111475 82765
rect 108475 79773 108483 82757
rect 111467 79773 111475 82757
rect 108475 79765 111475 79773
rect 111665 82757 114665 82765
rect 111665 79773 111673 82757
rect 114657 79773 114665 82757
rect 111665 79765 114665 79773
rect 114855 82757 117855 82765
rect 114855 79773 114863 82757
rect 117847 79773 117855 82757
rect 114855 79765 117855 79773
rect 118045 82757 121045 82765
rect 118045 79773 118053 82757
rect 121037 79773 121045 82757
rect 118045 79765 121045 79773
rect 121235 82757 124235 82765
rect 121235 79773 121243 82757
rect 124227 79773 124235 82757
rect 121235 79765 124235 79773
rect 124425 82757 127425 82765
rect 124425 79773 124433 82757
rect 127417 79773 127425 82757
rect 124425 79765 127425 79773
rect 127615 82757 130615 82765
rect 127615 79773 127623 82757
rect 130607 79773 130615 82757
rect 127615 79765 130615 79773
rect 130805 82757 133805 82765
rect 130805 79773 130813 82757
rect 133797 79773 133805 82757
rect 130805 79765 133805 79773
rect 133995 82757 136995 82765
rect 133995 79773 134003 82757
rect 136987 79773 136995 82757
rect 133995 79765 136995 79773
rect 15 79567 3015 79575
rect 15 76583 23 79567
rect 3007 76583 3015 79567
rect 15 76575 3015 76583
rect 3205 79567 6205 79575
rect 3205 76583 3213 79567
rect 6197 76583 6205 79567
rect 3205 76575 6205 76583
rect 6395 79567 9395 79575
rect 6395 76583 6403 79567
rect 9387 76583 9395 79567
rect 6395 76575 9395 76583
rect 9585 79567 12585 79575
rect 9585 76583 9593 79567
rect 12577 76583 12585 79567
rect 9585 76575 12585 76583
rect 12775 79567 15775 79575
rect 12775 76583 12783 79567
rect 15767 76583 15775 79567
rect 12775 76575 15775 76583
rect 15965 79567 18965 79575
rect 15965 76583 15973 79567
rect 18957 76583 18965 79567
rect 15965 76575 18965 76583
rect 19155 79567 22155 79575
rect 19155 76583 19163 79567
rect 22147 76583 22155 79567
rect 19155 76575 22155 76583
rect 22345 79567 25345 79575
rect 22345 76583 22353 79567
rect 25337 76583 25345 79567
rect 22345 76575 25345 76583
rect 25535 79567 28535 79575
rect 25535 76583 25543 79567
rect 28527 76583 28535 79567
rect 25535 76575 28535 76583
rect 28725 79567 31725 79575
rect 28725 76583 28733 79567
rect 31717 76583 31725 79567
rect 28725 76575 31725 76583
rect 31915 79567 34915 79575
rect 31915 76583 31923 79567
rect 34907 76583 34915 79567
rect 31915 76575 34915 76583
rect 35105 79567 38105 79575
rect 35105 76583 35113 79567
rect 38097 76583 38105 79567
rect 35105 76575 38105 76583
rect 38295 79567 41295 79575
rect 38295 76583 38303 79567
rect 41287 76583 41295 79567
rect 38295 76575 41295 76583
rect 41485 79567 44485 79575
rect 41485 76583 41493 79567
rect 44477 76583 44485 79567
rect 41485 76575 44485 76583
rect 44675 79567 47675 79575
rect 44675 76583 44683 79567
rect 47667 76583 47675 79567
rect 44675 76575 47675 76583
rect 47865 79567 50865 79575
rect 47865 76583 47873 79567
rect 50857 76583 50865 79567
rect 47865 76575 50865 76583
rect 51055 79567 54055 79575
rect 51055 76583 51063 79567
rect 54047 76583 54055 79567
rect 51055 76575 54055 76583
rect 54245 79567 57245 79575
rect 54245 76583 54253 79567
rect 57237 76583 57245 79567
rect 54245 76575 57245 76583
rect 57435 79567 60435 79575
rect 57435 76583 57443 79567
rect 60427 76583 60435 79567
rect 57435 76575 60435 76583
rect 60625 79567 63625 79575
rect 60625 76583 60633 79567
rect 63617 76583 63625 79567
rect 60625 76575 63625 76583
rect 63815 79567 66815 79575
rect 63815 76583 63823 79567
rect 66807 76583 66815 79567
rect 63815 76575 66815 76583
rect 67005 79567 70005 79575
rect 67005 76583 67013 79567
rect 69997 76583 70005 79567
rect 67005 76575 70005 76583
rect 70195 79567 73195 79575
rect 70195 76583 70203 79567
rect 73187 76583 73195 79567
rect 70195 76575 73195 76583
rect 73385 79567 76385 79575
rect 73385 76583 73393 79567
rect 76377 76583 76385 79567
rect 73385 76575 76385 76583
rect 76575 79567 79575 79575
rect 76575 76583 76583 79567
rect 79567 76583 79575 79567
rect 76575 76575 79575 76583
rect 79765 79567 82765 79575
rect 79765 76583 79773 79567
rect 82757 76583 82765 79567
rect 79765 76575 82765 76583
rect 82955 79567 85955 79575
rect 82955 76583 82963 79567
rect 85947 76583 85955 79567
rect 82955 76575 85955 76583
rect 86145 79567 89145 79575
rect 86145 76583 86153 79567
rect 89137 76583 89145 79567
rect 86145 76575 89145 76583
rect 89335 79567 92335 79575
rect 89335 76583 89343 79567
rect 92327 76583 92335 79567
rect 89335 76575 92335 76583
rect 92525 79567 95525 79575
rect 92525 76583 92533 79567
rect 95517 76583 95525 79567
rect 92525 76575 95525 76583
rect 95715 79567 98715 79575
rect 95715 76583 95723 79567
rect 98707 76583 98715 79567
rect 95715 76575 98715 76583
rect 98905 79567 101905 79575
rect 98905 76583 98913 79567
rect 101897 76583 101905 79567
rect 98905 76575 101905 76583
rect 102095 79567 105095 79575
rect 102095 76583 102103 79567
rect 105087 76583 105095 79567
rect 102095 76575 105095 76583
rect 105285 79567 108285 79575
rect 105285 76583 105293 79567
rect 108277 76583 108285 79567
rect 105285 76575 108285 76583
rect 108475 79567 111475 79575
rect 108475 76583 108483 79567
rect 111467 76583 111475 79567
rect 108475 76575 111475 76583
rect 111665 79567 114665 79575
rect 111665 76583 111673 79567
rect 114657 76583 114665 79567
rect 111665 76575 114665 76583
rect 114855 79567 117855 79575
rect 114855 76583 114863 79567
rect 117847 76583 117855 79567
rect 114855 76575 117855 76583
rect 118045 79567 121045 79575
rect 118045 76583 118053 79567
rect 121037 76583 121045 79567
rect 118045 76575 121045 76583
rect 121235 79567 124235 79575
rect 121235 76583 121243 79567
rect 124227 76583 124235 79567
rect 121235 76575 124235 76583
rect 124425 79567 127425 79575
rect 124425 76583 124433 79567
rect 127417 76583 127425 79567
rect 124425 76575 127425 76583
rect 127615 79567 130615 79575
rect 127615 76583 127623 79567
rect 130607 76583 130615 79567
rect 127615 76575 130615 76583
rect 130805 79567 133805 79575
rect 130805 76583 130813 79567
rect 133797 76583 133805 79567
rect 130805 76575 133805 76583
rect 133995 79567 136995 79575
rect 133995 76583 134003 79567
rect 136987 76583 136995 79567
rect 133995 76575 136995 76583
rect 15 76377 3015 76385
rect 15 73393 23 76377
rect 3007 73393 3015 76377
rect 15 73385 3015 73393
rect 3205 76377 6205 76385
rect 3205 73393 3213 76377
rect 6197 73393 6205 76377
rect 3205 73385 6205 73393
rect 6395 76377 9395 76385
rect 6395 73393 6403 76377
rect 9387 73393 9395 76377
rect 6395 73385 9395 73393
rect 9585 76377 12585 76385
rect 9585 73393 9593 76377
rect 12577 73393 12585 76377
rect 9585 73385 12585 73393
rect 12775 76377 15775 76385
rect 12775 73393 12783 76377
rect 15767 73393 15775 76377
rect 12775 73385 15775 73393
rect 15965 76377 18965 76385
rect 15965 73393 15973 76377
rect 18957 73393 18965 76377
rect 15965 73385 18965 73393
rect 19155 76377 22155 76385
rect 19155 73393 19163 76377
rect 22147 73393 22155 76377
rect 19155 73385 22155 73393
rect 22345 76377 25345 76385
rect 22345 73393 22353 76377
rect 25337 73393 25345 76377
rect 22345 73385 25345 73393
rect 25535 76377 28535 76385
rect 25535 73393 25543 76377
rect 28527 73393 28535 76377
rect 25535 73385 28535 73393
rect 28725 76377 31725 76385
rect 28725 73393 28733 76377
rect 31717 73393 31725 76377
rect 28725 73385 31725 73393
rect 31915 76377 34915 76385
rect 31915 73393 31923 76377
rect 34907 73393 34915 76377
rect 31915 73385 34915 73393
rect 35105 76377 38105 76385
rect 35105 73393 35113 76377
rect 38097 73393 38105 76377
rect 35105 73385 38105 73393
rect 38295 76377 41295 76385
rect 38295 73393 38303 76377
rect 41287 73393 41295 76377
rect 38295 73385 41295 73393
rect 41485 76377 44485 76385
rect 41485 73393 41493 76377
rect 44477 73393 44485 76377
rect 41485 73385 44485 73393
rect 44675 76377 47675 76385
rect 44675 73393 44683 76377
rect 47667 73393 47675 76377
rect 44675 73385 47675 73393
rect 47865 76377 50865 76385
rect 47865 73393 47873 76377
rect 50857 73393 50865 76377
rect 47865 73385 50865 73393
rect 51055 76377 54055 76385
rect 51055 73393 51063 76377
rect 54047 73393 54055 76377
rect 51055 73385 54055 73393
rect 54245 76377 57245 76385
rect 54245 73393 54253 76377
rect 57237 73393 57245 76377
rect 54245 73385 57245 73393
rect 57435 76377 60435 76385
rect 57435 73393 57443 76377
rect 60427 73393 60435 76377
rect 57435 73385 60435 73393
rect 60625 76377 63625 76385
rect 60625 73393 60633 76377
rect 63617 73393 63625 76377
rect 60625 73385 63625 73393
rect 63815 76377 66815 76385
rect 63815 73393 63823 76377
rect 66807 73393 66815 76377
rect 63815 73385 66815 73393
rect 67005 76377 70005 76385
rect 67005 73393 67013 76377
rect 69997 73393 70005 76377
rect 67005 73385 70005 73393
rect 70195 76377 73195 76385
rect 70195 73393 70203 76377
rect 73187 73393 73195 76377
rect 70195 73385 73195 73393
rect 73385 76377 76385 76385
rect 73385 73393 73393 76377
rect 76377 73393 76385 76377
rect 73385 73385 76385 73393
rect 76575 76377 79575 76385
rect 76575 73393 76583 76377
rect 79567 73393 79575 76377
rect 76575 73385 79575 73393
rect 79765 76377 82765 76385
rect 79765 73393 79773 76377
rect 82757 73393 82765 76377
rect 79765 73385 82765 73393
rect 82955 76377 85955 76385
rect 82955 73393 82963 76377
rect 85947 73393 85955 76377
rect 82955 73385 85955 73393
rect 86145 76377 89145 76385
rect 86145 73393 86153 76377
rect 89137 73393 89145 76377
rect 86145 73385 89145 73393
rect 89335 76377 92335 76385
rect 89335 73393 89343 76377
rect 92327 73393 92335 76377
rect 89335 73385 92335 73393
rect 92525 76377 95525 76385
rect 92525 73393 92533 76377
rect 95517 73393 95525 76377
rect 92525 73385 95525 73393
rect 95715 76377 98715 76385
rect 95715 73393 95723 76377
rect 98707 73393 98715 76377
rect 95715 73385 98715 73393
rect 98905 76377 101905 76385
rect 98905 73393 98913 76377
rect 101897 73393 101905 76377
rect 98905 73385 101905 73393
rect 102095 76377 105095 76385
rect 102095 73393 102103 76377
rect 105087 73393 105095 76377
rect 102095 73385 105095 73393
rect 105285 76377 108285 76385
rect 105285 73393 105293 76377
rect 108277 73393 108285 76377
rect 105285 73385 108285 73393
rect 108475 76377 111475 76385
rect 108475 73393 108483 76377
rect 111467 73393 111475 76377
rect 108475 73385 111475 73393
rect 111665 76377 114665 76385
rect 111665 73393 111673 76377
rect 114657 73393 114665 76377
rect 111665 73385 114665 73393
rect 114855 76377 117855 76385
rect 114855 73393 114863 76377
rect 117847 73393 117855 76377
rect 114855 73385 117855 73393
rect 118045 76377 121045 76385
rect 118045 73393 118053 76377
rect 121037 73393 121045 76377
rect 118045 73385 121045 73393
rect 121235 76377 124235 76385
rect 121235 73393 121243 76377
rect 124227 73393 124235 76377
rect 121235 73385 124235 73393
rect 124425 76377 127425 76385
rect 124425 73393 124433 76377
rect 127417 73393 127425 76377
rect 124425 73385 127425 73393
rect 127615 76377 130615 76385
rect 127615 73393 127623 76377
rect 130607 73393 130615 76377
rect 127615 73385 130615 73393
rect 130805 76377 133805 76385
rect 130805 73393 130813 76377
rect 133797 73393 133805 76377
rect 130805 73385 133805 73393
rect 133995 76377 136995 76385
rect 133995 73393 134003 76377
rect 136987 73393 136995 76377
rect 133995 73385 136995 73393
rect 15 73187 3015 73195
rect 15 70203 23 73187
rect 3007 70203 3015 73187
rect 15 70195 3015 70203
rect 3205 73187 6205 73195
rect 3205 70203 3213 73187
rect 6197 70203 6205 73187
rect 3205 70195 6205 70203
rect 6395 73187 9395 73195
rect 6395 70203 6403 73187
rect 9387 70203 9395 73187
rect 6395 70195 9395 70203
rect 9585 73187 12585 73195
rect 9585 70203 9593 73187
rect 12577 70203 12585 73187
rect 9585 70195 12585 70203
rect 12775 73187 15775 73195
rect 12775 70203 12783 73187
rect 15767 70203 15775 73187
rect 12775 70195 15775 70203
rect 15965 73187 18965 73195
rect 15965 70203 15973 73187
rect 18957 70203 18965 73187
rect 15965 70195 18965 70203
rect 19155 73187 22155 73195
rect 19155 70203 19163 73187
rect 22147 70203 22155 73187
rect 19155 70195 22155 70203
rect 22345 73187 25345 73195
rect 22345 70203 22353 73187
rect 25337 70203 25345 73187
rect 22345 70195 25345 70203
rect 25535 73187 28535 73195
rect 25535 70203 25543 73187
rect 28527 70203 28535 73187
rect 25535 70195 28535 70203
rect 28725 73187 31725 73195
rect 28725 70203 28733 73187
rect 31717 70203 31725 73187
rect 28725 70195 31725 70203
rect 31915 73187 34915 73195
rect 31915 70203 31923 73187
rect 34907 70203 34915 73187
rect 31915 70195 34915 70203
rect 35105 73187 38105 73195
rect 35105 70203 35113 73187
rect 38097 70203 38105 73187
rect 35105 70195 38105 70203
rect 38295 73187 41295 73195
rect 38295 70203 38303 73187
rect 41287 70203 41295 73187
rect 38295 70195 41295 70203
rect 41485 73187 44485 73195
rect 41485 70203 41493 73187
rect 44477 70203 44485 73187
rect 41485 70195 44485 70203
rect 44675 73187 47675 73195
rect 44675 70203 44683 73187
rect 47667 70203 47675 73187
rect 44675 70195 47675 70203
rect 47865 73187 50865 73195
rect 47865 70203 47873 73187
rect 50857 70203 50865 73187
rect 47865 70195 50865 70203
rect 51055 73187 54055 73195
rect 51055 70203 51063 73187
rect 54047 70203 54055 73187
rect 51055 70195 54055 70203
rect 54245 73187 57245 73195
rect 54245 70203 54253 73187
rect 57237 70203 57245 73187
rect 54245 70195 57245 70203
rect 57435 73187 60435 73195
rect 57435 70203 57443 73187
rect 60427 70203 60435 73187
rect 57435 70195 60435 70203
rect 60625 73187 63625 73195
rect 60625 70203 60633 73187
rect 63617 70203 63625 73187
rect 60625 70195 63625 70203
rect 63815 73187 66815 73195
rect 63815 70203 63823 73187
rect 66807 70203 66815 73187
rect 63815 70195 66815 70203
rect 67005 73187 70005 73195
rect 67005 70203 67013 73187
rect 69997 70203 70005 73187
rect 67005 70195 70005 70203
rect 70195 73187 73195 73195
rect 70195 70203 70203 73187
rect 73187 70203 73195 73187
rect 70195 70195 73195 70203
rect 73385 73187 76385 73195
rect 73385 70203 73393 73187
rect 76377 70203 76385 73187
rect 73385 70195 76385 70203
rect 76575 73187 79575 73195
rect 76575 70203 76583 73187
rect 79567 70203 79575 73187
rect 76575 70195 79575 70203
rect 79765 73187 82765 73195
rect 79765 70203 79773 73187
rect 82757 70203 82765 73187
rect 79765 70195 82765 70203
rect 82955 73187 85955 73195
rect 82955 70203 82963 73187
rect 85947 70203 85955 73187
rect 82955 70195 85955 70203
rect 86145 73187 89145 73195
rect 86145 70203 86153 73187
rect 89137 70203 89145 73187
rect 86145 70195 89145 70203
rect 89335 73187 92335 73195
rect 89335 70203 89343 73187
rect 92327 70203 92335 73187
rect 89335 70195 92335 70203
rect 92525 73187 95525 73195
rect 92525 70203 92533 73187
rect 95517 70203 95525 73187
rect 92525 70195 95525 70203
rect 95715 73187 98715 73195
rect 95715 70203 95723 73187
rect 98707 70203 98715 73187
rect 95715 70195 98715 70203
rect 98905 73187 101905 73195
rect 98905 70203 98913 73187
rect 101897 70203 101905 73187
rect 98905 70195 101905 70203
rect 102095 73187 105095 73195
rect 102095 70203 102103 73187
rect 105087 70203 105095 73187
rect 102095 70195 105095 70203
rect 105285 73187 108285 73195
rect 105285 70203 105293 73187
rect 108277 70203 108285 73187
rect 105285 70195 108285 70203
rect 108475 73187 111475 73195
rect 108475 70203 108483 73187
rect 111467 70203 111475 73187
rect 108475 70195 111475 70203
rect 111665 73187 114665 73195
rect 111665 70203 111673 73187
rect 114657 70203 114665 73187
rect 111665 70195 114665 70203
rect 114855 73187 117855 73195
rect 114855 70203 114863 73187
rect 117847 70203 117855 73187
rect 114855 70195 117855 70203
rect 118045 73187 121045 73195
rect 118045 70203 118053 73187
rect 121037 70203 121045 73187
rect 118045 70195 121045 70203
rect 121235 73187 124235 73195
rect 121235 70203 121243 73187
rect 124227 70203 124235 73187
rect 121235 70195 124235 70203
rect 124425 73187 127425 73195
rect 124425 70203 124433 73187
rect 127417 70203 127425 73187
rect 124425 70195 127425 70203
rect 127615 73187 130615 73195
rect 127615 70203 127623 73187
rect 130607 70203 130615 73187
rect 127615 70195 130615 70203
rect 130805 73187 133805 73195
rect 130805 70203 130813 73187
rect 133797 70203 133805 73187
rect 130805 70195 133805 70203
rect 133995 73187 136995 73195
rect 133995 70203 134003 73187
rect 136987 70203 136995 73187
rect 133995 70195 136995 70203
rect 15 69997 3015 70005
rect 15 67013 23 69997
rect 3007 67013 3015 69997
rect 15 67005 3015 67013
rect 3205 69997 6205 70005
rect 3205 67013 3213 69997
rect 6197 67013 6205 69997
rect 3205 67005 6205 67013
rect 6395 69997 9395 70005
rect 6395 67013 6403 69997
rect 9387 67013 9395 69997
rect 6395 67005 9395 67013
rect 9585 69997 12585 70005
rect 9585 67013 9593 69997
rect 12577 67013 12585 69997
rect 9585 67005 12585 67013
rect 12775 69997 15775 70005
rect 12775 67013 12783 69997
rect 15767 67013 15775 69997
rect 12775 67005 15775 67013
rect 15965 69997 18965 70005
rect 15965 67013 15973 69997
rect 18957 67013 18965 69997
rect 15965 67005 18965 67013
rect 19155 69997 22155 70005
rect 19155 67013 19163 69997
rect 22147 67013 22155 69997
rect 19155 67005 22155 67013
rect 22345 69997 25345 70005
rect 22345 67013 22353 69997
rect 25337 67013 25345 69997
rect 22345 67005 25345 67013
rect 25535 69997 28535 70005
rect 25535 67013 25543 69997
rect 28527 67013 28535 69997
rect 25535 67005 28535 67013
rect 28725 69997 31725 70005
rect 28725 67013 28733 69997
rect 31717 67013 31725 69997
rect 28725 67005 31725 67013
rect 31915 69997 34915 70005
rect 31915 67013 31923 69997
rect 34907 67013 34915 69997
rect 31915 67005 34915 67013
rect 35105 69997 38105 70005
rect 35105 67013 35113 69997
rect 38097 67013 38105 69997
rect 35105 67005 38105 67013
rect 38295 69997 41295 70005
rect 38295 67013 38303 69997
rect 41287 67013 41295 69997
rect 38295 67005 41295 67013
rect 41485 69997 44485 70005
rect 41485 67013 41493 69997
rect 44477 67013 44485 69997
rect 41485 67005 44485 67013
rect 44675 69997 47675 70005
rect 44675 67013 44683 69997
rect 47667 67013 47675 69997
rect 44675 67005 47675 67013
rect 47865 69997 50865 70005
rect 47865 67013 47873 69997
rect 50857 67013 50865 69997
rect 47865 67005 50865 67013
rect 51055 69997 54055 70005
rect 51055 67013 51063 69997
rect 54047 67013 54055 69997
rect 51055 67005 54055 67013
rect 54245 69997 57245 70005
rect 54245 67013 54253 69997
rect 57237 67013 57245 69997
rect 54245 67005 57245 67013
rect 57435 69997 60435 70005
rect 57435 67013 57443 69997
rect 60427 67013 60435 69997
rect 57435 67005 60435 67013
rect 60625 69997 63625 70005
rect 60625 67013 60633 69997
rect 63617 67013 63625 69997
rect 60625 67005 63625 67013
rect 63815 69997 66815 70005
rect 63815 67013 63823 69997
rect 66807 67013 66815 69997
rect 63815 67005 66815 67013
rect 67005 69997 70005 70005
rect 67005 67013 67013 69997
rect 69997 67013 70005 69997
rect 67005 67005 70005 67013
rect 70195 69997 73195 70005
rect 70195 67013 70203 69997
rect 73187 67013 73195 69997
rect 70195 67005 73195 67013
rect 73385 69997 76385 70005
rect 73385 67013 73393 69997
rect 76377 67013 76385 69997
rect 73385 67005 76385 67013
rect 76575 69997 79575 70005
rect 76575 67013 76583 69997
rect 79567 67013 79575 69997
rect 76575 67005 79575 67013
rect 79765 69997 82765 70005
rect 79765 67013 79773 69997
rect 82757 67013 82765 69997
rect 79765 67005 82765 67013
rect 82955 69997 85955 70005
rect 82955 67013 82963 69997
rect 85947 67013 85955 69997
rect 82955 67005 85955 67013
rect 86145 69997 89145 70005
rect 86145 67013 86153 69997
rect 89137 67013 89145 69997
rect 86145 67005 89145 67013
rect 89335 69997 92335 70005
rect 89335 67013 89343 69997
rect 92327 67013 92335 69997
rect 89335 67005 92335 67013
rect 92525 69997 95525 70005
rect 92525 67013 92533 69997
rect 95517 67013 95525 69997
rect 92525 67005 95525 67013
rect 95715 69997 98715 70005
rect 95715 67013 95723 69997
rect 98707 67013 98715 69997
rect 95715 67005 98715 67013
rect 98905 69997 101905 70005
rect 98905 67013 98913 69997
rect 101897 67013 101905 69997
rect 98905 67005 101905 67013
rect 102095 69997 105095 70005
rect 102095 67013 102103 69997
rect 105087 67013 105095 69997
rect 102095 67005 105095 67013
rect 105285 69997 108285 70005
rect 105285 67013 105293 69997
rect 108277 67013 108285 69997
rect 105285 67005 108285 67013
rect 108475 69997 111475 70005
rect 108475 67013 108483 69997
rect 111467 67013 111475 69997
rect 108475 67005 111475 67013
rect 111665 69997 114665 70005
rect 111665 67013 111673 69997
rect 114657 67013 114665 69997
rect 111665 67005 114665 67013
rect 114855 69997 117855 70005
rect 114855 67013 114863 69997
rect 117847 67013 117855 69997
rect 114855 67005 117855 67013
rect 118045 69997 121045 70005
rect 118045 67013 118053 69997
rect 121037 67013 121045 69997
rect 118045 67005 121045 67013
rect 121235 69997 124235 70005
rect 121235 67013 121243 69997
rect 124227 67013 124235 69997
rect 121235 67005 124235 67013
rect 124425 69997 127425 70005
rect 124425 67013 124433 69997
rect 127417 67013 127425 69997
rect 124425 67005 127425 67013
rect 127615 69997 130615 70005
rect 127615 67013 127623 69997
rect 130607 67013 130615 69997
rect 127615 67005 130615 67013
rect 130805 69997 133805 70005
rect 130805 67013 130813 69997
rect 133797 67013 133805 69997
rect 130805 67005 133805 67013
rect 133995 69997 136995 70005
rect 133995 67013 134003 69997
rect 136987 67013 136995 69997
rect 133995 67005 136995 67013
rect 15 66807 3015 66815
rect 15 63823 23 66807
rect 3007 63823 3015 66807
rect 15 63815 3015 63823
rect 3205 66807 6205 66815
rect 3205 63823 3213 66807
rect 6197 63823 6205 66807
rect 3205 63815 6205 63823
rect 6395 66807 9395 66815
rect 6395 63823 6403 66807
rect 9387 63823 9395 66807
rect 6395 63815 9395 63823
rect 9585 66807 12585 66815
rect 9585 63823 9593 66807
rect 12577 63823 12585 66807
rect 9585 63815 12585 63823
rect 12775 66807 15775 66815
rect 12775 63823 12783 66807
rect 15767 63823 15775 66807
rect 12775 63815 15775 63823
rect 15965 66807 18965 66815
rect 15965 63823 15973 66807
rect 18957 63823 18965 66807
rect 15965 63815 18965 63823
rect 19155 66807 22155 66815
rect 19155 63823 19163 66807
rect 22147 63823 22155 66807
rect 19155 63815 22155 63823
rect 22345 66807 25345 66815
rect 22345 63823 22353 66807
rect 25337 63823 25345 66807
rect 22345 63815 25345 63823
rect 25535 66807 28535 66815
rect 25535 63823 25543 66807
rect 28527 63823 28535 66807
rect 25535 63815 28535 63823
rect 28725 66807 31725 66815
rect 28725 63823 28733 66807
rect 31717 63823 31725 66807
rect 28725 63815 31725 63823
rect 31915 66807 34915 66815
rect 31915 63823 31923 66807
rect 34907 63823 34915 66807
rect 31915 63815 34915 63823
rect 35105 66807 38105 66815
rect 35105 63823 35113 66807
rect 38097 63823 38105 66807
rect 35105 63815 38105 63823
rect 38295 66807 41295 66815
rect 38295 63823 38303 66807
rect 41287 63823 41295 66807
rect 38295 63815 41295 63823
rect 41485 66807 44485 66815
rect 41485 63823 41493 66807
rect 44477 63823 44485 66807
rect 41485 63815 44485 63823
rect 44675 66807 47675 66815
rect 44675 63823 44683 66807
rect 47667 63823 47675 66807
rect 44675 63815 47675 63823
rect 47865 66807 50865 66815
rect 47865 63823 47873 66807
rect 50857 63823 50865 66807
rect 47865 63815 50865 63823
rect 51055 66807 54055 66815
rect 51055 63823 51063 66807
rect 54047 63823 54055 66807
rect 51055 63815 54055 63823
rect 54245 66807 57245 66815
rect 54245 63823 54253 66807
rect 57237 63823 57245 66807
rect 54245 63815 57245 63823
rect 57435 66807 60435 66815
rect 57435 63823 57443 66807
rect 60427 63823 60435 66807
rect 57435 63815 60435 63823
rect 60625 66807 63625 66815
rect 60625 63823 60633 66807
rect 63617 63823 63625 66807
rect 60625 63815 63625 63823
rect 63815 66807 66815 66815
rect 63815 63823 63823 66807
rect 66807 63823 66815 66807
rect 63815 63815 66815 63823
rect 67005 66807 70005 66815
rect 67005 63823 67013 66807
rect 69997 63823 70005 66807
rect 67005 63815 70005 63823
rect 70195 66807 73195 66815
rect 70195 63823 70203 66807
rect 73187 63823 73195 66807
rect 70195 63815 73195 63823
rect 73385 66807 76385 66815
rect 73385 63823 73393 66807
rect 76377 63823 76385 66807
rect 73385 63815 76385 63823
rect 76575 66807 79575 66815
rect 76575 63823 76583 66807
rect 79567 63823 79575 66807
rect 76575 63815 79575 63823
rect 79765 66807 82765 66815
rect 79765 63823 79773 66807
rect 82757 63823 82765 66807
rect 79765 63815 82765 63823
rect 82955 66807 85955 66815
rect 82955 63823 82963 66807
rect 85947 63823 85955 66807
rect 82955 63815 85955 63823
rect 86145 66807 89145 66815
rect 86145 63823 86153 66807
rect 89137 63823 89145 66807
rect 86145 63815 89145 63823
rect 89335 66807 92335 66815
rect 89335 63823 89343 66807
rect 92327 63823 92335 66807
rect 89335 63815 92335 63823
rect 92525 66807 95525 66815
rect 92525 63823 92533 66807
rect 95517 63823 95525 66807
rect 92525 63815 95525 63823
rect 95715 66807 98715 66815
rect 95715 63823 95723 66807
rect 98707 63823 98715 66807
rect 95715 63815 98715 63823
rect 98905 66807 101905 66815
rect 98905 63823 98913 66807
rect 101897 63823 101905 66807
rect 98905 63815 101905 63823
rect 102095 66807 105095 66815
rect 102095 63823 102103 66807
rect 105087 63823 105095 66807
rect 102095 63815 105095 63823
rect 105285 66807 108285 66815
rect 105285 63823 105293 66807
rect 108277 63823 108285 66807
rect 105285 63815 108285 63823
rect 108475 66807 111475 66815
rect 108475 63823 108483 66807
rect 111467 63823 111475 66807
rect 108475 63815 111475 63823
rect 111665 66807 114665 66815
rect 111665 63823 111673 66807
rect 114657 63823 114665 66807
rect 111665 63815 114665 63823
rect 114855 66807 117855 66815
rect 114855 63823 114863 66807
rect 117847 63823 117855 66807
rect 114855 63815 117855 63823
rect 118045 66807 121045 66815
rect 118045 63823 118053 66807
rect 121037 63823 121045 66807
rect 118045 63815 121045 63823
rect 121235 66807 124235 66815
rect 121235 63823 121243 66807
rect 124227 63823 124235 66807
rect 121235 63815 124235 63823
rect 124425 66807 127425 66815
rect 124425 63823 124433 66807
rect 127417 63823 127425 66807
rect 124425 63815 127425 63823
rect 127615 66807 130615 66815
rect 127615 63823 127623 66807
rect 130607 63823 130615 66807
rect 127615 63815 130615 63823
rect 130805 66807 133805 66815
rect 130805 63823 130813 66807
rect 133797 63823 133805 66807
rect 130805 63815 133805 63823
rect 133995 66807 136995 66815
rect 133995 63823 134003 66807
rect 136987 63823 136995 66807
rect 133995 63815 136995 63823
rect 15 63617 3015 63625
rect 15 60633 23 63617
rect 3007 60633 3015 63617
rect 15 60625 3015 60633
rect 3205 63617 6205 63625
rect 3205 60633 3213 63617
rect 6197 60633 6205 63617
rect 3205 60625 6205 60633
rect 6395 63617 9395 63625
rect 6395 60633 6403 63617
rect 9387 60633 9395 63617
rect 6395 60625 9395 60633
rect 9585 63617 12585 63625
rect 9585 60633 9593 63617
rect 12577 60633 12585 63617
rect 9585 60625 12585 60633
rect 12775 63617 15775 63625
rect 12775 60633 12783 63617
rect 15767 60633 15775 63617
rect 12775 60625 15775 60633
rect 15965 63617 18965 63625
rect 15965 60633 15973 63617
rect 18957 60633 18965 63617
rect 15965 60625 18965 60633
rect 19155 63617 22155 63625
rect 19155 60633 19163 63617
rect 22147 60633 22155 63617
rect 19155 60625 22155 60633
rect 22345 63617 25345 63625
rect 22345 60633 22353 63617
rect 25337 60633 25345 63617
rect 22345 60625 25345 60633
rect 25535 63617 28535 63625
rect 25535 60633 25543 63617
rect 28527 60633 28535 63617
rect 25535 60625 28535 60633
rect 28725 63617 31725 63625
rect 28725 60633 28733 63617
rect 31717 60633 31725 63617
rect 28725 60625 31725 60633
rect 31915 63617 34915 63625
rect 31915 60633 31923 63617
rect 34907 60633 34915 63617
rect 31915 60625 34915 60633
rect 35105 63617 38105 63625
rect 35105 60633 35113 63617
rect 38097 60633 38105 63617
rect 35105 60625 38105 60633
rect 38295 63617 41295 63625
rect 38295 60633 38303 63617
rect 41287 60633 41295 63617
rect 38295 60625 41295 60633
rect 41485 63617 44485 63625
rect 41485 60633 41493 63617
rect 44477 60633 44485 63617
rect 41485 60625 44485 60633
rect 44675 63617 47675 63625
rect 44675 60633 44683 63617
rect 47667 60633 47675 63617
rect 44675 60625 47675 60633
rect 47865 63617 50865 63625
rect 47865 60633 47873 63617
rect 50857 60633 50865 63617
rect 47865 60625 50865 60633
rect 51055 63617 54055 63625
rect 51055 60633 51063 63617
rect 54047 60633 54055 63617
rect 51055 60625 54055 60633
rect 54245 63617 57245 63625
rect 54245 60633 54253 63617
rect 57237 60633 57245 63617
rect 54245 60625 57245 60633
rect 57435 63617 60435 63625
rect 57435 60633 57443 63617
rect 60427 60633 60435 63617
rect 57435 60625 60435 60633
rect 60625 63617 63625 63625
rect 60625 60633 60633 63617
rect 63617 60633 63625 63617
rect 60625 60625 63625 60633
rect 63815 63617 66815 63625
rect 63815 60633 63823 63617
rect 66807 60633 66815 63617
rect 63815 60625 66815 60633
rect 67005 63617 70005 63625
rect 67005 60633 67013 63617
rect 69997 60633 70005 63617
rect 67005 60625 70005 60633
rect 70195 63617 73195 63625
rect 70195 60633 70203 63617
rect 73187 60633 73195 63617
rect 70195 60625 73195 60633
rect 73385 63617 76385 63625
rect 73385 60633 73393 63617
rect 76377 60633 76385 63617
rect 73385 60625 76385 60633
rect 76575 63617 79575 63625
rect 76575 60633 76583 63617
rect 79567 60633 79575 63617
rect 76575 60625 79575 60633
rect 79765 63617 82765 63625
rect 79765 60633 79773 63617
rect 82757 60633 82765 63617
rect 79765 60625 82765 60633
rect 82955 63617 85955 63625
rect 82955 60633 82963 63617
rect 85947 60633 85955 63617
rect 82955 60625 85955 60633
rect 86145 63617 89145 63625
rect 86145 60633 86153 63617
rect 89137 60633 89145 63617
rect 86145 60625 89145 60633
rect 89335 63617 92335 63625
rect 89335 60633 89343 63617
rect 92327 60633 92335 63617
rect 89335 60625 92335 60633
rect 92525 63617 95525 63625
rect 92525 60633 92533 63617
rect 95517 60633 95525 63617
rect 92525 60625 95525 60633
rect 95715 63617 98715 63625
rect 95715 60633 95723 63617
rect 98707 60633 98715 63617
rect 95715 60625 98715 60633
rect 98905 63617 101905 63625
rect 98905 60633 98913 63617
rect 101897 60633 101905 63617
rect 98905 60625 101905 60633
rect 102095 63617 105095 63625
rect 102095 60633 102103 63617
rect 105087 60633 105095 63617
rect 102095 60625 105095 60633
rect 105285 63617 108285 63625
rect 105285 60633 105293 63617
rect 108277 60633 108285 63617
rect 105285 60625 108285 60633
rect 108475 63617 111475 63625
rect 108475 60633 108483 63617
rect 111467 60633 111475 63617
rect 108475 60625 111475 60633
rect 111665 63617 114665 63625
rect 111665 60633 111673 63617
rect 114657 60633 114665 63617
rect 111665 60625 114665 60633
rect 114855 63617 117855 63625
rect 114855 60633 114863 63617
rect 117847 60633 117855 63617
rect 114855 60625 117855 60633
rect 118045 63617 121045 63625
rect 118045 60633 118053 63617
rect 121037 60633 121045 63617
rect 118045 60625 121045 60633
rect 121235 63617 124235 63625
rect 121235 60633 121243 63617
rect 124227 60633 124235 63617
rect 121235 60625 124235 60633
rect 124425 63617 127425 63625
rect 124425 60633 124433 63617
rect 127417 60633 127425 63617
rect 124425 60625 127425 60633
rect 127615 63617 130615 63625
rect 127615 60633 127623 63617
rect 130607 60633 130615 63617
rect 127615 60625 130615 60633
rect 130805 63617 133805 63625
rect 130805 60633 130813 63617
rect 133797 60633 133805 63617
rect 130805 60625 133805 60633
rect 133995 63617 136995 63625
rect 133995 60633 134003 63617
rect 136987 60633 136995 63617
rect 133995 60625 136995 60633
rect 15 60427 3015 60435
rect 15 57443 23 60427
rect 3007 57443 3015 60427
rect 15 57435 3015 57443
rect 3205 60427 6205 60435
rect 3205 57443 3213 60427
rect 6197 57443 6205 60427
rect 3205 57435 6205 57443
rect 6395 60427 9395 60435
rect 6395 57443 6403 60427
rect 9387 57443 9395 60427
rect 6395 57435 9395 57443
rect 9585 60427 12585 60435
rect 9585 57443 9593 60427
rect 12577 57443 12585 60427
rect 9585 57435 12585 57443
rect 12775 60427 15775 60435
rect 12775 57443 12783 60427
rect 15767 57443 15775 60427
rect 12775 57435 15775 57443
rect 15965 60427 18965 60435
rect 15965 57443 15973 60427
rect 18957 57443 18965 60427
rect 15965 57435 18965 57443
rect 19155 60427 22155 60435
rect 19155 57443 19163 60427
rect 22147 57443 22155 60427
rect 19155 57435 22155 57443
rect 22345 60427 25345 60435
rect 22345 57443 22353 60427
rect 25337 57443 25345 60427
rect 22345 57435 25345 57443
rect 25535 60427 28535 60435
rect 25535 57443 25543 60427
rect 28527 57443 28535 60427
rect 25535 57435 28535 57443
rect 28725 60427 31725 60435
rect 28725 57443 28733 60427
rect 31717 57443 31725 60427
rect 28725 57435 31725 57443
rect 31915 60427 34915 60435
rect 31915 57443 31923 60427
rect 34907 57443 34915 60427
rect 31915 57435 34915 57443
rect 35105 60427 38105 60435
rect 35105 57443 35113 60427
rect 38097 57443 38105 60427
rect 35105 57435 38105 57443
rect 38295 60427 41295 60435
rect 38295 57443 38303 60427
rect 41287 57443 41295 60427
rect 38295 57435 41295 57443
rect 41485 60427 44485 60435
rect 41485 57443 41493 60427
rect 44477 57443 44485 60427
rect 41485 57435 44485 57443
rect 44675 60427 47675 60435
rect 44675 57443 44683 60427
rect 47667 57443 47675 60427
rect 44675 57435 47675 57443
rect 47865 60427 50865 60435
rect 47865 57443 47873 60427
rect 50857 57443 50865 60427
rect 47865 57435 50865 57443
rect 51055 60427 54055 60435
rect 51055 57443 51063 60427
rect 54047 57443 54055 60427
rect 51055 57435 54055 57443
rect 54245 60427 57245 60435
rect 54245 57443 54253 60427
rect 57237 57443 57245 60427
rect 54245 57435 57245 57443
rect 57435 60427 60435 60435
rect 57435 57443 57443 60427
rect 60427 57443 60435 60427
rect 57435 57435 60435 57443
rect 60625 60427 63625 60435
rect 60625 57443 60633 60427
rect 63617 57443 63625 60427
rect 60625 57435 63625 57443
rect 63815 60427 66815 60435
rect 63815 57443 63823 60427
rect 66807 57443 66815 60427
rect 63815 57435 66815 57443
rect 67005 60427 70005 60435
rect 67005 57443 67013 60427
rect 69997 57443 70005 60427
rect 67005 57435 70005 57443
rect 70195 60427 73195 60435
rect 70195 57443 70203 60427
rect 73187 57443 73195 60427
rect 70195 57435 73195 57443
rect 73385 60427 76385 60435
rect 73385 57443 73393 60427
rect 76377 57443 76385 60427
rect 73385 57435 76385 57443
rect 76575 60427 79575 60435
rect 76575 57443 76583 60427
rect 79567 57443 79575 60427
rect 76575 57435 79575 57443
rect 79765 60427 82765 60435
rect 79765 57443 79773 60427
rect 82757 57443 82765 60427
rect 79765 57435 82765 57443
rect 82955 60427 85955 60435
rect 82955 57443 82963 60427
rect 85947 57443 85955 60427
rect 82955 57435 85955 57443
rect 86145 60427 89145 60435
rect 86145 57443 86153 60427
rect 89137 57443 89145 60427
rect 86145 57435 89145 57443
rect 89335 60427 92335 60435
rect 89335 57443 89343 60427
rect 92327 57443 92335 60427
rect 89335 57435 92335 57443
rect 92525 60427 95525 60435
rect 92525 57443 92533 60427
rect 95517 57443 95525 60427
rect 92525 57435 95525 57443
rect 95715 60427 98715 60435
rect 95715 57443 95723 60427
rect 98707 57443 98715 60427
rect 95715 57435 98715 57443
rect 98905 60427 101905 60435
rect 98905 57443 98913 60427
rect 101897 57443 101905 60427
rect 98905 57435 101905 57443
rect 102095 60427 105095 60435
rect 102095 57443 102103 60427
rect 105087 57443 105095 60427
rect 102095 57435 105095 57443
rect 105285 60427 108285 60435
rect 105285 57443 105293 60427
rect 108277 57443 108285 60427
rect 105285 57435 108285 57443
rect 108475 60427 111475 60435
rect 108475 57443 108483 60427
rect 111467 57443 111475 60427
rect 108475 57435 111475 57443
rect 111665 60427 114665 60435
rect 111665 57443 111673 60427
rect 114657 57443 114665 60427
rect 111665 57435 114665 57443
rect 114855 60427 117855 60435
rect 114855 57443 114863 60427
rect 117847 57443 117855 60427
rect 114855 57435 117855 57443
rect 118045 60427 121045 60435
rect 118045 57443 118053 60427
rect 121037 57443 121045 60427
rect 118045 57435 121045 57443
rect 121235 60427 124235 60435
rect 121235 57443 121243 60427
rect 124227 57443 124235 60427
rect 121235 57435 124235 57443
rect 124425 60427 127425 60435
rect 124425 57443 124433 60427
rect 127417 57443 127425 60427
rect 124425 57435 127425 57443
rect 127615 60427 130615 60435
rect 127615 57443 127623 60427
rect 130607 57443 130615 60427
rect 127615 57435 130615 57443
rect 130805 60427 133805 60435
rect 130805 57443 130813 60427
rect 133797 57443 133805 60427
rect 130805 57435 133805 57443
rect 133995 60427 136995 60435
rect 133995 57443 134003 60427
rect 136987 57443 136995 60427
rect 133995 57435 136995 57443
rect 15 57237 3015 57245
rect 15 54253 23 57237
rect 3007 54253 3015 57237
rect 15 54245 3015 54253
rect 3205 57237 6205 57245
rect 3205 54253 3213 57237
rect 6197 54253 6205 57237
rect 3205 54245 6205 54253
rect 6395 57237 9395 57245
rect 6395 54253 6403 57237
rect 9387 54253 9395 57237
rect 6395 54245 9395 54253
rect 9585 57237 12585 57245
rect 9585 54253 9593 57237
rect 12577 54253 12585 57237
rect 9585 54245 12585 54253
rect 12775 57237 15775 57245
rect 12775 54253 12783 57237
rect 15767 54253 15775 57237
rect 12775 54245 15775 54253
rect 15965 57237 18965 57245
rect 15965 54253 15973 57237
rect 18957 54253 18965 57237
rect 15965 54245 18965 54253
rect 19155 57237 22155 57245
rect 19155 54253 19163 57237
rect 22147 54253 22155 57237
rect 19155 54245 22155 54253
rect 22345 57237 25345 57245
rect 22345 54253 22353 57237
rect 25337 54253 25345 57237
rect 22345 54245 25345 54253
rect 25535 57237 28535 57245
rect 25535 54253 25543 57237
rect 28527 54253 28535 57237
rect 25535 54245 28535 54253
rect 28725 57237 31725 57245
rect 28725 54253 28733 57237
rect 31717 54253 31725 57237
rect 28725 54245 31725 54253
rect 31915 57237 34915 57245
rect 31915 54253 31923 57237
rect 34907 54253 34915 57237
rect 31915 54245 34915 54253
rect 35105 57237 38105 57245
rect 35105 54253 35113 57237
rect 38097 54253 38105 57237
rect 35105 54245 38105 54253
rect 38295 57237 41295 57245
rect 38295 54253 38303 57237
rect 41287 54253 41295 57237
rect 38295 54245 41295 54253
rect 41485 57237 44485 57245
rect 41485 54253 41493 57237
rect 44477 54253 44485 57237
rect 41485 54245 44485 54253
rect 44675 57237 47675 57245
rect 44675 54253 44683 57237
rect 47667 54253 47675 57237
rect 44675 54245 47675 54253
rect 47865 57237 50865 57245
rect 47865 54253 47873 57237
rect 50857 54253 50865 57237
rect 47865 54245 50865 54253
rect 51055 57237 54055 57245
rect 51055 54253 51063 57237
rect 54047 54253 54055 57237
rect 51055 54245 54055 54253
rect 54245 57237 57245 57245
rect 54245 54253 54253 57237
rect 57237 54253 57245 57237
rect 54245 54245 57245 54253
rect 57435 57237 60435 57245
rect 57435 54253 57443 57237
rect 60427 54253 60435 57237
rect 57435 54245 60435 54253
rect 60625 57237 63625 57245
rect 60625 54253 60633 57237
rect 63617 54253 63625 57237
rect 60625 54245 63625 54253
rect 63815 57237 66815 57245
rect 63815 54253 63823 57237
rect 66807 54253 66815 57237
rect 63815 54245 66815 54253
rect 67005 57237 70005 57245
rect 67005 54253 67013 57237
rect 69997 54253 70005 57237
rect 67005 54245 70005 54253
rect 70195 57237 73195 57245
rect 70195 54253 70203 57237
rect 73187 54253 73195 57237
rect 70195 54245 73195 54253
rect 73385 57237 76385 57245
rect 73385 54253 73393 57237
rect 76377 54253 76385 57237
rect 73385 54245 76385 54253
rect 76575 57237 79575 57245
rect 76575 54253 76583 57237
rect 79567 54253 79575 57237
rect 76575 54245 79575 54253
rect 79765 57237 82765 57245
rect 79765 54253 79773 57237
rect 82757 54253 82765 57237
rect 79765 54245 82765 54253
rect 82955 57237 85955 57245
rect 82955 54253 82963 57237
rect 85947 54253 85955 57237
rect 82955 54245 85955 54253
rect 86145 57237 89145 57245
rect 86145 54253 86153 57237
rect 89137 54253 89145 57237
rect 86145 54245 89145 54253
rect 89335 57237 92335 57245
rect 89335 54253 89343 57237
rect 92327 54253 92335 57237
rect 89335 54245 92335 54253
rect 92525 57237 95525 57245
rect 92525 54253 92533 57237
rect 95517 54253 95525 57237
rect 92525 54245 95525 54253
rect 95715 57237 98715 57245
rect 95715 54253 95723 57237
rect 98707 54253 98715 57237
rect 95715 54245 98715 54253
rect 98905 57237 101905 57245
rect 98905 54253 98913 57237
rect 101897 54253 101905 57237
rect 98905 54245 101905 54253
rect 102095 57237 105095 57245
rect 102095 54253 102103 57237
rect 105087 54253 105095 57237
rect 102095 54245 105095 54253
rect 105285 57237 108285 57245
rect 105285 54253 105293 57237
rect 108277 54253 108285 57237
rect 105285 54245 108285 54253
rect 108475 57237 111475 57245
rect 108475 54253 108483 57237
rect 111467 54253 111475 57237
rect 108475 54245 111475 54253
rect 111665 57237 114665 57245
rect 111665 54253 111673 57237
rect 114657 54253 114665 57237
rect 111665 54245 114665 54253
rect 114855 57237 117855 57245
rect 114855 54253 114863 57237
rect 117847 54253 117855 57237
rect 114855 54245 117855 54253
rect 118045 57237 121045 57245
rect 118045 54253 118053 57237
rect 121037 54253 121045 57237
rect 118045 54245 121045 54253
rect 121235 57237 124235 57245
rect 121235 54253 121243 57237
rect 124227 54253 124235 57237
rect 121235 54245 124235 54253
rect 124425 57237 127425 57245
rect 124425 54253 124433 57237
rect 127417 54253 127425 57237
rect 124425 54245 127425 54253
rect 127615 57237 130615 57245
rect 127615 54253 127623 57237
rect 130607 54253 130615 57237
rect 127615 54245 130615 54253
rect 130805 57237 133805 57245
rect 130805 54253 130813 57237
rect 133797 54253 133805 57237
rect 130805 54245 133805 54253
rect 133995 57237 136995 57245
rect 133995 54253 134003 57237
rect 136987 54253 136995 57237
rect 133995 54245 136995 54253
rect 15 54047 3015 54055
rect 15 51063 23 54047
rect 3007 51063 3015 54047
rect 15 51055 3015 51063
rect 3205 54047 6205 54055
rect 3205 51063 3213 54047
rect 6197 51063 6205 54047
rect 3205 51055 6205 51063
rect 6395 54047 9395 54055
rect 6395 51063 6403 54047
rect 9387 51063 9395 54047
rect 6395 51055 9395 51063
rect 9585 54047 12585 54055
rect 9585 51063 9593 54047
rect 12577 51063 12585 54047
rect 9585 51055 12585 51063
rect 12775 54047 15775 54055
rect 12775 51063 12783 54047
rect 15767 51063 15775 54047
rect 12775 51055 15775 51063
rect 15965 54047 18965 54055
rect 15965 51063 15973 54047
rect 18957 51063 18965 54047
rect 15965 51055 18965 51063
rect 19155 54047 22155 54055
rect 19155 51063 19163 54047
rect 22147 51063 22155 54047
rect 19155 51055 22155 51063
rect 22345 54047 25345 54055
rect 22345 51063 22353 54047
rect 25337 51063 25345 54047
rect 22345 51055 25345 51063
rect 25535 54047 28535 54055
rect 25535 51063 25543 54047
rect 28527 51063 28535 54047
rect 25535 51055 28535 51063
rect 28725 54047 31725 54055
rect 28725 51063 28733 54047
rect 31717 51063 31725 54047
rect 28725 51055 31725 51063
rect 31915 54047 34915 54055
rect 31915 51063 31923 54047
rect 34907 51063 34915 54047
rect 31915 51055 34915 51063
rect 35105 54047 38105 54055
rect 35105 51063 35113 54047
rect 38097 51063 38105 54047
rect 35105 51055 38105 51063
rect 38295 54047 41295 54055
rect 38295 51063 38303 54047
rect 41287 51063 41295 54047
rect 38295 51055 41295 51063
rect 41485 54047 44485 54055
rect 41485 51063 41493 54047
rect 44477 51063 44485 54047
rect 41485 51055 44485 51063
rect 44675 54047 47675 54055
rect 44675 51063 44683 54047
rect 47667 51063 47675 54047
rect 44675 51055 47675 51063
rect 47865 54047 50865 54055
rect 47865 51063 47873 54047
rect 50857 51063 50865 54047
rect 47865 51055 50865 51063
rect 51055 54047 54055 54055
rect 51055 51063 51063 54047
rect 54047 51063 54055 54047
rect 51055 51055 54055 51063
rect 54245 54047 57245 54055
rect 54245 51063 54253 54047
rect 57237 51063 57245 54047
rect 54245 51055 57245 51063
rect 57435 54047 60435 54055
rect 57435 51063 57443 54047
rect 60427 51063 60435 54047
rect 57435 51055 60435 51063
rect 60625 54047 63625 54055
rect 60625 51063 60633 54047
rect 63617 51063 63625 54047
rect 60625 51055 63625 51063
rect 63815 54047 66815 54055
rect 63815 51063 63823 54047
rect 66807 51063 66815 54047
rect 63815 51055 66815 51063
rect 67005 54047 70005 54055
rect 67005 51063 67013 54047
rect 69997 51063 70005 54047
rect 67005 51055 70005 51063
rect 70195 54047 73195 54055
rect 70195 51063 70203 54047
rect 73187 51063 73195 54047
rect 70195 51055 73195 51063
rect 73385 54047 76385 54055
rect 73385 51063 73393 54047
rect 76377 51063 76385 54047
rect 73385 51055 76385 51063
rect 76575 54047 79575 54055
rect 76575 51063 76583 54047
rect 79567 51063 79575 54047
rect 76575 51055 79575 51063
rect 79765 54047 82765 54055
rect 79765 51063 79773 54047
rect 82757 51063 82765 54047
rect 79765 51055 82765 51063
rect 82955 54047 85955 54055
rect 82955 51063 82963 54047
rect 85947 51063 85955 54047
rect 82955 51055 85955 51063
rect 86145 54047 89145 54055
rect 86145 51063 86153 54047
rect 89137 51063 89145 54047
rect 86145 51055 89145 51063
rect 89335 54047 92335 54055
rect 89335 51063 89343 54047
rect 92327 51063 92335 54047
rect 89335 51055 92335 51063
rect 92525 54047 95525 54055
rect 92525 51063 92533 54047
rect 95517 51063 95525 54047
rect 92525 51055 95525 51063
rect 95715 54047 98715 54055
rect 95715 51063 95723 54047
rect 98707 51063 98715 54047
rect 95715 51055 98715 51063
rect 98905 54047 101905 54055
rect 98905 51063 98913 54047
rect 101897 51063 101905 54047
rect 98905 51055 101905 51063
rect 102095 54047 105095 54055
rect 102095 51063 102103 54047
rect 105087 51063 105095 54047
rect 102095 51055 105095 51063
rect 105285 54047 108285 54055
rect 105285 51063 105293 54047
rect 108277 51063 108285 54047
rect 105285 51055 108285 51063
rect 108475 54047 111475 54055
rect 108475 51063 108483 54047
rect 111467 51063 111475 54047
rect 108475 51055 111475 51063
rect 111665 54047 114665 54055
rect 111665 51063 111673 54047
rect 114657 51063 114665 54047
rect 111665 51055 114665 51063
rect 114855 54047 117855 54055
rect 114855 51063 114863 54047
rect 117847 51063 117855 54047
rect 114855 51055 117855 51063
rect 118045 54047 121045 54055
rect 118045 51063 118053 54047
rect 121037 51063 121045 54047
rect 118045 51055 121045 51063
rect 121235 54047 124235 54055
rect 121235 51063 121243 54047
rect 124227 51063 124235 54047
rect 121235 51055 124235 51063
rect 124425 54047 127425 54055
rect 124425 51063 124433 54047
rect 127417 51063 127425 54047
rect 124425 51055 127425 51063
rect 127615 54047 130615 54055
rect 127615 51063 127623 54047
rect 130607 51063 130615 54047
rect 127615 51055 130615 51063
rect 130805 54047 133805 54055
rect 130805 51063 130813 54047
rect 133797 51063 133805 54047
rect 130805 51055 133805 51063
rect 133995 54047 136995 54055
rect 133995 51063 134003 54047
rect 136987 51063 136995 54047
rect 133995 51055 136995 51063
rect 15 50857 3015 50865
rect 15 47873 23 50857
rect 3007 47873 3015 50857
rect 15 47865 3015 47873
rect 3205 50857 6205 50865
rect 3205 47873 3213 50857
rect 6197 47873 6205 50857
rect 3205 47865 6205 47873
rect 6395 50857 9395 50865
rect 6395 47873 6403 50857
rect 9387 47873 9395 50857
rect 6395 47865 9395 47873
rect 9585 50857 12585 50865
rect 9585 47873 9593 50857
rect 12577 47873 12585 50857
rect 9585 47865 12585 47873
rect 12775 50857 15775 50865
rect 12775 47873 12783 50857
rect 15767 47873 15775 50857
rect 12775 47865 15775 47873
rect 15965 50857 18965 50865
rect 15965 47873 15973 50857
rect 18957 47873 18965 50857
rect 15965 47865 18965 47873
rect 19155 50857 22155 50865
rect 19155 47873 19163 50857
rect 22147 47873 22155 50857
rect 19155 47865 22155 47873
rect 22345 50857 25345 50865
rect 22345 47873 22353 50857
rect 25337 47873 25345 50857
rect 22345 47865 25345 47873
rect 25535 50857 28535 50865
rect 25535 47873 25543 50857
rect 28527 47873 28535 50857
rect 25535 47865 28535 47873
rect 28725 50857 31725 50865
rect 28725 47873 28733 50857
rect 31717 47873 31725 50857
rect 28725 47865 31725 47873
rect 31915 50857 34915 50865
rect 31915 47873 31923 50857
rect 34907 47873 34915 50857
rect 31915 47865 34915 47873
rect 35105 50857 38105 50865
rect 35105 47873 35113 50857
rect 38097 47873 38105 50857
rect 35105 47865 38105 47873
rect 38295 50857 41295 50865
rect 38295 47873 38303 50857
rect 41287 47873 41295 50857
rect 38295 47865 41295 47873
rect 41485 50857 44485 50865
rect 41485 47873 41493 50857
rect 44477 47873 44485 50857
rect 41485 47865 44485 47873
rect 44675 50857 47675 50865
rect 44675 47873 44683 50857
rect 47667 47873 47675 50857
rect 44675 47865 47675 47873
rect 47865 50857 50865 50865
rect 47865 47873 47873 50857
rect 50857 47873 50865 50857
rect 47865 47865 50865 47873
rect 51055 50857 54055 50865
rect 51055 47873 51063 50857
rect 54047 47873 54055 50857
rect 51055 47865 54055 47873
rect 54245 50857 57245 50865
rect 54245 47873 54253 50857
rect 57237 47873 57245 50857
rect 54245 47865 57245 47873
rect 57435 50857 60435 50865
rect 57435 47873 57443 50857
rect 60427 47873 60435 50857
rect 57435 47865 60435 47873
rect 60625 50857 63625 50865
rect 60625 47873 60633 50857
rect 63617 47873 63625 50857
rect 60625 47865 63625 47873
rect 63815 50857 66815 50865
rect 63815 47873 63823 50857
rect 66807 47873 66815 50857
rect 63815 47865 66815 47873
rect 67005 50857 70005 50865
rect 67005 47873 67013 50857
rect 69997 47873 70005 50857
rect 67005 47865 70005 47873
rect 70195 50857 73195 50865
rect 70195 47873 70203 50857
rect 73187 47873 73195 50857
rect 70195 47865 73195 47873
rect 73385 50857 76385 50865
rect 73385 47873 73393 50857
rect 76377 47873 76385 50857
rect 73385 47865 76385 47873
rect 76575 50857 79575 50865
rect 76575 47873 76583 50857
rect 79567 47873 79575 50857
rect 76575 47865 79575 47873
rect 79765 50857 82765 50865
rect 79765 47873 79773 50857
rect 82757 47873 82765 50857
rect 79765 47865 82765 47873
rect 82955 50857 85955 50865
rect 82955 47873 82963 50857
rect 85947 47873 85955 50857
rect 82955 47865 85955 47873
rect 86145 50857 89145 50865
rect 86145 47873 86153 50857
rect 89137 47873 89145 50857
rect 86145 47865 89145 47873
rect 89335 50857 92335 50865
rect 89335 47873 89343 50857
rect 92327 47873 92335 50857
rect 89335 47865 92335 47873
rect 92525 50857 95525 50865
rect 92525 47873 92533 50857
rect 95517 47873 95525 50857
rect 92525 47865 95525 47873
rect 95715 50857 98715 50865
rect 95715 47873 95723 50857
rect 98707 47873 98715 50857
rect 95715 47865 98715 47873
rect 98905 50857 101905 50865
rect 98905 47873 98913 50857
rect 101897 47873 101905 50857
rect 98905 47865 101905 47873
rect 102095 50857 105095 50865
rect 102095 47873 102103 50857
rect 105087 47873 105095 50857
rect 102095 47865 105095 47873
rect 105285 50857 108285 50865
rect 105285 47873 105293 50857
rect 108277 47873 108285 50857
rect 105285 47865 108285 47873
rect 108475 50857 111475 50865
rect 108475 47873 108483 50857
rect 111467 47873 111475 50857
rect 108475 47865 111475 47873
rect 111665 50857 114665 50865
rect 111665 47873 111673 50857
rect 114657 47873 114665 50857
rect 111665 47865 114665 47873
rect 114855 50857 117855 50865
rect 114855 47873 114863 50857
rect 117847 47873 117855 50857
rect 114855 47865 117855 47873
rect 118045 50857 121045 50865
rect 118045 47873 118053 50857
rect 121037 47873 121045 50857
rect 118045 47865 121045 47873
rect 121235 50857 124235 50865
rect 121235 47873 121243 50857
rect 124227 47873 124235 50857
rect 121235 47865 124235 47873
rect 124425 50857 127425 50865
rect 124425 47873 124433 50857
rect 127417 47873 127425 50857
rect 124425 47865 127425 47873
rect 127615 50857 130615 50865
rect 127615 47873 127623 50857
rect 130607 47873 130615 50857
rect 127615 47865 130615 47873
rect 130805 50857 133805 50865
rect 130805 47873 130813 50857
rect 133797 47873 133805 50857
rect 130805 47865 133805 47873
rect 133995 50857 136995 50865
rect 133995 47873 134003 50857
rect 136987 47873 136995 50857
rect 133995 47865 136995 47873
rect 15 47667 3015 47675
rect 15 44683 23 47667
rect 3007 44683 3015 47667
rect 15 44675 3015 44683
rect 3205 47667 6205 47675
rect 3205 44683 3213 47667
rect 6197 44683 6205 47667
rect 3205 44675 6205 44683
rect 6395 47667 9395 47675
rect 6395 44683 6403 47667
rect 9387 44683 9395 47667
rect 6395 44675 9395 44683
rect 9585 47667 12585 47675
rect 9585 44683 9593 47667
rect 12577 44683 12585 47667
rect 9585 44675 12585 44683
rect 12775 47667 15775 47675
rect 12775 44683 12783 47667
rect 15767 44683 15775 47667
rect 12775 44675 15775 44683
rect 15965 47667 18965 47675
rect 15965 44683 15973 47667
rect 18957 44683 18965 47667
rect 15965 44675 18965 44683
rect 19155 47667 22155 47675
rect 19155 44683 19163 47667
rect 22147 44683 22155 47667
rect 19155 44675 22155 44683
rect 22345 47667 25345 47675
rect 22345 44683 22353 47667
rect 25337 44683 25345 47667
rect 22345 44675 25345 44683
rect 25535 47667 28535 47675
rect 25535 44683 25543 47667
rect 28527 44683 28535 47667
rect 25535 44675 28535 44683
rect 28725 47667 31725 47675
rect 28725 44683 28733 47667
rect 31717 44683 31725 47667
rect 28725 44675 31725 44683
rect 31915 47667 34915 47675
rect 31915 44683 31923 47667
rect 34907 44683 34915 47667
rect 31915 44675 34915 44683
rect 35105 47667 38105 47675
rect 35105 44683 35113 47667
rect 38097 44683 38105 47667
rect 35105 44675 38105 44683
rect 38295 47667 41295 47675
rect 38295 44683 38303 47667
rect 41287 44683 41295 47667
rect 38295 44675 41295 44683
rect 41485 47667 44485 47675
rect 41485 44683 41493 47667
rect 44477 44683 44485 47667
rect 41485 44675 44485 44683
rect 44675 47667 47675 47675
rect 44675 44683 44683 47667
rect 47667 44683 47675 47667
rect 44675 44675 47675 44683
rect 47865 47667 50865 47675
rect 47865 44683 47873 47667
rect 50857 44683 50865 47667
rect 47865 44675 50865 44683
rect 51055 47667 54055 47675
rect 51055 44683 51063 47667
rect 54047 44683 54055 47667
rect 51055 44675 54055 44683
rect 54245 47667 57245 47675
rect 54245 44683 54253 47667
rect 57237 44683 57245 47667
rect 54245 44675 57245 44683
rect 57435 47667 60435 47675
rect 57435 44683 57443 47667
rect 60427 44683 60435 47667
rect 57435 44675 60435 44683
rect 60625 47667 63625 47675
rect 60625 44683 60633 47667
rect 63617 44683 63625 47667
rect 60625 44675 63625 44683
rect 63815 47667 66815 47675
rect 63815 44683 63823 47667
rect 66807 44683 66815 47667
rect 63815 44675 66815 44683
rect 67005 47667 70005 47675
rect 67005 44683 67013 47667
rect 69997 44683 70005 47667
rect 67005 44675 70005 44683
rect 70195 47667 73195 47675
rect 70195 44683 70203 47667
rect 73187 44683 73195 47667
rect 70195 44675 73195 44683
rect 73385 47667 76385 47675
rect 73385 44683 73393 47667
rect 76377 44683 76385 47667
rect 73385 44675 76385 44683
rect 76575 47667 79575 47675
rect 76575 44683 76583 47667
rect 79567 44683 79575 47667
rect 76575 44675 79575 44683
rect 79765 47667 82765 47675
rect 79765 44683 79773 47667
rect 82757 44683 82765 47667
rect 79765 44675 82765 44683
rect 82955 47667 85955 47675
rect 82955 44683 82963 47667
rect 85947 44683 85955 47667
rect 82955 44675 85955 44683
rect 86145 47667 89145 47675
rect 86145 44683 86153 47667
rect 89137 44683 89145 47667
rect 86145 44675 89145 44683
rect 89335 47667 92335 47675
rect 89335 44683 89343 47667
rect 92327 44683 92335 47667
rect 89335 44675 92335 44683
rect 92525 47667 95525 47675
rect 92525 44683 92533 47667
rect 95517 44683 95525 47667
rect 92525 44675 95525 44683
rect 95715 47667 98715 47675
rect 95715 44683 95723 47667
rect 98707 44683 98715 47667
rect 95715 44675 98715 44683
rect 98905 47667 101905 47675
rect 98905 44683 98913 47667
rect 101897 44683 101905 47667
rect 98905 44675 101905 44683
rect 102095 47667 105095 47675
rect 102095 44683 102103 47667
rect 105087 44683 105095 47667
rect 102095 44675 105095 44683
rect 105285 47667 108285 47675
rect 105285 44683 105293 47667
rect 108277 44683 108285 47667
rect 105285 44675 108285 44683
rect 108475 47667 111475 47675
rect 108475 44683 108483 47667
rect 111467 44683 111475 47667
rect 108475 44675 111475 44683
rect 111665 47667 114665 47675
rect 111665 44683 111673 47667
rect 114657 44683 114665 47667
rect 111665 44675 114665 44683
rect 114855 47667 117855 47675
rect 114855 44683 114863 47667
rect 117847 44683 117855 47667
rect 114855 44675 117855 44683
rect 118045 47667 121045 47675
rect 118045 44683 118053 47667
rect 121037 44683 121045 47667
rect 118045 44675 121045 44683
rect 121235 47667 124235 47675
rect 121235 44683 121243 47667
rect 124227 44683 124235 47667
rect 121235 44675 124235 44683
rect 124425 47667 127425 47675
rect 124425 44683 124433 47667
rect 127417 44683 127425 47667
rect 124425 44675 127425 44683
rect 127615 47667 130615 47675
rect 127615 44683 127623 47667
rect 130607 44683 130615 47667
rect 127615 44675 130615 44683
rect 130805 47667 133805 47675
rect 130805 44683 130813 47667
rect 133797 44683 133805 47667
rect 130805 44675 133805 44683
rect 133995 47667 136995 47675
rect 133995 44683 134003 47667
rect 136987 44683 136995 47667
rect 133995 44675 136995 44683
rect 15 44477 3015 44485
rect 15 41493 23 44477
rect 3007 41493 3015 44477
rect 15 41485 3015 41493
rect 3205 44477 6205 44485
rect 3205 41493 3213 44477
rect 6197 41493 6205 44477
rect 3205 41485 6205 41493
rect 6395 44477 9395 44485
rect 6395 41493 6403 44477
rect 9387 41493 9395 44477
rect 6395 41485 9395 41493
rect 9585 44477 12585 44485
rect 9585 41493 9593 44477
rect 12577 41493 12585 44477
rect 9585 41485 12585 41493
rect 12775 44477 15775 44485
rect 12775 41493 12783 44477
rect 15767 41493 15775 44477
rect 12775 41485 15775 41493
rect 15965 44477 18965 44485
rect 15965 41493 15973 44477
rect 18957 41493 18965 44477
rect 15965 41485 18965 41493
rect 19155 44477 22155 44485
rect 19155 41493 19163 44477
rect 22147 41493 22155 44477
rect 19155 41485 22155 41493
rect 22345 44477 25345 44485
rect 22345 41493 22353 44477
rect 25337 41493 25345 44477
rect 22345 41485 25345 41493
rect 25535 44477 28535 44485
rect 25535 41493 25543 44477
rect 28527 41493 28535 44477
rect 25535 41485 28535 41493
rect 28725 44477 31725 44485
rect 28725 41493 28733 44477
rect 31717 41493 31725 44477
rect 28725 41485 31725 41493
rect 31915 44477 34915 44485
rect 31915 41493 31923 44477
rect 34907 41493 34915 44477
rect 31915 41485 34915 41493
rect 35105 44477 38105 44485
rect 35105 41493 35113 44477
rect 38097 41493 38105 44477
rect 35105 41485 38105 41493
rect 38295 44477 41295 44485
rect 38295 41493 38303 44477
rect 41287 41493 41295 44477
rect 38295 41485 41295 41493
rect 41485 44477 44485 44485
rect 41485 41493 41493 44477
rect 44477 41493 44485 44477
rect 41485 41485 44485 41493
rect 44675 44477 47675 44485
rect 44675 41493 44683 44477
rect 47667 41493 47675 44477
rect 44675 41485 47675 41493
rect 47865 44477 50865 44485
rect 47865 41493 47873 44477
rect 50857 41493 50865 44477
rect 47865 41485 50865 41493
rect 51055 44477 54055 44485
rect 51055 41493 51063 44477
rect 54047 41493 54055 44477
rect 51055 41485 54055 41493
rect 54245 44477 57245 44485
rect 54245 41493 54253 44477
rect 57237 41493 57245 44477
rect 54245 41485 57245 41493
rect 57435 44477 60435 44485
rect 57435 41493 57443 44477
rect 60427 41493 60435 44477
rect 57435 41485 60435 41493
rect 60625 44477 63625 44485
rect 60625 41493 60633 44477
rect 63617 41493 63625 44477
rect 60625 41485 63625 41493
rect 63815 44477 66815 44485
rect 63815 41493 63823 44477
rect 66807 41493 66815 44477
rect 63815 41485 66815 41493
rect 67005 44477 70005 44485
rect 67005 41493 67013 44477
rect 69997 41493 70005 44477
rect 67005 41485 70005 41493
rect 70195 44477 73195 44485
rect 70195 41493 70203 44477
rect 73187 41493 73195 44477
rect 70195 41485 73195 41493
rect 73385 44477 76385 44485
rect 73385 41493 73393 44477
rect 76377 41493 76385 44477
rect 73385 41485 76385 41493
rect 76575 44477 79575 44485
rect 76575 41493 76583 44477
rect 79567 41493 79575 44477
rect 76575 41485 79575 41493
rect 79765 44477 82765 44485
rect 79765 41493 79773 44477
rect 82757 41493 82765 44477
rect 79765 41485 82765 41493
rect 82955 44477 85955 44485
rect 82955 41493 82963 44477
rect 85947 41493 85955 44477
rect 82955 41485 85955 41493
rect 86145 44477 89145 44485
rect 86145 41493 86153 44477
rect 89137 41493 89145 44477
rect 86145 41485 89145 41493
rect 89335 44477 92335 44485
rect 89335 41493 89343 44477
rect 92327 41493 92335 44477
rect 89335 41485 92335 41493
rect 92525 44477 95525 44485
rect 92525 41493 92533 44477
rect 95517 41493 95525 44477
rect 92525 41485 95525 41493
rect 95715 44477 98715 44485
rect 95715 41493 95723 44477
rect 98707 41493 98715 44477
rect 95715 41485 98715 41493
rect 98905 44477 101905 44485
rect 98905 41493 98913 44477
rect 101897 41493 101905 44477
rect 98905 41485 101905 41493
rect 102095 44477 105095 44485
rect 102095 41493 102103 44477
rect 105087 41493 105095 44477
rect 102095 41485 105095 41493
rect 105285 44477 108285 44485
rect 105285 41493 105293 44477
rect 108277 41493 108285 44477
rect 105285 41485 108285 41493
rect 108475 44477 111475 44485
rect 108475 41493 108483 44477
rect 111467 41493 111475 44477
rect 108475 41485 111475 41493
rect 111665 44477 114665 44485
rect 111665 41493 111673 44477
rect 114657 41493 114665 44477
rect 111665 41485 114665 41493
rect 114855 44477 117855 44485
rect 114855 41493 114863 44477
rect 117847 41493 117855 44477
rect 114855 41485 117855 41493
rect 118045 44477 121045 44485
rect 118045 41493 118053 44477
rect 121037 41493 121045 44477
rect 118045 41485 121045 41493
rect 121235 44477 124235 44485
rect 121235 41493 121243 44477
rect 124227 41493 124235 44477
rect 121235 41485 124235 41493
rect 124425 44477 127425 44485
rect 124425 41493 124433 44477
rect 127417 41493 127425 44477
rect 124425 41485 127425 41493
rect 127615 44477 130615 44485
rect 127615 41493 127623 44477
rect 130607 41493 130615 44477
rect 127615 41485 130615 41493
rect 130805 44477 133805 44485
rect 130805 41493 130813 44477
rect 133797 41493 133805 44477
rect 130805 41485 133805 41493
rect 133995 44477 136995 44485
rect 133995 41493 134003 44477
rect 136987 41493 136995 44477
rect 133995 41485 136995 41493
rect 15 41287 3015 41295
rect 15 38303 23 41287
rect 3007 38303 3015 41287
rect 15 38295 3015 38303
rect 3205 41287 6205 41295
rect 3205 38303 3213 41287
rect 6197 38303 6205 41287
rect 3205 38295 6205 38303
rect 6395 41287 9395 41295
rect 6395 38303 6403 41287
rect 9387 38303 9395 41287
rect 6395 38295 9395 38303
rect 9585 41287 12585 41295
rect 9585 38303 9593 41287
rect 12577 38303 12585 41287
rect 9585 38295 12585 38303
rect 12775 41287 15775 41295
rect 12775 38303 12783 41287
rect 15767 38303 15775 41287
rect 12775 38295 15775 38303
rect 15965 41287 18965 41295
rect 15965 38303 15973 41287
rect 18957 38303 18965 41287
rect 15965 38295 18965 38303
rect 19155 41287 22155 41295
rect 19155 38303 19163 41287
rect 22147 38303 22155 41287
rect 19155 38295 22155 38303
rect 22345 41287 25345 41295
rect 22345 38303 22353 41287
rect 25337 38303 25345 41287
rect 22345 38295 25345 38303
rect 25535 41287 28535 41295
rect 25535 38303 25543 41287
rect 28527 38303 28535 41287
rect 25535 38295 28535 38303
rect 28725 41287 31725 41295
rect 28725 38303 28733 41287
rect 31717 38303 31725 41287
rect 28725 38295 31725 38303
rect 31915 41287 34915 41295
rect 31915 38303 31923 41287
rect 34907 38303 34915 41287
rect 31915 38295 34915 38303
rect 35105 41287 38105 41295
rect 35105 38303 35113 41287
rect 38097 38303 38105 41287
rect 35105 38295 38105 38303
rect 38295 41287 41295 41295
rect 38295 38303 38303 41287
rect 41287 38303 41295 41287
rect 38295 38295 41295 38303
rect 41485 41287 44485 41295
rect 41485 38303 41493 41287
rect 44477 38303 44485 41287
rect 41485 38295 44485 38303
rect 44675 41287 47675 41295
rect 44675 38303 44683 41287
rect 47667 38303 47675 41287
rect 44675 38295 47675 38303
rect 47865 41287 50865 41295
rect 47865 38303 47873 41287
rect 50857 38303 50865 41287
rect 47865 38295 50865 38303
rect 51055 41287 54055 41295
rect 51055 38303 51063 41287
rect 54047 38303 54055 41287
rect 51055 38295 54055 38303
rect 54245 41287 57245 41295
rect 54245 38303 54253 41287
rect 57237 38303 57245 41287
rect 54245 38295 57245 38303
rect 57435 41287 60435 41295
rect 57435 38303 57443 41287
rect 60427 38303 60435 41287
rect 57435 38295 60435 38303
rect 60625 41287 63625 41295
rect 60625 38303 60633 41287
rect 63617 38303 63625 41287
rect 60625 38295 63625 38303
rect 63815 41287 66815 41295
rect 63815 38303 63823 41287
rect 66807 38303 66815 41287
rect 63815 38295 66815 38303
rect 67005 41287 70005 41295
rect 67005 38303 67013 41287
rect 69997 38303 70005 41287
rect 67005 38295 70005 38303
rect 70195 41287 73195 41295
rect 70195 38303 70203 41287
rect 73187 38303 73195 41287
rect 70195 38295 73195 38303
rect 73385 41287 76385 41295
rect 73385 38303 73393 41287
rect 76377 38303 76385 41287
rect 73385 38295 76385 38303
rect 76575 41287 79575 41295
rect 76575 38303 76583 41287
rect 79567 38303 79575 41287
rect 76575 38295 79575 38303
rect 79765 41287 82765 41295
rect 79765 38303 79773 41287
rect 82757 38303 82765 41287
rect 79765 38295 82765 38303
rect 82955 41287 85955 41295
rect 82955 38303 82963 41287
rect 85947 38303 85955 41287
rect 82955 38295 85955 38303
rect 86145 41287 89145 41295
rect 86145 38303 86153 41287
rect 89137 38303 89145 41287
rect 86145 38295 89145 38303
rect 89335 41287 92335 41295
rect 89335 38303 89343 41287
rect 92327 38303 92335 41287
rect 89335 38295 92335 38303
rect 92525 41287 95525 41295
rect 92525 38303 92533 41287
rect 95517 38303 95525 41287
rect 92525 38295 95525 38303
rect 95715 41287 98715 41295
rect 95715 38303 95723 41287
rect 98707 38303 98715 41287
rect 95715 38295 98715 38303
rect 98905 41287 101905 41295
rect 98905 38303 98913 41287
rect 101897 38303 101905 41287
rect 98905 38295 101905 38303
rect 102095 41287 105095 41295
rect 102095 38303 102103 41287
rect 105087 38303 105095 41287
rect 102095 38295 105095 38303
rect 105285 41287 108285 41295
rect 105285 38303 105293 41287
rect 108277 38303 108285 41287
rect 105285 38295 108285 38303
rect 108475 41287 111475 41295
rect 108475 38303 108483 41287
rect 111467 38303 111475 41287
rect 108475 38295 111475 38303
rect 111665 41287 114665 41295
rect 111665 38303 111673 41287
rect 114657 38303 114665 41287
rect 111665 38295 114665 38303
rect 114855 41287 117855 41295
rect 114855 38303 114863 41287
rect 117847 38303 117855 41287
rect 114855 38295 117855 38303
rect 118045 41287 121045 41295
rect 118045 38303 118053 41287
rect 121037 38303 121045 41287
rect 118045 38295 121045 38303
rect 121235 41287 124235 41295
rect 121235 38303 121243 41287
rect 124227 38303 124235 41287
rect 121235 38295 124235 38303
rect 124425 41287 127425 41295
rect 124425 38303 124433 41287
rect 127417 38303 127425 41287
rect 124425 38295 127425 38303
rect 127615 41287 130615 41295
rect 127615 38303 127623 41287
rect 130607 38303 130615 41287
rect 127615 38295 130615 38303
rect 130805 41287 133805 41295
rect 130805 38303 130813 41287
rect 133797 38303 133805 41287
rect 130805 38295 133805 38303
rect 133995 41287 136995 41295
rect 133995 38303 134003 41287
rect 136987 38303 136995 41287
rect 133995 38295 136995 38303
rect 15 38097 3015 38105
rect 15 35113 23 38097
rect 3007 35113 3015 38097
rect 15 35105 3015 35113
rect 3205 38097 6205 38105
rect 3205 35113 3213 38097
rect 6197 35113 6205 38097
rect 3205 35105 6205 35113
rect 6395 38097 9395 38105
rect 6395 35113 6403 38097
rect 9387 35113 9395 38097
rect 6395 35105 9395 35113
rect 9585 38097 12585 38105
rect 9585 35113 9593 38097
rect 12577 35113 12585 38097
rect 9585 35105 12585 35113
rect 12775 38097 15775 38105
rect 12775 35113 12783 38097
rect 15767 35113 15775 38097
rect 12775 35105 15775 35113
rect 15965 38097 18965 38105
rect 15965 35113 15973 38097
rect 18957 35113 18965 38097
rect 15965 35105 18965 35113
rect 19155 38097 22155 38105
rect 19155 35113 19163 38097
rect 22147 35113 22155 38097
rect 19155 35105 22155 35113
rect 22345 38097 25345 38105
rect 22345 35113 22353 38097
rect 25337 35113 25345 38097
rect 22345 35105 25345 35113
rect 25535 38097 28535 38105
rect 25535 35113 25543 38097
rect 28527 35113 28535 38097
rect 25535 35105 28535 35113
rect 28725 38097 31725 38105
rect 28725 35113 28733 38097
rect 31717 35113 31725 38097
rect 28725 35105 31725 35113
rect 31915 38097 34915 38105
rect 31915 35113 31923 38097
rect 34907 35113 34915 38097
rect 31915 35105 34915 35113
rect 35105 38097 38105 38105
rect 35105 35113 35113 38097
rect 38097 35113 38105 38097
rect 35105 35105 38105 35113
rect 38295 38097 41295 38105
rect 38295 35113 38303 38097
rect 41287 35113 41295 38097
rect 38295 35105 41295 35113
rect 41485 38097 44485 38105
rect 41485 35113 41493 38097
rect 44477 35113 44485 38097
rect 41485 35105 44485 35113
rect 44675 38097 47675 38105
rect 44675 35113 44683 38097
rect 47667 35113 47675 38097
rect 44675 35105 47675 35113
rect 47865 38097 50865 38105
rect 47865 35113 47873 38097
rect 50857 35113 50865 38097
rect 47865 35105 50865 35113
rect 51055 38097 54055 38105
rect 51055 35113 51063 38097
rect 54047 35113 54055 38097
rect 51055 35105 54055 35113
rect 54245 38097 57245 38105
rect 54245 35113 54253 38097
rect 57237 35113 57245 38097
rect 54245 35105 57245 35113
rect 57435 38097 60435 38105
rect 57435 35113 57443 38097
rect 60427 35113 60435 38097
rect 57435 35105 60435 35113
rect 60625 38097 63625 38105
rect 60625 35113 60633 38097
rect 63617 35113 63625 38097
rect 60625 35105 63625 35113
rect 63815 38097 66815 38105
rect 63815 35113 63823 38097
rect 66807 35113 66815 38097
rect 63815 35105 66815 35113
rect 67005 38097 70005 38105
rect 67005 35113 67013 38097
rect 69997 35113 70005 38097
rect 67005 35105 70005 35113
rect 70195 38097 73195 38105
rect 70195 35113 70203 38097
rect 73187 35113 73195 38097
rect 70195 35105 73195 35113
rect 73385 38097 76385 38105
rect 73385 35113 73393 38097
rect 76377 35113 76385 38097
rect 73385 35105 76385 35113
rect 76575 38097 79575 38105
rect 76575 35113 76583 38097
rect 79567 35113 79575 38097
rect 76575 35105 79575 35113
rect 79765 38097 82765 38105
rect 79765 35113 79773 38097
rect 82757 35113 82765 38097
rect 79765 35105 82765 35113
rect 82955 38097 85955 38105
rect 82955 35113 82963 38097
rect 85947 35113 85955 38097
rect 82955 35105 85955 35113
rect 86145 38097 89145 38105
rect 86145 35113 86153 38097
rect 89137 35113 89145 38097
rect 86145 35105 89145 35113
rect 89335 38097 92335 38105
rect 89335 35113 89343 38097
rect 92327 35113 92335 38097
rect 89335 35105 92335 35113
rect 92525 38097 95525 38105
rect 92525 35113 92533 38097
rect 95517 35113 95525 38097
rect 92525 35105 95525 35113
rect 95715 38097 98715 38105
rect 95715 35113 95723 38097
rect 98707 35113 98715 38097
rect 95715 35105 98715 35113
rect 98905 38097 101905 38105
rect 98905 35113 98913 38097
rect 101897 35113 101905 38097
rect 98905 35105 101905 35113
rect 102095 38097 105095 38105
rect 102095 35113 102103 38097
rect 105087 35113 105095 38097
rect 102095 35105 105095 35113
rect 105285 38097 108285 38105
rect 105285 35113 105293 38097
rect 108277 35113 108285 38097
rect 105285 35105 108285 35113
rect 108475 38097 111475 38105
rect 108475 35113 108483 38097
rect 111467 35113 111475 38097
rect 108475 35105 111475 35113
rect 111665 38097 114665 38105
rect 111665 35113 111673 38097
rect 114657 35113 114665 38097
rect 111665 35105 114665 35113
rect 114855 38097 117855 38105
rect 114855 35113 114863 38097
rect 117847 35113 117855 38097
rect 114855 35105 117855 35113
rect 118045 38097 121045 38105
rect 118045 35113 118053 38097
rect 121037 35113 121045 38097
rect 118045 35105 121045 35113
rect 121235 38097 124235 38105
rect 121235 35113 121243 38097
rect 124227 35113 124235 38097
rect 121235 35105 124235 35113
rect 124425 38097 127425 38105
rect 124425 35113 124433 38097
rect 127417 35113 127425 38097
rect 124425 35105 127425 35113
rect 127615 38097 130615 38105
rect 127615 35113 127623 38097
rect 130607 35113 130615 38097
rect 127615 35105 130615 35113
rect 130805 38097 133805 38105
rect 130805 35113 130813 38097
rect 133797 35113 133805 38097
rect 130805 35105 133805 35113
rect 133995 38097 136995 38105
rect 133995 35113 134003 38097
rect 136987 35113 136995 38097
rect 133995 35105 136995 35113
rect 15 34907 3015 34915
rect 15 31923 23 34907
rect 3007 31923 3015 34907
rect 15 31915 3015 31923
rect 3205 34907 6205 34915
rect 3205 31923 3213 34907
rect 6197 31923 6205 34907
rect 3205 31915 6205 31923
rect 6395 34907 9395 34915
rect 6395 31923 6403 34907
rect 9387 31923 9395 34907
rect 6395 31915 9395 31923
rect 9585 34907 12585 34915
rect 9585 31923 9593 34907
rect 12577 31923 12585 34907
rect 9585 31915 12585 31923
rect 12775 34907 15775 34915
rect 12775 31923 12783 34907
rect 15767 31923 15775 34907
rect 12775 31915 15775 31923
rect 15965 34907 18965 34915
rect 15965 31923 15973 34907
rect 18957 31923 18965 34907
rect 15965 31915 18965 31923
rect 19155 34907 22155 34915
rect 19155 31923 19163 34907
rect 22147 31923 22155 34907
rect 19155 31915 22155 31923
rect 22345 34907 25345 34915
rect 22345 31923 22353 34907
rect 25337 31923 25345 34907
rect 22345 31915 25345 31923
rect 25535 34907 28535 34915
rect 25535 31923 25543 34907
rect 28527 31923 28535 34907
rect 25535 31915 28535 31923
rect 28725 34907 31725 34915
rect 28725 31923 28733 34907
rect 31717 31923 31725 34907
rect 28725 31915 31725 31923
rect 31915 34907 34915 34915
rect 31915 31923 31923 34907
rect 34907 31923 34915 34907
rect 31915 31915 34915 31923
rect 35105 34907 38105 34915
rect 35105 31923 35113 34907
rect 38097 31923 38105 34907
rect 35105 31915 38105 31923
rect 38295 34907 41295 34915
rect 38295 31923 38303 34907
rect 41287 31923 41295 34907
rect 38295 31915 41295 31923
rect 41485 34907 44485 34915
rect 41485 31923 41493 34907
rect 44477 31923 44485 34907
rect 41485 31915 44485 31923
rect 44675 34907 47675 34915
rect 44675 31923 44683 34907
rect 47667 31923 47675 34907
rect 44675 31915 47675 31923
rect 47865 34907 50865 34915
rect 47865 31923 47873 34907
rect 50857 31923 50865 34907
rect 47865 31915 50865 31923
rect 51055 34907 54055 34915
rect 51055 31923 51063 34907
rect 54047 31923 54055 34907
rect 51055 31915 54055 31923
rect 54245 34907 57245 34915
rect 54245 31923 54253 34907
rect 57237 31923 57245 34907
rect 54245 31915 57245 31923
rect 57435 34907 60435 34915
rect 57435 31923 57443 34907
rect 60427 31923 60435 34907
rect 57435 31915 60435 31923
rect 60625 34907 63625 34915
rect 60625 31923 60633 34907
rect 63617 31923 63625 34907
rect 60625 31915 63625 31923
rect 63815 34907 66815 34915
rect 63815 31923 63823 34907
rect 66807 31923 66815 34907
rect 63815 31915 66815 31923
rect 67005 34907 70005 34915
rect 67005 31923 67013 34907
rect 69997 31923 70005 34907
rect 67005 31915 70005 31923
rect 70195 34907 73195 34915
rect 70195 31923 70203 34907
rect 73187 31923 73195 34907
rect 70195 31915 73195 31923
rect 73385 34907 76385 34915
rect 73385 31923 73393 34907
rect 76377 31923 76385 34907
rect 73385 31915 76385 31923
rect 76575 34907 79575 34915
rect 76575 31923 76583 34907
rect 79567 31923 79575 34907
rect 76575 31915 79575 31923
rect 79765 34907 82765 34915
rect 79765 31923 79773 34907
rect 82757 31923 82765 34907
rect 79765 31915 82765 31923
rect 82955 34907 85955 34915
rect 82955 31923 82963 34907
rect 85947 31923 85955 34907
rect 82955 31915 85955 31923
rect 86145 34907 89145 34915
rect 86145 31923 86153 34907
rect 89137 31923 89145 34907
rect 86145 31915 89145 31923
rect 89335 34907 92335 34915
rect 89335 31923 89343 34907
rect 92327 31923 92335 34907
rect 89335 31915 92335 31923
rect 92525 34907 95525 34915
rect 92525 31923 92533 34907
rect 95517 31923 95525 34907
rect 92525 31915 95525 31923
rect 95715 34907 98715 34915
rect 95715 31923 95723 34907
rect 98707 31923 98715 34907
rect 95715 31915 98715 31923
rect 98905 34907 101905 34915
rect 98905 31923 98913 34907
rect 101897 31923 101905 34907
rect 98905 31915 101905 31923
rect 102095 34907 105095 34915
rect 102095 31923 102103 34907
rect 105087 31923 105095 34907
rect 102095 31915 105095 31923
rect 105285 34907 108285 34915
rect 105285 31923 105293 34907
rect 108277 31923 108285 34907
rect 105285 31915 108285 31923
rect 108475 34907 111475 34915
rect 108475 31923 108483 34907
rect 111467 31923 111475 34907
rect 108475 31915 111475 31923
rect 111665 34907 114665 34915
rect 111665 31923 111673 34907
rect 114657 31923 114665 34907
rect 111665 31915 114665 31923
rect 114855 34907 117855 34915
rect 114855 31923 114863 34907
rect 117847 31923 117855 34907
rect 114855 31915 117855 31923
rect 118045 34907 121045 34915
rect 118045 31923 118053 34907
rect 121037 31923 121045 34907
rect 118045 31915 121045 31923
rect 121235 34907 124235 34915
rect 121235 31923 121243 34907
rect 124227 31923 124235 34907
rect 121235 31915 124235 31923
rect 124425 34907 127425 34915
rect 124425 31923 124433 34907
rect 127417 31923 127425 34907
rect 124425 31915 127425 31923
rect 127615 34907 130615 34915
rect 127615 31923 127623 34907
rect 130607 31923 130615 34907
rect 127615 31915 130615 31923
rect 130805 34907 133805 34915
rect 130805 31923 130813 34907
rect 133797 31923 133805 34907
rect 130805 31915 133805 31923
rect 133995 34907 136995 34915
rect 133995 31923 134003 34907
rect 136987 31923 136995 34907
rect 133995 31915 136995 31923
rect 15 31717 3015 31725
rect 15 28733 23 31717
rect 3007 28733 3015 31717
rect 15 28725 3015 28733
rect 3205 31717 6205 31725
rect 3205 28733 3213 31717
rect 6197 28733 6205 31717
rect 3205 28725 6205 28733
rect 6395 31717 9395 31725
rect 6395 28733 6403 31717
rect 9387 28733 9395 31717
rect 6395 28725 9395 28733
rect 9585 31717 12585 31725
rect 9585 28733 9593 31717
rect 12577 28733 12585 31717
rect 9585 28725 12585 28733
rect 12775 31717 15775 31725
rect 12775 28733 12783 31717
rect 15767 28733 15775 31717
rect 12775 28725 15775 28733
rect 15965 31717 18965 31725
rect 15965 28733 15973 31717
rect 18957 28733 18965 31717
rect 15965 28725 18965 28733
rect 19155 31717 22155 31725
rect 19155 28733 19163 31717
rect 22147 28733 22155 31717
rect 19155 28725 22155 28733
rect 22345 31717 25345 31725
rect 22345 28733 22353 31717
rect 25337 28733 25345 31717
rect 22345 28725 25345 28733
rect 25535 31717 28535 31725
rect 25535 28733 25543 31717
rect 28527 28733 28535 31717
rect 25535 28725 28535 28733
rect 28725 31717 31725 31725
rect 28725 28733 28733 31717
rect 31717 28733 31725 31717
rect 28725 28725 31725 28733
rect 31915 31717 34915 31725
rect 31915 28733 31923 31717
rect 34907 28733 34915 31717
rect 31915 28725 34915 28733
rect 35105 31717 38105 31725
rect 35105 28733 35113 31717
rect 38097 28733 38105 31717
rect 35105 28725 38105 28733
rect 38295 31717 41295 31725
rect 38295 28733 38303 31717
rect 41287 28733 41295 31717
rect 38295 28725 41295 28733
rect 41485 31717 44485 31725
rect 41485 28733 41493 31717
rect 44477 28733 44485 31717
rect 41485 28725 44485 28733
rect 44675 31717 47675 31725
rect 44675 28733 44683 31717
rect 47667 28733 47675 31717
rect 44675 28725 47675 28733
rect 47865 31717 50865 31725
rect 47865 28733 47873 31717
rect 50857 28733 50865 31717
rect 47865 28725 50865 28733
rect 51055 31717 54055 31725
rect 51055 28733 51063 31717
rect 54047 28733 54055 31717
rect 51055 28725 54055 28733
rect 54245 31717 57245 31725
rect 54245 28733 54253 31717
rect 57237 28733 57245 31717
rect 54245 28725 57245 28733
rect 57435 31717 60435 31725
rect 57435 28733 57443 31717
rect 60427 28733 60435 31717
rect 57435 28725 60435 28733
rect 60625 31717 63625 31725
rect 60625 28733 60633 31717
rect 63617 28733 63625 31717
rect 60625 28725 63625 28733
rect 63815 31717 66815 31725
rect 63815 28733 63823 31717
rect 66807 28733 66815 31717
rect 63815 28725 66815 28733
rect 67005 31717 70005 31725
rect 67005 28733 67013 31717
rect 69997 28733 70005 31717
rect 67005 28725 70005 28733
rect 70195 31717 73195 31725
rect 70195 28733 70203 31717
rect 73187 28733 73195 31717
rect 70195 28725 73195 28733
rect 73385 31717 76385 31725
rect 73385 28733 73393 31717
rect 76377 28733 76385 31717
rect 73385 28725 76385 28733
rect 76575 31717 79575 31725
rect 76575 28733 76583 31717
rect 79567 28733 79575 31717
rect 76575 28725 79575 28733
rect 79765 31717 82765 31725
rect 79765 28733 79773 31717
rect 82757 28733 82765 31717
rect 79765 28725 82765 28733
rect 82955 31717 85955 31725
rect 82955 28733 82963 31717
rect 85947 28733 85955 31717
rect 82955 28725 85955 28733
rect 86145 31717 89145 31725
rect 86145 28733 86153 31717
rect 89137 28733 89145 31717
rect 86145 28725 89145 28733
rect 89335 31717 92335 31725
rect 89335 28733 89343 31717
rect 92327 28733 92335 31717
rect 89335 28725 92335 28733
rect 92525 31717 95525 31725
rect 92525 28733 92533 31717
rect 95517 28733 95525 31717
rect 92525 28725 95525 28733
rect 95715 31717 98715 31725
rect 95715 28733 95723 31717
rect 98707 28733 98715 31717
rect 95715 28725 98715 28733
rect 98905 31717 101905 31725
rect 98905 28733 98913 31717
rect 101897 28733 101905 31717
rect 98905 28725 101905 28733
rect 102095 31717 105095 31725
rect 102095 28733 102103 31717
rect 105087 28733 105095 31717
rect 102095 28725 105095 28733
rect 105285 31717 108285 31725
rect 105285 28733 105293 31717
rect 108277 28733 108285 31717
rect 105285 28725 108285 28733
rect 108475 31717 111475 31725
rect 108475 28733 108483 31717
rect 111467 28733 111475 31717
rect 108475 28725 111475 28733
rect 111665 31717 114665 31725
rect 111665 28733 111673 31717
rect 114657 28733 114665 31717
rect 111665 28725 114665 28733
rect 114855 31717 117855 31725
rect 114855 28733 114863 31717
rect 117847 28733 117855 31717
rect 114855 28725 117855 28733
rect 118045 31717 121045 31725
rect 118045 28733 118053 31717
rect 121037 28733 121045 31717
rect 118045 28725 121045 28733
rect 121235 31717 124235 31725
rect 121235 28733 121243 31717
rect 124227 28733 124235 31717
rect 121235 28725 124235 28733
rect 124425 31717 127425 31725
rect 124425 28733 124433 31717
rect 127417 28733 127425 31717
rect 124425 28725 127425 28733
rect 127615 31717 130615 31725
rect 127615 28733 127623 31717
rect 130607 28733 130615 31717
rect 127615 28725 130615 28733
rect 130805 31717 133805 31725
rect 130805 28733 130813 31717
rect 133797 28733 133805 31717
rect 130805 28725 133805 28733
rect 133995 31717 136995 31725
rect 133995 28733 134003 31717
rect 136987 28733 136995 31717
rect 133995 28725 136995 28733
rect 15 28527 3015 28535
rect 15 25543 23 28527
rect 3007 25543 3015 28527
rect 15 25535 3015 25543
rect 3205 28527 6205 28535
rect 3205 25543 3213 28527
rect 6197 25543 6205 28527
rect 3205 25535 6205 25543
rect 6395 28527 9395 28535
rect 6395 25543 6403 28527
rect 9387 25543 9395 28527
rect 6395 25535 9395 25543
rect 9585 28527 12585 28535
rect 9585 25543 9593 28527
rect 12577 25543 12585 28527
rect 9585 25535 12585 25543
rect 12775 28527 15775 28535
rect 12775 25543 12783 28527
rect 15767 25543 15775 28527
rect 12775 25535 15775 25543
rect 15965 28527 18965 28535
rect 15965 25543 15973 28527
rect 18957 25543 18965 28527
rect 15965 25535 18965 25543
rect 19155 28527 22155 28535
rect 19155 25543 19163 28527
rect 22147 25543 22155 28527
rect 19155 25535 22155 25543
rect 22345 28527 25345 28535
rect 22345 25543 22353 28527
rect 25337 25543 25345 28527
rect 22345 25535 25345 25543
rect 25535 28527 28535 28535
rect 25535 25543 25543 28527
rect 28527 25543 28535 28527
rect 25535 25535 28535 25543
rect 28725 28527 31725 28535
rect 28725 25543 28733 28527
rect 31717 25543 31725 28527
rect 28725 25535 31725 25543
rect 31915 28527 34915 28535
rect 31915 25543 31923 28527
rect 34907 25543 34915 28527
rect 31915 25535 34915 25543
rect 35105 28527 38105 28535
rect 35105 25543 35113 28527
rect 38097 25543 38105 28527
rect 35105 25535 38105 25543
rect 38295 28527 41295 28535
rect 38295 25543 38303 28527
rect 41287 25543 41295 28527
rect 38295 25535 41295 25543
rect 41485 28527 44485 28535
rect 41485 25543 41493 28527
rect 44477 25543 44485 28527
rect 41485 25535 44485 25543
rect 44675 28527 47675 28535
rect 44675 25543 44683 28527
rect 47667 25543 47675 28527
rect 44675 25535 47675 25543
rect 47865 28527 50865 28535
rect 47865 25543 47873 28527
rect 50857 25543 50865 28527
rect 47865 25535 50865 25543
rect 51055 28527 54055 28535
rect 51055 25543 51063 28527
rect 54047 25543 54055 28527
rect 51055 25535 54055 25543
rect 54245 28527 57245 28535
rect 54245 25543 54253 28527
rect 57237 25543 57245 28527
rect 54245 25535 57245 25543
rect 57435 28527 60435 28535
rect 57435 25543 57443 28527
rect 60427 25543 60435 28527
rect 57435 25535 60435 25543
rect 60625 28527 63625 28535
rect 60625 25543 60633 28527
rect 63617 25543 63625 28527
rect 60625 25535 63625 25543
rect 63815 28527 66815 28535
rect 63815 25543 63823 28527
rect 66807 25543 66815 28527
rect 63815 25535 66815 25543
rect 67005 28527 70005 28535
rect 67005 25543 67013 28527
rect 69997 25543 70005 28527
rect 67005 25535 70005 25543
rect 70195 28527 73195 28535
rect 70195 25543 70203 28527
rect 73187 25543 73195 28527
rect 70195 25535 73195 25543
rect 73385 28527 76385 28535
rect 73385 25543 73393 28527
rect 76377 25543 76385 28527
rect 73385 25535 76385 25543
rect 76575 28527 79575 28535
rect 76575 25543 76583 28527
rect 79567 25543 79575 28527
rect 76575 25535 79575 25543
rect 79765 28527 82765 28535
rect 79765 25543 79773 28527
rect 82757 25543 82765 28527
rect 79765 25535 82765 25543
rect 82955 28527 85955 28535
rect 82955 25543 82963 28527
rect 85947 25543 85955 28527
rect 82955 25535 85955 25543
rect 86145 28527 89145 28535
rect 86145 25543 86153 28527
rect 89137 25543 89145 28527
rect 86145 25535 89145 25543
rect 89335 28527 92335 28535
rect 89335 25543 89343 28527
rect 92327 25543 92335 28527
rect 89335 25535 92335 25543
rect 92525 28527 95525 28535
rect 92525 25543 92533 28527
rect 95517 25543 95525 28527
rect 92525 25535 95525 25543
rect 95715 28527 98715 28535
rect 95715 25543 95723 28527
rect 98707 25543 98715 28527
rect 95715 25535 98715 25543
rect 98905 28527 101905 28535
rect 98905 25543 98913 28527
rect 101897 25543 101905 28527
rect 98905 25535 101905 25543
rect 102095 28527 105095 28535
rect 102095 25543 102103 28527
rect 105087 25543 105095 28527
rect 102095 25535 105095 25543
rect 105285 28527 108285 28535
rect 105285 25543 105293 28527
rect 108277 25543 108285 28527
rect 105285 25535 108285 25543
rect 108475 28527 111475 28535
rect 108475 25543 108483 28527
rect 111467 25543 111475 28527
rect 108475 25535 111475 25543
rect 111665 28527 114665 28535
rect 111665 25543 111673 28527
rect 114657 25543 114665 28527
rect 111665 25535 114665 25543
rect 114855 28527 117855 28535
rect 114855 25543 114863 28527
rect 117847 25543 117855 28527
rect 114855 25535 117855 25543
rect 118045 28527 121045 28535
rect 118045 25543 118053 28527
rect 121037 25543 121045 28527
rect 118045 25535 121045 25543
rect 121235 28527 124235 28535
rect 121235 25543 121243 28527
rect 124227 25543 124235 28527
rect 121235 25535 124235 25543
rect 124425 28527 127425 28535
rect 124425 25543 124433 28527
rect 127417 25543 127425 28527
rect 124425 25535 127425 25543
rect 127615 28527 130615 28535
rect 127615 25543 127623 28527
rect 130607 25543 130615 28527
rect 127615 25535 130615 25543
rect 130805 28527 133805 28535
rect 130805 25543 130813 28527
rect 133797 25543 133805 28527
rect 130805 25535 133805 25543
rect 133995 28527 136995 28535
rect 133995 25543 134003 28527
rect 136987 25543 136995 28527
rect 133995 25535 136995 25543
rect 15 25337 3015 25345
rect 15 22353 23 25337
rect 3007 22353 3015 25337
rect 15 22345 3015 22353
rect 3205 25337 6205 25345
rect 3205 22353 3213 25337
rect 6197 22353 6205 25337
rect 3205 22345 6205 22353
rect 6395 25337 9395 25345
rect 6395 22353 6403 25337
rect 9387 22353 9395 25337
rect 6395 22345 9395 22353
rect 9585 25337 12585 25345
rect 9585 22353 9593 25337
rect 12577 22353 12585 25337
rect 9585 22345 12585 22353
rect 12775 25337 15775 25345
rect 12775 22353 12783 25337
rect 15767 22353 15775 25337
rect 12775 22345 15775 22353
rect 15965 25337 18965 25345
rect 15965 22353 15973 25337
rect 18957 22353 18965 25337
rect 15965 22345 18965 22353
rect 19155 25337 22155 25345
rect 19155 22353 19163 25337
rect 22147 22353 22155 25337
rect 19155 22345 22155 22353
rect 22345 25337 25345 25345
rect 22345 22353 22353 25337
rect 25337 22353 25345 25337
rect 22345 22345 25345 22353
rect 25535 25337 28535 25345
rect 25535 22353 25543 25337
rect 28527 22353 28535 25337
rect 25535 22345 28535 22353
rect 28725 25337 31725 25345
rect 28725 22353 28733 25337
rect 31717 22353 31725 25337
rect 28725 22345 31725 22353
rect 31915 25337 34915 25345
rect 31915 22353 31923 25337
rect 34907 22353 34915 25337
rect 31915 22345 34915 22353
rect 35105 25337 38105 25345
rect 35105 22353 35113 25337
rect 38097 22353 38105 25337
rect 35105 22345 38105 22353
rect 38295 25337 41295 25345
rect 38295 22353 38303 25337
rect 41287 22353 41295 25337
rect 38295 22345 41295 22353
rect 41485 25337 44485 25345
rect 41485 22353 41493 25337
rect 44477 22353 44485 25337
rect 41485 22345 44485 22353
rect 44675 25337 47675 25345
rect 44675 22353 44683 25337
rect 47667 22353 47675 25337
rect 44675 22345 47675 22353
rect 47865 25337 50865 25345
rect 47865 22353 47873 25337
rect 50857 22353 50865 25337
rect 47865 22345 50865 22353
rect 51055 25337 54055 25345
rect 51055 22353 51063 25337
rect 54047 22353 54055 25337
rect 51055 22345 54055 22353
rect 54245 25337 57245 25345
rect 54245 22353 54253 25337
rect 57237 22353 57245 25337
rect 54245 22345 57245 22353
rect 57435 25337 60435 25345
rect 57435 22353 57443 25337
rect 60427 22353 60435 25337
rect 57435 22345 60435 22353
rect 60625 25337 63625 25345
rect 60625 22353 60633 25337
rect 63617 22353 63625 25337
rect 60625 22345 63625 22353
rect 63815 25337 66815 25345
rect 63815 22353 63823 25337
rect 66807 22353 66815 25337
rect 63815 22345 66815 22353
rect 67005 25337 70005 25345
rect 67005 22353 67013 25337
rect 69997 22353 70005 25337
rect 67005 22345 70005 22353
rect 70195 25337 73195 25345
rect 70195 22353 70203 25337
rect 73187 22353 73195 25337
rect 70195 22345 73195 22353
rect 73385 25337 76385 25345
rect 73385 22353 73393 25337
rect 76377 22353 76385 25337
rect 73385 22345 76385 22353
rect 76575 25337 79575 25345
rect 76575 22353 76583 25337
rect 79567 22353 79575 25337
rect 76575 22345 79575 22353
rect 79765 25337 82765 25345
rect 79765 22353 79773 25337
rect 82757 22353 82765 25337
rect 79765 22345 82765 22353
rect 82955 25337 85955 25345
rect 82955 22353 82963 25337
rect 85947 22353 85955 25337
rect 82955 22345 85955 22353
rect 86145 25337 89145 25345
rect 86145 22353 86153 25337
rect 89137 22353 89145 25337
rect 86145 22345 89145 22353
rect 89335 25337 92335 25345
rect 89335 22353 89343 25337
rect 92327 22353 92335 25337
rect 89335 22345 92335 22353
rect 92525 25337 95525 25345
rect 92525 22353 92533 25337
rect 95517 22353 95525 25337
rect 92525 22345 95525 22353
rect 95715 25337 98715 25345
rect 95715 22353 95723 25337
rect 98707 22353 98715 25337
rect 95715 22345 98715 22353
rect 98905 25337 101905 25345
rect 98905 22353 98913 25337
rect 101897 22353 101905 25337
rect 98905 22345 101905 22353
rect 102095 25337 105095 25345
rect 102095 22353 102103 25337
rect 105087 22353 105095 25337
rect 102095 22345 105095 22353
rect 105285 25337 108285 25345
rect 105285 22353 105293 25337
rect 108277 22353 108285 25337
rect 105285 22345 108285 22353
rect 108475 25337 111475 25345
rect 108475 22353 108483 25337
rect 111467 22353 111475 25337
rect 108475 22345 111475 22353
rect 111665 25337 114665 25345
rect 111665 22353 111673 25337
rect 114657 22353 114665 25337
rect 111665 22345 114665 22353
rect 114855 25337 117855 25345
rect 114855 22353 114863 25337
rect 117847 22353 117855 25337
rect 114855 22345 117855 22353
rect 118045 25337 121045 25345
rect 118045 22353 118053 25337
rect 121037 22353 121045 25337
rect 118045 22345 121045 22353
rect 121235 25337 124235 25345
rect 121235 22353 121243 25337
rect 124227 22353 124235 25337
rect 121235 22345 124235 22353
rect 124425 25337 127425 25345
rect 124425 22353 124433 25337
rect 127417 22353 127425 25337
rect 124425 22345 127425 22353
rect 127615 25337 130615 25345
rect 127615 22353 127623 25337
rect 130607 22353 130615 25337
rect 127615 22345 130615 22353
rect 130805 25337 133805 25345
rect 130805 22353 130813 25337
rect 133797 22353 133805 25337
rect 130805 22345 133805 22353
rect 133995 25337 136995 25345
rect 133995 22353 134003 25337
rect 136987 22353 136995 25337
rect 133995 22345 136995 22353
rect 15 22147 3015 22155
rect 15 19163 23 22147
rect 3007 19163 3015 22147
rect 15 19155 3015 19163
rect 3205 22147 6205 22155
rect 3205 19163 3213 22147
rect 6197 19163 6205 22147
rect 3205 19155 6205 19163
rect 6395 22147 9395 22155
rect 6395 19163 6403 22147
rect 9387 19163 9395 22147
rect 6395 19155 9395 19163
rect 9585 22147 12585 22155
rect 9585 19163 9593 22147
rect 12577 19163 12585 22147
rect 9585 19155 12585 19163
rect 12775 22147 15775 22155
rect 12775 19163 12783 22147
rect 15767 19163 15775 22147
rect 12775 19155 15775 19163
rect 15965 22147 18965 22155
rect 15965 19163 15973 22147
rect 18957 19163 18965 22147
rect 15965 19155 18965 19163
rect 19155 22147 22155 22155
rect 19155 19163 19163 22147
rect 22147 19163 22155 22147
rect 19155 19155 22155 19163
rect 22345 22147 25345 22155
rect 22345 19163 22353 22147
rect 25337 19163 25345 22147
rect 22345 19155 25345 19163
rect 25535 22147 28535 22155
rect 25535 19163 25543 22147
rect 28527 19163 28535 22147
rect 25535 19155 28535 19163
rect 28725 22147 31725 22155
rect 28725 19163 28733 22147
rect 31717 19163 31725 22147
rect 28725 19155 31725 19163
rect 31915 22147 34915 22155
rect 31915 19163 31923 22147
rect 34907 19163 34915 22147
rect 31915 19155 34915 19163
rect 35105 22147 38105 22155
rect 35105 19163 35113 22147
rect 38097 19163 38105 22147
rect 35105 19155 38105 19163
rect 38295 22147 41295 22155
rect 38295 19163 38303 22147
rect 41287 19163 41295 22147
rect 38295 19155 41295 19163
rect 41485 22147 44485 22155
rect 41485 19163 41493 22147
rect 44477 19163 44485 22147
rect 41485 19155 44485 19163
rect 44675 22147 47675 22155
rect 44675 19163 44683 22147
rect 47667 19163 47675 22147
rect 44675 19155 47675 19163
rect 47865 22147 50865 22155
rect 47865 19163 47873 22147
rect 50857 19163 50865 22147
rect 47865 19155 50865 19163
rect 51055 22147 54055 22155
rect 51055 19163 51063 22147
rect 54047 19163 54055 22147
rect 51055 19155 54055 19163
rect 54245 22147 57245 22155
rect 54245 19163 54253 22147
rect 57237 19163 57245 22147
rect 54245 19155 57245 19163
rect 57435 22147 60435 22155
rect 57435 19163 57443 22147
rect 60427 19163 60435 22147
rect 57435 19155 60435 19163
rect 60625 22147 63625 22155
rect 60625 19163 60633 22147
rect 63617 19163 63625 22147
rect 60625 19155 63625 19163
rect 63815 22147 66815 22155
rect 63815 19163 63823 22147
rect 66807 19163 66815 22147
rect 63815 19155 66815 19163
rect 67005 22147 70005 22155
rect 67005 19163 67013 22147
rect 69997 19163 70005 22147
rect 67005 19155 70005 19163
rect 70195 22147 73195 22155
rect 70195 19163 70203 22147
rect 73187 19163 73195 22147
rect 70195 19155 73195 19163
rect 73385 22147 76385 22155
rect 73385 19163 73393 22147
rect 76377 19163 76385 22147
rect 73385 19155 76385 19163
rect 76575 22147 79575 22155
rect 76575 19163 76583 22147
rect 79567 19163 79575 22147
rect 76575 19155 79575 19163
rect 79765 22147 82765 22155
rect 79765 19163 79773 22147
rect 82757 19163 82765 22147
rect 79765 19155 82765 19163
rect 82955 22147 85955 22155
rect 82955 19163 82963 22147
rect 85947 19163 85955 22147
rect 82955 19155 85955 19163
rect 86145 22147 89145 22155
rect 86145 19163 86153 22147
rect 89137 19163 89145 22147
rect 86145 19155 89145 19163
rect 89335 22147 92335 22155
rect 89335 19163 89343 22147
rect 92327 19163 92335 22147
rect 89335 19155 92335 19163
rect 92525 22147 95525 22155
rect 92525 19163 92533 22147
rect 95517 19163 95525 22147
rect 92525 19155 95525 19163
rect 95715 22147 98715 22155
rect 95715 19163 95723 22147
rect 98707 19163 98715 22147
rect 95715 19155 98715 19163
rect 98905 22147 101905 22155
rect 98905 19163 98913 22147
rect 101897 19163 101905 22147
rect 98905 19155 101905 19163
rect 102095 22147 105095 22155
rect 102095 19163 102103 22147
rect 105087 19163 105095 22147
rect 102095 19155 105095 19163
rect 105285 22147 108285 22155
rect 105285 19163 105293 22147
rect 108277 19163 108285 22147
rect 105285 19155 108285 19163
rect 108475 22147 111475 22155
rect 108475 19163 108483 22147
rect 111467 19163 111475 22147
rect 108475 19155 111475 19163
rect 111665 22147 114665 22155
rect 111665 19163 111673 22147
rect 114657 19163 114665 22147
rect 111665 19155 114665 19163
rect 114855 22147 117855 22155
rect 114855 19163 114863 22147
rect 117847 19163 117855 22147
rect 114855 19155 117855 19163
rect 118045 22147 121045 22155
rect 118045 19163 118053 22147
rect 121037 19163 121045 22147
rect 118045 19155 121045 19163
rect 121235 22147 124235 22155
rect 121235 19163 121243 22147
rect 124227 19163 124235 22147
rect 121235 19155 124235 19163
rect 124425 22147 127425 22155
rect 124425 19163 124433 22147
rect 127417 19163 127425 22147
rect 124425 19155 127425 19163
rect 127615 22147 130615 22155
rect 127615 19163 127623 22147
rect 130607 19163 130615 22147
rect 127615 19155 130615 19163
rect 130805 22147 133805 22155
rect 130805 19163 130813 22147
rect 133797 19163 133805 22147
rect 130805 19155 133805 19163
rect 133995 22147 136995 22155
rect 133995 19163 134003 22147
rect 136987 19163 136995 22147
rect 133995 19155 136995 19163
rect 15 18957 3015 18965
rect 15 15973 23 18957
rect 3007 15973 3015 18957
rect 15 15965 3015 15973
rect 3205 18957 6205 18965
rect 3205 15973 3213 18957
rect 6197 15973 6205 18957
rect 3205 15965 6205 15973
rect 6395 18957 9395 18965
rect 6395 15973 6403 18957
rect 9387 15973 9395 18957
rect 6395 15965 9395 15973
rect 9585 18957 12585 18965
rect 9585 15973 9593 18957
rect 12577 15973 12585 18957
rect 9585 15965 12585 15973
rect 12775 18957 15775 18965
rect 12775 15973 12783 18957
rect 15767 15973 15775 18957
rect 12775 15965 15775 15973
rect 15965 18957 18965 18965
rect 15965 15973 15973 18957
rect 18957 15973 18965 18957
rect 15965 15965 18965 15973
rect 19155 18957 22155 18965
rect 19155 15973 19163 18957
rect 22147 15973 22155 18957
rect 19155 15965 22155 15973
rect 22345 18957 25345 18965
rect 22345 15973 22353 18957
rect 25337 15973 25345 18957
rect 22345 15965 25345 15973
rect 25535 18957 28535 18965
rect 25535 15973 25543 18957
rect 28527 15973 28535 18957
rect 25535 15965 28535 15973
rect 28725 18957 31725 18965
rect 28725 15973 28733 18957
rect 31717 15973 31725 18957
rect 28725 15965 31725 15973
rect 31915 18957 34915 18965
rect 31915 15973 31923 18957
rect 34907 15973 34915 18957
rect 31915 15965 34915 15973
rect 35105 18957 38105 18965
rect 35105 15973 35113 18957
rect 38097 15973 38105 18957
rect 35105 15965 38105 15973
rect 38295 18957 41295 18965
rect 38295 15973 38303 18957
rect 41287 15973 41295 18957
rect 38295 15965 41295 15973
rect 41485 18957 44485 18965
rect 41485 15973 41493 18957
rect 44477 15973 44485 18957
rect 41485 15965 44485 15973
rect 44675 18957 47675 18965
rect 44675 15973 44683 18957
rect 47667 15973 47675 18957
rect 44675 15965 47675 15973
rect 47865 18957 50865 18965
rect 47865 15973 47873 18957
rect 50857 15973 50865 18957
rect 47865 15965 50865 15973
rect 51055 18957 54055 18965
rect 51055 15973 51063 18957
rect 54047 15973 54055 18957
rect 51055 15965 54055 15973
rect 54245 18957 57245 18965
rect 54245 15973 54253 18957
rect 57237 15973 57245 18957
rect 54245 15965 57245 15973
rect 57435 18957 60435 18965
rect 57435 15973 57443 18957
rect 60427 15973 60435 18957
rect 57435 15965 60435 15973
rect 60625 18957 63625 18965
rect 60625 15973 60633 18957
rect 63617 15973 63625 18957
rect 60625 15965 63625 15973
rect 63815 18957 66815 18965
rect 63815 15973 63823 18957
rect 66807 15973 66815 18957
rect 63815 15965 66815 15973
rect 67005 18957 70005 18965
rect 67005 15973 67013 18957
rect 69997 15973 70005 18957
rect 67005 15965 70005 15973
rect 70195 18957 73195 18965
rect 70195 15973 70203 18957
rect 73187 15973 73195 18957
rect 70195 15965 73195 15973
rect 73385 18957 76385 18965
rect 73385 15973 73393 18957
rect 76377 15973 76385 18957
rect 73385 15965 76385 15973
rect 76575 18957 79575 18965
rect 76575 15973 76583 18957
rect 79567 15973 79575 18957
rect 76575 15965 79575 15973
rect 79765 18957 82765 18965
rect 79765 15973 79773 18957
rect 82757 15973 82765 18957
rect 79765 15965 82765 15973
rect 82955 18957 85955 18965
rect 82955 15973 82963 18957
rect 85947 15973 85955 18957
rect 82955 15965 85955 15973
rect 86145 18957 89145 18965
rect 86145 15973 86153 18957
rect 89137 15973 89145 18957
rect 86145 15965 89145 15973
rect 89335 18957 92335 18965
rect 89335 15973 89343 18957
rect 92327 15973 92335 18957
rect 89335 15965 92335 15973
rect 92525 18957 95525 18965
rect 92525 15973 92533 18957
rect 95517 15973 95525 18957
rect 92525 15965 95525 15973
rect 95715 18957 98715 18965
rect 95715 15973 95723 18957
rect 98707 15973 98715 18957
rect 95715 15965 98715 15973
rect 98905 18957 101905 18965
rect 98905 15973 98913 18957
rect 101897 15973 101905 18957
rect 98905 15965 101905 15973
rect 102095 18957 105095 18965
rect 102095 15973 102103 18957
rect 105087 15973 105095 18957
rect 102095 15965 105095 15973
rect 105285 18957 108285 18965
rect 105285 15973 105293 18957
rect 108277 15973 108285 18957
rect 105285 15965 108285 15973
rect 108475 18957 111475 18965
rect 108475 15973 108483 18957
rect 111467 15973 111475 18957
rect 108475 15965 111475 15973
rect 111665 18957 114665 18965
rect 111665 15973 111673 18957
rect 114657 15973 114665 18957
rect 111665 15965 114665 15973
rect 114855 18957 117855 18965
rect 114855 15973 114863 18957
rect 117847 15973 117855 18957
rect 114855 15965 117855 15973
rect 118045 18957 121045 18965
rect 118045 15973 118053 18957
rect 121037 15973 121045 18957
rect 118045 15965 121045 15973
rect 121235 18957 124235 18965
rect 121235 15973 121243 18957
rect 124227 15973 124235 18957
rect 121235 15965 124235 15973
rect 124425 18957 127425 18965
rect 124425 15973 124433 18957
rect 127417 15973 127425 18957
rect 124425 15965 127425 15973
rect 127615 18957 130615 18965
rect 127615 15973 127623 18957
rect 130607 15973 130615 18957
rect 127615 15965 130615 15973
rect 130805 18957 133805 18965
rect 130805 15973 130813 18957
rect 133797 15973 133805 18957
rect 130805 15965 133805 15973
rect 133995 18957 136995 18965
rect 133995 15973 134003 18957
rect 136987 15973 136995 18957
rect 133995 15965 136995 15973
rect 15 15767 3015 15775
rect 15 12783 23 15767
rect 3007 12783 3015 15767
rect 15 12775 3015 12783
rect 3205 15767 6205 15775
rect 3205 12783 3213 15767
rect 6197 12783 6205 15767
rect 3205 12775 6205 12783
rect 6395 15767 9395 15775
rect 6395 12783 6403 15767
rect 9387 12783 9395 15767
rect 6395 12775 9395 12783
rect 9585 15767 12585 15775
rect 9585 12783 9593 15767
rect 12577 12783 12585 15767
rect 9585 12775 12585 12783
rect 12775 15767 15775 15775
rect 12775 12783 12783 15767
rect 15767 12783 15775 15767
rect 12775 12775 15775 12783
rect 15965 15767 18965 15775
rect 15965 12783 15973 15767
rect 18957 12783 18965 15767
rect 15965 12775 18965 12783
rect 19155 15767 22155 15775
rect 19155 12783 19163 15767
rect 22147 12783 22155 15767
rect 19155 12775 22155 12783
rect 22345 15767 25345 15775
rect 22345 12783 22353 15767
rect 25337 12783 25345 15767
rect 22345 12775 25345 12783
rect 25535 15767 28535 15775
rect 25535 12783 25543 15767
rect 28527 12783 28535 15767
rect 25535 12775 28535 12783
rect 28725 15767 31725 15775
rect 28725 12783 28733 15767
rect 31717 12783 31725 15767
rect 28725 12775 31725 12783
rect 31915 15767 34915 15775
rect 31915 12783 31923 15767
rect 34907 12783 34915 15767
rect 31915 12775 34915 12783
rect 35105 15767 38105 15775
rect 35105 12783 35113 15767
rect 38097 12783 38105 15767
rect 35105 12775 38105 12783
rect 38295 15767 41295 15775
rect 38295 12783 38303 15767
rect 41287 12783 41295 15767
rect 38295 12775 41295 12783
rect 41485 15767 44485 15775
rect 41485 12783 41493 15767
rect 44477 12783 44485 15767
rect 41485 12775 44485 12783
rect 44675 15767 47675 15775
rect 44675 12783 44683 15767
rect 47667 12783 47675 15767
rect 44675 12775 47675 12783
rect 47865 15767 50865 15775
rect 47865 12783 47873 15767
rect 50857 12783 50865 15767
rect 47865 12775 50865 12783
rect 51055 15767 54055 15775
rect 51055 12783 51063 15767
rect 54047 12783 54055 15767
rect 51055 12775 54055 12783
rect 54245 15767 57245 15775
rect 54245 12783 54253 15767
rect 57237 12783 57245 15767
rect 54245 12775 57245 12783
rect 57435 15767 60435 15775
rect 57435 12783 57443 15767
rect 60427 12783 60435 15767
rect 57435 12775 60435 12783
rect 60625 15767 63625 15775
rect 60625 12783 60633 15767
rect 63617 12783 63625 15767
rect 60625 12775 63625 12783
rect 63815 15767 66815 15775
rect 63815 12783 63823 15767
rect 66807 12783 66815 15767
rect 63815 12775 66815 12783
rect 67005 15767 70005 15775
rect 67005 12783 67013 15767
rect 69997 12783 70005 15767
rect 67005 12775 70005 12783
rect 70195 15767 73195 15775
rect 70195 12783 70203 15767
rect 73187 12783 73195 15767
rect 70195 12775 73195 12783
rect 73385 15767 76385 15775
rect 73385 12783 73393 15767
rect 76377 12783 76385 15767
rect 73385 12775 76385 12783
rect 76575 15767 79575 15775
rect 76575 12783 76583 15767
rect 79567 12783 79575 15767
rect 76575 12775 79575 12783
rect 79765 15767 82765 15775
rect 79765 12783 79773 15767
rect 82757 12783 82765 15767
rect 79765 12775 82765 12783
rect 82955 15767 85955 15775
rect 82955 12783 82963 15767
rect 85947 12783 85955 15767
rect 82955 12775 85955 12783
rect 86145 15767 89145 15775
rect 86145 12783 86153 15767
rect 89137 12783 89145 15767
rect 86145 12775 89145 12783
rect 89335 15767 92335 15775
rect 89335 12783 89343 15767
rect 92327 12783 92335 15767
rect 89335 12775 92335 12783
rect 92525 15767 95525 15775
rect 92525 12783 92533 15767
rect 95517 12783 95525 15767
rect 92525 12775 95525 12783
rect 95715 15767 98715 15775
rect 95715 12783 95723 15767
rect 98707 12783 98715 15767
rect 95715 12775 98715 12783
rect 98905 15767 101905 15775
rect 98905 12783 98913 15767
rect 101897 12783 101905 15767
rect 98905 12775 101905 12783
rect 102095 15767 105095 15775
rect 102095 12783 102103 15767
rect 105087 12783 105095 15767
rect 102095 12775 105095 12783
rect 105285 15767 108285 15775
rect 105285 12783 105293 15767
rect 108277 12783 108285 15767
rect 105285 12775 108285 12783
rect 108475 15767 111475 15775
rect 108475 12783 108483 15767
rect 111467 12783 111475 15767
rect 108475 12775 111475 12783
rect 111665 15767 114665 15775
rect 111665 12783 111673 15767
rect 114657 12783 114665 15767
rect 111665 12775 114665 12783
rect 114855 15767 117855 15775
rect 114855 12783 114863 15767
rect 117847 12783 117855 15767
rect 114855 12775 117855 12783
rect 118045 15767 121045 15775
rect 118045 12783 118053 15767
rect 121037 12783 121045 15767
rect 118045 12775 121045 12783
rect 121235 15767 124235 15775
rect 121235 12783 121243 15767
rect 124227 12783 124235 15767
rect 121235 12775 124235 12783
rect 124425 15767 127425 15775
rect 124425 12783 124433 15767
rect 127417 12783 127425 15767
rect 124425 12775 127425 12783
rect 127615 15767 130615 15775
rect 127615 12783 127623 15767
rect 130607 12783 130615 15767
rect 127615 12775 130615 12783
rect 130805 15767 133805 15775
rect 130805 12783 130813 15767
rect 133797 12783 133805 15767
rect 130805 12775 133805 12783
rect 133995 15767 136995 15775
rect 133995 12783 134003 15767
rect 136987 12783 136995 15767
rect 133995 12775 136995 12783
rect 15 12577 3015 12585
rect 15 9593 23 12577
rect 3007 9593 3015 12577
rect 15 9585 3015 9593
rect 3205 12577 6205 12585
rect 3205 9593 3213 12577
rect 6197 9593 6205 12577
rect 3205 9585 6205 9593
rect 6395 12577 9395 12585
rect 6395 9593 6403 12577
rect 9387 9593 9395 12577
rect 6395 9585 9395 9593
rect 9585 12577 12585 12585
rect 9585 9593 9593 12577
rect 12577 9593 12585 12577
rect 9585 9585 12585 9593
rect 12775 12577 15775 12585
rect 12775 9593 12783 12577
rect 15767 9593 15775 12577
rect 12775 9585 15775 9593
rect 15965 12577 18965 12585
rect 15965 9593 15973 12577
rect 18957 9593 18965 12577
rect 15965 9585 18965 9593
rect 19155 12577 22155 12585
rect 19155 9593 19163 12577
rect 22147 9593 22155 12577
rect 19155 9585 22155 9593
rect 22345 12577 25345 12585
rect 22345 9593 22353 12577
rect 25337 9593 25345 12577
rect 22345 9585 25345 9593
rect 25535 12577 28535 12585
rect 25535 9593 25543 12577
rect 28527 9593 28535 12577
rect 25535 9585 28535 9593
rect 28725 12577 31725 12585
rect 28725 9593 28733 12577
rect 31717 9593 31725 12577
rect 28725 9585 31725 9593
rect 31915 12577 34915 12585
rect 31915 9593 31923 12577
rect 34907 9593 34915 12577
rect 31915 9585 34915 9593
rect 35105 12577 38105 12585
rect 35105 9593 35113 12577
rect 38097 9593 38105 12577
rect 35105 9585 38105 9593
rect 38295 12577 41295 12585
rect 38295 9593 38303 12577
rect 41287 9593 41295 12577
rect 38295 9585 41295 9593
rect 41485 12577 44485 12585
rect 41485 9593 41493 12577
rect 44477 9593 44485 12577
rect 41485 9585 44485 9593
rect 44675 12577 47675 12585
rect 44675 9593 44683 12577
rect 47667 9593 47675 12577
rect 44675 9585 47675 9593
rect 47865 12577 50865 12585
rect 47865 9593 47873 12577
rect 50857 9593 50865 12577
rect 47865 9585 50865 9593
rect 51055 12577 54055 12585
rect 51055 9593 51063 12577
rect 54047 9593 54055 12577
rect 51055 9585 54055 9593
rect 54245 12577 57245 12585
rect 54245 9593 54253 12577
rect 57237 9593 57245 12577
rect 54245 9585 57245 9593
rect 57435 12577 60435 12585
rect 57435 9593 57443 12577
rect 60427 9593 60435 12577
rect 57435 9585 60435 9593
rect 60625 12577 63625 12585
rect 60625 9593 60633 12577
rect 63617 9593 63625 12577
rect 60625 9585 63625 9593
rect 63815 12577 66815 12585
rect 63815 9593 63823 12577
rect 66807 9593 66815 12577
rect 63815 9585 66815 9593
rect 67005 12577 70005 12585
rect 67005 9593 67013 12577
rect 69997 9593 70005 12577
rect 67005 9585 70005 9593
rect 70195 12577 73195 12585
rect 70195 9593 70203 12577
rect 73187 9593 73195 12577
rect 70195 9585 73195 9593
rect 73385 12577 76385 12585
rect 73385 9593 73393 12577
rect 76377 9593 76385 12577
rect 73385 9585 76385 9593
rect 76575 12577 79575 12585
rect 76575 9593 76583 12577
rect 79567 9593 79575 12577
rect 76575 9585 79575 9593
rect 79765 12577 82765 12585
rect 79765 9593 79773 12577
rect 82757 9593 82765 12577
rect 79765 9585 82765 9593
rect 82955 12577 85955 12585
rect 82955 9593 82963 12577
rect 85947 9593 85955 12577
rect 82955 9585 85955 9593
rect 86145 12577 89145 12585
rect 86145 9593 86153 12577
rect 89137 9593 89145 12577
rect 86145 9585 89145 9593
rect 89335 12577 92335 12585
rect 89335 9593 89343 12577
rect 92327 9593 92335 12577
rect 89335 9585 92335 9593
rect 92525 12577 95525 12585
rect 92525 9593 92533 12577
rect 95517 9593 95525 12577
rect 92525 9585 95525 9593
rect 95715 12577 98715 12585
rect 95715 9593 95723 12577
rect 98707 9593 98715 12577
rect 95715 9585 98715 9593
rect 98905 12577 101905 12585
rect 98905 9593 98913 12577
rect 101897 9593 101905 12577
rect 98905 9585 101905 9593
rect 102095 12577 105095 12585
rect 102095 9593 102103 12577
rect 105087 9593 105095 12577
rect 102095 9585 105095 9593
rect 105285 12577 108285 12585
rect 105285 9593 105293 12577
rect 108277 9593 108285 12577
rect 105285 9585 108285 9593
rect 108475 12577 111475 12585
rect 108475 9593 108483 12577
rect 111467 9593 111475 12577
rect 108475 9585 111475 9593
rect 111665 12577 114665 12585
rect 111665 9593 111673 12577
rect 114657 9593 114665 12577
rect 111665 9585 114665 9593
rect 114855 12577 117855 12585
rect 114855 9593 114863 12577
rect 117847 9593 117855 12577
rect 114855 9585 117855 9593
rect 118045 12577 121045 12585
rect 118045 9593 118053 12577
rect 121037 9593 121045 12577
rect 118045 9585 121045 9593
rect 121235 12577 124235 12585
rect 121235 9593 121243 12577
rect 124227 9593 124235 12577
rect 121235 9585 124235 9593
rect 124425 12577 127425 12585
rect 124425 9593 124433 12577
rect 127417 9593 127425 12577
rect 124425 9585 127425 9593
rect 127615 12577 130615 12585
rect 127615 9593 127623 12577
rect 130607 9593 130615 12577
rect 127615 9585 130615 9593
rect 130805 12577 133805 12585
rect 130805 9593 130813 12577
rect 133797 9593 133805 12577
rect 130805 9585 133805 9593
rect 133995 12577 136995 12585
rect 133995 9593 134003 12577
rect 136987 9593 136995 12577
rect 133995 9585 136995 9593
rect 15 9387 3015 9395
rect 15 6403 23 9387
rect 3007 6403 3015 9387
rect 15 6395 3015 6403
rect 3205 9387 6205 9395
rect 3205 6403 3213 9387
rect 6197 6403 6205 9387
rect 3205 6395 6205 6403
rect 6395 9387 9395 9395
rect 6395 6403 6403 9387
rect 9387 6403 9395 9387
rect 6395 6395 9395 6403
rect 9585 9387 12585 9395
rect 9585 6403 9593 9387
rect 12577 6403 12585 9387
rect 9585 6395 12585 6403
rect 12775 9387 15775 9395
rect 12775 6403 12783 9387
rect 15767 6403 15775 9387
rect 12775 6395 15775 6403
rect 15965 9387 18965 9395
rect 15965 6403 15973 9387
rect 18957 6403 18965 9387
rect 15965 6395 18965 6403
rect 19155 9387 22155 9395
rect 19155 6403 19163 9387
rect 22147 6403 22155 9387
rect 19155 6395 22155 6403
rect 22345 9387 25345 9395
rect 22345 6403 22353 9387
rect 25337 6403 25345 9387
rect 22345 6395 25345 6403
rect 25535 9387 28535 9395
rect 25535 6403 25543 9387
rect 28527 6403 28535 9387
rect 25535 6395 28535 6403
rect 28725 9387 31725 9395
rect 28725 6403 28733 9387
rect 31717 6403 31725 9387
rect 28725 6395 31725 6403
rect 31915 9387 34915 9395
rect 31915 6403 31923 9387
rect 34907 6403 34915 9387
rect 31915 6395 34915 6403
rect 35105 9387 38105 9395
rect 35105 6403 35113 9387
rect 38097 6403 38105 9387
rect 35105 6395 38105 6403
rect 38295 9387 41295 9395
rect 38295 6403 38303 9387
rect 41287 6403 41295 9387
rect 38295 6395 41295 6403
rect 41485 9387 44485 9395
rect 41485 6403 41493 9387
rect 44477 6403 44485 9387
rect 41485 6395 44485 6403
rect 44675 9387 47675 9395
rect 44675 6403 44683 9387
rect 47667 6403 47675 9387
rect 44675 6395 47675 6403
rect 47865 9387 50865 9395
rect 47865 6403 47873 9387
rect 50857 6403 50865 9387
rect 47865 6395 50865 6403
rect 51055 9387 54055 9395
rect 51055 6403 51063 9387
rect 54047 6403 54055 9387
rect 51055 6395 54055 6403
rect 54245 9387 57245 9395
rect 54245 6403 54253 9387
rect 57237 6403 57245 9387
rect 54245 6395 57245 6403
rect 57435 9387 60435 9395
rect 57435 6403 57443 9387
rect 60427 6403 60435 9387
rect 57435 6395 60435 6403
rect 60625 9387 63625 9395
rect 60625 6403 60633 9387
rect 63617 6403 63625 9387
rect 60625 6395 63625 6403
rect 63815 9387 66815 9395
rect 63815 6403 63823 9387
rect 66807 6403 66815 9387
rect 63815 6395 66815 6403
rect 67005 9387 70005 9395
rect 67005 6403 67013 9387
rect 69997 6403 70005 9387
rect 67005 6395 70005 6403
rect 70195 9387 73195 9395
rect 70195 6403 70203 9387
rect 73187 6403 73195 9387
rect 70195 6395 73195 6403
rect 73385 9387 76385 9395
rect 73385 6403 73393 9387
rect 76377 6403 76385 9387
rect 73385 6395 76385 6403
rect 76575 9387 79575 9395
rect 76575 6403 76583 9387
rect 79567 6403 79575 9387
rect 76575 6395 79575 6403
rect 79765 9387 82765 9395
rect 79765 6403 79773 9387
rect 82757 6403 82765 9387
rect 79765 6395 82765 6403
rect 82955 9387 85955 9395
rect 82955 6403 82963 9387
rect 85947 6403 85955 9387
rect 82955 6395 85955 6403
rect 86145 9387 89145 9395
rect 86145 6403 86153 9387
rect 89137 6403 89145 9387
rect 86145 6395 89145 6403
rect 89335 9387 92335 9395
rect 89335 6403 89343 9387
rect 92327 6403 92335 9387
rect 89335 6395 92335 6403
rect 92525 9387 95525 9395
rect 92525 6403 92533 9387
rect 95517 6403 95525 9387
rect 92525 6395 95525 6403
rect 95715 9387 98715 9395
rect 95715 6403 95723 9387
rect 98707 6403 98715 9387
rect 95715 6395 98715 6403
rect 98905 9387 101905 9395
rect 98905 6403 98913 9387
rect 101897 6403 101905 9387
rect 98905 6395 101905 6403
rect 102095 9387 105095 9395
rect 102095 6403 102103 9387
rect 105087 6403 105095 9387
rect 102095 6395 105095 6403
rect 105285 9387 108285 9395
rect 105285 6403 105293 9387
rect 108277 6403 108285 9387
rect 105285 6395 108285 6403
rect 108475 9387 111475 9395
rect 108475 6403 108483 9387
rect 111467 6403 111475 9387
rect 108475 6395 111475 6403
rect 111665 9387 114665 9395
rect 111665 6403 111673 9387
rect 114657 6403 114665 9387
rect 111665 6395 114665 6403
rect 114855 9387 117855 9395
rect 114855 6403 114863 9387
rect 117847 6403 117855 9387
rect 114855 6395 117855 6403
rect 118045 9387 121045 9395
rect 118045 6403 118053 9387
rect 121037 6403 121045 9387
rect 118045 6395 121045 6403
rect 121235 9387 124235 9395
rect 121235 6403 121243 9387
rect 124227 6403 124235 9387
rect 121235 6395 124235 6403
rect 124425 9387 127425 9395
rect 124425 6403 124433 9387
rect 127417 6403 127425 9387
rect 124425 6395 127425 6403
rect 127615 9387 130615 9395
rect 127615 6403 127623 9387
rect 130607 6403 130615 9387
rect 127615 6395 130615 6403
rect 130805 9387 133805 9395
rect 130805 6403 130813 9387
rect 133797 6403 133805 9387
rect 130805 6395 133805 6403
rect 133995 9387 136995 9395
rect 133995 6403 134003 9387
rect 136987 6403 136995 9387
rect 133995 6395 136995 6403
rect 15 6197 3015 6205
rect 15 3213 23 6197
rect 3007 3213 3015 6197
rect 15 3205 3015 3213
rect 3205 6197 6205 6205
rect 3205 3213 3213 6197
rect 6197 3213 6205 6197
rect 3205 3205 6205 3213
rect 6395 6197 9395 6205
rect 6395 3213 6403 6197
rect 9387 3213 9395 6197
rect 6395 3205 9395 3213
rect 9585 6197 12585 6205
rect 9585 3213 9593 6197
rect 12577 3213 12585 6197
rect 9585 3205 12585 3213
rect 12775 6197 15775 6205
rect 12775 3213 12783 6197
rect 15767 3213 15775 6197
rect 12775 3205 15775 3213
rect 15965 6197 18965 6205
rect 15965 3213 15973 6197
rect 18957 3213 18965 6197
rect 15965 3205 18965 3213
rect 19155 6197 22155 6205
rect 19155 3213 19163 6197
rect 22147 3213 22155 6197
rect 19155 3205 22155 3213
rect 22345 6197 25345 6205
rect 22345 3213 22353 6197
rect 25337 3213 25345 6197
rect 22345 3205 25345 3213
rect 25535 6197 28535 6205
rect 25535 3213 25543 6197
rect 28527 3213 28535 6197
rect 25535 3205 28535 3213
rect 28725 6197 31725 6205
rect 28725 3213 28733 6197
rect 31717 3213 31725 6197
rect 28725 3205 31725 3213
rect 31915 6197 34915 6205
rect 31915 3213 31923 6197
rect 34907 3213 34915 6197
rect 31915 3205 34915 3213
rect 35105 6197 38105 6205
rect 35105 3213 35113 6197
rect 38097 3213 38105 6197
rect 35105 3205 38105 3213
rect 38295 6197 41295 6205
rect 38295 3213 38303 6197
rect 41287 3213 41295 6197
rect 38295 3205 41295 3213
rect 41485 6197 44485 6205
rect 41485 3213 41493 6197
rect 44477 3213 44485 6197
rect 41485 3205 44485 3213
rect 44675 6197 47675 6205
rect 44675 3213 44683 6197
rect 47667 3213 47675 6197
rect 44675 3205 47675 3213
rect 47865 6197 50865 6205
rect 47865 3213 47873 6197
rect 50857 3213 50865 6197
rect 47865 3205 50865 3213
rect 51055 6197 54055 6205
rect 51055 3213 51063 6197
rect 54047 3213 54055 6197
rect 51055 3205 54055 3213
rect 54245 6197 57245 6205
rect 54245 3213 54253 6197
rect 57237 3213 57245 6197
rect 54245 3205 57245 3213
rect 57435 6197 60435 6205
rect 57435 3213 57443 6197
rect 60427 3213 60435 6197
rect 57435 3205 60435 3213
rect 60625 6197 63625 6205
rect 60625 3213 60633 6197
rect 63617 3213 63625 6197
rect 60625 3205 63625 3213
rect 63815 6197 66815 6205
rect 63815 3213 63823 6197
rect 66807 3213 66815 6197
rect 63815 3205 66815 3213
rect 67005 6197 70005 6205
rect 67005 3213 67013 6197
rect 69997 3213 70005 6197
rect 67005 3205 70005 3213
rect 70195 6197 73195 6205
rect 70195 3213 70203 6197
rect 73187 3213 73195 6197
rect 70195 3205 73195 3213
rect 73385 6197 76385 6205
rect 73385 3213 73393 6197
rect 76377 3213 76385 6197
rect 73385 3205 76385 3213
rect 76575 6197 79575 6205
rect 76575 3213 76583 6197
rect 79567 3213 79575 6197
rect 76575 3205 79575 3213
rect 79765 6197 82765 6205
rect 79765 3213 79773 6197
rect 82757 3213 82765 6197
rect 79765 3205 82765 3213
rect 82955 6197 85955 6205
rect 82955 3213 82963 6197
rect 85947 3213 85955 6197
rect 82955 3205 85955 3213
rect 86145 6197 89145 6205
rect 86145 3213 86153 6197
rect 89137 3213 89145 6197
rect 86145 3205 89145 3213
rect 89335 6197 92335 6205
rect 89335 3213 89343 6197
rect 92327 3213 92335 6197
rect 89335 3205 92335 3213
rect 92525 6197 95525 6205
rect 92525 3213 92533 6197
rect 95517 3213 95525 6197
rect 92525 3205 95525 3213
rect 95715 6197 98715 6205
rect 95715 3213 95723 6197
rect 98707 3213 98715 6197
rect 95715 3205 98715 3213
rect 98905 6197 101905 6205
rect 98905 3213 98913 6197
rect 101897 3213 101905 6197
rect 98905 3205 101905 3213
rect 102095 6197 105095 6205
rect 102095 3213 102103 6197
rect 105087 3213 105095 6197
rect 102095 3205 105095 3213
rect 105285 6197 108285 6205
rect 105285 3213 105293 6197
rect 108277 3213 108285 6197
rect 105285 3205 108285 3213
rect 108475 6197 111475 6205
rect 108475 3213 108483 6197
rect 111467 3213 111475 6197
rect 108475 3205 111475 3213
rect 111665 6197 114665 6205
rect 111665 3213 111673 6197
rect 114657 3213 114665 6197
rect 111665 3205 114665 3213
rect 114855 6197 117855 6205
rect 114855 3213 114863 6197
rect 117847 3213 117855 6197
rect 114855 3205 117855 3213
rect 118045 6197 121045 6205
rect 118045 3213 118053 6197
rect 121037 3213 121045 6197
rect 118045 3205 121045 3213
rect 121235 6197 124235 6205
rect 121235 3213 121243 6197
rect 124227 3213 124235 6197
rect 121235 3205 124235 3213
rect 124425 6197 127425 6205
rect 124425 3213 124433 6197
rect 127417 3213 127425 6197
rect 124425 3205 127425 3213
rect 127615 6197 130615 6205
rect 127615 3213 127623 6197
rect 130607 3213 130615 6197
rect 127615 3205 130615 3213
rect 130805 6197 133805 6205
rect 130805 3213 130813 6197
rect 133797 3213 133805 6197
rect 130805 3205 133805 3213
rect 133995 6197 136995 6205
rect 133995 3213 134003 6197
rect 136987 3213 136995 6197
rect 133995 3205 136995 3213
rect 15 3007 3015 3015
rect 15 23 23 3007
rect 3007 23 3015 3007
rect 15 15 3015 23
rect 3205 3007 6205 3015
rect 3205 23 3213 3007
rect 6197 23 6205 3007
rect 3205 15 6205 23
rect 6395 3007 9395 3015
rect 6395 23 6403 3007
rect 9387 23 9395 3007
rect 6395 15 9395 23
rect 9585 3007 12585 3015
rect 9585 23 9593 3007
rect 12577 23 12585 3007
rect 9585 15 12585 23
rect 12775 3007 15775 3015
rect 12775 23 12783 3007
rect 15767 23 15775 3007
rect 12775 15 15775 23
rect 15965 3007 18965 3015
rect 15965 23 15973 3007
rect 18957 23 18965 3007
rect 15965 15 18965 23
rect 19155 3007 22155 3015
rect 19155 23 19163 3007
rect 22147 23 22155 3007
rect 19155 15 22155 23
rect 22345 3007 25345 3015
rect 22345 23 22353 3007
rect 25337 23 25345 3007
rect 22345 15 25345 23
rect 25535 3007 28535 3015
rect 25535 23 25543 3007
rect 28527 23 28535 3007
rect 25535 15 28535 23
rect 28725 3007 31725 3015
rect 28725 23 28733 3007
rect 31717 23 31725 3007
rect 28725 15 31725 23
rect 31915 3007 34915 3015
rect 31915 23 31923 3007
rect 34907 23 34915 3007
rect 31915 15 34915 23
rect 35105 3007 38105 3015
rect 35105 23 35113 3007
rect 38097 23 38105 3007
rect 35105 15 38105 23
rect 38295 3007 41295 3015
rect 38295 23 38303 3007
rect 41287 23 41295 3007
rect 38295 15 41295 23
rect 41485 3007 44485 3015
rect 41485 23 41493 3007
rect 44477 23 44485 3007
rect 41485 15 44485 23
rect 44675 3007 47675 3015
rect 44675 23 44683 3007
rect 47667 23 47675 3007
rect 44675 15 47675 23
rect 47865 3007 50865 3015
rect 47865 23 47873 3007
rect 50857 23 50865 3007
rect 47865 15 50865 23
rect 51055 3007 54055 3015
rect 51055 23 51063 3007
rect 54047 23 54055 3007
rect 51055 15 54055 23
rect 54245 3007 57245 3015
rect 54245 23 54253 3007
rect 57237 23 57245 3007
rect 54245 15 57245 23
rect 57435 3007 60435 3015
rect 57435 23 57443 3007
rect 60427 23 60435 3007
rect 57435 15 60435 23
rect 60625 3007 63625 3015
rect 60625 23 60633 3007
rect 63617 23 63625 3007
rect 60625 15 63625 23
rect 63815 3007 66815 3015
rect 63815 23 63823 3007
rect 66807 23 66815 3007
rect 63815 15 66815 23
rect 67005 3007 70005 3015
rect 67005 23 67013 3007
rect 69997 23 70005 3007
rect 67005 15 70005 23
rect 70195 3007 73195 3015
rect 70195 23 70203 3007
rect 73187 23 73195 3007
rect 70195 15 73195 23
rect 73385 3007 76385 3015
rect 73385 23 73393 3007
rect 76377 23 76385 3007
rect 73385 15 76385 23
rect 76575 3007 79575 3015
rect 76575 23 76583 3007
rect 79567 23 79575 3007
rect 76575 15 79575 23
rect 79765 3007 82765 3015
rect 79765 23 79773 3007
rect 82757 23 82765 3007
rect 79765 15 82765 23
rect 82955 3007 85955 3015
rect 82955 23 82963 3007
rect 85947 23 85955 3007
rect 82955 15 85955 23
rect 86145 3007 89145 3015
rect 86145 23 86153 3007
rect 89137 23 89145 3007
rect 86145 15 89145 23
rect 89335 3007 92335 3015
rect 89335 23 89343 3007
rect 92327 23 92335 3007
rect 89335 15 92335 23
rect 92525 3007 95525 3015
rect 92525 23 92533 3007
rect 95517 23 95525 3007
rect 92525 15 95525 23
rect 95715 3007 98715 3015
rect 95715 23 95723 3007
rect 98707 23 98715 3007
rect 95715 15 98715 23
rect 98905 3007 101905 3015
rect 98905 23 98913 3007
rect 101897 23 101905 3007
rect 98905 15 101905 23
rect 102095 3007 105095 3015
rect 102095 23 102103 3007
rect 105087 23 105095 3007
rect 102095 15 105095 23
rect 105285 3007 108285 3015
rect 105285 23 105293 3007
rect 108277 23 108285 3007
rect 105285 15 108285 23
rect 108475 3007 111475 3015
rect 108475 23 108483 3007
rect 111467 23 111475 3007
rect 108475 15 111475 23
rect 111665 3007 114665 3015
rect 111665 23 111673 3007
rect 114657 23 114665 3007
rect 111665 15 114665 23
rect 114855 3007 117855 3015
rect 114855 23 114863 3007
rect 117847 23 117855 3007
rect 114855 15 117855 23
rect 118045 3007 121045 3015
rect 118045 23 118053 3007
rect 121037 23 121045 3007
rect 118045 15 121045 23
rect 121235 3007 124235 3015
rect 121235 23 121243 3007
rect 124227 23 124235 3007
rect 121235 15 124235 23
rect 124425 3007 127425 3015
rect 124425 23 124433 3007
rect 127417 23 127425 3007
rect 124425 15 127425 23
rect 127615 3007 130615 3015
rect 127615 23 127623 3007
rect 130607 23 130615 3007
rect 127615 15 130615 23
rect 130805 3007 133805 3015
rect 130805 23 130813 3007
rect 133797 23 133805 3007
rect 130805 15 133805 23
rect 133995 3007 136995 3015
rect 133995 23 134003 3007
rect 136987 23 136995 3007
rect 133995 15 136995 23
<< mimcapcontact >>
rect 23 162713 3007 165697
rect 3213 162713 6197 165697
rect 6403 162713 9387 165697
rect 9593 162713 12577 165697
rect 12783 162713 15767 165697
rect 15973 162713 18957 165697
rect 19163 162713 22147 165697
rect 22353 162713 25337 165697
rect 25543 162713 28527 165697
rect 28733 162713 31717 165697
rect 31923 162713 34907 165697
rect 35113 162713 38097 165697
rect 38303 162713 41287 165697
rect 41493 162713 44477 165697
rect 44683 162713 47667 165697
rect 47873 162713 50857 165697
rect 51063 162713 54047 165697
rect 54253 162713 57237 165697
rect 57443 162713 60427 165697
rect 60633 162713 63617 165697
rect 63823 162713 66807 165697
rect 67013 162713 69997 165697
rect 70203 162713 73187 165697
rect 73393 162713 76377 165697
rect 76583 162713 79567 165697
rect 79773 162713 82757 165697
rect 82963 162713 85947 165697
rect 86153 162713 89137 165697
rect 89343 162713 92327 165697
rect 92533 162713 95517 165697
rect 95723 162713 98707 165697
rect 98913 162713 101897 165697
rect 102103 162713 105087 165697
rect 105293 162713 108277 165697
rect 108483 162713 111467 165697
rect 111673 162713 114657 165697
rect 114863 162713 117847 165697
rect 118053 162713 121037 165697
rect 121243 162713 124227 165697
rect 124433 162713 127417 165697
rect 127623 162713 130607 165697
rect 130813 162713 133797 165697
rect 134003 162713 136987 165697
rect 23 159523 3007 162507
rect 3213 159523 6197 162507
rect 6403 159523 9387 162507
rect 9593 159523 12577 162507
rect 12783 159523 15767 162507
rect 15973 159523 18957 162507
rect 19163 159523 22147 162507
rect 22353 159523 25337 162507
rect 25543 159523 28527 162507
rect 28733 159523 31717 162507
rect 31923 159523 34907 162507
rect 35113 159523 38097 162507
rect 38303 159523 41287 162507
rect 41493 159523 44477 162507
rect 44683 159523 47667 162507
rect 47873 159523 50857 162507
rect 51063 159523 54047 162507
rect 54253 159523 57237 162507
rect 57443 159523 60427 162507
rect 60633 159523 63617 162507
rect 63823 159523 66807 162507
rect 67013 159523 69997 162507
rect 70203 159523 73187 162507
rect 73393 159523 76377 162507
rect 76583 159523 79567 162507
rect 79773 159523 82757 162507
rect 82963 159523 85947 162507
rect 86153 159523 89137 162507
rect 89343 159523 92327 162507
rect 92533 159523 95517 162507
rect 95723 159523 98707 162507
rect 98913 159523 101897 162507
rect 102103 159523 105087 162507
rect 105293 159523 108277 162507
rect 108483 159523 111467 162507
rect 111673 159523 114657 162507
rect 114863 159523 117847 162507
rect 118053 159523 121037 162507
rect 121243 159523 124227 162507
rect 124433 159523 127417 162507
rect 127623 159523 130607 162507
rect 130813 159523 133797 162507
rect 134003 159523 136987 162507
rect 23 156333 3007 159317
rect 3213 156333 6197 159317
rect 6403 156333 9387 159317
rect 9593 156333 12577 159317
rect 12783 156333 15767 159317
rect 15973 156333 18957 159317
rect 19163 156333 22147 159317
rect 22353 156333 25337 159317
rect 25543 156333 28527 159317
rect 28733 156333 31717 159317
rect 31923 156333 34907 159317
rect 35113 156333 38097 159317
rect 38303 156333 41287 159317
rect 41493 156333 44477 159317
rect 44683 156333 47667 159317
rect 47873 156333 50857 159317
rect 51063 156333 54047 159317
rect 54253 156333 57237 159317
rect 57443 156333 60427 159317
rect 60633 156333 63617 159317
rect 63823 156333 66807 159317
rect 67013 156333 69997 159317
rect 70203 156333 73187 159317
rect 73393 156333 76377 159317
rect 76583 156333 79567 159317
rect 79773 156333 82757 159317
rect 82963 156333 85947 159317
rect 86153 156333 89137 159317
rect 89343 156333 92327 159317
rect 92533 156333 95517 159317
rect 95723 156333 98707 159317
rect 98913 156333 101897 159317
rect 102103 156333 105087 159317
rect 105293 156333 108277 159317
rect 108483 156333 111467 159317
rect 111673 156333 114657 159317
rect 114863 156333 117847 159317
rect 118053 156333 121037 159317
rect 121243 156333 124227 159317
rect 124433 156333 127417 159317
rect 127623 156333 130607 159317
rect 130813 156333 133797 159317
rect 134003 156333 136987 159317
rect 23 153143 3007 156127
rect 3213 153143 6197 156127
rect 6403 153143 9387 156127
rect 9593 153143 12577 156127
rect 12783 153143 15767 156127
rect 15973 153143 18957 156127
rect 19163 153143 22147 156127
rect 22353 153143 25337 156127
rect 25543 153143 28527 156127
rect 28733 153143 31717 156127
rect 31923 153143 34907 156127
rect 35113 153143 38097 156127
rect 38303 153143 41287 156127
rect 41493 153143 44477 156127
rect 44683 153143 47667 156127
rect 47873 153143 50857 156127
rect 51063 153143 54047 156127
rect 54253 153143 57237 156127
rect 57443 153143 60427 156127
rect 60633 153143 63617 156127
rect 63823 153143 66807 156127
rect 67013 153143 69997 156127
rect 70203 153143 73187 156127
rect 73393 153143 76377 156127
rect 76583 153143 79567 156127
rect 79773 153143 82757 156127
rect 82963 153143 85947 156127
rect 86153 153143 89137 156127
rect 89343 153143 92327 156127
rect 92533 153143 95517 156127
rect 95723 153143 98707 156127
rect 98913 153143 101897 156127
rect 102103 153143 105087 156127
rect 105293 153143 108277 156127
rect 108483 153143 111467 156127
rect 111673 153143 114657 156127
rect 114863 153143 117847 156127
rect 118053 153143 121037 156127
rect 121243 153143 124227 156127
rect 124433 153143 127417 156127
rect 127623 153143 130607 156127
rect 130813 153143 133797 156127
rect 134003 153143 136987 156127
rect 23 149953 3007 152937
rect 3213 149953 6197 152937
rect 6403 149953 9387 152937
rect 9593 149953 12577 152937
rect 12783 149953 15767 152937
rect 15973 149953 18957 152937
rect 19163 149953 22147 152937
rect 22353 149953 25337 152937
rect 25543 149953 28527 152937
rect 28733 149953 31717 152937
rect 31923 149953 34907 152937
rect 35113 149953 38097 152937
rect 38303 149953 41287 152937
rect 41493 149953 44477 152937
rect 44683 149953 47667 152937
rect 47873 149953 50857 152937
rect 51063 149953 54047 152937
rect 54253 149953 57237 152937
rect 57443 149953 60427 152937
rect 60633 149953 63617 152937
rect 63823 149953 66807 152937
rect 67013 149953 69997 152937
rect 70203 149953 73187 152937
rect 73393 149953 76377 152937
rect 76583 149953 79567 152937
rect 79773 149953 82757 152937
rect 82963 149953 85947 152937
rect 86153 149953 89137 152937
rect 89343 149953 92327 152937
rect 92533 149953 95517 152937
rect 95723 149953 98707 152937
rect 98913 149953 101897 152937
rect 102103 149953 105087 152937
rect 105293 149953 108277 152937
rect 108483 149953 111467 152937
rect 111673 149953 114657 152937
rect 114863 149953 117847 152937
rect 118053 149953 121037 152937
rect 121243 149953 124227 152937
rect 124433 149953 127417 152937
rect 127623 149953 130607 152937
rect 130813 149953 133797 152937
rect 134003 149953 136987 152937
rect 23 146763 3007 149747
rect 3213 146763 6197 149747
rect 6403 146763 9387 149747
rect 9593 146763 12577 149747
rect 12783 146763 15767 149747
rect 15973 146763 18957 149747
rect 19163 146763 22147 149747
rect 22353 146763 25337 149747
rect 25543 146763 28527 149747
rect 28733 146763 31717 149747
rect 31923 146763 34907 149747
rect 35113 146763 38097 149747
rect 38303 146763 41287 149747
rect 41493 146763 44477 149747
rect 44683 146763 47667 149747
rect 47873 146763 50857 149747
rect 51063 146763 54047 149747
rect 54253 146763 57237 149747
rect 57443 146763 60427 149747
rect 60633 146763 63617 149747
rect 63823 146763 66807 149747
rect 67013 146763 69997 149747
rect 70203 146763 73187 149747
rect 73393 146763 76377 149747
rect 76583 146763 79567 149747
rect 79773 146763 82757 149747
rect 82963 146763 85947 149747
rect 86153 146763 89137 149747
rect 89343 146763 92327 149747
rect 92533 146763 95517 149747
rect 95723 146763 98707 149747
rect 98913 146763 101897 149747
rect 102103 146763 105087 149747
rect 105293 146763 108277 149747
rect 108483 146763 111467 149747
rect 111673 146763 114657 149747
rect 114863 146763 117847 149747
rect 118053 146763 121037 149747
rect 121243 146763 124227 149747
rect 124433 146763 127417 149747
rect 127623 146763 130607 149747
rect 130813 146763 133797 149747
rect 134003 146763 136987 149747
rect 23 143573 3007 146557
rect 3213 143573 6197 146557
rect 6403 143573 9387 146557
rect 9593 143573 12577 146557
rect 12783 143573 15767 146557
rect 15973 143573 18957 146557
rect 19163 143573 22147 146557
rect 22353 143573 25337 146557
rect 25543 143573 28527 146557
rect 28733 143573 31717 146557
rect 31923 143573 34907 146557
rect 35113 143573 38097 146557
rect 38303 143573 41287 146557
rect 41493 143573 44477 146557
rect 44683 143573 47667 146557
rect 47873 143573 50857 146557
rect 51063 143573 54047 146557
rect 54253 143573 57237 146557
rect 57443 143573 60427 146557
rect 60633 143573 63617 146557
rect 63823 143573 66807 146557
rect 67013 143573 69997 146557
rect 70203 143573 73187 146557
rect 73393 143573 76377 146557
rect 76583 143573 79567 146557
rect 79773 143573 82757 146557
rect 82963 143573 85947 146557
rect 86153 143573 89137 146557
rect 89343 143573 92327 146557
rect 92533 143573 95517 146557
rect 95723 143573 98707 146557
rect 98913 143573 101897 146557
rect 102103 143573 105087 146557
rect 105293 143573 108277 146557
rect 108483 143573 111467 146557
rect 111673 143573 114657 146557
rect 114863 143573 117847 146557
rect 118053 143573 121037 146557
rect 121243 143573 124227 146557
rect 124433 143573 127417 146557
rect 127623 143573 130607 146557
rect 130813 143573 133797 146557
rect 134003 143573 136987 146557
rect 23 140383 3007 143367
rect 3213 140383 6197 143367
rect 6403 140383 9387 143367
rect 9593 140383 12577 143367
rect 12783 140383 15767 143367
rect 15973 140383 18957 143367
rect 19163 140383 22147 143367
rect 22353 140383 25337 143367
rect 25543 140383 28527 143367
rect 28733 140383 31717 143367
rect 31923 140383 34907 143367
rect 35113 140383 38097 143367
rect 38303 140383 41287 143367
rect 41493 140383 44477 143367
rect 44683 140383 47667 143367
rect 47873 140383 50857 143367
rect 51063 140383 54047 143367
rect 54253 140383 57237 143367
rect 57443 140383 60427 143367
rect 60633 140383 63617 143367
rect 63823 140383 66807 143367
rect 67013 140383 69997 143367
rect 70203 140383 73187 143367
rect 73393 140383 76377 143367
rect 76583 140383 79567 143367
rect 79773 140383 82757 143367
rect 82963 140383 85947 143367
rect 86153 140383 89137 143367
rect 89343 140383 92327 143367
rect 92533 140383 95517 143367
rect 95723 140383 98707 143367
rect 98913 140383 101897 143367
rect 102103 140383 105087 143367
rect 105293 140383 108277 143367
rect 108483 140383 111467 143367
rect 111673 140383 114657 143367
rect 114863 140383 117847 143367
rect 118053 140383 121037 143367
rect 121243 140383 124227 143367
rect 124433 140383 127417 143367
rect 127623 140383 130607 143367
rect 130813 140383 133797 143367
rect 134003 140383 136987 143367
rect 9593 137193 12577 140177
rect 12783 137193 15767 140177
rect 15973 137193 18957 140177
rect 19163 137193 22147 140177
rect 22353 137193 25337 140177
rect 25543 137193 28527 140177
rect 28733 137193 31717 140177
rect 31923 137193 34907 140177
rect 35113 137193 38097 140177
rect 38303 137193 41287 140177
rect 41493 137193 44477 140177
rect 44683 137193 47667 140177
rect 47873 137193 50857 140177
rect 51063 137193 54047 140177
rect 54253 137193 57237 140177
rect 57443 137193 60427 140177
rect 60633 137193 63617 140177
rect 63823 137193 66807 140177
rect 67013 137193 69997 140177
rect 70203 137193 73187 140177
rect 73393 137193 76377 140177
rect 76583 137193 79567 140177
rect 79773 137193 82757 140177
rect 82963 137193 85947 140177
rect 86153 137193 89137 140177
rect 89343 137193 92327 140177
rect 92533 137193 95517 140177
rect 95723 137193 98707 140177
rect 98913 137193 101897 140177
rect 102103 137193 105087 140177
rect 105293 137193 108277 140177
rect 108483 137193 111467 140177
rect 111673 137193 114657 140177
rect 114863 137193 117847 140177
rect 118053 137193 121037 140177
rect 121243 137193 124227 140177
rect 124433 137193 127417 140177
rect 127623 137193 130607 140177
rect 130813 137193 133797 140177
rect 134003 137193 136987 140177
rect 9593 134003 12577 136987
rect 12783 134003 15767 136987
rect 15973 134003 18957 136987
rect 19163 134003 22147 136987
rect 22353 134003 25337 136987
rect 25543 134003 28527 136987
rect 28733 134003 31717 136987
rect 31923 134003 34907 136987
rect 35113 134003 38097 136987
rect 38303 134003 41287 136987
rect 41493 134003 44477 136987
rect 44683 134003 47667 136987
rect 47873 134003 50857 136987
rect 51063 134003 54047 136987
rect 54253 134003 57237 136987
rect 57443 134003 60427 136987
rect 60633 134003 63617 136987
rect 63823 134003 66807 136987
rect 67013 134003 69997 136987
rect 70203 134003 73187 136987
rect 73393 134003 76377 136987
rect 76583 134003 79567 136987
rect 79773 134003 82757 136987
rect 82963 134003 85947 136987
rect 86153 134003 89137 136987
rect 89343 134003 92327 136987
rect 92533 134003 95517 136987
rect 95723 134003 98707 136987
rect 98913 134003 101897 136987
rect 102103 134003 105087 136987
rect 105293 134003 108277 136987
rect 108483 134003 111467 136987
rect 111673 134003 114657 136987
rect 114863 134003 117847 136987
rect 118053 134003 121037 136987
rect 121243 134003 124227 136987
rect 124433 134003 127417 136987
rect 127623 134003 130607 136987
rect 130813 134003 133797 136987
rect 134003 134003 136987 136987
rect 9593 130813 12577 133797
rect 12783 130813 15767 133797
rect 15973 130813 18957 133797
rect 19163 130813 22147 133797
rect 22353 130813 25337 133797
rect 25543 130813 28527 133797
rect 28733 130813 31717 133797
rect 31923 130813 34907 133797
rect 35113 130813 38097 133797
rect 38303 130813 41287 133797
rect 41493 130813 44477 133797
rect 44683 130813 47667 133797
rect 47873 130813 50857 133797
rect 51063 130813 54047 133797
rect 54253 130813 57237 133797
rect 57443 130813 60427 133797
rect 60633 130813 63617 133797
rect 63823 130813 66807 133797
rect 67013 130813 69997 133797
rect 70203 130813 73187 133797
rect 73393 130813 76377 133797
rect 76583 130813 79567 133797
rect 79773 130813 82757 133797
rect 82963 130813 85947 133797
rect 86153 130813 89137 133797
rect 89343 130813 92327 133797
rect 92533 130813 95517 133797
rect 95723 130813 98707 133797
rect 98913 130813 101897 133797
rect 102103 130813 105087 133797
rect 105293 130813 108277 133797
rect 108483 130813 111467 133797
rect 111673 130813 114657 133797
rect 114863 130813 117847 133797
rect 118053 130813 121037 133797
rect 121243 130813 124227 133797
rect 124433 130813 127417 133797
rect 127623 130813 130607 133797
rect 130813 130813 133797 133797
rect 134003 130813 136987 133797
rect 9593 127623 12577 130607
rect 12783 127623 15767 130607
rect 15973 127623 18957 130607
rect 19163 127623 22147 130607
rect 22353 127623 25337 130607
rect 25543 127623 28527 130607
rect 28733 127623 31717 130607
rect 31923 127623 34907 130607
rect 35113 127623 38097 130607
rect 38303 127623 41287 130607
rect 41493 127623 44477 130607
rect 44683 127623 47667 130607
rect 47873 127623 50857 130607
rect 51063 127623 54047 130607
rect 54253 127623 57237 130607
rect 57443 127623 60427 130607
rect 60633 127623 63617 130607
rect 63823 127623 66807 130607
rect 67013 127623 69997 130607
rect 70203 127623 73187 130607
rect 73393 127623 76377 130607
rect 76583 127623 79567 130607
rect 79773 127623 82757 130607
rect 82963 127623 85947 130607
rect 86153 127623 89137 130607
rect 89343 127623 92327 130607
rect 92533 127623 95517 130607
rect 95723 127623 98707 130607
rect 98913 127623 101897 130607
rect 102103 127623 105087 130607
rect 105293 127623 108277 130607
rect 108483 127623 111467 130607
rect 111673 127623 114657 130607
rect 114863 127623 117847 130607
rect 118053 127623 121037 130607
rect 121243 127623 124227 130607
rect 124433 127623 127417 130607
rect 127623 127623 130607 130607
rect 130813 127623 133797 130607
rect 134003 127623 136987 130607
rect 9593 124433 12577 127417
rect 12783 124433 15767 127417
rect 15973 124433 18957 127417
rect 19163 124433 22147 127417
rect 22353 124433 25337 127417
rect 25543 124433 28527 127417
rect 28733 124433 31717 127417
rect 31923 124433 34907 127417
rect 35113 124433 38097 127417
rect 38303 124433 41287 127417
rect 41493 124433 44477 127417
rect 44683 124433 47667 127417
rect 47873 124433 50857 127417
rect 51063 124433 54047 127417
rect 54253 124433 57237 127417
rect 57443 124433 60427 127417
rect 60633 124433 63617 127417
rect 63823 124433 66807 127417
rect 67013 124433 69997 127417
rect 70203 124433 73187 127417
rect 73393 124433 76377 127417
rect 76583 124433 79567 127417
rect 79773 124433 82757 127417
rect 82963 124433 85947 127417
rect 86153 124433 89137 127417
rect 89343 124433 92327 127417
rect 92533 124433 95517 127417
rect 95723 124433 98707 127417
rect 98913 124433 101897 127417
rect 102103 124433 105087 127417
rect 105293 124433 108277 127417
rect 108483 124433 111467 127417
rect 111673 124433 114657 127417
rect 114863 124433 117847 127417
rect 118053 124433 121037 127417
rect 121243 124433 124227 127417
rect 124433 124433 127417 127417
rect 127623 124433 130607 127417
rect 130813 124433 133797 127417
rect 134003 124433 136987 127417
rect 9593 121243 12577 124227
rect 12783 121243 15767 124227
rect 15973 121243 18957 124227
rect 19163 121243 22147 124227
rect 22353 121243 25337 124227
rect 25543 121243 28527 124227
rect 28733 121243 31717 124227
rect 31923 121243 34907 124227
rect 35113 121243 38097 124227
rect 38303 121243 41287 124227
rect 41493 121243 44477 124227
rect 44683 121243 47667 124227
rect 47873 121243 50857 124227
rect 51063 121243 54047 124227
rect 54253 121243 57237 124227
rect 57443 121243 60427 124227
rect 60633 121243 63617 124227
rect 63823 121243 66807 124227
rect 67013 121243 69997 124227
rect 70203 121243 73187 124227
rect 73393 121243 76377 124227
rect 76583 121243 79567 124227
rect 79773 121243 82757 124227
rect 82963 121243 85947 124227
rect 86153 121243 89137 124227
rect 89343 121243 92327 124227
rect 92533 121243 95517 124227
rect 95723 121243 98707 124227
rect 98913 121243 101897 124227
rect 102103 121243 105087 124227
rect 105293 121243 108277 124227
rect 108483 121243 111467 124227
rect 111673 121243 114657 124227
rect 114863 121243 117847 124227
rect 118053 121243 121037 124227
rect 121243 121243 124227 124227
rect 124433 121243 127417 124227
rect 127623 121243 130607 124227
rect 130813 121243 133797 124227
rect 134003 121243 136987 124227
rect 23 118053 3007 121037
rect 3213 118053 6197 121037
rect 6403 118053 9387 121037
rect 9593 118053 12577 121037
rect 12783 118053 15767 121037
rect 15973 118053 18957 121037
rect 19163 118053 22147 121037
rect 22353 118053 25337 121037
rect 25543 118053 28527 121037
rect 28733 118053 31717 121037
rect 31923 118053 34907 121037
rect 35113 118053 38097 121037
rect 38303 118053 41287 121037
rect 41493 118053 44477 121037
rect 44683 118053 47667 121037
rect 47873 118053 50857 121037
rect 51063 118053 54047 121037
rect 54253 118053 57237 121037
rect 57443 118053 60427 121037
rect 60633 118053 63617 121037
rect 63823 118053 66807 121037
rect 67013 118053 69997 121037
rect 70203 118053 73187 121037
rect 73393 118053 76377 121037
rect 76583 118053 79567 121037
rect 79773 118053 82757 121037
rect 82963 118053 85947 121037
rect 86153 118053 89137 121037
rect 89343 118053 92327 121037
rect 92533 118053 95517 121037
rect 95723 118053 98707 121037
rect 98913 118053 101897 121037
rect 102103 118053 105087 121037
rect 105293 118053 108277 121037
rect 108483 118053 111467 121037
rect 111673 118053 114657 121037
rect 114863 118053 117847 121037
rect 118053 118053 121037 121037
rect 121243 118053 124227 121037
rect 124433 118053 127417 121037
rect 127623 118053 130607 121037
rect 130813 118053 133797 121037
rect 134003 118053 136987 121037
rect 23 114863 3007 117847
rect 3213 114863 6197 117847
rect 6403 114863 9387 117847
rect 9593 114863 12577 117847
rect 12783 114863 15767 117847
rect 15973 114863 18957 117847
rect 19163 114863 22147 117847
rect 22353 114863 25337 117847
rect 25543 114863 28527 117847
rect 28733 114863 31717 117847
rect 31923 114863 34907 117847
rect 35113 114863 38097 117847
rect 38303 114863 41287 117847
rect 41493 114863 44477 117847
rect 44683 114863 47667 117847
rect 47873 114863 50857 117847
rect 51063 114863 54047 117847
rect 54253 114863 57237 117847
rect 57443 114863 60427 117847
rect 60633 114863 63617 117847
rect 63823 114863 66807 117847
rect 67013 114863 69997 117847
rect 70203 114863 73187 117847
rect 73393 114863 76377 117847
rect 76583 114863 79567 117847
rect 79773 114863 82757 117847
rect 82963 114863 85947 117847
rect 86153 114863 89137 117847
rect 89343 114863 92327 117847
rect 92533 114863 95517 117847
rect 95723 114863 98707 117847
rect 98913 114863 101897 117847
rect 102103 114863 105087 117847
rect 105293 114863 108277 117847
rect 108483 114863 111467 117847
rect 111673 114863 114657 117847
rect 114863 114863 117847 117847
rect 118053 114863 121037 117847
rect 121243 114863 124227 117847
rect 124433 114863 127417 117847
rect 127623 114863 130607 117847
rect 130813 114863 133797 117847
rect 134003 114863 136987 117847
rect 23 111673 3007 114657
rect 3213 111673 6197 114657
rect 6403 111673 9387 114657
rect 9593 111673 12577 114657
rect 12783 111673 15767 114657
rect 15973 111673 18957 114657
rect 19163 111673 22147 114657
rect 22353 111673 25337 114657
rect 25543 111673 28527 114657
rect 28733 111673 31717 114657
rect 31923 111673 34907 114657
rect 35113 111673 38097 114657
rect 38303 111673 41287 114657
rect 41493 111673 44477 114657
rect 44683 111673 47667 114657
rect 47873 111673 50857 114657
rect 51063 111673 54047 114657
rect 54253 111673 57237 114657
rect 57443 111673 60427 114657
rect 60633 111673 63617 114657
rect 63823 111673 66807 114657
rect 67013 111673 69997 114657
rect 70203 111673 73187 114657
rect 73393 111673 76377 114657
rect 76583 111673 79567 114657
rect 79773 111673 82757 114657
rect 82963 111673 85947 114657
rect 86153 111673 89137 114657
rect 89343 111673 92327 114657
rect 92533 111673 95517 114657
rect 95723 111673 98707 114657
rect 98913 111673 101897 114657
rect 102103 111673 105087 114657
rect 105293 111673 108277 114657
rect 108483 111673 111467 114657
rect 111673 111673 114657 114657
rect 114863 111673 117847 114657
rect 118053 111673 121037 114657
rect 121243 111673 124227 114657
rect 124433 111673 127417 114657
rect 127623 111673 130607 114657
rect 130813 111673 133797 114657
rect 134003 111673 136987 114657
rect 23 108483 3007 111467
rect 3213 108483 6197 111467
rect 6403 108483 9387 111467
rect 9593 108483 12577 111467
rect 12783 108483 15767 111467
rect 15973 108483 18957 111467
rect 19163 108483 22147 111467
rect 22353 108483 25337 111467
rect 25543 108483 28527 111467
rect 28733 108483 31717 111467
rect 31923 108483 34907 111467
rect 35113 108483 38097 111467
rect 38303 108483 41287 111467
rect 41493 108483 44477 111467
rect 44683 108483 47667 111467
rect 47873 108483 50857 111467
rect 51063 108483 54047 111467
rect 54253 108483 57237 111467
rect 57443 108483 60427 111467
rect 60633 108483 63617 111467
rect 63823 108483 66807 111467
rect 67013 108483 69997 111467
rect 70203 108483 73187 111467
rect 73393 108483 76377 111467
rect 76583 108483 79567 111467
rect 79773 108483 82757 111467
rect 82963 108483 85947 111467
rect 86153 108483 89137 111467
rect 89343 108483 92327 111467
rect 92533 108483 95517 111467
rect 95723 108483 98707 111467
rect 98913 108483 101897 111467
rect 102103 108483 105087 111467
rect 105293 108483 108277 111467
rect 108483 108483 111467 111467
rect 111673 108483 114657 111467
rect 114863 108483 117847 111467
rect 118053 108483 121037 111467
rect 121243 108483 124227 111467
rect 124433 108483 127417 111467
rect 127623 108483 130607 111467
rect 130813 108483 133797 111467
rect 134003 108483 136987 111467
rect 23 105293 3007 108277
rect 3213 105293 6197 108277
rect 6403 105293 9387 108277
rect 9593 105293 12577 108277
rect 12783 105293 15767 108277
rect 15973 105293 18957 108277
rect 19163 105293 22147 108277
rect 22353 105293 25337 108277
rect 25543 105293 28527 108277
rect 28733 105293 31717 108277
rect 31923 105293 34907 108277
rect 35113 105293 38097 108277
rect 38303 105293 41287 108277
rect 41493 105293 44477 108277
rect 44683 105293 47667 108277
rect 47873 105293 50857 108277
rect 51063 105293 54047 108277
rect 54253 105293 57237 108277
rect 57443 105293 60427 108277
rect 60633 105293 63617 108277
rect 63823 105293 66807 108277
rect 67013 105293 69997 108277
rect 70203 105293 73187 108277
rect 73393 105293 76377 108277
rect 76583 105293 79567 108277
rect 79773 105293 82757 108277
rect 82963 105293 85947 108277
rect 86153 105293 89137 108277
rect 89343 105293 92327 108277
rect 92533 105293 95517 108277
rect 95723 105293 98707 108277
rect 98913 105293 101897 108277
rect 102103 105293 105087 108277
rect 105293 105293 108277 108277
rect 108483 105293 111467 108277
rect 111673 105293 114657 108277
rect 114863 105293 117847 108277
rect 118053 105293 121037 108277
rect 121243 105293 124227 108277
rect 124433 105293 127417 108277
rect 127623 105293 130607 108277
rect 130813 105293 133797 108277
rect 134003 105293 136987 108277
rect 23 102103 3007 105087
rect 3213 102103 6197 105087
rect 6403 102103 9387 105087
rect 9593 102103 12577 105087
rect 12783 102103 15767 105087
rect 15973 102103 18957 105087
rect 19163 102103 22147 105087
rect 22353 102103 25337 105087
rect 25543 102103 28527 105087
rect 28733 102103 31717 105087
rect 31923 102103 34907 105087
rect 35113 102103 38097 105087
rect 38303 102103 41287 105087
rect 41493 102103 44477 105087
rect 44683 102103 47667 105087
rect 47873 102103 50857 105087
rect 51063 102103 54047 105087
rect 54253 102103 57237 105087
rect 57443 102103 60427 105087
rect 60633 102103 63617 105087
rect 63823 102103 66807 105087
rect 67013 102103 69997 105087
rect 70203 102103 73187 105087
rect 73393 102103 76377 105087
rect 76583 102103 79567 105087
rect 79773 102103 82757 105087
rect 82963 102103 85947 105087
rect 86153 102103 89137 105087
rect 89343 102103 92327 105087
rect 92533 102103 95517 105087
rect 95723 102103 98707 105087
rect 98913 102103 101897 105087
rect 102103 102103 105087 105087
rect 105293 102103 108277 105087
rect 108483 102103 111467 105087
rect 111673 102103 114657 105087
rect 114863 102103 117847 105087
rect 118053 102103 121037 105087
rect 121243 102103 124227 105087
rect 124433 102103 127417 105087
rect 127623 102103 130607 105087
rect 130813 102103 133797 105087
rect 134003 102103 136987 105087
rect 23 98913 3007 101897
rect 3213 98913 6197 101897
rect 6403 98913 9387 101897
rect 9593 98913 12577 101897
rect 12783 98913 15767 101897
rect 15973 98913 18957 101897
rect 19163 98913 22147 101897
rect 22353 98913 25337 101897
rect 25543 98913 28527 101897
rect 28733 98913 31717 101897
rect 31923 98913 34907 101897
rect 35113 98913 38097 101897
rect 38303 98913 41287 101897
rect 41493 98913 44477 101897
rect 44683 98913 47667 101897
rect 47873 98913 50857 101897
rect 51063 98913 54047 101897
rect 54253 98913 57237 101897
rect 57443 98913 60427 101897
rect 60633 98913 63617 101897
rect 63823 98913 66807 101897
rect 67013 98913 69997 101897
rect 70203 98913 73187 101897
rect 73393 98913 76377 101897
rect 76583 98913 79567 101897
rect 79773 98913 82757 101897
rect 82963 98913 85947 101897
rect 86153 98913 89137 101897
rect 89343 98913 92327 101897
rect 92533 98913 95517 101897
rect 95723 98913 98707 101897
rect 98913 98913 101897 101897
rect 102103 98913 105087 101897
rect 105293 98913 108277 101897
rect 108483 98913 111467 101897
rect 111673 98913 114657 101897
rect 114863 98913 117847 101897
rect 118053 98913 121037 101897
rect 121243 98913 124227 101897
rect 124433 98913 127417 101897
rect 127623 98913 130607 101897
rect 130813 98913 133797 101897
rect 134003 98913 136987 101897
rect 9593 95723 12577 98707
rect 12783 95723 15767 98707
rect 15973 95723 18957 98707
rect 19163 95723 22147 98707
rect 22353 95723 25337 98707
rect 25543 95723 28527 98707
rect 28733 95723 31717 98707
rect 31923 95723 34907 98707
rect 35113 95723 38097 98707
rect 38303 95723 41287 98707
rect 41493 95723 44477 98707
rect 44683 95723 47667 98707
rect 47873 95723 50857 98707
rect 51063 95723 54047 98707
rect 54253 95723 57237 98707
rect 57443 95723 60427 98707
rect 60633 95723 63617 98707
rect 63823 95723 66807 98707
rect 67013 95723 69997 98707
rect 70203 95723 73187 98707
rect 73393 95723 76377 98707
rect 76583 95723 79567 98707
rect 79773 95723 82757 98707
rect 82963 95723 85947 98707
rect 86153 95723 89137 98707
rect 89343 95723 92327 98707
rect 92533 95723 95517 98707
rect 95723 95723 98707 98707
rect 98913 95723 101897 98707
rect 102103 95723 105087 98707
rect 105293 95723 108277 98707
rect 108483 95723 111467 98707
rect 111673 95723 114657 98707
rect 114863 95723 117847 98707
rect 118053 95723 121037 98707
rect 121243 95723 124227 98707
rect 124433 95723 127417 98707
rect 127623 95723 130607 98707
rect 130813 95723 133797 98707
rect 134003 95723 136987 98707
rect 9593 92533 12577 95517
rect 12783 92533 15767 95517
rect 15973 92533 18957 95517
rect 19163 92533 22147 95517
rect 22353 92533 25337 95517
rect 25543 92533 28527 95517
rect 28733 92533 31717 95517
rect 31923 92533 34907 95517
rect 35113 92533 38097 95517
rect 38303 92533 41287 95517
rect 41493 92533 44477 95517
rect 44683 92533 47667 95517
rect 47873 92533 50857 95517
rect 51063 92533 54047 95517
rect 54253 92533 57237 95517
rect 57443 92533 60427 95517
rect 60633 92533 63617 95517
rect 63823 92533 66807 95517
rect 67013 92533 69997 95517
rect 70203 92533 73187 95517
rect 73393 92533 76377 95517
rect 76583 92533 79567 95517
rect 79773 92533 82757 95517
rect 82963 92533 85947 95517
rect 86153 92533 89137 95517
rect 89343 92533 92327 95517
rect 92533 92533 95517 95517
rect 95723 92533 98707 95517
rect 98913 92533 101897 95517
rect 102103 92533 105087 95517
rect 105293 92533 108277 95517
rect 108483 92533 111467 95517
rect 111673 92533 114657 95517
rect 114863 92533 117847 95517
rect 118053 92533 121037 95517
rect 121243 92533 124227 95517
rect 124433 92533 127417 95517
rect 127623 92533 130607 95517
rect 130813 92533 133797 95517
rect 134003 92533 136987 95517
rect 9593 89343 12577 92327
rect 12783 89343 15767 92327
rect 15973 89343 18957 92327
rect 19163 89343 22147 92327
rect 22353 89343 25337 92327
rect 25543 89343 28527 92327
rect 28733 89343 31717 92327
rect 31923 89343 34907 92327
rect 35113 89343 38097 92327
rect 38303 89343 41287 92327
rect 41493 89343 44477 92327
rect 44683 89343 47667 92327
rect 47873 89343 50857 92327
rect 51063 89343 54047 92327
rect 54253 89343 57237 92327
rect 57443 89343 60427 92327
rect 60633 89343 63617 92327
rect 63823 89343 66807 92327
rect 67013 89343 69997 92327
rect 70203 89343 73187 92327
rect 73393 89343 76377 92327
rect 76583 89343 79567 92327
rect 79773 89343 82757 92327
rect 82963 89343 85947 92327
rect 86153 89343 89137 92327
rect 89343 89343 92327 92327
rect 92533 89343 95517 92327
rect 95723 89343 98707 92327
rect 98913 89343 101897 92327
rect 102103 89343 105087 92327
rect 105293 89343 108277 92327
rect 108483 89343 111467 92327
rect 111673 89343 114657 92327
rect 114863 89343 117847 92327
rect 118053 89343 121037 92327
rect 121243 89343 124227 92327
rect 124433 89343 127417 92327
rect 127623 89343 130607 92327
rect 130813 89343 133797 92327
rect 134003 89343 136987 92327
rect 9593 86153 12577 89137
rect 12783 86153 15767 89137
rect 15973 86153 18957 89137
rect 19163 86153 22147 89137
rect 22353 86153 25337 89137
rect 25543 86153 28527 89137
rect 28733 86153 31717 89137
rect 31923 86153 34907 89137
rect 35113 86153 38097 89137
rect 38303 86153 41287 89137
rect 41493 86153 44477 89137
rect 44683 86153 47667 89137
rect 47873 86153 50857 89137
rect 51063 86153 54047 89137
rect 54253 86153 57237 89137
rect 57443 86153 60427 89137
rect 60633 86153 63617 89137
rect 63823 86153 66807 89137
rect 67013 86153 69997 89137
rect 70203 86153 73187 89137
rect 73393 86153 76377 89137
rect 76583 86153 79567 89137
rect 79773 86153 82757 89137
rect 82963 86153 85947 89137
rect 86153 86153 89137 89137
rect 89343 86153 92327 89137
rect 92533 86153 95517 89137
rect 95723 86153 98707 89137
rect 98913 86153 101897 89137
rect 102103 86153 105087 89137
rect 105293 86153 108277 89137
rect 108483 86153 111467 89137
rect 111673 86153 114657 89137
rect 114863 86153 117847 89137
rect 118053 86153 121037 89137
rect 121243 86153 124227 89137
rect 124433 86153 127417 89137
rect 127623 86153 130607 89137
rect 130813 86153 133797 89137
rect 134003 86153 136987 89137
rect 9593 82963 12577 85947
rect 12783 82963 15767 85947
rect 15973 82963 18957 85947
rect 19163 82963 22147 85947
rect 22353 82963 25337 85947
rect 25543 82963 28527 85947
rect 28733 82963 31717 85947
rect 31923 82963 34907 85947
rect 35113 82963 38097 85947
rect 38303 82963 41287 85947
rect 41493 82963 44477 85947
rect 44683 82963 47667 85947
rect 47873 82963 50857 85947
rect 51063 82963 54047 85947
rect 54253 82963 57237 85947
rect 57443 82963 60427 85947
rect 60633 82963 63617 85947
rect 63823 82963 66807 85947
rect 67013 82963 69997 85947
rect 70203 82963 73187 85947
rect 73393 82963 76377 85947
rect 76583 82963 79567 85947
rect 79773 82963 82757 85947
rect 82963 82963 85947 85947
rect 86153 82963 89137 85947
rect 89343 82963 92327 85947
rect 92533 82963 95517 85947
rect 95723 82963 98707 85947
rect 98913 82963 101897 85947
rect 102103 82963 105087 85947
rect 105293 82963 108277 85947
rect 108483 82963 111467 85947
rect 111673 82963 114657 85947
rect 114863 82963 117847 85947
rect 118053 82963 121037 85947
rect 121243 82963 124227 85947
rect 124433 82963 127417 85947
rect 127623 82963 130607 85947
rect 130813 82963 133797 85947
rect 134003 82963 136987 85947
rect 9593 79773 12577 82757
rect 12783 79773 15767 82757
rect 15973 79773 18957 82757
rect 19163 79773 22147 82757
rect 22353 79773 25337 82757
rect 25543 79773 28527 82757
rect 28733 79773 31717 82757
rect 31923 79773 34907 82757
rect 35113 79773 38097 82757
rect 38303 79773 41287 82757
rect 41493 79773 44477 82757
rect 44683 79773 47667 82757
rect 47873 79773 50857 82757
rect 51063 79773 54047 82757
rect 54253 79773 57237 82757
rect 57443 79773 60427 82757
rect 60633 79773 63617 82757
rect 63823 79773 66807 82757
rect 67013 79773 69997 82757
rect 70203 79773 73187 82757
rect 73393 79773 76377 82757
rect 76583 79773 79567 82757
rect 79773 79773 82757 82757
rect 82963 79773 85947 82757
rect 86153 79773 89137 82757
rect 89343 79773 92327 82757
rect 92533 79773 95517 82757
rect 95723 79773 98707 82757
rect 98913 79773 101897 82757
rect 102103 79773 105087 82757
rect 105293 79773 108277 82757
rect 108483 79773 111467 82757
rect 111673 79773 114657 82757
rect 114863 79773 117847 82757
rect 118053 79773 121037 82757
rect 121243 79773 124227 82757
rect 124433 79773 127417 82757
rect 127623 79773 130607 82757
rect 130813 79773 133797 82757
rect 134003 79773 136987 82757
rect 23 76583 3007 79567
rect 3213 76583 6197 79567
rect 6403 76583 9387 79567
rect 9593 76583 12577 79567
rect 12783 76583 15767 79567
rect 15973 76583 18957 79567
rect 19163 76583 22147 79567
rect 22353 76583 25337 79567
rect 25543 76583 28527 79567
rect 28733 76583 31717 79567
rect 31923 76583 34907 79567
rect 35113 76583 38097 79567
rect 38303 76583 41287 79567
rect 41493 76583 44477 79567
rect 44683 76583 47667 79567
rect 47873 76583 50857 79567
rect 51063 76583 54047 79567
rect 54253 76583 57237 79567
rect 57443 76583 60427 79567
rect 60633 76583 63617 79567
rect 63823 76583 66807 79567
rect 67013 76583 69997 79567
rect 70203 76583 73187 79567
rect 73393 76583 76377 79567
rect 76583 76583 79567 79567
rect 79773 76583 82757 79567
rect 82963 76583 85947 79567
rect 86153 76583 89137 79567
rect 89343 76583 92327 79567
rect 92533 76583 95517 79567
rect 95723 76583 98707 79567
rect 98913 76583 101897 79567
rect 102103 76583 105087 79567
rect 105293 76583 108277 79567
rect 108483 76583 111467 79567
rect 111673 76583 114657 79567
rect 114863 76583 117847 79567
rect 118053 76583 121037 79567
rect 121243 76583 124227 79567
rect 124433 76583 127417 79567
rect 127623 76583 130607 79567
rect 130813 76583 133797 79567
rect 134003 76583 136987 79567
rect 23 73393 3007 76377
rect 3213 73393 6197 76377
rect 6403 73393 9387 76377
rect 9593 73393 12577 76377
rect 12783 73393 15767 76377
rect 15973 73393 18957 76377
rect 19163 73393 22147 76377
rect 22353 73393 25337 76377
rect 25543 73393 28527 76377
rect 28733 73393 31717 76377
rect 31923 73393 34907 76377
rect 35113 73393 38097 76377
rect 38303 73393 41287 76377
rect 41493 73393 44477 76377
rect 44683 73393 47667 76377
rect 47873 73393 50857 76377
rect 51063 73393 54047 76377
rect 54253 73393 57237 76377
rect 57443 73393 60427 76377
rect 60633 73393 63617 76377
rect 63823 73393 66807 76377
rect 67013 73393 69997 76377
rect 70203 73393 73187 76377
rect 73393 73393 76377 76377
rect 76583 73393 79567 76377
rect 79773 73393 82757 76377
rect 82963 73393 85947 76377
rect 86153 73393 89137 76377
rect 89343 73393 92327 76377
rect 92533 73393 95517 76377
rect 95723 73393 98707 76377
rect 98913 73393 101897 76377
rect 102103 73393 105087 76377
rect 105293 73393 108277 76377
rect 108483 73393 111467 76377
rect 111673 73393 114657 76377
rect 114863 73393 117847 76377
rect 118053 73393 121037 76377
rect 121243 73393 124227 76377
rect 124433 73393 127417 76377
rect 127623 73393 130607 76377
rect 130813 73393 133797 76377
rect 134003 73393 136987 76377
rect 23 70203 3007 73187
rect 3213 70203 6197 73187
rect 6403 70203 9387 73187
rect 9593 70203 12577 73187
rect 12783 70203 15767 73187
rect 15973 70203 18957 73187
rect 19163 70203 22147 73187
rect 22353 70203 25337 73187
rect 25543 70203 28527 73187
rect 28733 70203 31717 73187
rect 31923 70203 34907 73187
rect 35113 70203 38097 73187
rect 38303 70203 41287 73187
rect 41493 70203 44477 73187
rect 44683 70203 47667 73187
rect 47873 70203 50857 73187
rect 51063 70203 54047 73187
rect 54253 70203 57237 73187
rect 57443 70203 60427 73187
rect 60633 70203 63617 73187
rect 63823 70203 66807 73187
rect 67013 70203 69997 73187
rect 70203 70203 73187 73187
rect 73393 70203 76377 73187
rect 76583 70203 79567 73187
rect 79773 70203 82757 73187
rect 82963 70203 85947 73187
rect 86153 70203 89137 73187
rect 89343 70203 92327 73187
rect 92533 70203 95517 73187
rect 95723 70203 98707 73187
rect 98913 70203 101897 73187
rect 102103 70203 105087 73187
rect 105293 70203 108277 73187
rect 108483 70203 111467 73187
rect 111673 70203 114657 73187
rect 114863 70203 117847 73187
rect 118053 70203 121037 73187
rect 121243 70203 124227 73187
rect 124433 70203 127417 73187
rect 127623 70203 130607 73187
rect 130813 70203 133797 73187
rect 134003 70203 136987 73187
rect 23 67013 3007 69997
rect 3213 67013 6197 69997
rect 6403 67013 9387 69997
rect 9593 67013 12577 69997
rect 12783 67013 15767 69997
rect 15973 67013 18957 69997
rect 19163 67013 22147 69997
rect 22353 67013 25337 69997
rect 25543 67013 28527 69997
rect 28733 67013 31717 69997
rect 31923 67013 34907 69997
rect 35113 67013 38097 69997
rect 38303 67013 41287 69997
rect 41493 67013 44477 69997
rect 44683 67013 47667 69997
rect 47873 67013 50857 69997
rect 51063 67013 54047 69997
rect 54253 67013 57237 69997
rect 57443 67013 60427 69997
rect 60633 67013 63617 69997
rect 63823 67013 66807 69997
rect 67013 67013 69997 69997
rect 70203 67013 73187 69997
rect 73393 67013 76377 69997
rect 76583 67013 79567 69997
rect 79773 67013 82757 69997
rect 82963 67013 85947 69997
rect 86153 67013 89137 69997
rect 89343 67013 92327 69997
rect 92533 67013 95517 69997
rect 95723 67013 98707 69997
rect 98913 67013 101897 69997
rect 102103 67013 105087 69997
rect 105293 67013 108277 69997
rect 108483 67013 111467 69997
rect 111673 67013 114657 69997
rect 114863 67013 117847 69997
rect 118053 67013 121037 69997
rect 121243 67013 124227 69997
rect 124433 67013 127417 69997
rect 127623 67013 130607 69997
rect 130813 67013 133797 69997
rect 134003 67013 136987 69997
rect 23 63823 3007 66807
rect 3213 63823 6197 66807
rect 6403 63823 9387 66807
rect 9593 63823 12577 66807
rect 12783 63823 15767 66807
rect 15973 63823 18957 66807
rect 19163 63823 22147 66807
rect 22353 63823 25337 66807
rect 25543 63823 28527 66807
rect 28733 63823 31717 66807
rect 31923 63823 34907 66807
rect 35113 63823 38097 66807
rect 38303 63823 41287 66807
rect 41493 63823 44477 66807
rect 44683 63823 47667 66807
rect 47873 63823 50857 66807
rect 51063 63823 54047 66807
rect 54253 63823 57237 66807
rect 57443 63823 60427 66807
rect 60633 63823 63617 66807
rect 63823 63823 66807 66807
rect 67013 63823 69997 66807
rect 70203 63823 73187 66807
rect 73393 63823 76377 66807
rect 76583 63823 79567 66807
rect 79773 63823 82757 66807
rect 82963 63823 85947 66807
rect 86153 63823 89137 66807
rect 89343 63823 92327 66807
rect 92533 63823 95517 66807
rect 95723 63823 98707 66807
rect 98913 63823 101897 66807
rect 102103 63823 105087 66807
rect 105293 63823 108277 66807
rect 108483 63823 111467 66807
rect 111673 63823 114657 66807
rect 114863 63823 117847 66807
rect 118053 63823 121037 66807
rect 121243 63823 124227 66807
rect 124433 63823 127417 66807
rect 127623 63823 130607 66807
rect 130813 63823 133797 66807
rect 134003 63823 136987 66807
rect 23 60633 3007 63617
rect 3213 60633 6197 63617
rect 6403 60633 9387 63617
rect 9593 60633 12577 63617
rect 12783 60633 15767 63617
rect 15973 60633 18957 63617
rect 19163 60633 22147 63617
rect 22353 60633 25337 63617
rect 25543 60633 28527 63617
rect 28733 60633 31717 63617
rect 31923 60633 34907 63617
rect 35113 60633 38097 63617
rect 38303 60633 41287 63617
rect 41493 60633 44477 63617
rect 44683 60633 47667 63617
rect 47873 60633 50857 63617
rect 51063 60633 54047 63617
rect 54253 60633 57237 63617
rect 57443 60633 60427 63617
rect 60633 60633 63617 63617
rect 63823 60633 66807 63617
rect 67013 60633 69997 63617
rect 70203 60633 73187 63617
rect 73393 60633 76377 63617
rect 76583 60633 79567 63617
rect 79773 60633 82757 63617
rect 82963 60633 85947 63617
rect 86153 60633 89137 63617
rect 89343 60633 92327 63617
rect 92533 60633 95517 63617
rect 95723 60633 98707 63617
rect 98913 60633 101897 63617
rect 102103 60633 105087 63617
rect 105293 60633 108277 63617
rect 108483 60633 111467 63617
rect 111673 60633 114657 63617
rect 114863 60633 117847 63617
rect 118053 60633 121037 63617
rect 121243 60633 124227 63617
rect 124433 60633 127417 63617
rect 127623 60633 130607 63617
rect 130813 60633 133797 63617
rect 134003 60633 136987 63617
rect 23 57443 3007 60427
rect 3213 57443 6197 60427
rect 6403 57443 9387 60427
rect 9593 57443 12577 60427
rect 12783 57443 15767 60427
rect 15973 57443 18957 60427
rect 19163 57443 22147 60427
rect 22353 57443 25337 60427
rect 25543 57443 28527 60427
rect 28733 57443 31717 60427
rect 31923 57443 34907 60427
rect 35113 57443 38097 60427
rect 38303 57443 41287 60427
rect 41493 57443 44477 60427
rect 44683 57443 47667 60427
rect 47873 57443 50857 60427
rect 51063 57443 54047 60427
rect 54253 57443 57237 60427
rect 57443 57443 60427 60427
rect 60633 57443 63617 60427
rect 63823 57443 66807 60427
rect 67013 57443 69997 60427
rect 70203 57443 73187 60427
rect 73393 57443 76377 60427
rect 76583 57443 79567 60427
rect 79773 57443 82757 60427
rect 82963 57443 85947 60427
rect 86153 57443 89137 60427
rect 89343 57443 92327 60427
rect 92533 57443 95517 60427
rect 95723 57443 98707 60427
rect 98913 57443 101897 60427
rect 102103 57443 105087 60427
rect 105293 57443 108277 60427
rect 108483 57443 111467 60427
rect 111673 57443 114657 60427
rect 114863 57443 117847 60427
rect 118053 57443 121037 60427
rect 121243 57443 124227 60427
rect 124433 57443 127417 60427
rect 127623 57443 130607 60427
rect 130813 57443 133797 60427
rect 134003 57443 136987 60427
rect 23 54253 3007 57237
rect 3213 54253 6197 57237
rect 6403 54253 9387 57237
rect 9593 54253 12577 57237
rect 12783 54253 15767 57237
rect 15973 54253 18957 57237
rect 19163 54253 22147 57237
rect 22353 54253 25337 57237
rect 25543 54253 28527 57237
rect 28733 54253 31717 57237
rect 31923 54253 34907 57237
rect 35113 54253 38097 57237
rect 38303 54253 41287 57237
rect 41493 54253 44477 57237
rect 44683 54253 47667 57237
rect 47873 54253 50857 57237
rect 51063 54253 54047 57237
rect 54253 54253 57237 57237
rect 57443 54253 60427 57237
rect 60633 54253 63617 57237
rect 63823 54253 66807 57237
rect 67013 54253 69997 57237
rect 70203 54253 73187 57237
rect 73393 54253 76377 57237
rect 76583 54253 79567 57237
rect 79773 54253 82757 57237
rect 82963 54253 85947 57237
rect 86153 54253 89137 57237
rect 89343 54253 92327 57237
rect 92533 54253 95517 57237
rect 95723 54253 98707 57237
rect 98913 54253 101897 57237
rect 102103 54253 105087 57237
rect 105293 54253 108277 57237
rect 108483 54253 111467 57237
rect 111673 54253 114657 57237
rect 114863 54253 117847 57237
rect 118053 54253 121037 57237
rect 121243 54253 124227 57237
rect 124433 54253 127417 57237
rect 127623 54253 130607 57237
rect 130813 54253 133797 57237
rect 134003 54253 136987 57237
rect 23 51063 3007 54047
rect 3213 51063 6197 54047
rect 6403 51063 9387 54047
rect 9593 51063 12577 54047
rect 12783 51063 15767 54047
rect 15973 51063 18957 54047
rect 19163 51063 22147 54047
rect 22353 51063 25337 54047
rect 25543 51063 28527 54047
rect 28733 51063 31717 54047
rect 31923 51063 34907 54047
rect 35113 51063 38097 54047
rect 38303 51063 41287 54047
rect 41493 51063 44477 54047
rect 44683 51063 47667 54047
rect 47873 51063 50857 54047
rect 51063 51063 54047 54047
rect 54253 51063 57237 54047
rect 57443 51063 60427 54047
rect 60633 51063 63617 54047
rect 63823 51063 66807 54047
rect 67013 51063 69997 54047
rect 70203 51063 73187 54047
rect 73393 51063 76377 54047
rect 76583 51063 79567 54047
rect 79773 51063 82757 54047
rect 82963 51063 85947 54047
rect 86153 51063 89137 54047
rect 89343 51063 92327 54047
rect 92533 51063 95517 54047
rect 95723 51063 98707 54047
rect 98913 51063 101897 54047
rect 102103 51063 105087 54047
rect 105293 51063 108277 54047
rect 108483 51063 111467 54047
rect 111673 51063 114657 54047
rect 114863 51063 117847 54047
rect 118053 51063 121037 54047
rect 121243 51063 124227 54047
rect 124433 51063 127417 54047
rect 127623 51063 130607 54047
rect 130813 51063 133797 54047
rect 134003 51063 136987 54047
rect 23 47873 3007 50857
rect 3213 47873 6197 50857
rect 6403 47873 9387 50857
rect 9593 47873 12577 50857
rect 12783 47873 15767 50857
rect 15973 47873 18957 50857
rect 19163 47873 22147 50857
rect 22353 47873 25337 50857
rect 25543 47873 28527 50857
rect 28733 47873 31717 50857
rect 31923 47873 34907 50857
rect 35113 47873 38097 50857
rect 38303 47873 41287 50857
rect 41493 47873 44477 50857
rect 44683 47873 47667 50857
rect 47873 47873 50857 50857
rect 51063 47873 54047 50857
rect 54253 47873 57237 50857
rect 57443 47873 60427 50857
rect 60633 47873 63617 50857
rect 63823 47873 66807 50857
rect 67013 47873 69997 50857
rect 70203 47873 73187 50857
rect 73393 47873 76377 50857
rect 76583 47873 79567 50857
rect 79773 47873 82757 50857
rect 82963 47873 85947 50857
rect 86153 47873 89137 50857
rect 89343 47873 92327 50857
rect 92533 47873 95517 50857
rect 95723 47873 98707 50857
rect 98913 47873 101897 50857
rect 102103 47873 105087 50857
rect 105293 47873 108277 50857
rect 108483 47873 111467 50857
rect 111673 47873 114657 50857
rect 114863 47873 117847 50857
rect 118053 47873 121037 50857
rect 121243 47873 124227 50857
rect 124433 47873 127417 50857
rect 127623 47873 130607 50857
rect 130813 47873 133797 50857
rect 134003 47873 136987 50857
rect 23 44683 3007 47667
rect 3213 44683 6197 47667
rect 6403 44683 9387 47667
rect 9593 44683 12577 47667
rect 12783 44683 15767 47667
rect 15973 44683 18957 47667
rect 19163 44683 22147 47667
rect 22353 44683 25337 47667
rect 25543 44683 28527 47667
rect 28733 44683 31717 47667
rect 31923 44683 34907 47667
rect 35113 44683 38097 47667
rect 38303 44683 41287 47667
rect 41493 44683 44477 47667
rect 44683 44683 47667 47667
rect 47873 44683 50857 47667
rect 51063 44683 54047 47667
rect 54253 44683 57237 47667
rect 57443 44683 60427 47667
rect 60633 44683 63617 47667
rect 63823 44683 66807 47667
rect 67013 44683 69997 47667
rect 70203 44683 73187 47667
rect 73393 44683 76377 47667
rect 76583 44683 79567 47667
rect 79773 44683 82757 47667
rect 82963 44683 85947 47667
rect 86153 44683 89137 47667
rect 89343 44683 92327 47667
rect 92533 44683 95517 47667
rect 95723 44683 98707 47667
rect 98913 44683 101897 47667
rect 102103 44683 105087 47667
rect 105293 44683 108277 47667
rect 108483 44683 111467 47667
rect 111673 44683 114657 47667
rect 114863 44683 117847 47667
rect 118053 44683 121037 47667
rect 121243 44683 124227 47667
rect 124433 44683 127417 47667
rect 127623 44683 130607 47667
rect 130813 44683 133797 47667
rect 134003 44683 136987 47667
rect 23 41493 3007 44477
rect 3213 41493 6197 44477
rect 6403 41493 9387 44477
rect 9593 41493 12577 44477
rect 12783 41493 15767 44477
rect 15973 41493 18957 44477
rect 19163 41493 22147 44477
rect 22353 41493 25337 44477
rect 25543 41493 28527 44477
rect 28733 41493 31717 44477
rect 31923 41493 34907 44477
rect 35113 41493 38097 44477
rect 38303 41493 41287 44477
rect 41493 41493 44477 44477
rect 44683 41493 47667 44477
rect 47873 41493 50857 44477
rect 51063 41493 54047 44477
rect 54253 41493 57237 44477
rect 57443 41493 60427 44477
rect 60633 41493 63617 44477
rect 63823 41493 66807 44477
rect 67013 41493 69997 44477
rect 70203 41493 73187 44477
rect 73393 41493 76377 44477
rect 76583 41493 79567 44477
rect 79773 41493 82757 44477
rect 82963 41493 85947 44477
rect 86153 41493 89137 44477
rect 89343 41493 92327 44477
rect 92533 41493 95517 44477
rect 95723 41493 98707 44477
rect 98913 41493 101897 44477
rect 102103 41493 105087 44477
rect 105293 41493 108277 44477
rect 108483 41493 111467 44477
rect 111673 41493 114657 44477
rect 114863 41493 117847 44477
rect 118053 41493 121037 44477
rect 121243 41493 124227 44477
rect 124433 41493 127417 44477
rect 127623 41493 130607 44477
rect 130813 41493 133797 44477
rect 134003 41493 136987 44477
rect 23 38303 3007 41287
rect 3213 38303 6197 41287
rect 6403 38303 9387 41287
rect 9593 38303 12577 41287
rect 12783 38303 15767 41287
rect 15973 38303 18957 41287
rect 19163 38303 22147 41287
rect 22353 38303 25337 41287
rect 25543 38303 28527 41287
rect 28733 38303 31717 41287
rect 31923 38303 34907 41287
rect 35113 38303 38097 41287
rect 38303 38303 41287 41287
rect 41493 38303 44477 41287
rect 44683 38303 47667 41287
rect 47873 38303 50857 41287
rect 51063 38303 54047 41287
rect 54253 38303 57237 41287
rect 57443 38303 60427 41287
rect 60633 38303 63617 41287
rect 63823 38303 66807 41287
rect 67013 38303 69997 41287
rect 70203 38303 73187 41287
rect 73393 38303 76377 41287
rect 76583 38303 79567 41287
rect 79773 38303 82757 41287
rect 82963 38303 85947 41287
rect 86153 38303 89137 41287
rect 89343 38303 92327 41287
rect 92533 38303 95517 41287
rect 95723 38303 98707 41287
rect 98913 38303 101897 41287
rect 102103 38303 105087 41287
rect 105293 38303 108277 41287
rect 108483 38303 111467 41287
rect 111673 38303 114657 41287
rect 114863 38303 117847 41287
rect 118053 38303 121037 41287
rect 121243 38303 124227 41287
rect 124433 38303 127417 41287
rect 127623 38303 130607 41287
rect 130813 38303 133797 41287
rect 134003 38303 136987 41287
rect 23 35113 3007 38097
rect 3213 35113 6197 38097
rect 6403 35113 9387 38097
rect 9593 35113 12577 38097
rect 12783 35113 15767 38097
rect 15973 35113 18957 38097
rect 19163 35113 22147 38097
rect 22353 35113 25337 38097
rect 25543 35113 28527 38097
rect 28733 35113 31717 38097
rect 31923 35113 34907 38097
rect 35113 35113 38097 38097
rect 38303 35113 41287 38097
rect 41493 35113 44477 38097
rect 44683 35113 47667 38097
rect 47873 35113 50857 38097
rect 51063 35113 54047 38097
rect 54253 35113 57237 38097
rect 57443 35113 60427 38097
rect 60633 35113 63617 38097
rect 63823 35113 66807 38097
rect 67013 35113 69997 38097
rect 70203 35113 73187 38097
rect 73393 35113 76377 38097
rect 76583 35113 79567 38097
rect 79773 35113 82757 38097
rect 82963 35113 85947 38097
rect 86153 35113 89137 38097
rect 89343 35113 92327 38097
rect 92533 35113 95517 38097
rect 95723 35113 98707 38097
rect 98913 35113 101897 38097
rect 102103 35113 105087 38097
rect 105293 35113 108277 38097
rect 108483 35113 111467 38097
rect 111673 35113 114657 38097
rect 114863 35113 117847 38097
rect 118053 35113 121037 38097
rect 121243 35113 124227 38097
rect 124433 35113 127417 38097
rect 127623 35113 130607 38097
rect 130813 35113 133797 38097
rect 134003 35113 136987 38097
rect 23 31923 3007 34907
rect 3213 31923 6197 34907
rect 6403 31923 9387 34907
rect 9593 31923 12577 34907
rect 12783 31923 15767 34907
rect 15973 31923 18957 34907
rect 19163 31923 22147 34907
rect 22353 31923 25337 34907
rect 25543 31923 28527 34907
rect 28733 31923 31717 34907
rect 31923 31923 34907 34907
rect 35113 31923 38097 34907
rect 38303 31923 41287 34907
rect 41493 31923 44477 34907
rect 44683 31923 47667 34907
rect 47873 31923 50857 34907
rect 51063 31923 54047 34907
rect 54253 31923 57237 34907
rect 57443 31923 60427 34907
rect 60633 31923 63617 34907
rect 63823 31923 66807 34907
rect 67013 31923 69997 34907
rect 70203 31923 73187 34907
rect 73393 31923 76377 34907
rect 76583 31923 79567 34907
rect 79773 31923 82757 34907
rect 82963 31923 85947 34907
rect 86153 31923 89137 34907
rect 89343 31923 92327 34907
rect 92533 31923 95517 34907
rect 95723 31923 98707 34907
rect 98913 31923 101897 34907
rect 102103 31923 105087 34907
rect 105293 31923 108277 34907
rect 108483 31923 111467 34907
rect 111673 31923 114657 34907
rect 114863 31923 117847 34907
rect 118053 31923 121037 34907
rect 121243 31923 124227 34907
rect 124433 31923 127417 34907
rect 127623 31923 130607 34907
rect 130813 31923 133797 34907
rect 134003 31923 136987 34907
rect 23 28733 3007 31717
rect 3213 28733 6197 31717
rect 6403 28733 9387 31717
rect 9593 28733 12577 31717
rect 12783 28733 15767 31717
rect 15973 28733 18957 31717
rect 19163 28733 22147 31717
rect 22353 28733 25337 31717
rect 25543 28733 28527 31717
rect 28733 28733 31717 31717
rect 31923 28733 34907 31717
rect 35113 28733 38097 31717
rect 38303 28733 41287 31717
rect 41493 28733 44477 31717
rect 44683 28733 47667 31717
rect 47873 28733 50857 31717
rect 51063 28733 54047 31717
rect 54253 28733 57237 31717
rect 57443 28733 60427 31717
rect 60633 28733 63617 31717
rect 63823 28733 66807 31717
rect 67013 28733 69997 31717
rect 70203 28733 73187 31717
rect 73393 28733 76377 31717
rect 76583 28733 79567 31717
rect 79773 28733 82757 31717
rect 82963 28733 85947 31717
rect 86153 28733 89137 31717
rect 89343 28733 92327 31717
rect 92533 28733 95517 31717
rect 95723 28733 98707 31717
rect 98913 28733 101897 31717
rect 102103 28733 105087 31717
rect 105293 28733 108277 31717
rect 108483 28733 111467 31717
rect 111673 28733 114657 31717
rect 114863 28733 117847 31717
rect 118053 28733 121037 31717
rect 121243 28733 124227 31717
rect 124433 28733 127417 31717
rect 127623 28733 130607 31717
rect 130813 28733 133797 31717
rect 134003 28733 136987 31717
rect 23 25543 3007 28527
rect 3213 25543 6197 28527
rect 6403 25543 9387 28527
rect 9593 25543 12577 28527
rect 12783 25543 15767 28527
rect 15973 25543 18957 28527
rect 19163 25543 22147 28527
rect 22353 25543 25337 28527
rect 25543 25543 28527 28527
rect 28733 25543 31717 28527
rect 31923 25543 34907 28527
rect 35113 25543 38097 28527
rect 38303 25543 41287 28527
rect 41493 25543 44477 28527
rect 44683 25543 47667 28527
rect 47873 25543 50857 28527
rect 51063 25543 54047 28527
rect 54253 25543 57237 28527
rect 57443 25543 60427 28527
rect 60633 25543 63617 28527
rect 63823 25543 66807 28527
rect 67013 25543 69997 28527
rect 70203 25543 73187 28527
rect 73393 25543 76377 28527
rect 76583 25543 79567 28527
rect 79773 25543 82757 28527
rect 82963 25543 85947 28527
rect 86153 25543 89137 28527
rect 89343 25543 92327 28527
rect 92533 25543 95517 28527
rect 95723 25543 98707 28527
rect 98913 25543 101897 28527
rect 102103 25543 105087 28527
rect 105293 25543 108277 28527
rect 108483 25543 111467 28527
rect 111673 25543 114657 28527
rect 114863 25543 117847 28527
rect 118053 25543 121037 28527
rect 121243 25543 124227 28527
rect 124433 25543 127417 28527
rect 127623 25543 130607 28527
rect 130813 25543 133797 28527
rect 134003 25543 136987 28527
rect 23 22353 3007 25337
rect 3213 22353 6197 25337
rect 6403 22353 9387 25337
rect 9593 22353 12577 25337
rect 12783 22353 15767 25337
rect 15973 22353 18957 25337
rect 19163 22353 22147 25337
rect 22353 22353 25337 25337
rect 25543 22353 28527 25337
rect 28733 22353 31717 25337
rect 31923 22353 34907 25337
rect 35113 22353 38097 25337
rect 38303 22353 41287 25337
rect 41493 22353 44477 25337
rect 44683 22353 47667 25337
rect 47873 22353 50857 25337
rect 51063 22353 54047 25337
rect 54253 22353 57237 25337
rect 57443 22353 60427 25337
rect 60633 22353 63617 25337
rect 63823 22353 66807 25337
rect 67013 22353 69997 25337
rect 70203 22353 73187 25337
rect 73393 22353 76377 25337
rect 76583 22353 79567 25337
rect 79773 22353 82757 25337
rect 82963 22353 85947 25337
rect 86153 22353 89137 25337
rect 89343 22353 92327 25337
rect 92533 22353 95517 25337
rect 95723 22353 98707 25337
rect 98913 22353 101897 25337
rect 102103 22353 105087 25337
rect 105293 22353 108277 25337
rect 108483 22353 111467 25337
rect 111673 22353 114657 25337
rect 114863 22353 117847 25337
rect 118053 22353 121037 25337
rect 121243 22353 124227 25337
rect 124433 22353 127417 25337
rect 127623 22353 130607 25337
rect 130813 22353 133797 25337
rect 134003 22353 136987 25337
rect 23 19163 3007 22147
rect 3213 19163 6197 22147
rect 6403 19163 9387 22147
rect 9593 19163 12577 22147
rect 12783 19163 15767 22147
rect 15973 19163 18957 22147
rect 19163 19163 22147 22147
rect 22353 19163 25337 22147
rect 25543 19163 28527 22147
rect 28733 19163 31717 22147
rect 31923 19163 34907 22147
rect 35113 19163 38097 22147
rect 38303 19163 41287 22147
rect 41493 19163 44477 22147
rect 44683 19163 47667 22147
rect 47873 19163 50857 22147
rect 51063 19163 54047 22147
rect 54253 19163 57237 22147
rect 57443 19163 60427 22147
rect 60633 19163 63617 22147
rect 63823 19163 66807 22147
rect 67013 19163 69997 22147
rect 70203 19163 73187 22147
rect 73393 19163 76377 22147
rect 76583 19163 79567 22147
rect 79773 19163 82757 22147
rect 82963 19163 85947 22147
rect 86153 19163 89137 22147
rect 89343 19163 92327 22147
rect 92533 19163 95517 22147
rect 95723 19163 98707 22147
rect 98913 19163 101897 22147
rect 102103 19163 105087 22147
rect 105293 19163 108277 22147
rect 108483 19163 111467 22147
rect 111673 19163 114657 22147
rect 114863 19163 117847 22147
rect 118053 19163 121037 22147
rect 121243 19163 124227 22147
rect 124433 19163 127417 22147
rect 127623 19163 130607 22147
rect 130813 19163 133797 22147
rect 134003 19163 136987 22147
rect 23 15973 3007 18957
rect 3213 15973 6197 18957
rect 6403 15973 9387 18957
rect 9593 15973 12577 18957
rect 12783 15973 15767 18957
rect 15973 15973 18957 18957
rect 19163 15973 22147 18957
rect 22353 15973 25337 18957
rect 25543 15973 28527 18957
rect 28733 15973 31717 18957
rect 31923 15973 34907 18957
rect 35113 15973 38097 18957
rect 38303 15973 41287 18957
rect 41493 15973 44477 18957
rect 44683 15973 47667 18957
rect 47873 15973 50857 18957
rect 51063 15973 54047 18957
rect 54253 15973 57237 18957
rect 57443 15973 60427 18957
rect 60633 15973 63617 18957
rect 63823 15973 66807 18957
rect 67013 15973 69997 18957
rect 70203 15973 73187 18957
rect 73393 15973 76377 18957
rect 76583 15973 79567 18957
rect 79773 15973 82757 18957
rect 82963 15973 85947 18957
rect 86153 15973 89137 18957
rect 89343 15973 92327 18957
rect 92533 15973 95517 18957
rect 95723 15973 98707 18957
rect 98913 15973 101897 18957
rect 102103 15973 105087 18957
rect 105293 15973 108277 18957
rect 108483 15973 111467 18957
rect 111673 15973 114657 18957
rect 114863 15973 117847 18957
rect 118053 15973 121037 18957
rect 121243 15973 124227 18957
rect 124433 15973 127417 18957
rect 127623 15973 130607 18957
rect 130813 15973 133797 18957
rect 134003 15973 136987 18957
rect 23 12783 3007 15767
rect 3213 12783 6197 15767
rect 6403 12783 9387 15767
rect 9593 12783 12577 15767
rect 12783 12783 15767 15767
rect 15973 12783 18957 15767
rect 19163 12783 22147 15767
rect 22353 12783 25337 15767
rect 25543 12783 28527 15767
rect 28733 12783 31717 15767
rect 31923 12783 34907 15767
rect 35113 12783 38097 15767
rect 38303 12783 41287 15767
rect 41493 12783 44477 15767
rect 44683 12783 47667 15767
rect 47873 12783 50857 15767
rect 51063 12783 54047 15767
rect 54253 12783 57237 15767
rect 57443 12783 60427 15767
rect 60633 12783 63617 15767
rect 63823 12783 66807 15767
rect 67013 12783 69997 15767
rect 70203 12783 73187 15767
rect 73393 12783 76377 15767
rect 76583 12783 79567 15767
rect 79773 12783 82757 15767
rect 82963 12783 85947 15767
rect 86153 12783 89137 15767
rect 89343 12783 92327 15767
rect 92533 12783 95517 15767
rect 95723 12783 98707 15767
rect 98913 12783 101897 15767
rect 102103 12783 105087 15767
rect 105293 12783 108277 15767
rect 108483 12783 111467 15767
rect 111673 12783 114657 15767
rect 114863 12783 117847 15767
rect 118053 12783 121037 15767
rect 121243 12783 124227 15767
rect 124433 12783 127417 15767
rect 127623 12783 130607 15767
rect 130813 12783 133797 15767
rect 134003 12783 136987 15767
rect 23 9593 3007 12577
rect 3213 9593 6197 12577
rect 6403 9593 9387 12577
rect 9593 9593 12577 12577
rect 12783 9593 15767 12577
rect 15973 9593 18957 12577
rect 19163 9593 22147 12577
rect 22353 9593 25337 12577
rect 25543 9593 28527 12577
rect 28733 9593 31717 12577
rect 31923 9593 34907 12577
rect 35113 9593 38097 12577
rect 38303 9593 41287 12577
rect 41493 9593 44477 12577
rect 44683 9593 47667 12577
rect 47873 9593 50857 12577
rect 51063 9593 54047 12577
rect 54253 9593 57237 12577
rect 57443 9593 60427 12577
rect 60633 9593 63617 12577
rect 63823 9593 66807 12577
rect 67013 9593 69997 12577
rect 70203 9593 73187 12577
rect 73393 9593 76377 12577
rect 76583 9593 79567 12577
rect 79773 9593 82757 12577
rect 82963 9593 85947 12577
rect 86153 9593 89137 12577
rect 89343 9593 92327 12577
rect 92533 9593 95517 12577
rect 95723 9593 98707 12577
rect 98913 9593 101897 12577
rect 102103 9593 105087 12577
rect 105293 9593 108277 12577
rect 108483 9593 111467 12577
rect 111673 9593 114657 12577
rect 114863 9593 117847 12577
rect 118053 9593 121037 12577
rect 121243 9593 124227 12577
rect 124433 9593 127417 12577
rect 127623 9593 130607 12577
rect 130813 9593 133797 12577
rect 134003 9593 136987 12577
rect 23 6403 3007 9387
rect 3213 6403 6197 9387
rect 6403 6403 9387 9387
rect 9593 6403 12577 9387
rect 12783 6403 15767 9387
rect 15973 6403 18957 9387
rect 19163 6403 22147 9387
rect 22353 6403 25337 9387
rect 25543 6403 28527 9387
rect 28733 6403 31717 9387
rect 31923 6403 34907 9387
rect 35113 6403 38097 9387
rect 38303 6403 41287 9387
rect 41493 6403 44477 9387
rect 44683 6403 47667 9387
rect 47873 6403 50857 9387
rect 51063 6403 54047 9387
rect 54253 6403 57237 9387
rect 57443 6403 60427 9387
rect 60633 6403 63617 9387
rect 63823 6403 66807 9387
rect 67013 6403 69997 9387
rect 70203 6403 73187 9387
rect 73393 6403 76377 9387
rect 76583 6403 79567 9387
rect 79773 6403 82757 9387
rect 82963 6403 85947 9387
rect 86153 6403 89137 9387
rect 89343 6403 92327 9387
rect 92533 6403 95517 9387
rect 95723 6403 98707 9387
rect 98913 6403 101897 9387
rect 102103 6403 105087 9387
rect 105293 6403 108277 9387
rect 108483 6403 111467 9387
rect 111673 6403 114657 9387
rect 114863 6403 117847 9387
rect 118053 6403 121037 9387
rect 121243 6403 124227 9387
rect 124433 6403 127417 9387
rect 127623 6403 130607 9387
rect 130813 6403 133797 9387
rect 134003 6403 136987 9387
rect 23 3213 3007 6197
rect 3213 3213 6197 6197
rect 6403 3213 9387 6197
rect 9593 3213 12577 6197
rect 12783 3213 15767 6197
rect 15973 3213 18957 6197
rect 19163 3213 22147 6197
rect 22353 3213 25337 6197
rect 25543 3213 28527 6197
rect 28733 3213 31717 6197
rect 31923 3213 34907 6197
rect 35113 3213 38097 6197
rect 38303 3213 41287 6197
rect 41493 3213 44477 6197
rect 44683 3213 47667 6197
rect 47873 3213 50857 6197
rect 51063 3213 54047 6197
rect 54253 3213 57237 6197
rect 57443 3213 60427 6197
rect 60633 3213 63617 6197
rect 63823 3213 66807 6197
rect 67013 3213 69997 6197
rect 70203 3213 73187 6197
rect 73393 3213 76377 6197
rect 76583 3213 79567 6197
rect 79773 3213 82757 6197
rect 82963 3213 85947 6197
rect 86153 3213 89137 6197
rect 89343 3213 92327 6197
rect 92533 3213 95517 6197
rect 95723 3213 98707 6197
rect 98913 3213 101897 6197
rect 102103 3213 105087 6197
rect 105293 3213 108277 6197
rect 108483 3213 111467 6197
rect 111673 3213 114657 6197
rect 114863 3213 117847 6197
rect 118053 3213 121037 6197
rect 121243 3213 124227 6197
rect 124433 3213 127417 6197
rect 127623 3213 130607 6197
rect 130813 3213 133797 6197
rect 134003 3213 136987 6197
rect 23 23 3007 3007
rect 3213 23 6197 3007
rect 6403 23 9387 3007
rect 9593 23 12577 3007
rect 12783 23 15767 3007
rect 15973 23 18957 3007
rect 19163 23 22147 3007
rect 22353 23 25337 3007
rect 25543 23 28527 3007
rect 28733 23 31717 3007
rect 31923 23 34907 3007
rect 35113 23 38097 3007
rect 38303 23 41287 3007
rect 41493 23 44477 3007
rect 44683 23 47667 3007
rect 47873 23 50857 3007
rect 51063 23 54047 3007
rect 54253 23 57237 3007
rect 57443 23 60427 3007
rect 60633 23 63617 3007
rect 63823 23 66807 3007
rect 67013 23 69997 3007
rect 70203 23 73187 3007
rect 73393 23 76377 3007
rect 76583 23 79567 3007
rect 79773 23 82757 3007
rect 82963 23 85947 3007
rect 86153 23 89137 3007
rect 89343 23 92327 3007
rect 92533 23 95517 3007
rect 95723 23 98707 3007
rect 98913 23 101897 3007
rect 102103 23 105087 3007
rect 105293 23 108277 3007
rect 108483 23 111467 3007
rect 111673 23 114657 3007
rect 114863 23 117847 3007
rect 118053 23 121037 3007
rect 121243 23 124227 3007
rect 124433 23 127417 3007
rect 127623 23 130607 3007
rect 130813 23 133797 3007
rect 134003 23 136987 3007
<< metal4 >>
rect 1000 166980 68990 168000
rect 1000 166020 1020 166980
rect 68970 166020 68990 166980
rect 1000 166000 68990 166020
rect 71180 166980 135980 167000
rect 71180 166020 71200 166980
rect 135960 166020 135980 166980
rect 71180 165880 135980 166020
rect 1000 165720 2000 165880
rect 4190 165720 5190 165880
rect 7380 165720 8380 165880
rect 10570 165720 11570 165880
rect 13760 165720 14760 165880
rect 16950 165720 17950 165880
rect 20140 165720 21140 165880
rect 23330 165720 24330 165880
rect 26520 165720 27520 165880
rect 29710 165720 30710 165880
rect 32900 165720 33900 165880
rect 36090 165720 37090 165880
rect 39280 165720 40280 165880
rect 42470 165720 43470 165880
rect 45660 165720 46660 165880
rect 48850 165720 49850 165880
rect 52040 165720 53040 165880
rect 55230 165720 56230 165880
rect 58420 165720 59420 165880
rect 61610 165720 62610 165880
rect 64800 165720 65800 165880
rect 67990 165720 68990 165880
rect 71180 165720 72180 165880
rect 74370 165720 75370 165880
rect 77560 165720 78560 165880
rect 80750 165720 81750 165880
rect 83940 165720 84940 165880
rect 87130 165720 88130 165880
rect 90320 165720 91320 165880
rect 93510 165720 94510 165880
rect 96700 165720 97700 165880
rect 99890 165720 100890 165880
rect 103080 165720 104080 165880
rect 106270 165720 107270 165880
rect 109460 165720 110460 165880
rect 112650 165720 113650 165880
rect 115840 165720 116840 165880
rect 119030 165720 120030 165880
rect 122220 165720 123220 165880
rect 125410 165720 126410 165880
rect 128600 165720 129600 165880
rect 131790 165720 132790 165880
rect 134980 165720 135980 165880
rect 0 165697 3030 165720
rect 0 162713 23 165697
rect 3007 164690 3030 165697
rect 3190 165697 6220 165720
rect 3190 164690 3213 165697
rect 3007 163690 3213 164690
rect 3007 162713 3030 163690
rect 0 162690 3030 162713
rect 3190 162713 3213 163690
rect 6197 164690 6220 165697
rect 6380 165697 9410 165720
rect 6380 164690 6403 165697
rect 6197 163690 6403 164690
rect 6197 162713 6220 163690
rect 3190 162690 6220 162713
rect 6380 162713 6403 163690
rect 9387 164690 9410 165697
rect 9570 165697 12600 165720
rect 9570 164690 9593 165697
rect 9387 163690 9593 164690
rect 9387 162713 9410 163690
rect 6380 162690 9410 162713
rect 9570 162713 9593 163690
rect 12577 164690 12600 165697
rect 12760 165697 15790 165720
rect 12760 164690 12783 165697
rect 12577 163690 12783 164690
rect 12577 162713 12600 163690
rect 9570 162690 12600 162713
rect 12760 162713 12783 163690
rect 15767 164690 15790 165697
rect 15950 165697 18980 165720
rect 15950 164690 15973 165697
rect 15767 163690 15973 164690
rect 15767 162713 15790 163690
rect 12760 162690 15790 162713
rect 15950 162713 15973 163690
rect 18957 164690 18980 165697
rect 19140 165697 22170 165720
rect 19140 164690 19163 165697
rect 18957 163690 19163 164690
rect 18957 162713 18980 163690
rect 15950 162690 18980 162713
rect 19140 162713 19163 163690
rect 22147 164690 22170 165697
rect 22330 165697 25360 165720
rect 22330 164690 22353 165697
rect 22147 163690 22353 164690
rect 22147 162713 22170 163690
rect 19140 162690 22170 162713
rect 22330 162713 22353 163690
rect 25337 164690 25360 165697
rect 25520 165697 28550 165720
rect 25520 164690 25543 165697
rect 25337 163690 25543 164690
rect 25337 162713 25360 163690
rect 22330 162690 25360 162713
rect 25520 162713 25543 163690
rect 28527 164690 28550 165697
rect 28710 165697 31740 165720
rect 28710 164690 28733 165697
rect 28527 163690 28733 164690
rect 28527 162713 28550 163690
rect 25520 162690 28550 162713
rect 28710 162713 28733 163690
rect 31717 164690 31740 165697
rect 31900 165697 34930 165720
rect 31900 164690 31923 165697
rect 31717 163690 31923 164690
rect 31717 162713 31740 163690
rect 28710 162690 31740 162713
rect 31900 162713 31923 163690
rect 34907 164690 34930 165697
rect 35090 165697 38120 165720
rect 35090 164690 35113 165697
rect 34907 163690 35113 164690
rect 34907 162713 34930 163690
rect 31900 162690 34930 162713
rect 35090 162713 35113 163690
rect 38097 164690 38120 165697
rect 38280 165697 41310 165720
rect 38280 164690 38303 165697
rect 38097 163690 38303 164690
rect 38097 162713 38120 163690
rect 35090 162690 38120 162713
rect 38280 162713 38303 163690
rect 41287 164690 41310 165697
rect 41470 165697 44500 165720
rect 41470 164690 41493 165697
rect 41287 163690 41493 164690
rect 41287 162713 41310 163690
rect 38280 162690 41310 162713
rect 41470 162713 41493 163690
rect 44477 164690 44500 165697
rect 44660 165697 47690 165720
rect 44660 164690 44683 165697
rect 44477 163690 44683 164690
rect 44477 162713 44500 163690
rect 41470 162690 44500 162713
rect 44660 162713 44683 163690
rect 47667 164690 47690 165697
rect 47850 165697 50880 165720
rect 47850 164690 47873 165697
rect 47667 163690 47873 164690
rect 47667 162713 47690 163690
rect 44660 162690 47690 162713
rect 47850 162713 47873 163690
rect 50857 164690 50880 165697
rect 51040 165697 54070 165720
rect 51040 164690 51063 165697
rect 50857 163690 51063 164690
rect 50857 162713 50880 163690
rect 47850 162690 50880 162713
rect 51040 162713 51063 163690
rect 54047 164690 54070 165697
rect 54230 165697 57260 165720
rect 54230 164690 54253 165697
rect 54047 163690 54253 164690
rect 54047 162713 54070 163690
rect 51040 162690 54070 162713
rect 54230 162713 54253 163690
rect 57237 164690 57260 165697
rect 57420 165697 60450 165720
rect 57420 164690 57443 165697
rect 57237 163690 57443 164690
rect 57237 162713 57260 163690
rect 54230 162690 57260 162713
rect 57420 162713 57443 163690
rect 60427 164690 60450 165697
rect 60610 165697 63640 165720
rect 60610 164690 60633 165697
rect 60427 163690 60633 164690
rect 60427 162713 60450 163690
rect 57420 162690 60450 162713
rect 60610 162713 60633 163690
rect 63617 164690 63640 165697
rect 63800 165697 66830 165720
rect 63800 164690 63823 165697
rect 63617 163690 63823 164690
rect 63617 162713 63640 163690
rect 60610 162690 63640 162713
rect 63800 162713 63823 163690
rect 66807 164690 66830 165697
rect 66990 165697 70020 165720
rect 66990 164690 67013 165697
rect 66807 163690 67013 164690
rect 66807 162713 66830 163690
rect 63800 162690 66830 162713
rect 66990 162713 67013 163690
rect 69997 164690 70020 165697
rect 70180 165697 73210 165720
rect 70180 164690 70203 165697
rect 69997 163690 70203 164690
rect 69997 162713 70020 163690
rect 66990 162690 70020 162713
rect 70180 162713 70203 163690
rect 73187 164690 73210 165697
rect 73370 165697 76400 165720
rect 73370 164690 73393 165697
rect 73187 163690 73393 164690
rect 73187 162713 73210 163690
rect 70180 162690 73210 162713
rect 73370 162713 73393 163690
rect 76377 164690 76400 165697
rect 76560 165697 79590 165720
rect 76560 164690 76583 165697
rect 76377 163690 76583 164690
rect 76377 162713 76400 163690
rect 73370 162690 76400 162713
rect 76560 162713 76583 163690
rect 79567 164690 79590 165697
rect 79750 165697 82780 165720
rect 79750 164690 79773 165697
rect 79567 163690 79773 164690
rect 79567 162713 79590 163690
rect 76560 162690 79590 162713
rect 79750 162713 79773 163690
rect 82757 164690 82780 165697
rect 82940 165697 85970 165720
rect 82940 164690 82963 165697
rect 82757 163690 82963 164690
rect 82757 162713 82780 163690
rect 79750 162690 82780 162713
rect 82940 162713 82963 163690
rect 85947 164690 85970 165697
rect 86130 165697 89160 165720
rect 86130 164690 86153 165697
rect 85947 163690 86153 164690
rect 85947 162713 85970 163690
rect 82940 162690 85970 162713
rect 86130 162713 86153 163690
rect 89137 164690 89160 165697
rect 89320 165697 92350 165720
rect 89320 164690 89343 165697
rect 89137 163690 89343 164690
rect 89137 162713 89160 163690
rect 86130 162690 89160 162713
rect 89320 162713 89343 163690
rect 92327 164690 92350 165697
rect 92510 165697 95540 165720
rect 92510 164690 92533 165697
rect 92327 163690 92533 164690
rect 92327 162713 92350 163690
rect 89320 162690 92350 162713
rect 92510 162713 92533 163690
rect 95517 164690 95540 165697
rect 95700 165697 98730 165720
rect 95700 164690 95723 165697
rect 95517 163690 95723 164690
rect 95517 162713 95540 163690
rect 92510 162690 95540 162713
rect 95700 162713 95723 163690
rect 98707 164690 98730 165697
rect 98890 165697 101920 165720
rect 98890 164690 98913 165697
rect 98707 163690 98913 164690
rect 98707 162713 98730 163690
rect 95700 162690 98730 162713
rect 98890 162713 98913 163690
rect 101897 164690 101920 165697
rect 102080 165697 105110 165720
rect 102080 164690 102103 165697
rect 101897 163690 102103 164690
rect 101897 162713 101920 163690
rect 98890 162690 101920 162713
rect 102080 162713 102103 163690
rect 105087 164690 105110 165697
rect 105270 165697 108300 165720
rect 105270 164690 105293 165697
rect 105087 163690 105293 164690
rect 105087 162713 105110 163690
rect 102080 162690 105110 162713
rect 105270 162713 105293 163690
rect 108277 164690 108300 165697
rect 108460 165697 111490 165720
rect 108460 164690 108483 165697
rect 108277 163690 108483 164690
rect 108277 162713 108300 163690
rect 105270 162690 108300 162713
rect 108460 162713 108483 163690
rect 111467 164690 111490 165697
rect 111650 165697 114680 165720
rect 111650 164690 111673 165697
rect 111467 163690 111673 164690
rect 111467 162713 111490 163690
rect 108460 162690 111490 162713
rect 111650 162713 111673 163690
rect 114657 164690 114680 165697
rect 114840 165697 117870 165720
rect 114840 164690 114863 165697
rect 114657 163690 114863 164690
rect 114657 162713 114680 163690
rect 111650 162690 114680 162713
rect 114840 162713 114863 163690
rect 117847 164690 117870 165697
rect 118030 165697 121060 165720
rect 118030 164690 118053 165697
rect 117847 163690 118053 164690
rect 117847 162713 117870 163690
rect 114840 162690 117870 162713
rect 118030 162713 118053 163690
rect 121037 164690 121060 165697
rect 121220 165697 124250 165720
rect 121220 164690 121243 165697
rect 121037 163690 121243 164690
rect 121037 162713 121060 163690
rect 118030 162690 121060 162713
rect 121220 162713 121243 163690
rect 124227 164690 124250 165697
rect 124410 165697 127440 165720
rect 124410 164690 124433 165697
rect 124227 163690 124433 164690
rect 124227 162713 124250 163690
rect 121220 162690 124250 162713
rect 124410 162713 124433 163690
rect 127417 164690 127440 165697
rect 127600 165697 130630 165720
rect 127600 164690 127623 165697
rect 127417 163690 127623 164690
rect 127417 162713 127440 163690
rect 124410 162690 127440 162713
rect 127600 162713 127623 163690
rect 130607 164690 130630 165697
rect 130790 165697 133820 165720
rect 130790 164690 130813 165697
rect 130607 163690 130813 164690
rect 130607 162713 130630 163690
rect 127600 162690 130630 162713
rect 130790 162713 130813 163690
rect 133797 164690 133820 165697
rect 133980 165697 137010 165720
rect 133980 164690 134003 165697
rect 133797 163690 134003 164690
rect 133797 162713 133820 163690
rect 130790 162690 133820 162713
rect 133980 162713 134003 163690
rect 136987 164690 137010 165697
rect 136987 163690 137170 164690
rect 136987 162713 137010 163690
rect 133980 162690 137010 162713
rect 1000 162530 2000 162690
rect 4190 162530 5190 162690
rect 7380 162530 8380 162690
rect 10570 162530 11570 162690
rect 13760 162530 14760 162690
rect 16950 162530 17950 162690
rect 20140 162530 21140 162690
rect 23330 162530 24330 162690
rect 26520 162530 27520 162690
rect 29710 162530 30710 162690
rect 32900 162530 33900 162690
rect 36090 162530 37090 162690
rect 39280 162530 40280 162690
rect 42470 162530 43470 162690
rect 45660 162530 46660 162690
rect 48850 162530 49850 162690
rect 52040 162530 53040 162690
rect 55230 162530 56230 162690
rect 58420 162530 59420 162690
rect 61610 162530 62610 162690
rect 64800 162530 65800 162690
rect 67990 162530 68990 162690
rect 71180 162530 72180 162690
rect 74370 162530 75370 162690
rect 77560 162530 78560 162690
rect 80750 162530 81750 162690
rect 83940 162530 84940 162690
rect 87130 162530 88130 162690
rect 90320 162530 91320 162690
rect 93510 162530 94510 162690
rect 96700 162530 97700 162690
rect 99890 162530 100890 162690
rect 103080 162530 104080 162690
rect 106270 162530 107270 162690
rect 109460 162530 110460 162690
rect 112650 162530 113650 162690
rect 115840 162530 116840 162690
rect 119030 162530 120030 162690
rect 122220 162530 123220 162690
rect 125410 162530 126410 162690
rect 128600 162530 129600 162690
rect 131790 162530 132790 162690
rect 134980 162530 135980 162690
rect 0 162507 3030 162530
rect 0 159523 23 162507
rect 3007 161500 3030 162507
rect 3190 162507 6220 162530
rect 3190 161500 3213 162507
rect 3007 160500 3213 161500
rect 3007 159523 3030 160500
rect 0 159500 3030 159523
rect 3190 159523 3213 160500
rect 6197 161500 6220 162507
rect 6380 162507 9410 162530
rect 6380 161500 6403 162507
rect 6197 160500 6403 161500
rect 6197 159523 6220 160500
rect 3190 159500 6220 159523
rect 6380 159523 6403 160500
rect 9387 161500 9410 162507
rect 9570 162507 12600 162530
rect 9570 161500 9593 162507
rect 9387 160500 9593 161500
rect 9387 159523 9410 160500
rect 6380 159500 9410 159523
rect 9570 159523 9593 160500
rect 12577 161500 12600 162507
rect 12760 162507 15790 162530
rect 12760 161500 12783 162507
rect 12577 160500 12783 161500
rect 12577 159523 12600 160500
rect 9570 159500 12600 159523
rect 12760 159523 12783 160500
rect 15767 161500 15790 162507
rect 15950 162507 18980 162530
rect 15950 161500 15973 162507
rect 15767 160500 15973 161500
rect 15767 159523 15790 160500
rect 12760 159500 15790 159523
rect 15950 159523 15973 160500
rect 18957 161500 18980 162507
rect 19140 162507 22170 162530
rect 19140 161500 19163 162507
rect 18957 160500 19163 161500
rect 18957 159523 18980 160500
rect 15950 159500 18980 159523
rect 19140 159523 19163 160500
rect 22147 161500 22170 162507
rect 22330 162507 25360 162530
rect 22330 161500 22353 162507
rect 22147 160500 22353 161500
rect 22147 159523 22170 160500
rect 19140 159500 22170 159523
rect 22330 159523 22353 160500
rect 25337 161500 25360 162507
rect 25520 162507 28550 162530
rect 25520 161500 25543 162507
rect 25337 160500 25543 161500
rect 25337 159523 25360 160500
rect 22330 159500 25360 159523
rect 25520 159523 25543 160500
rect 28527 161500 28550 162507
rect 28710 162507 31740 162530
rect 28710 161500 28733 162507
rect 28527 160500 28733 161500
rect 28527 159523 28550 160500
rect 25520 159500 28550 159523
rect 28710 159523 28733 160500
rect 31717 161500 31740 162507
rect 31900 162507 34930 162530
rect 31900 161500 31923 162507
rect 31717 160500 31923 161500
rect 31717 159523 31740 160500
rect 28710 159500 31740 159523
rect 31900 159523 31923 160500
rect 34907 161500 34930 162507
rect 35090 162507 38120 162530
rect 35090 161500 35113 162507
rect 34907 160500 35113 161500
rect 34907 159523 34930 160500
rect 31900 159500 34930 159523
rect 35090 159523 35113 160500
rect 38097 161500 38120 162507
rect 38280 162507 41310 162530
rect 38280 161500 38303 162507
rect 38097 160500 38303 161500
rect 38097 159523 38120 160500
rect 35090 159500 38120 159523
rect 38280 159523 38303 160500
rect 41287 161500 41310 162507
rect 41470 162507 44500 162530
rect 41470 161500 41493 162507
rect 41287 160500 41493 161500
rect 41287 159523 41310 160500
rect 38280 159500 41310 159523
rect 41470 159523 41493 160500
rect 44477 161500 44500 162507
rect 44660 162507 47690 162530
rect 44660 161500 44683 162507
rect 44477 160500 44683 161500
rect 44477 159523 44500 160500
rect 41470 159500 44500 159523
rect 44660 159523 44683 160500
rect 47667 161500 47690 162507
rect 47850 162507 50880 162530
rect 47850 161500 47873 162507
rect 47667 160500 47873 161500
rect 47667 159523 47690 160500
rect 44660 159500 47690 159523
rect 47850 159523 47873 160500
rect 50857 161500 50880 162507
rect 51040 162507 54070 162530
rect 51040 161500 51063 162507
rect 50857 160500 51063 161500
rect 50857 159523 50880 160500
rect 47850 159500 50880 159523
rect 51040 159523 51063 160500
rect 54047 161500 54070 162507
rect 54230 162507 57260 162530
rect 54230 161500 54253 162507
rect 54047 160500 54253 161500
rect 54047 159523 54070 160500
rect 51040 159500 54070 159523
rect 54230 159523 54253 160500
rect 57237 161500 57260 162507
rect 57420 162507 60450 162530
rect 57420 161500 57443 162507
rect 57237 160500 57443 161500
rect 57237 159523 57260 160500
rect 54230 159500 57260 159523
rect 57420 159523 57443 160500
rect 60427 161500 60450 162507
rect 60610 162507 63640 162530
rect 60610 161500 60633 162507
rect 60427 160500 60633 161500
rect 60427 159523 60450 160500
rect 57420 159500 60450 159523
rect 60610 159523 60633 160500
rect 63617 161500 63640 162507
rect 63800 162507 66830 162530
rect 63800 161500 63823 162507
rect 63617 160500 63823 161500
rect 63617 159523 63640 160500
rect 60610 159500 63640 159523
rect 63800 159523 63823 160500
rect 66807 161500 66830 162507
rect 66990 162507 70020 162530
rect 66990 161500 67013 162507
rect 66807 160500 67013 161500
rect 66807 159523 66830 160500
rect 63800 159500 66830 159523
rect 66990 159523 67013 160500
rect 69997 161500 70020 162507
rect 70180 162507 73210 162530
rect 70180 161500 70203 162507
rect 69997 160500 70203 161500
rect 69997 159523 70020 160500
rect 66990 159500 70020 159523
rect 70180 159523 70203 160500
rect 73187 161500 73210 162507
rect 73370 162507 76400 162530
rect 73370 161500 73393 162507
rect 73187 160500 73393 161500
rect 73187 159523 73210 160500
rect 70180 159500 73210 159523
rect 73370 159523 73393 160500
rect 76377 161500 76400 162507
rect 76560 162507 79590 162530
rect 76560 161500 76583 162507
rect 76377 160500 76583 161500
rect 76377 159523 76400 160500
rect 73370 159500 76400 159523
rect 76560 159523 76583 160500
rect 79567 161500 79590 162507
rect 79750 162507 82780 162530
rect 79750 161500 79773 162507
rect 79567 160500 79773 161500
rect 79567 159523 79590 160500
rect 76560 159500 79590 159523
rect 79750 159523 79773 160500
rect 82757 161500 82780 162507
rect 82940 162507 85970 162530
rect 82940 161500 82963 162507
rect 82757 160500 82963 161500
rect 82757 159523 82780 160500
rect 79750 159500 82780 159523
rect 82940 159523 82963 160500
rect 85947 161500 85970 162507
rect 86130 162507 89160 162530
rect 86130 161500 86153 162507
rect 85947 160500 86153 161500
rect 85947 159523 85970 160500
rect 82940 159500 85970 159523
rect 86130 159523 86153 160500
rect 89137 161500 89160 162507
rect 89320 162507 92350 162530
rect 89320 161500 89343 162507
rect 89137 160500 89343 161500
rect 89137 159523 89160 160500
rect 86130 159500 89160 159523
rect 89320 159523 89343 160500
rect 92327 161500 92350 162507
rect 92510 162507 95540 162530
rect 92510 161500 92533 162507
rect 92327 160500 92533 161500
rect 92327 159523 92350 160500
rect 89320 159500 92350 159523
rect 92510 159523 92533 160500
rect 95517 161500 95540 162507
rect 95700 162507 98730 162530
rect 95700 161500 95723 162507
rect 95517 160500 95723 161500
rect 95517 159523 95540 160500
rect 92510 159500 95540 159523
rect 95700 159523 95723 160500
rect 98707 161500 98730 162507
rect 98890 162507 101920 162530
rect 98890 161500 98913 162507
rect 98707 160500 98913 161500
rect 98707 159523 98730 160500
rect 95700 159500 98730 159523
rect 98890 159523 98913 160500
rect 101897 161500 101920 162507
rect 102080 162507 105110 162530
rect 102080 161500 102103 162507
rect 101897 160500 102103 161500
rect 101897 159523 101920 160500
rect 98890 159500 101920 159523
rect 102080 159523 102103 160500
rect 105087 161500 105110 162507
rect 105270 162507 108300 162530
rect 105270 161500 105293 162507
rect 105087 160500 105293 161500
rect 105087 159523 105110 160500
rect 102080 159500 105110 159523
rect 105270 159523 105293 160500
rect 108277 161500 108300 162507
rect 108460 162507 111490 162530
rect 108460 161500 108483 162507
rect 108277 160500 108483 161500
rect 108277 159523 108300 160500
rect 105270 159500 108300 159523
rect 108460 159523 108483 160500
rect 111467 161500 111490 162507
rect 111650 162507 114680 162530
rect 111650 161500 111673 162507
rect 111467 160500 111673 161500
rect 111467 159523 111490 160500
rect 108460 159500 111490 159523
rect 111650 159523 111673 160500
rect 114657 161500 114680 162507
rect 114840 162507 117870 162530
rect 114840 161500 114863 162507
rect 114657 160500 114863 161500
rect 114657 159523 114680 160500
rect 111650 159500 114680 159523
rect 114840 159523 114863 160500
rect 117847 161500 117870 162507
rect 118030 162507 121060 162530
rect 118030 161500 118053 162507
rect 117847 160500 118053 161500
rect 117847 159523 117870 160500
rect 114840 159500 117870 159523
rect 118030 159523 118053 160500
rect 121037 161500 121060 162507
rect 121220 162507 124250 162530
rect 121220 161500 121243 162507
rect 121037 160500 121243 161500
rect 121037 159523 121060 160500
rect 118030 159500 121060 159523
rect 121220 159523 121243 160500
rect 124227 161500 124250 162507
rect 124410 162507 127440 162530
rect 124410 161500 124433 162507
rect 124227 160500 124433 161500
rect 124227 159523 124250 160500
rect 121220 159500 124250 159523
rect 124410 159523 124433 160500
rect 127417 161500 127440 162507
rect 127600 162507 130630 162530
rect 127600 161500 127623 162507
rect 127417 160500 127623 161500
rect 127417 159523 127440 160500
rect 124410 159500 127440 159523
rect 127600 159523 127623 160500
rect 130607 161500 130630 162507
rect 130790 162507 133820 162530
rect 130790 161500 130813 162507
rect 130607 160500 130813 161500
rect 130607 159523 130630 160500
rect 127600 159500 130630 159523
rect 130790 159523 130813 160500
rect 133797 161500 133820 162507
rect 133980 162507 137010 162530
rect 133980 161500 134003 162507
rect 133797 160500 134003 161500
rect 133797 159523 133820 160500
rect 130790 159500 133820 159523
rect 133980 159523 134003 160500
rect 136987 161500 137010 162507
rect 136987 160500 137170 161500
rect 136987 159523 137010 160500
rect 133980 159500 137010 159523
rect 1000 159340 2000 159500
rect 4190 159340 5190 159500
rect 7380 159340 8380 159500
rect 10570 159340 11570 159500
rect 13760 159340 14760 159500
rect 16950 159340 17950 159500
rect 20140 159340 21140 159500
rect 23330 159340 24330 159500
rect 26520 159340 27520 159500
rect 29710 159340 30710 159500
rect 32900 159340 33900 159500
rect 36090 159340 37090 159500
rect 39280 159340 40280 159500
rect 42470 159340 43470 159500
rect 45660 159340 46660 159500
rect 48850 159340 49850 159500
rect 52040 159340 53040 159500
rect 55230 159340 56230 159500
rect 58420 159340 59420 159500
rect 61610 159340 62610 159500
rect 64800 159340 65800 159500
rect 67990 159340 68990 159500
rect 71180 159340 72180 159500
rect 74370 159340 75370 159500
rect 77560 159340 78560 159500
rect 80750 159340 81750 159500
rect 83940 159340 84940 159500
rect 87130 159340 88130 159500
rect 90320 159340 91320 159500
rect 93510 159340 94510 159500
rect 96700 159340 97700 159500
rect 99890 159340 100890 159500
rect 103080 159340 104080 159500
rect 106270 159340 107270 159500
rect 109460 159340 110460 159500
rect 112650 159340 113650 159500
rect 115840 159340 116840 159500
rect 119030 159340 120030 159500
rect 122220 159340 123220 159500
rect 125410 159340 126410 159500
rect 128600 159340 129600 159500
rect 131790 159340 132790 159500
rect 134980 159340 135980 159500
rect 0 159317 3030 159340
rect 0 156333 23 159317
rect 3007 158310 3030 159317
rect 3190 159317 6220 159340
rect 3190 158310 3213 159317
rect 3007 157310 3213 158310
rect 3007 156333 3030 157310
rect 0 156310 3030 156333
rect 3190 156333 3213 157310
rect 6197 158310 6220 159317
rect 6380 159317 9410 159340
rect 6380 158310 6403 159317
rect 6197 157310 6403 158310
rect 6197 156333 6220 157310
rect 3190 156310 6220 156333
rect 6380 156333 6403 157310
rect 9387 158310 9410 159317
rect 9570 159317 12600 159340
rect 9570 158310 9593 159317
rect 9387 157310 9593 158310
rect 9387 156333 9410 157310
rect 6380 156310 9410 156333
rect 9570 156333 9593 157310
rect 12577 158310 12600 159317
rect 12760 159317 15790 159340
rect 12760 158310 12783 159317
rect 12577 157310 12783 158310
rect 12577 156333 12600 157310
rect 9570 156310 12600 156333
rect 12760 156333 12783 157310
rect 15767 158310 15790 159317
rect 15950 159317 18980 159340
rect 15950 158310 15973 159317
rect 15767 157310 15973 158310
rect 15767 156333 15790 157310
rect 12760 156310 15790 156333
rect 15950 156333 15973 157310
rect 18957 158310 18980 159317
rect 19140 159317 22170 159340
rect 19140 158310 19163 159317
rect 18957 157310 19163 158310
rect 18957 156333 18980 157310
rect 15950 156310 18980 156333
rect 19140 156333 19163 157310
rect 22147 158310 22170 159317
rect 22330 159317 25360 159340
rect 22330 158310 22353 159317
rect 22147 157310 22353 158310
rect 22147 156333 22170 157310
rect 19140 156310 22170 156333
rect 22330 156333 22353 157310
rect 25337 158310 25360 159317
rect 25520 159317 28550 159340
rect 25520 158310 25543 159317
rect 25337 157310 25543 158310
rect 25337 156333 25360 157310
rect 22330 156310 25360 156333
rect 25520 156333 25543 157310
rect 28527 158310 28550 159317
rect 28710 159317 31740 159340
rect 28710 158310 28733 159317
rect 28527 157310 28733 158310
rect 28527 156333 28550 157310
rect 25520 156310 28550 156333
rect 28710 156333 28733 157310
rect 31717 158310 31740 159317
rect 31900 159317 34930 159340
rect 31900 158310 31923 159317
rect 31717 157310 31923 158310
rect 31717 156333 31740 157310
rect 28710 156310 31740 156333
rect 31900 156333 31923 157310
rect 34907 158310 34930 159317
rect 35090 159317 38120 159340
rect 35090 158310 35113 159317
rect 34907 157310 35113 158310
rect 34907 156333 34930 157310
rect 31900 156310 34930 156333
rect 35090 156333 35113 157310
rect 38097 158310 38120 159317
rect 38280 159317 41310 159340
rect 38280 158310 38303 159317
rect 38097 157310 38303 158310
rect 38097 156333 38120 157310
rect 35090 156310 38120 156333
rect 38280 156333 38303 157310
rect 41287 158310 41310 159317
rect 41470 159317 44500 159340
rect 41470 158310 41493 159317
rect 41287 157310 41493 158310
rect 41287 156333 41310 157310
rect 38280 156310 41310 156333
rect 41470 156333 41493 157310
rect 44477 158310 44500 159317
rect 44660 159317 47690 159340
rect 44660 158310 44683 159317
rect 44477 157310 44683 158310
rect 44477 156333 44500 157310
rect 41470 156310 44500 156333
rect 44660 156333 44683 157310
rect 47667 158310 47690 159317
rect 47850 159317 50880 159340
rect 47850 158310 47873 159317
rect 47667 157310 47873 158310
rect 47667 156333 47690 157310
rect 44660 156310 47690 156333
rect 47850 156333 47873 157310
rect 50857 158310 50880 159317
rect 51040 159317 54070 159340
rect 51040 158310 51063 159317
rect 50857 157310 51063 158310
rect 50857 156333 50880 157310
rect 47850 156310 50880 156333
rect 51040 156333 51063 157310
rect 54047 158310 54070 159317
rect 54230 159317 57260 159340
rect 54230 158310 54253 159317
rect 54047 157310 54253 158310
rect 54047 156333 54070 157310
rect 51040 156310 54070 156333
rect 54230 156333 54253 157310
rect 57237 158310 57260 159317
rect 57420 159317 60450 159340
rect 57420 158310 57443 159317
rect 57237 157310 57443 158310
rect 57237 156333 57260 157310
rect 54230 156310 57260 156333
rect 57420 156333 57443 157310
rect 60427 158310 60450 159317
rect 60610 159317 63640 159340
rect 60610 158310 60633 159317
rect 60427 157310 60633 158310
rect 60427 156333 60450 157310
rect 57420 156310 60450 156333
rect 60610 156333 60633 157310
rect 63617 158310 63640 159317
rect 63800 159317 66830 159340
rect 63800 158310 63823 159317
rect 63617 157310 63823 158310
rect 63617 156333 63640 157310
rect 60610 156310 63640 156333
rect 63800 156333 63823 157310
rect 66807 158310 66830 159317
rect 66990 159317 70020 159340
rect 66990 158310 67013 159317
rect 66807 157310 67013 158310
rect 66807 156333 66830 157310
rect 63800 156310 66830 156333
rect 66990 156333 67013 157310
rect 69997 158310 70020 159317
rect 70180 159317 73210 159340
rect 70180 158310 70203 159317
rect 69997 157310 70203 158310
rect 69997 156333 70020 157310
rect 66990 156310 70020 156333
rect 70180 156333 70203 157310
rect 73187 158310 73210 159317
rect 73370 159317 76400 159340
rect 73370 158310 73393 159317
rect 73187 157310 73393 158310
rect 73187 156333 73210 157310
rect 70180 156310 73210 156333
rect 73370 156333 73393 157310
rect 76377 158310 76400 159317
rect 76560 159317 79590 159340
rect 76560 158310 76583 159317
rect 76377 157310 76583 158310
rect 76377 156333 76400 157310
rect 73370 156310 76400 156333
rect 76560 156333 76583 157310
rect 79567 158310 79590 159317
rect 79750 159317 82780 159340
rect 79750 158310 79773 159317
rect 79567 157310 79773 158310
rect 79567 156333 79590 157310
rect 76560 156310 79590 156333
rect 79750 156333 79773 157310
rect 82757 158310 82780 159317
rect 82940 159317 85970 159340
rect 82940 158310 82963 159317
rect 82757 157310 82963 158310
rect 82757 156333 82780 157310
rect 79750 156310 82780 156333
rect 82940 156333 82963 157310
rect 85947 158310 85970 159317
rect 86130 159317 89160 159340
rect 86130 158310 86153 159317
rect 85947 157310 86153 158310
rect 85947 156333 85970 157310
rect 82940 156310 85970 156333
rect 86130 156333 86153 157310
rect 89137 158310 89160 159317
rect 89320 159317 92350 159340
rect 89320 158310 89343 159317
rect 89137 157310 89343 158310
rect 89137 156333 89160 157310
rect 86130 156310 89160 156333
rect 89320 156333 89343 157310
rect 92327 158310 92350 159317
rect 92510 159317 95540 159340
rect 92510 158310 92533 159317
rect 92327 157310 92533 158310
rect 92327 156333 92350 157310
rect 89320 156310 92350 156333
rect 92510 156333 92533 157310
rect 95517 158310 95540 159317
rect 95700 159317 98730 159340
rect 95700 158310 95723 159317
rect 95517 157310 95723 158310
rect 95517 156333 95540 157310
rect 92510 156310 95540 156333
rect 95700 156333 95723 157310
rect 98707 158310 98730 159317
rect 98890 159317 101920 159340
rect 98890 158310 98913 159317
rect 98707 157310 98913 158310
rect 98707 156333 98730 157310
rect 95700 156310 98730 156333
rect 98890 156333 98913 157310
rect 101897 158310 101920 159317
rect 102080 159317 105110 159340
rect 102080 158310 102103 159317
rect 101897 157310 102103 158310
rect 101897 156333 101920 157310
rect 98890 156310 101920 156333
rect 102080 156333 102103 157310
rect 105087 158310 105110 159317
rect 105270 159317 108300 159340
rect 105270 158310 105293 159317
rect 105087 157310 105293 158310
rect 105087 156333 105110 157310
rect 102080 156310 105110 156333
rect 105270 156333 105293 157310
rect 108277 158310 108300 159317
rect 108460 159317 111490 159340
rect 108460 158310 108483 159317
rect 108277 157310 108483 158310
rect 108277 156333 108300 157310
rect 105270 156310 108300 156333
rect 108460 156333 108483 157310
rect 111467 158310 111490 159317
rect 111650 159317 114680 159340
rect 111650 158310 111673 159317
rect 111467 157310 111673 158310
rect 111467 156333 111490 157310
rect 108460 156310 111490 156333
rect 111650 156333 111673 157310
rect 114657 158310 114680 159317
rect 114840 159317 117870 159340
rect 114840 158310 114863 159317
rect 114657 157310 114863 158310
rect 114657 156333 114680 157310
rect 111650 156310 114680 156333
rect 114840 156333 114863 157310
rect 117847 158310 117870 159317
rect 118030 159317 121060 159340
rect 118030 158310 118053 159317
rect 117847 157310 118053 158310
rect 117847 156333 117870 157310
rect 114840 156310 117870 156333
rect 118030 156333 118053 157310
rect 121037 158310 121060 159317
rect 121220 159317 124250 159340
rect 121220 158310 121243 159317
rect 121037 157310 121243 158310
rect 121037 156333 121060 157310
rect 118030 156310 121060 156333
rect 121220 156333 121243 157310
rect 124227 158310 124250 159317
rect 124410 159317 127440 159340
rect 124410 158310 124433 159317
rect 124227 157310 124433 158310
rect 124227 156333 124250 157310
rect 121220 156310 124250 156333
rect 124410 156333 124433 157310
rect 127417 158310 127440 159317
rect 127600 159317 130630 159340
rect 127600 158310 127623 159317
rect 127417 157310 127623 158310
rect 127417 156333 127440 157310
rect 124410 156310 127440 156333
rect 127600 156333 127623 157310
rect 130607 158310 130630 159317
rect 130790 159317 133820 159340
rect 130790 158310 130813 159317
rect 130607 157310 130813 158310
rect 130607 156333 130630 157310
rect 127600 156310 130630 156333
rect 130790 156333 130813 157310
rect 133797 158310 133820 159317
rect 133980 159317 137010 159340
rect 133980 158310 134003 159317
rect 133797 157310 134003 158310
rect 133797 156333 133820 157310
rect 130790 156310 133820 156333
rect 133980 156333 134003 157310
rect 136987 158310 137010 159317
rect 136987 157310 137170 158310
rect 136987 156333 137010 157310
rect 133980 156310 137010 156333
rect 1000 156150 2000 156310
rect 4190 156150 5190 156310
rect 7380 156150 8380 156310
rect 10570 156150 11570 156310
rect 13760 156150 14760 156310
rect 16950 156150 17950 156310
rect 20140 156150 21140 156310
rect 23330 156150 24330 156310
rect 26520 156150 27520 156310
rect 29710 156150 30710 156310
rect 32900 156150 33900 156310
rect 36090 156150 37090 156310
rect 39280 156150 40280 156310
rect 42470 156150 43470 156310
rect 45660 156150 46660 156310
rect 48850 156150 49850 156310
rect 52040 156150 53040 156310
rect 55230 156150 56230 156310
rect 58420 156150 59420 156310
rect 61610 156150 62610 156310
rect 64800 156150 65800 156310
rect 67990 156150 68990 156310
rect 71180 156150 72180 156310
rect 74370 156150 75370 156310
rect 77560 156150 78560 156310
rect 80750 156150 81750 156310
rect 83940 156150 84940 156310
rect 87130 156150 88130 156310
rect 90320 156150 91320 156310
rect 93510 156150 94510 156310
rect 96700 156150 97700 156310
rect 99890 156150 100890 156310
rect 103080 156150 104080 156310
rect 106270 156150 107270 156310
rect 109460 156150 110460 156310
rect 112650 156150 113650 156310
rect 115840 156150 116840 156310
rect 119030 156150 120030 156310
rect 122220 156150 123220 156310
rect 125410 156150 126410 156310
rect 128600 156150 129600 156310
rect 131790 156150 132790 156310
rect 134980 156150 135980 156310
rect 0 156127 3030 156150
rect 0 153143 23 156127
rect 3007 155120 3030 156127
rect 3190 156127 6220 156150
rect 3190 155120 3213 156127
rect 3007 154120 3213 155120
rect 3007 153143 3030 154120
rect 0 153120 3030 153143
rect 3190 153143 3213 154120
rect 6197 155120 6220 156127
rect 6380 156127 9410 156150
rect 6380 155120 6403 156127
rect 6197 154120 6403 155120
rect 6197 153143 6220 154120
rect 3190 153120 6220 153143
rect 6380 153143 6403 154120
rect 9387 155120 9410 156127
rect 9570 156127 12600 156150
rect 9570 155120 9593 156127
rect 9387 154120 9593 155120
rect 9387 153143 9410 154120
rect 6380 153120 9410 153143
rect 9570 153143 9593 154120
rect 12577 155120 12600 156127
rect 12760 156127 15790 156150
rect 12760 155120 12783 156127
rect 12577 154120 12783 155120
rect 12577 153143 12600 154120
rect 9570 153120 12600 153143
rect 12760 153143 12783 154120
rect 15767 155120 15790 156127
rect 15950 156127 18980 156150
rect 15950 155120 15973 156127
rect 15767 154120 15973 155120
rect 15767 153143 15790 154120
rect 12760 153120 15790 153143
rect 15950 153143 15973 154120
rect 18957 155120 18980 156127
rect 19140 156127 22170 156150
rect 19140 155120 19163 156127
rect 18957 154120 19163 155120
rect 18957 153143 18980 154120
rect 15950 153120 18980 153143
rect 19140 153143 19163 154120
rect 22147 155120 22170 156127
rect 22330 156127 25360 156150
rect 22330 155120 22353 156127
rect 22147 154120 22353 155120
rect 22147 153143 22170 154120
rect 19140 153120 22170 153143
rect 22330 153143 22353 154120
rect 25337 155120 25360 156127
rect 25520 156127 28550 156150
rect 25520 155120 25543 156127
rect 25337 154120 25543 155120
rect 25337 153143 25360 154120
rect 22330 153120 25360 153143
rect 25520 153143 25543 154120
rect 28527 155120 28550 156127
rect 28710 156127 31740 156150
rect 28710 155120 28733 156127
rect 28527 154120 28733 155120
rect 28527 153143 28550 154120
rect 25520 153120 28550 153143
rect 28710 153143 28733 154120
rect 31717 155120 31740 156127
rect 31900 156127 34930 156150
rect 31900 155120 31923 156127
rect 31717 154120 31923 155120
rect 31717 153143 31740 154120
rect 28710 153120 31740 153143
rect 31900 153143 31923 154120
rect 34907 155120 34930 156127
rect 35090 156127 38120 156150
rect 35090 155120 35113 156127
rect 34907 154120 35113 155120
rect 34907 153143 34930 154120
rect 31900 153120 34930 153143
rect 35090 153143 35113 154120
rect 38097 155120 38120 156127
rect 38280 156127 41310 156150
rect 38280 155120 38303 156127
rect 38097 154120 38303 155120
rect 38097 153143 38120 154120
rect 35090 153120 38120 153143
rect 38280 153143 38303 154120
rect 41287 155120 41310 156127
rect 41470 156127 44500 156150
rect 41470 155120 41493 156127
rect 41287 154120 41493 155120
rect 41287 153143 41310 154120
rect 38280 153120 41310 153143
rect 41470 153143 41493 154120
rect 44477 155120 44500 156127
rect 44660 156127 47690 156150
rect 44660 155120 44683 156127
rect 44477 154120 44683 155120
rect 44477 153143 44500 154120
rect 41470 153120 44500 153143
rect 44660 153143 44683 154120
rect 47667 155120 47690 156127
rect 47850 156127 50880 156150
rect 47850 155120 47873 156127
rect 47667 154120 47873 155120
rect 47667 153143 47690 154120
rect 44660 153120 47690 153143
rect 47850 153143 47873 154120
rect 50857 155120 50880 156127
rect 51040 156127 54070 156150
rect 51040 155120 51063 156127
rect 50857 154120 51063 155120
rect 50857 153143 50880 154120
rect 47850 153120 50880 153143
rect 51040 153143 51063 154120
rect 54047 155120 54070 156127
rect 54230 156127 57260 156150
rect 54230 155120 54253 156127
rect 54047 154120 54253 155120
rect 54047 153143 54070 154120
rect 51040 153120 54070 153143
rect 54230 153143 54253 154120
rect 57237 155120 57260 156127
rect 57420 156127 60450 156150
rect 57420 155120 57443 156127
rect 57237 154120 57443 155120
rect 57237 153143 57260 154120
rect 54230 153120 57260 153143
rect 57420 153143 57443 154120
rect 60427 155120 60450 156127
rect 60610 156127 63640 156150
rect 60610 155120 60633 156127
rect 60427 154120 60633 155120
rect 60427 153143 60450 154120
rect 57420 153120 60450 153143
rect 60610 153143 60633 154120
rect 63617 155120 63640 156127
rect 63800 156127 66830 156150
rect 63800 155120 63823 156127
rect 63617 154120 63823 155120
rect 63617 153143 63640 154120
rect 60610 153120 63640 153143
rect 63800 153143 63823 154120
rect 66807 155120 66830 156127
rect 66990 156127 70020 156150
rect 66990 155120 67013 156127
rect 66807 154120 67013 155120
rect 66807 153143 66830 154120
rect 63800 153120 66830 153143
rect 66990 153143 67013 154120
rect 69997 155120 70020 156127
rect 70180 156127 73210 156150
rect 70180 155120 70203 156127
rect 69997 154120 70203 155120
rect 69997 153143 70020 154120
rect 66990 153120 70020 153143
rect 70180 153143 70203 154120
rect 73187 155120 73210 156127
rect 73370 156127 76400 156150
rect 73370 155120 73393 156127
rect 73187 154120 73393 155120
rect 73187 153143 73210 154120
rect 70180 153120 73210 153143
rect 73370 153143 73393 154120
rect 76377 155120 76400 156127
rect 76560 156127 79590 156150
rect 76560 155120 76583 156127
rect 76377 154120 76583 155120
rect 76377 153143 76400 154120
rect 73370 153120 76400 153143
rect 76560 153143 76583 154120
rect 79567 155120 79590 156127
rect 79750 156127 82780 156150
rect 79750 155120 79773 156127
rect 79567 154120 79773 155120
rect 79567 153143 79590 154120
rect 76560 153120 79590 153143
rect 79750 153143 79773 154120
rect 82757 155120 82780 156127
rect 82940 156127 85970 156150
rect 82940 155120 82963 156127
rect 82757 154120 82963 155120
rect 82757 153143 82780 154120
rect 79750 153120 82780 153143
rect 82940 153143 82963 154120
rect 85947 155120 85970 156127
rect 86130 156127 89160 156150
rect 86130 155120 86153 156127
rect 85947 154120 86153 155120
rect 85947 153143 85970 154120
rect 82940 153120 85970 153143
rect 86130 153143 86153 154120
rect 89137 155120 89160 156127
rect 89320 156127 92350 156150
rect 89320 155120 89343 156127
rect 89137 154120 89343 155120
rect 89137 153143 89160 154120
rect 86130 153120 89160 153143
rect 89320 153143 89343 154120
rect 92327 155120 92350 156127
rect 92510 156127 95540 156150
rect 92510 155120 92533 156127
rect 92327 154120 92533 155120
rect 92327 153143 92350 154120
rect 89320 153120 92350 153143
rect 92510 153143 92533 154120
rect 95517 155120 95540 156127
rect 95700 156127 98730 156150
rect 95700 155120 95723 156127
rect 95517 154120 95723 155120
rect 95517 153143 95540 154120
rect 92510 153120 95540 153143
rect 95700 153143 95723 154120
rect 98707 155120 98730 156127
rect 98890 156127 101920 156150
rect 98890 155120 98913 156127
rect 98707 154120 98913 155120
rect 98707 153143 98730 154120
rect 95700 153120 98730 153143
rect 98890 153143 98913 154120
rect 101897 155120 101920 156127
rect 102080 156127 105110 156150
rect 102080 155120 102103 156127
rect 101897 154120 102103 155120
rect 101897 153143 101920 154120
rect 98890 153120 101920 153143
rect 102080 153143 102103 154120
rect 105087 155120 105110 156127
rect 105270 156127 108300 156150
rect 105270 155120 105293 156127
rect 105087 154120 105293 155120
rect 105087 153143 105110 154120
rect 102080 153120 105110 153143
rect 105270 153143 105293 154120
rect 108277 155120 108300 156127
rect 108460 156127 111490 156150
rect 108460 155120 108483 156127
rect 108277 154120 108483 155120
rect 108277 153143 108300 154120
rect 105270 153120 108300 153143
rect 108460 153143 108483 154120
rect 111467 155120 111490 156127
rect 111650 156127 114680 156150
rect 111650 155120 111673 156127
rect 111467 154120 111673 155120
rect 111467 153143 111490 154120
rect 108460 153120 111490 153143
rect 111650 153143 111673 154120
rect 114657 155120 114680 156127
rect 114840 156127 117870 156150
rect 114840 155120 114863 156127
rect 114657 154120 114863 155120
rect 114657 153143 114680 154120
rect 111650 153120 114680 153143
rect 114840 153143 114863 154120
rect 117847 155120 117870 156127
rect 118030 156127 121060 156150
rect 118030 155120 118053 156127
rect 117847 154120 118053 155120
rect 117847 153143 117870 154120
rect 114840 153120 117870 153143
rect 118030 153143 118053 154120
rect 121037 155120 121060 156127
rect 121220 156127 124250 156150
rect 121220 155120 121243 156127
rect 121037 154120 121243 155120
rect 121037 153143 121060 154120
rect 118030 153120 121060 153143
rect 121220 153143 121243 154120
rect 124227 155120 124250 156127
rect 124410 156127 127440 156150
rect 124410 155120 124433 156127
rect 124227 154120 124433 155120
rect 124227 153143 124250 154120
rect 121220 153120 124250 153143
rect 124410 153143 124433 154120
rect 127417 155120 127440 156127
rect 127600 156127 130630 156150
rect 127600 155120 127623 156127
rect 127417 154120 127623 155120
rect 127417 153143 127440 154120
rect 124410 153120 127440 153143
rect 127600 153143 127623 154120
rect 130607 155120 130630 156127
rect 130790 156127 133820 156150
rect 130790 155120 130813 156127
rect 130607 154120 130813 155120
rect 130607 153143 130630 154120
rect 127600 153120 130630 153143
rect 130790 153143 130813 154120
rect 133797 155120 133820 156127
rect 133980 156127 137010 156150
rect 133980 155120 134003 156127
rect 133797 154120 134003 155120
rect 133797 153143 133820 154120
rect 130790 153120 133820 153143
rect 133980 153143 134003 154120
rect 136987 155120 137010 156127
rect 136987 154120 137170 155120
rect 136987 153143 137010 154120
rect 133980 153120 137010 153143
rect 1000 152960 2000 153120
rect 4190 152960 5190 153120
rect 7380 152960 8380 153120
rect 10570 152960 11570 153120
rect 13760 152960 14760 153120
rect 16950 152960 17950 153120
rect 20140 152960 21140 153120
rect 23330 152960 24330 153120
rect 26520 152960 27520 153120
rect 29710 152960 30710 153120
rect 32900 152960 33900 153120
rect 36090 152960 37090 153120
rect 39280 152960 40280 153120
rect 42470 152960 43470 153120
rect 45660 152960 46660 153120
rect 48850 152960 49850 153120
rect 52040 152960 53040 153120
rect 55230 152960 56230 153120
rect 58420 152960 59420 153120
rect 61610 152960 62610 153120
rect 64800 152960 65800 153120
rect 67990 152960 68990 153120
rect 71180 152960 72180 153120
rect 74370 152960 75370 153120
rect 77560 152960 78560 153120
rect 80750 152960 81750 153120
rect 83940 152960 84940 153120
rect 87130 152960 88130 153120
rect 90320 152960 91320 153120
rect 93510 152960 94510 153120
rect 96700 152960 97700 153120
rect 99890 152960 100890 153120
rect 103080 152960 104080 153120
rect 106270 152960 107270 153120
rect 109460 152960 110460 153120
rect 112650 152960 113650 153120
rect 115840 152960 116840 153120
rect 119030 152960 120030 153120
rect 122220 152960 123220 153120
rect 125410 152960 126410 153120
rect 128600 152960 129600 153120
rect 131790 152960 132790 153120
rect 134980 152960 135980 153120
rect 0 152937 3030 152960
rect 0 149953 23 152937
rect 3007 151930 3030 152937
rect 3190 152937 6220 152960
rect 3190 151930 3213 152937
rect 3007 150930 3213 151930
rect 3007 149953 3030 150930
rect 0 149930 3030 149953
rect 3190 149953 3213 150930
rect 6197 151930 6220 152937
rect 6380 152937 9410 152960
rect 6380 151930 6403 152937
rect 6197 150930 6403 151930
rect 6197 149953 6220 150930
rect 3190 149930 6220 149953
rect 6380 149953 6403 150930
rect 9387 151930 9410 152937
rect 9570 152937 12600 152960
rect 9570 151930 9593 152937
rect 9387 150930 9593 151930
rect 9387 149953 9410 150930
rect 6380 149930 9410 149953
rect 9570 149953 9593 150930
rect 12577 151930 12600 152937
rect 12760 152937 15790 152960
rect 12760 151930 12783 152937
rect 12577 150930 12783 151930
rect 12577 149953 12600 150930
rect 9570 149930 12600 149953
rect 12760 149953 12783 150930
rect 15767 151930 15790 152937
rect 15950 152937 18980 152960
rect 15950 151930 15973 152937
rect 15767 150930 15973 151930
rect 15767 149953 15790 150930
rect 12760 149930 15790 149953
rect 15950 149953 15973 150930
rect 18957 151930 18980 152937
rect 19140 152937 22170 152960
rect 19140 151930 19163 152937
rect 18957 150930 19163 151930
rect 18957 149953 18980 150930
rect 15950 149930 18980 149953
rect 19140 149953 19163 150930
rect 22147 151930 22170 152937
rect 22330 152937 25360 152960
rect 22330 151930 22353 152937
rect 22147 150930 22353 151930
rect 22147 149953 22170 150930
rect 19140 149930 22170 149953
rect 22330 149953 22353 150930
rect 25337 151930 25360 152937
rect 25520 152937 28550 152960
rect 25520 151930 25543 152937
rect 25337 150930 25543 151930
rect 25337 149953 25360 150930
rect 22330 149930 25360 149953
rect 25520 149953 25543 150930
rect 28527 151930 28550 152937
rect 28710 152937 31740 152960
rect 28710 151930 28733 152937
rect 28527 150930 28733 151930
rect 28527 149953 28550 150930
rect 25520 149930 28550 149953
rect 28710 149953 28733 150930
rect 31717 151930 31740 152937
rect 31900 152937 34930 152960
rect 31900 151930 31923 152937
rect 31717 150930 31923 151930
rect 31717 149953 31740 150930
rect 28710 149930 31740 149953
rect 31900 149953 31923 150930
rect 34907 151930 34930 152937
rect 35090 152937 38120 152960
rect 35090 151930 35113 152937
rect 34907 150930 35113 151930
rect 34907 149953 34930 150930
rect 31900 149930 34930 149953
rect 35090 149953 35113 150930
rect 38097 151930 38120 152937
rect 38280 152937 41310 152960
rect 38280 151930 38303 152937
rect 38097 150930 38303 151930
rect 38097 149953 38120 150930
rect 35090 149930 38120 149953
rect 38280 149953 38303 150930
rect 41287 151930 41310 152937
rect 41470 152937 44500 152960
rect 41470 151930 41493 152937
rect 41287 150930 41493 151930
rect 41287 149953 41310 150930
rect 38280 149930 41310 149953
rect 41470 149953 41493 150930
rect 44477 151930 44500 152937
rect 44660 152937 47690 152960
rect 44660 151930 44683 152937
rect 44477 150930 44683 151930
rect 44477 149953 44500 150930
rect 41470 149930 44500 149953
rect 44660 149953 44683 150930
rect 47667 151930 47690 152937
rect 47850 152937 50880 152960
rect 47850 151930 47873 152937
rect 47667 150930 47873 151930
rect 47667 149953 47690 150930
rect 44660 149930 47690 149953
rect 47850 149953 47873 150930
rect 50857 151930 50880 152937
rect 51040 152937 54070 152960
rect 51040 151930 51063 152937
rect 50857 150930 51063 151930
rect 50857 149953 50880 150930
rect 47850 149930 50880 149953
rect 51040 149953 51063 150930
rect 54047 151930 54070 152937
rect 54230 152937 57260 152960
rect 54230 151930 54253 152937
rect 54047 150930 54253 151930
rect 54047 149953 54070 150930
rect 51040 149930 54070 149953
rect 54230 149953 54253 150930
rect 57237 151930 57260 152937
rect 57420 152937 60450 152960
rect 57420 151930 57443 152937
rect 57237 150930 57443 151930
rect 57237 149953 57260 150930
rect 54230 149930 57260 149953
rect 57420 149953 57443 150930
rect 60427 151930 60450 152937
rect 60610 152937 63640 152960
rect 60610 151930 60633 152937
rect 60427 150930 60633 151930
rect 60427 149953 60450 150930
rect 57420 149930 60450 149953
rect 60610 149953 60633 150930
rect 63617 151930 63640 152937
rect 63800 152937 66830 152960
rect 63800 151930 63823 152937
rect 63617 150930 63823 151930
rect 63617 149953 63640 150930
rect 60610 149930 63640 149953
rect 63800 149953 63823 150930
rect 66807 151930 66830 152937
rect 66990 152937 70020 152960
rect 66990 151930 67013 152937
rect 66807 150930 67013 151930
rect 66807 149953 66830 150930
rect 63800 149930 66830 149953
rect 66990 149953 67013 150930
rect 69997 151930 70020 152937
rect 70180 152937 73210 152960
rect 70180 151930 70203 152937
rect 69997 150930 70203 151930
rect 69997 149953 70020 150930
rect 66990 149930 70020 149953
rect 70180 149953 70203 150930
rect 73187 151930 73210 152937
rect 73370 152937 76400 152960
rect 73370 151930 73393 152937
rect 73187 150930 73393 151930
rect 73187 149953 73210 150930
rect 70180 149930 73210 149953
rect 73370 149953 73393 150930
rect 76377 151930 76400 152937
rect 76560 152937 79590 152960
rect 76560 151930 76583 152937
rect 76377 150930 76583 151930
rect 76377 149953 76400 150930
rect 73370 149930 76400 149953
rect 76560 149953 76583 150930
rect 79567 151930 79590 152937
rect 79750 152937 82780 152960
rect 79750 151930 79773 152937
rect 79567 150930 79773 151930
rect 79567 149953 79590 150930
rect 76560 149930 79590 149953
rect 79750 149953 79773 150930
rect 82757 151930 82780 152937
rect 82940 152937 85970 152960
rect 82940 151930 82963 152937
rect 82757 150930 82963 151930
rect 82757 149953 82780 150930
rect 79750 149930 82780 149953
rect 82940 149953 82963 150930
rect 85947 151930 85970 152937
rect 86130 152937 89160 152960
rect 86130 151930 86153 152937
rect 85947 150930 86153 151930
rect 85947 149953 85970 150930
rect 82940 149930 85970 149953
rect 86130 149953 86153 150930
rect 89137 151930 89160 152937
rect 89320 152937 92350 152960
rect 89320 151930 89343 152937
rect 89137 150930 89343 151930
rect 89137 149953 89160 150930
rect 86130 149930 89160 149953
rect 89320 149953 89343 150930
rect 92327 151930 92350 152937
rect 92510 152937 95540 152960
rect 92510 151930 92533 152937
rect 92327 150930 92533 151930
rect 92327 149953 92350 150930
rect 89320 149930 92350 149953
rect 92510 149953 92533 150930
rect 95517 151930 95540 152937
rect 95700 152937 98730 152960
rect 95700 151930 95723 152937
rect 95517 150930 95723 151930
rect 95517 149953 95540 150930
rect 92510 149930 95540 149953
rect 95700 149953 95723 150930
rect 98707 151930 98730 152937
rect 98890 152937 101920 152960
rect 98890 151930 98913 152937
rect 98707 150930 98913 151930
rect 98707 149953 98730 150930
rect 95700 149930 98730 149953
rect 98890 149953 98913 150930
rect 101897 151930 101920 152937
rect 102080 152937 105110 152960
rect 102080 151930 102103 152937
rect 101897 150930 102103 151930
rect 101897 149953 101920 150930
rect 98890 149930 101920 149953
rect 102080 149953 102103 150930
rect 105087 151930 105110 152937
rect 105270 152937 108300 152960
rect 105270 151930 105293 152937
rect 105087 150930 105293 151930
rect 105087 149953 105110 150930
rect 102080 149930 105110 149953
rect 105270 149953 105293 150930
rect 108277 151930 108300 152937
rect 108460 152937 111490 152960
rect 108460 151930 108483 152937
rect 108277 150930 108483 151930
rect 108277 149953 108300 150930
rect 105270 149930 108300 149953
rect 108460 149953 108483 150930
rect 111467 151930 111490 152937
rect 111650 152937 114680 152960
rect 111650 151930 111673 152937
rect 111467 150930 111673 151930
rect 111467 149953 111490 150930
rect 108460 149930 111490 149953
rect 111650 149953 111673 150930
rect 114657 151930 114680 152937
rect 114840 152937 117870 152960
rect 114840 151930 114863 152937
rect 114657 150930 114863 151930
rect 114657 149953 114680 150930
rect 111650 149930 114680 149953
rect 114840 149953 114863 150930
rect 117847 151930 117870 152937
rect 118030 152937 121060 152960
rect 118030 151930 118053 152937
rect 117847 150930 118053 151930
rect 117847 149953 117870 150930
rect 114840 149930 117870 149953
rect 118030 149953 118053 150930
rect 121037 151930 121060 152937
rect 121220 152937 124250 152960
rect 121220 151930 121243 152937
rect 121037 150930 121243 151930
rect 121037 149953 121060 150930
rect 118030 149930 121060 149953
rect 121220 149953 121243 150930
rect 124227 151930 124250 152937
rect 124410 152937 127440 152960
rect 124410 151930 124433 152937
rect 124227 150930 124433 151930
rect 124227 149953 124250 150930
rect 121220 149930 124250 149953
rect 124410 149953 124433 150930
rect 127417 151930 127440 152937
rect 127600 152937 130630 152960
rect 127600 151930 127623 152937
rect 127417 150930 127623 151930
rect 127417 149953 127440 150930
rect 124410 149930 127440 149953
rect 127600 149953 127623 150930
rect 130607 151930 130630 152937
rect 130790 152937 133820 152960
rect 130790 151930 130813 152937
rect 130607 150930 130813 151930
rect 130607 149953 130630 150930
rect 127600 149930 130630 149953
rect 130790 149953 130813 150930
rect 133797 151930 133820 152937
rect 133980 152937 137010 152960
rect 133980 151930 134003 152937
rect 133797 150930 134003 151930
rect 133797 149953 133820 150930
rect 130790 149930 133820 149953
rect 133980 149953 134003 150930
rect 136987 151930 137010 152937
rect 136987 150930 137170 151930
rect 136987 149953 137010 150930
rect 133980 149930 137010 149953
rect 1000 149770 2000 149930
rect 4190 149770 5190 149930
rect 7380 149770 8380 149930
rect 10570 149770 11570 149930
rect 13760 149770 14760 149930
rect 16950 149770 17950 149930
rect 20140 149770 21140 149930
rect 23330 149770 24330 149930
rect 26520 149770 27520 149930
rect 29710 149770 30710 149930
rect 32900 149770 33900 149930
rect 36090 149770 37090 149930
rect 39280 149770 40280 149930
rect 42470 149770 43470 149930
rect 45660 149770 46660 149930
rect 48850 149770 49850 149930
rect 52040 149770 53040 149930
rect 55230 149770 56230 149930
rect 58420 149770 59420 149930
rect 61610 149770 62610 149930
rect 64800 149770 65800 149930
rect 67990 149770 68990 149930
rect 71180 149770 72180 149930
rect 74370 149770 75370 149930
rect 77560 149770 78560 149930
rect 80750 149770 81750 149930
rect 83940 149770 84940 149930
rect 87130 149770 88130 149930
rect 90320 149770 91320 149930
rect 93510 149770 94510 149930
rect 96700 149770 97700 149930
rect 99890 149770 100890 149930
rect 103080 149770 104080 149930
rect 106270 149770 107270 149930
rect 109460 149770 110460 149930
rect 112650 149770 113650 149930
rect 115840 149770 116840 149930
rect 119030 149770 120030 149930
rect 122220 149770 123220 149930
rect 125410 149770 126410 149930
rect 128600 149770 129600 149930
rect 131790 149770 132790 149930
rect 134980 149770 135980 149930
rect 0 149747 3030 149770
rect 0 146763 23 149747
rect 3007 148740 3030 149747
rect 3190 149747 6220 149770
rect 3190 148740 3213 149747
rect 3007 147740 3213 148740
rect 3007 146763 3030 147740
rect 0 146740 3030 146763
rect 3190 146763 3213 147740
rect 6197 148740 6220 149747
rect 6380 149747 9410 149770
rect 6380 148740 6403 149747
rect 6197 147740 6403 148740
rect 6197 146763 6220 147740
rect 3190 146740 6220 146763
rect 6380 146763 6403 147740
rect 9387 148740 9410 149747
rect 9570 149747 12600 149770
rect 9570 148740 9593 149747
rect 9387 147740 9593 148740
rect 9387 146763 9410 147740
rect 6380 146740 9410 146763
rect 9570 146763 9593 147740
rect 12577 148740 12600 149747
rect 12760 149747 15790 149770
rect 12760 148740 12783 149747
rect 12577 147740 12783 148740
rect 12577 146763 12600 147740
rect 9570 146740 12600 146763
rect 12760 146763 12783 147740
rect 15767 148740 15790 149747
rect 15950 149747 18980 149770
rect 15950 148740 15973 149747
rect 15767 147740 15973 148740
rect 15767 146763 15790 147740
rect 12760 146740 15790 146763
rect 15950 146763 15973 147740
rect 18957 148740 18980 149747
rect 19140 149747 22170 149770
rect 19140 148740 19163 149747
rect 18957 147740 19163 148740
rect 18957 146763 18980 147740
rect 15950 146740 18980 146763
rect 19140 146763 19163 147740
rect 22147 148740 22170 149747
rect 22330 149747 25360 149770
rect 22330 148740 22353 149747
rect 22147 147740 22353 148740
rect 22147 146763 22170 147740
rect 19140 146740 22170 146763
rect 22330 146763 22353 147740
rect 25337 148740 25360 149747
rect 25520 149747 28550 149770
rect 25520 148740 25543 149747
rect 25337 147740 25543 148740
rect 25337 146763 25360 147740
rect 22330 146740 25360 146763
rect 25520 146763 25543 147740
rect 28527 148740 28550 149747
rect 28710 149747 31740 149770
rect 28710 148740 28733 149747
rect 28527 147740 28733 148740
rect 28527 146763 28550 147740
rect 25520 146740 28550 146763
rect 28710 146763 28733 147740
rect 31717 148740 31740 149747
rect 31900 149747 34930 149770
rect 31900 148740 31923 149747
rect 31717 147740 31923 148740
rect 31717 146763 31740 147740
rect 28710 146740 31740 146763
rect 31900 146763 31923 147740
rect 34907 148740 34930 149747
rect 35090 149747 38120 149770
rect 35090 148740 35113 149747
rect 34907 147740 35113 148740
rect 34907 146763 34930 147740
rect 31900 146740 34930 146763
rect 35090 146763 35113 147740
rect 38097 148740 38120 149747
rect 38280 149747 41310 149770
rect 38280 148740 38303 149747
rect 38097 147740 38303 148740
rect 38097 146763 38120 147740
rect 35090 146740 38120 146763
rect 38280 146763 38303 147740
rect 41287 148740 41310 149747
rect 41470 149747 44500 149770
rect 41470 148740 41493 149747
rect 41287 147740 41493 148740
rect 41287 146763 41310 147740
rect 38280 146740 41310 146763
rect 41470 146763 41493 147740
rect 44477 148740 44500 149747
rect 44660 149747 47690 149770
rect 44660 148740 44683 149747
rect 44477 147740 44683 148740
rect 44477 146763 44500 147740
rect 41470 146740 44500 146763
rect 44660 146763 44683 147740
rect 47667 148740 47690 149747
rect 47850 149747 50880 149770
rect 47850 148740 47873 149747
rect 47667 147740 47873 148740
rect 47667 146763 47690 147740
rect 44660 146740 47690 146763
rect 47850 146763 47873 147740
rect 50857 148740 50880 149747
rect 51040 149747 54070 149770
rect 51040 148740 51063 149747
rect 50857 147740 51063 148740
rect 50857 146763 50880 147740
rect 47850 146740 50880 146763
rect 51040 146763 51063 147740
rect 54047 148740 54070 149747
rect 54230 149747 57260 149770
rect 54230 148740 54253 149747
rect 54047 147740 54253 148740
rect 54047 146763 54070 147740
rect 51040 146740 54070 146763
rect 54230 146763 54253 147740
rect 57237 148740 57260 149747
rect 57420 149747 60450 149770
rect 57420 148740 57443 149747
rect 57237 147740 57443 148740
rect 57237 146763 57260 147740
rect 54230 146740 57260 146763
rect 57420 146763 57443 147740
rect 60427 148740 60450 149747
rect 60610 149747 63640 149770
rect 60610 148740 60633 149747
rect 60427 147740 60633 148740
rect 60427 146763 60450 147740
rect 57420 146740 60450 146763
rect 60610 146763 60633 147740
rect 63617 148740 63640 149747
rect 63800 149747 66830 149770
rect 63800 148740 63823 149747
rect 63617 147740 63823 148740
rect 63617 146763 63640 147740
rect 60610 146740 63640 146763
rect 63800 146763 63823 147740
rect 66807 148740 66830 149747
rect 66990 149747 70020 149770
rect 66990 148740 67013 149747
rect 66807 147740 67013 148740
rect 66807 146763 66830 147740
rect 63800 146740 66830 146763
rect 66990 146763 67013 147740
rect 69997 148740 70020 149747
rect 70180 149747 73210 149770
rect 70180 148740 70203 149747
rect 69997 147740 70203 148740
rect 69997 146763 70020 147740
rect 66990 146740 70020 146763
rect 70180 146763 70203 147740
rect 73187 148740 73210 149747
rect 73370 149747 76400 149770
rect 73370 148740 73393 149747
rect 73187 147740 73393 148740
rect 73187 146763 73210 147740
rect 70180 146740 73210 146763
rect 73370 146763 73393 147740
rect 76377 148740 76400 149747
rect 76560 149747 79590 149770
rect 76560 148740 76583 149747
rect 76377 147740 76583 148740
rect 76377 146763 76400 147740
rect 73370 146740 76400 146763
rect 76560 146763 76583 147740
rect 79567 148740 79590 149747
rect 79750 149747 82780 149770
rect 79750 148740 79773 149747
rect 79567 147740 79773 148740
rect 79567 146763 79590 147740
rect 76560 146740 79590 146763
rect 79750 146763 79773 147740
rect 82757 148740 82780 149747
rect 82940 149747 85970 149770
rect 82940 148740 82963 149747
rect 82757 147740 82963 148740
rect 82757 146763 82780 147740
rect 79750 146740 82780 146763
rect 82940 146763 82963 147740
rect 85947 148740 85970 149747
rect 86130 149747 89160 149770
rect 86130 148740 86153 149747
rect 85947 147740 86153 148740
rect 85947 146763 85970 147740
rect 82940 146740 85970 146763
rect 86130 146763 86153 147740
rect 89137 148740 89160 149747
rect 89320 149747 92350 149770
rect 89320 148740 89343 149747
rect 89137 147740 89343 148740
rect 89137 146763 89160 147740
rect 86130 146740 89160 146763
rect 89320 146763 89343 147740
rect 92327 148740 92350 149747
rect 92510 149747 95540 149770
rect 92510 148740 92533 149747
rect 92327 147740 92533 148740
rect 92327 146763 92350 147740
rect 89320 146740 92350 146763
rect 92510 146763 92533 147740
rect 95517 148740 95540 149747
rect 95700 149747 98730 149770
rect 95700 148740 95723 149747
rect 95517 147740 95723 148740
rect 95517 146763 95540 147740
rect 92510 146740 95540 146763
rect 95700 146763 95723 147740
rect 98707 148740 98730 149747
rect 98890 149747 101920 149770
rect 98890 148740 98913 149747
rect 98707 147740 98913 148740
rect 98707 146763 98730 147740
rect 95700 146740 98730 146763
rect 98890 146763 98913 147740
rect 101897 148740 101920 149747
rect 102080 149747 105110 149770
rect 102080 148740 102103 149747
rect 101897 147740 102103 148740
rect 101897 146763 101920 147740
rect 98890 146740 101920 146763
rect 102080 146763 102103 147740
rect 105087 148740 105110 149747
rect 105270 149747 108300 149770
rect 105270 148740 105293 149747
rect 105087 147740 105293 148740
rect 105087 146763 105110 147740
rect 102080 146740 105110 146763
rect 105270 146763 105293 147740
rect 108277 148740 108300 149747
rect 108460 149747 111490 149770
rect 108460 148740 108483 149747
rect 108277 147740 108483 148740
rect 108277 146763 108300 147740
rect 105270 146740 108300 146763
rect 108460 146763 108483 147740
rect 111467 148740 111490 149747
rect 111650 149747 114680 149770
rect 111650 148740 111673 149747
rect 111467 147740 111673 148740
rect 111467 146763 111490 147740
rect 108460 146740 111490 146763
rect 111650 146763 111673 147740
rect 114657 148740 114680 149747
rect 114840 149747 117870 149770
rect 114840 148740 114863 149747
rect 114657 147740 114863 148740
rect 114657 146763 114680 147740
rect 111650 146740 114680 146763
rect 114840 146763 114863 147740
rect 117847 148740 117870 149747
rect 118030 149747 121060 149770
rect 118030 148740 118053 149747
rect 117847 147740 118053 148740
rect 117847 146763 117870 147740
rect 114840 146740 117870 146763
rect 118030 146763 118053 147740
rect 121037 148740 121060 149747
rect 121220 149747 124250 149770
rect 121220 148740 121243 149747
rect 121037 147740 121243 148740
rect 121037 146763 121060 147740
rect 118030 146740 121060 146763
rect 121220 146763 121243 147740
rect 124227 148740 124250 149747
rect 124410 149747 127440 149770
rect 124410 148740 124433 149747
rect 124227 147740 124433 148740
rect 124227 146763 124250 147740
rect 121220 146740 124250 146763
rect 124410 146763 124433 147740
rect 127417 148740 127440 149747
rect 127600 149747 130630 149770
rect 127600 148740 127623 149747
rect 127417 147740 127623 148740
rect 127417 146763 127440 147740
rect 124410 146740 127440 146763
rect 127600 146763 127623 147740
rect 130607 148740 130630 149747
rect 130790 149747 133820 149770
rect 130790 148740 130813 149747
rect 130607 147740 130813 148740
rect 130607 146763 130630 147740
rect 127600 146740 130630 146763
rect 130790 146763 130813 147740
rect 133797 148740 133820 149747
rect 133980 149747 137010 149770
rect 133980 148740 134003 149747
rect 133797 147740 134003 148740
rect 133797 146763 133820 147740
rect 130790 146740 133820 146763
rect 133980 146763 134003 147740
rect 136987 148740 137010 149747
rect 136987 147740 137170 148740
rect 136987 146763 137010 147740
rect 133980 146740 137010 146763
rect 1000 146580 2000 146740
rect 4190 146580 5190 146740
rect 7380 146580 8380 146740
rect 10570 146580 11570 146740
rect 13760 146580 14760 146740
rect 16950 146580 17950 146740
rect 20140 146580 21140 146740
rect 23330 146580 24330 146740
rect 26520 146580 27520 146740
rect 29710 146580 30710 146740
rect 32900 146580 33900 146740
rect 36090 146580 37090 146740
rect 39280 146580 40280 146740
rect 42470 146580 43470 146740
rect 45660 146580 46660 146740
rect 48850 146580 49850 146740
rect 52040 146580 53040 146740
rect 55230 146580 56230 146740
rect 58420 146580 59420 146740
rect 61610 146580 62610 146740
rect 64800 146580 65800 146740
rect 67990 146580 68990 146740
rect 71180 146580 72180 146740
rect 74370 146580 75370 146740
rect 77560 146580 78560 146740
rect 80750 146580 81750 146740
rect 83940 146580 84940 146740
rect 87130 146580 88130 146740
rect 90320 146580 91320 146740
rect 93510 146580 94510 146740
rect 96700 146580 97700 146740
rect 99890 146580 100890 146740
rect 103080 146580 104080 146740
rect 106270 146580 107270 146740
rect 109460 146580 110460 146740
rect 112650 146580 113650 146740
rect 115840 146580 116840 146740
rect 119030 146580 120030 146740
rect 122220 146580 123220 146740
rect 125410 146580 126410 146740
rect 128600 146580 129600 146740
rect 131790 146580 132790 146740
rect 134980 146580 135980 146740
rect 0 146557 3030 146580
rect 0 143573 23 146557
rect 3007 145550 3030 146557
rect 3190 146557 6220 146580
rect 3190 145550 3213 146557
rect 3007 144550 3213 145550
rect 3007 143573 3030 144550
rect 0 143550 3030 143573
rect 3190 143573 3213 144550
rect 6197 145550 6220 146557
rect 6380 146557 9410 146580
rect 6380 145550 6403 146557
rect 6197 144550 6403 145550
rect 6197 143573 6220 144550
rect 3190 143550 6220 143573
rect 6380 143573 6403 144550
rect 9387 145550 9410 146557
rect 9570 146557 12600 146580
rect 9570 145550 9593 146557
rect 9387 144550 9593 145550
rect 9387 143573 9410 144550
rect 6380 143550 9410 143573
rect 9570 143573 9593 144550
rect 12577 145550 12600 146557
rect 12760 146557 15790 146580
rect 12760 145550 12783 146557
rect 12577 144550 12783 145550
rect 12577 143573 12600 144550
rect 9570 143550 12600 143573
rect 12760 143573 12783 144550
rect 15767 145550 15790 146557
rect 15950 146557 18980 146580
rect 15950 145550 15973 146557
rect 15767 144550 15973 145550
rect 15767 143573 15790 144550
rect 12760 143550 15790 143573
rect 15950 143573 15973 144550
rect 18957 145550 18980 146557
rect 19140 146557 22170 146580
rect 19140 145550 19163 146557
rect 18957 144550 19163 145550
rect 18957 143573 18980 144550
rect 15950 143550 18980 143573
rect 19140 143573 19163 144550
rect 22147 145550 22170 146557
rect 22330 146557 25360 146580
rect 22330 145550 22353 146557
rect 22147 144550 22353 145550
rect 22147 143573 22170 144550
rect 19140 143550 22170 143573
rect 22330 143573 22353 144550
rect 25337 145550 25360 146557
rect 25520 146557 28550 146580
rect 25520 145550 25543 146557
rect 25337 144550 25543 145550
rect 25337 143573 25360 144550
rect 22330 143550 25360 143573
rect 25520 143573 25543 144550
rect 28527 145550 28550 146557
rect 28710 146557 31740 146580
rect 28710 145550 28733 146557
rect 28527 144550 28733 145550
rect 28527 143573 28550 144550
rect 25520 143550 28550 143573
rect 28710 143573 28733 144550
rect 31717 145550 31740 146557
rect 31900 146557 34930 146580
rect 31900 145550 31923 146557
rect 31717 144550 31923 145550
rect 31717 143573 31740 144550
rect 28710 143550 31740 143573
rect 31900 143573 31923 144550
rect 34907 145550 34930 146557
rect 35090 146557 38120 146580
rect 35090 145550 35113 146557
rect 34907 144550 35113 145550
rect 34907 143573 34930 144550
rect 31900 143550 34930 143573
rect 35090 143573 35113 144550
rect 38097 145550 38120 146557
rect 38280 146557 41310 146580
rect 38280 145550 38303 146557
rect 38097 144550 38303 145550
rect 38097 143573 38120 144550
rect 35090 143550 38120 143573
rect 38280 143573 38303 144550
rect 41287 145550 41310 146557
rect 41470 146557 44500 146580
rect 41470 145550 41493 146557
rect 41287 144550 41493 145550
rect 41287 143573 41310 144550
rect 38280 143550 41310 143573
rect 41470 143573 41493 144550
rect 44477 145550 44500 146557
rect 44660 146557 47690 146580
rect 44660 145550 44683 146557
rect 44477 144550 44683 145550
rect 44477 143573 44500 144550
rect 41470 143550 44500 143573
rect 44660 143573 44683 144550
rect 47667 145550 47690 146557
rect 47850 146557 50880 146580
rect 47850 145550 47873 146557
rect 47667 144550 47873 145550
rect 47667 143573 47690 144550
rect 44660 143550 47690 143573
rect 47850 143573 47873 144550
rect 50857 145550 50880 146557
rect 51040 146557 54070 146580
rect 51040 145550 51063 146557
rect 50857 144550 51063 145550
rect 50857 143573 50880 144550
rect 47850 143550 50880 143573
rect 51040 143573 51063 144550
rect 54047 145550 54070 146557
rect 54230 146557 57260 146580
rect 54230 145550 54253 146557
rect 54047 144550 54253 145550
rect 54047 143573 54070 144550
rect 51040 143550 54070 143573
rect 54230 143573 54253 144550
rect 57237 145550 57260 146557
rect 57420 146557 60450 146580
rect 57420 145550 57443 146557
rect 57237 144550 57443 145550
rect 57237 143573 57260 144550
rect 54230 143550 57260 143573
rect 57420 143573 57443 144550
rect 60427 145550 60450 146557
rect 60610 146557 63640 146580
rect 60610 145550 60633 146557
rect 60427 144550 60633 145550
rect 60427 143573 60450 144550
rect 57420 143550 60450 143573
rect 60610 143573 60633 144550
rect 63617 145550 63640 146557
rect 63800 146557 66830 146580
rect 63800 145550 63823 146557
rect 63617 144550 63823 145550
rect 63617 143573 63640 144550
rect 60610 143550 63640 143573
rect 63800 143573 63823 144550
rect 66807 145550 66830 146557
rect 66990 146557 70020 146580
rect 66990 145550 67013 146557
rect 66807 144550 67013 145550
rect 66807 143573 66830 144550
rect 63800 143550 66830 143573
rect 66990 143573 67013 144550
rect 69997 145550 70020 146557
rect 70180 146557 73210 146580
rect 70180 145550 70203 146557
rect 69997 144550 70203 145550
rect 69997 143573 70020 144550
rect 66990 143550 70020 143573
rect 70180 143573 70203 144550
rect 73187 145550 73210 146557
rect 73370 146557 76400 146580
rect 73370 145550 73393 146557
rect 73187 144550 73393 145550
rect 73187 143573 73210 144550
rect 70180 143550 73210 143573
rect 73370 143573 73393 144550
rect 76377 145550 76400 146557
rect 76560 146557 79590 146580
rect 76560 145550 76583 146557
rect 76377 144550 76583 145550
rect 76377 143573 76400 144550
rect 73370 143550 76400 143573
rect 76560 143573 76583 144550
rect 79567 145550 79590 146557
rect 79750 146557 82780 146580
rect 79750 145550 79773 146557
rect 79567 144550 79773 145550
rect 79567 143573 79590 144550
rect 76560 143550 79590 143573
rect 79750 143573 79773 144550
rect 82757 145550 82780 146557
rect 82940 146557 85970 146580
rect 82940 145550 82963 146557
rect 82757 144550 82963 145550
rect 82757 143573 82780 144550
rect 79750 143550 82780 143573
rect 82940 143573 82963 144550
rect 85947 145550 85970 146557
rect 86130 146557 89160 146580
rect 86130 145550 86153 146557
rect 85947 144550 86153 145550
rect 85947 143573 85970 144550
rect 82940 143550 85970 143573
rect 86130 143573 86153 144550
rect 89137 145550 89160 146557
rect 89320 146557 92350 146580
rect 89320 145550 89343 146557
rect 89137 144550 89343 145550
rect 89137 143573 89160 144550
rect 86130 143550 89160 143573
rect 89320 143573 89343 144550
rect 92327 145550 92350 146557
rect 92510 146557 95540 146580
rect 92510 145550 92533 146557
rect 92327 144550 92533 145550
rect 92327 143573 92350 144550
rect 89320 143550 92350 143573
rect 92510 143573 92533 144550
rect 95517 145550 95540 146557
rect 95700 146557 98730 146580
rect 95700 145550 95723 146557
rect 95517 144550 95723 145550
rect 95517 143573 95540 144550
rect 92510 143550 95540 143573
rect 95700 143573 95723 144550
rect 98707 145550 98730 146557
rect 98890 146557 101920 146580
rect 98890 145550 98913 146557
rect 98707 144550 98913 145550
rect 98707 143573 98730 144550
rect 95700 143550 98730 143573
rect 98890 143573 98913 144550
rect 101897 145550 101920 146557
rect 102080 146557 105110 146580
rect 102080 145550 102103 146557
rect 101897 144550 102103 145550
rect 101897 143573 101920 144550
rect 98890 143550 101920 143573
rect 102080 143573 102103 144550
rect 105087 145550 105110 146557
rect 105270 146557 108300 146580
rect 105270 145550 105293 146557
rect 105087 144550 105293 145550
rect 105087 143573 105110 144550
rect 102080 143550 105110 143573
rect 105270 143573 105293 144550
rect 108277 145550 108300 146557
rect 108460 146557 111490 146580
rect 108460 145550 108483 146557
rect 108277 144550 108483 145550
rect 108277 143573 108300 144550
rect 105270 143550 108300 143573
rect 108460 143573 108483 144550
rect 111467 145550 111490 146557
rect 111650 146557 114680 146580
rect 111650 145550 111673 146557
rect 111467 144550 111673 145550
rect 111467 143573 111490 144550
rect 108460 143550 111490 143573
rect 111650 143573 111673 144550
rect 114657 145550 114680 146557
rect 114840 146557 117870 146580
rect 114840 145550 114863 146557
rect 114657 144550 114863 145550
rect 114657 143573 114680 144550
rect 111650 143550 114680 143573
rect 114840 143573 114863 144550
rect 117847 145550 117870 146557
rect 118030 146557 121060 146580
rect 118030 145550 118053 146557
rect 117847 144550 118053 145550
rect 117847 143573 117870 144550
rect 114840 143550 117870 143573
rect 118030 143573 118053 144550
rect 121037 145550 121060 146557
rect 121220 146557 124250 146580
rect 121220 145550 121243 146557
rect 121037 144550 121243 145550
rect 121037 143573 121060 144550
rect 118030 143550 121060 143573
rect 121220 143573 121243 144550
rect 124227 145550 124250 146557
rect 124410 146557 127440 146580
rect 124410 145550 124433 146557
rect 124227 144550 124433 145550
rect 124227 143573 124250 144550
rect 121220 143550 124250 143573
rect 124410 143573 124433 144550
rect 127417 145550 127440 146557
rect 127600 146557 130630 146580
rect 127600 145550 127623 146557
rect 127417 144550 127623 145550
rect 127417 143573 127440 144550
rect 124410 143550 127440 143573
rect 127600 143573 127623 144550
rect 130607 145550 130630 146557
rect 130790 146557 133820 146580
rect 130790 145550 130813 146557
rect 130607 144550 130813 145550
rect 130607 143573 130630 144550
rect 127600 143550 130630 143573
rect 130790 143573 130813 144550
rect 133797 145550 133820 146557
rect 133980 146557 137010 146580
rect 133980 145550 134003 146557
rect 133797 144550 134003 145550
rect 133797 143573 133820 144550
rect 130790 143550 133820 143573
rect 133980 143573 134003 144550
rect 136987 145550 137010 146557
rect 136987 144550 137170 145550
rect 136987 143573 137010 144550
rect 133980 143550 137010 143573
rect 1000 143390 2000 143550
rect 4190 143390 5190 143550
rect 7380 143390 8380 143550
rect 10570 143390 11570 143550
rect 13760 143390 14760 143550
rect 16950 143390 17950 143550
rect 20140 143390 21140 143550
rect 23330 143390 24330 143550
rect 26520 143390 27520 143550
rect 29710 143390 30710 143550
rect 32900 143390 33900 143550
rect 36090 143390 37090 143550
rect 39280 143390 40280 143550
rect 42470 143390 43470 143550
rect 45660 143390 46660 143550
rect 48850 143390 49850 143550
rect 52040 143390 53040 143550
rect 55230 143390 56230 143550
rect 58420 143390 59420 143550
rect 61610 143390 62610 143550
rect 64800 143390 65800 143550
rect 67990 143390 68990 143550
rect 71180 143390 72180 143550
rect 74370 143390 75370 143550
rect 77560 143390 78560 143550
rect 80750 143390 81750 143550
rect 83940 143390 84940 143550
rect 87130 143390 88130 143550
rect 90320 143390 91320 143550
rect 93510 143390 94510 143550
rect 96700 143390 97700 143550
rect 99890 143390 100890 143550
rect 103080 143390 104080 143550
rect 106270 143390 107270 143550
rect 109460 143390 110460 143550
rect 112650 143390 113650 143550
rect 115840 143390 116840 143550
rect 119030 143390 120030 143550
rect 122220 143390 123220 143550
rect 125410 143390 126410 143550
rect 128600 143390 129600 143550
rect 131790 143390 132790 143550
rect 134980 143390 135980 143550
rect 0 143367 3030 143390
rect 0 140383 23 143367
rect 3007 142360 3030 143367
rect 3190 143367 6220 143390
rect 3190 142360 3213 143367
rect 3007 141360 3213 142360
rect 3007 140383 3030 141360
rect 0 140360 3030 140383
rect 3190 140383 3213 141360
rect 6197 142360 6220 143367
rect 6380 143367 9410 143390
rect 6380 142360 6403 143367
rect 6197 141360 6403 142360
rect 6197 140383 6220 141360
rect 3190 140360 6220 140383
rect 6380 140383 6403 141360
rect 9387 142360 9410 143367
rect 9570 143367 12600 143390
rect 9570 142360 9593 143367
rect 9387 141360 9593 142360
rect 9387 140383 9410 141360
rect 6380 140360 9410 140383
rect 9570 140383 9593 141360
rect 12577 142360 12600 143367
rect 12760 143367 15790 143390
rect 12760 142360 12783 143367
rect 12577 141360 12783 142360
rect 12577 140383 12600 141360
rect 9570 140360 12600 140383
rect 12760 140383 12783 141360
rect 15767 142360 15790 143367
rect 15950 143367 18980 143390
rect 15950 142360 15973 143367
rect 15767 141360 15973 142360
rect 15767 140383 15790 141360
rect 12760 140360 15790 140383
rect 15950 140383 15973 141360
rect 18957 142360 18980 143367
rect 19140 143367 22170 143390
rect 19140 142360 19163 143367
rect 18957 141360 19163 142360
rect 18957 140383 18980 141360
rect 15950 140360 18980 140383
rect 19140 140383 19163 141360
rect 22147 142360 22170 143367
rect 22330 143367 25360 143390
rect 22330 142360 22353 143367
rect 22147 141360 22353 142360
rect 22147 140383 22170 141360
rect 19140 140360 22170 140383
rect 22330 140383 22353 141360
rect 25337 142360 25360 143367
rect 25520 143367 28550 143390
rect 25520 142360 25543 143367
rect 25337 141360 25543 142360
rect 25337 140383 25360 141360
rect 22330 140360 25360 140383
rect 25520 140383 25543 141360
rect 28527 142360 28550 143367
rect 28710 143367 31740 143390
rect 28710 142360 28733 143367
rect 28527 141360 28733 142360
rect 28527 140383 28550 141360
rect 25520 140360 28550 140383
rect 28710 140383 28733 141360
rect 31717 142360 31740 143367
rect 31900 143367 34930 143390
rect 31900 142360 31923 143367
rect 31717 141360 31923 142360
rect 31717 140383 31740 141360
rect 28710 140360 31740 140383
rect 31900 140383 31923 141360
rect 34907 142360 34930 143367
rect 35090 143367 38120 143390
rect 35090 142360 35113 143367
rect 34907 141360 35113 142360
rect 34907 140383 34930 141360
rect 31900 140360 34930 140383
rect 35090 140383 35113 141360
rect 38097 142360 38120 143367
rect 38280 143367 41310 143390
rect 38280 142360 38303 143367
rect 38097 141360 38303 142360
rect 38097 140383 38120 141360
rect 35090 140360 38120 140383
rect 38280 140383 38303 141360
rect 41287 142360 41310 143367
rect 41470 143367 44500 143390
rect 41470 142360 41493 143367
rect 41287 141360 41493 142360
rect 41287 140383 41310 141360
rect 38280 140360 41310 140383
rect 41470 140383 41493 141360
rect 44477 142360 44500 143367
rect 44660 143367 47690 143390
rect 44660 142360 44683 143367
rect 44477 141360 44683 142360
rect 44477 140383 44500 141360
rect 41470 140360 44500 140383
rect 44660 140383 44683 141360
rect 47667 142360 47690 143367
rect 47850 143367 50880 143390
rect 47850 142360 47873 143367
rect 47667 141360 47873 142360
rect 47667 140383 47690 141360
rect 44660 140360 47690 140383
rect 47850 140383 47873 141360
rect 50857 142360 50880 143367
rect 51040 143367 54070 143390
rect 51040 142360 51063 143367
rect 50857 141360 51063 142360
rect 50857 140383 50880 141360
rect 47850 140360 50880 140383
rect 51040 140383 51063 141360
rect 54047 142360 54070 143367
rect 54230 143367 57260 143390
rect 54230 142360 54253 143367
rect 54047 141360 54253 142360
rect 54047 140383 54070 141360
rect 51040 140360 54070 140383
rect 54230 140383 54253 141360
rect 57237 142360 57260 143367
rect 57420 143367 60450 143390
rect 57420 142360 57443 143367
rect 57237 141360 57443 142360
rect 57237 140383 57260 141360
rect 54230 140360 57260 140383
rect 57420 140383 57443 141360
rect 60427 142360 60450 143367
rect 60610 143367 63640 143390
rect 60610 142360 60633 143367
rect 60427 141360 60633 142360
rect 60427 140383 60450 141360
rect 57420 140360 60450 140383
rect 60610 140383 60633 141360
rect 63617 142360 63640 143367
rect 63800 143367 66830 143390
rect 63800 142360 63823 143367
rect 63617 141360 63823 142360
rect 63617 140383 63640 141360
rect 60610 140360 63640 140383
rect 63800 140383 63823 141360
rect 66807 142360 66830 143367
rect 66990 143367 70020 143390
rect 66990 142360 67013 143367
rect 66807 141360 67013 142360
rect 66807 140383 66830 141360
rect 63800 140360 66830 140383
rect 66990 140383 67013 141360
rect 69997 142360 70020 143367
rect 70180 143367 73210 143390
rect 70180 142360 70203 143367
rect 69997 141360 70203 142360
rect 69997 140383 70020 141360
rect 66990 140360 70020 140383
rect 70180 140383 70203 141360
rect 73187 142360 73210 143367
rect 73370 143367 76400 143390
rect 73370 142360 73393 143367
rect 73187 141360 73393 142360
rect 73187 140383 73210 141360
rect 70180 140360 73210 140383
rect 73370 140383 73393 141360
rect 76377 142360 76400 143367
rect 76560 143367 79590 143390
rect 76560 142360 76583 143367
rect 76377 141360 76583 142360
rect 76377 140383 76400 141360
rect 73370 140360 76400 140383
rect 76560 140383 76583 141360
rect 79567 142360 79590 143367
rect 79750 143367 82780 143390
rect 79750 142360 79773 143367
rect 79567 141360 79773 142360
rect 79567 140383 79590 141360
rect 76560 140360 79590 140383
rect 79750 140383 79773 141360
rect 82757 142360 82780 143367
rect 82940 143367 85970 143390
rect 82940 142360 82963 143367
rect 82757 141360 82963 142360
rect 82757 140383 82780 141360
rect 79750 140360 82780 140383
rect 82940 140383 82963 141360
rect 85947 142360 85970 143367
rect 86130 143367 89160 143390
rect 86130 142360 86153 143367
rect 85947 141360 86153 142360
rect 85947 140383 85970 141360
rect 82940 140360 85970 140383
rect 86130 140383 86153 141360
rect 89137 142360 89160 143367
rect 89320 143367 92350 143390
rect 89320 142360 89343 143367
rect 89137 141360 89343 142360
rect 89137 140383 89160 141360
rect 86130 140360 89160 140383
rect 89320 140383 89343 141360
rect 92327 142360 92350 143367
rect 92510 143367 95540 143390
rect 92510 142360 92533 143367
rect 92327 141360 92533 142360
rect 92327 140383 92350 141360
rect 89320 140360 92350 140383
rect 92510 140383 92533 141360
rect 95517 142360 95540 143367
rect 95700 143367 98730 143390
rect 95700 142360 95723 143367
rect 95517 141360 95723 142360
rect 95517 140383 95540 141360
rect 92510 140360 95540 140383
rect 95700 140383 95723 141360
rect 98707 142360 98730 143367
rect 98890 143367 101920 143390
rect 98890 142360 98913 143367
rect 98707 141360 98913 142360
rect 98707 140383 98730 141360
rect 95700 140360 98730 140383
rect 98890 140383 98913 141360
rect 101897 142360 101920 143367
rect 102080 143367 105110 143390
rect 102080 142360 102103 143367
rect 101897 141360 102103 142360
rect 101897 140383 101920 141360
rect 98890 140360 101920 140383
rect 102080 140383 102103 141360
rect 105087 142360 105110 143367
rect 105270 143367 108300 143390
rect 105270 142360 105293 143367
rect 105087 141360 105293 142360
rect 105087 140383 105110 141360
rect 102080 140360 105110 140383
rect 105270 140383 105293 141360
rect 108277 142360 108300 143367
rect 108460 143367 111490 143390
rect 108460 142360 108483 143367
rect 108277 141360 108483 142360
rect 108277 140383 108300 141360
rect 105270 140360 108300 140383
rect 108460 140383 108483 141360
rect 111467 142360 111490 143367
rect 111650 143367 114680 143390
rect 111650 142360 111673 143367
rect 111467 141360 111673 142360
rect 111467 140383 111490 141360
rect 108460 140360 111490 140383
rect 111650 140383 111673 141360
rect 114657 142360 114680 143367
rect 114840 143367 117870 143390
rect 114840 142360 114863 143367
rect 114657 141360 114863 142360
rect 114657 140383 114680 141360
rect 111650 140360 114680 140383
rect 114840 140383 114863 141360
rect 117847 142360 117870 143367
rect 118030 143367 121060 143390
rect 118030 142360 118053 143367
rect 117847 141360 118053 142360
rect 117847 140383 117870 141360
rect 114840 140360 117870 140383
rect 118030 140383 118053 141360
rect 121037 142360 121060 143367
rect 121220 143367 124250 143390
rect 121220 142360 121243 143367
rect 121037 141360 121243 142360
rect 121037 140383 121060 141360
rect 118030 140360 121060 140383
rect 121220 140383 121243 141360
rect 124227 142360 124250 143367
rect 124410 143367 127440 143390
rect 124410 142360 124433 143367
rect 124227 141360 124433 142360
rect 124227 140383 124250 141360
rect 121220 140360 124250 140383
rect 124410 140383 124433 141360
rect 127417 142360 127440 143367
rect 127600 143367 130630 143390
rect 127600 142360 127623 143367
rect 127417 141360 127623 142360
rect 127417 140383 127440 141360
rect 124410 140360 127440 140383
rect 127600 140383 127623 141360
rect 130607 142360 130630 143367
rect 130790 143367 133820 143390
rect 130790 142360 130813 143367
rect 130607 141360 130813 142360
rect 130607 140383 130630 141360
rect 127600 140360 130630 140383
rect 130790 140383 130813 141360
rect 133797 142360 133820 143367
rect 133980 143367 137010 143390
rect 133980 142360 134003 143367
rect 133797 141360 134003 142360
rect 133797 140383 133820 141360
rect 130790 140360 133820 140383
rect 133980 140383 134003 141360
rect 136987 142360 137010 143367
rect 136987 141360 137170 142360
rect 136987 140383 137010 141360
rect 133980 140360 137010 140383
rect 10570 140200 11570 140360
rect 13760 140200 14760 140360
rect 16950 140200 17950 140360
rect 20140 140200 21140 140360
rect 23330 140200 24330 140360
rect 26520 140200 27520 140360
rect 29710 140200 30710 140360
rect 32900 140200 33900 140360
rect 36090 140200 37090 140360
rect 39280 140200 40280 140360
rect 42470 140200 43470 140360
rect 45660 140200 46660 140360
rect 48850 140200 49850 140360
rect 52040 140200 53040 140360
rect 55230 140200 56230 140360
rect 58420 140200 59420 140360
rect 61610 140200 62610 140360
rect 64800 140200 65800 140360
rect 67990 140200 68990 140360
rect 71180 140200 72180 140360
rect 74370 140200 75370 140360
rect 77560 140200 78560 140360
rect 80750 140200 81750 140360
rect 83940 140200 84940 140360
rect 87130 140200 88130 140360
rect 90320 140200 91320 140360
rect 93510 140200 94510 140360
rect 96700 140200 97700 140360
rect 99890 140200 100890 140360
rect 103080 140200 104080 140360
rect 106270 140200 107270 140360
rect 109460 140200 110460 140360
rect 112650 140200 113650 140360
rect 115840 140200 116840 140360
rect 119030 140200 120030 140360
rect 122220 140200 123220 140360
rect 125410 140200 126410 140360
rect 128600 140200 129600 140360
rect 131790 140200 132790 140360
rect 134980 140200 135980 140360
rect 9570 140177 12600 140200
rect 0 140110 9370 140160
rect 0 121310 50 140110
rect 9320 121310 9370 140110
rect 9570 137193 9593 140177
rect 12577 139170 12600 140177
rect 12760 140177 15790 140200
rect 12760 139170 12783 140177
rect 12577 138170 12783 139170
rect 12577 137193 12600 138170
rect 9570 137170 12600 137193
rect 12760 137193 12783 138170
rect 15767 139170 15790 140177
rect 15950 140177 18980 140200
rect 15950 139170 15973 140177
rect 15767 138170 15973 139170
rect 15767 137193 15790 138170
rect 12760 137170 15790 137193
rect 15950 137193 15973 138170
rect 18957 139170 18980 140177
rect 19140 140177 22170 140200
rect 19140 139170 19163 140177
rect 18957 138170 19163 139170
rect 18957 137193 18980 138170
rect 15950 137170 18980 137193
rect 19140 137193 19163 138170
rect 22147 139170 22170 140177
rect 22330 140177 25360 140200
rect 22330 139170 22353 140177
rect 22147 138170 22353 139170
rect 22147 137193 22170 138170
rect 19140 137170 22170 137193
rect 22330 137193 22353 138170
rect 25337 139170 25360 140177
rect 25520 140177 28550 140200
rect 25520 139170 25543 140177
rect 25337 138170 25543 139170
rect 25337 137193 25360 138170
rect 22330 137170 25360 137193
rect 25520 137193 25543 138170
rect 28527 139170 28550 140177
rect 28710 140177 31740 140200
rect 28710 139170 28733 140177
rect 28527 138170 28733 139170
rect 28527 137193 28550 138170
rect 25520 137170 28550 137193
rect 28710 137193 28733 138170
rect 31717 139170 31740 140177
rect 31900 140177 34930 140200
rect 31900 139170 31923 140177
rect 31717 138170 31923 139170
rect 31717 137193 31740 138170
rect 28710 137170 31740 137193
rect 31900 137193 31923 138170
rect 34907 139170 34930 140177
rect 35090 140177 38120 140200
rect 35090 139170 35113 140177
rect 34907 138170 35113 139170
rect 34907 137193 34930 138170
rect 31900 137170 34930 137193
rect 35090 137193 35113 138170
rect 38097 139170 38120 140177
rect 38280 140177 41310 140200
rect 38280 139170 38303 140177
rect 38097 138170 38303 139170
rect 38097 137193 38120 138170
rect 35090 137170 38120 137193
rect 38280 137193 38303 138170
rect 41287 139170 41310 140177
rect 41470 140177 44500 140200
rect 41470 139170 41493 140177
rect 41287 138170 41493 139170
rect 41287 137193 41310 138170
rect 38280 137170 41310 137193
rect 41470 137193 41493 138170
rect 44477 139170 44500 140177
rect 44660 140177 47690 140200
rect 44660 139170 44683 140177
rect 44477 138170 44683 139170
rect 44477 137193 44500 138170
rect 41470 137170 44500 137193
rect 44660 137193 44683 138170
rect 47667 139170 47690 140177
rect 47850 140177 50880 140200
rect 47850 139170 47873 140177
rect 47667 138170 47873 139170
rect 47667 137193 47690 138170
rect 44660 137170 47690 137193
rect 47850 137193 47873 138170
rect 50857 139170 50880 140177
rect 51040 140177 54070 140200
rect 51040 139170 51063 140177
rect 50857 138170 51063 139170
rect 50857 137193 50880 138170
rect 47850 137170 50880 137193
rect 51040 137193 51063 138170
rect 54047 139170 54070 140177
rect 54230 140177 57260 140200
rect 54230 139170 54253 140177
rect 54047 138170 54253 139170
rect 54047 137193 54070 138170
rect 51040 137170 54070 137193
rect 54230 137193 54253 138170
rect 57237 139170 57260 140177
rect 57420 140177 60450 140200
rect 57420 139170 57443 140177
rect 57237 138170 57443 139170
rect 57237 137193 57260 138170
rect 54230 137170 57260 137193
rect 57420 137193 57443 138170
rect 60427 139170 60450 140177
rect 60610 140177 63640 140200
rect 60610 139170 60633 140177
rect 60427 138170 60633 139170
rect 60427 137193 60450 138170
rect 57420 137170 60450 137193
rect 60610 137193 60633 138170
rect 63617 139170 63640 140177
rect 63800 140177 66830 140200
rect 63800 139170 63823 140177
rect 63617 138170 63823 139170
rect 63617 137193 63640 138170
rect 60610 137170 63640 137193
rect 63800 137193 63823 138170
rect 66807 139170 66830 140177
rect 66990 140177 70020 140200
rect 66990 139170 67013 140177
rect 66807 138170 67013 139170
rect 66807 137193 66830 138170
rect 63800 137170 66830 137193
rect 66990 137193 67013 138170
rect 69997 139170 70020 140177
rect 70180 140177 73210 140200
rect 70180 139170 70203 140177
rect 69997 138170 70203 139170
rect 69997 137193 70020 138170
rect 66990 137170 70020 137193
rect 70180 137193 70203 138170
rect 73187 139170 73210 140177
rect 73370 140177 76400 140200
rect 73370 139170 73393 140177
rect 73187 138170 73393 139170
rect 73187 137193 73210 138170
rect 70180 137170 73210 137193
rect 73370 137193 73393 138170
rect 76377 139170 76400 140177
rect 76560 140177 79590 140200
rect 76560 139170 76583 140177
rect 76377 138170 76583 139170
rect 76377 137193 76400 138170
rect 73370 137170 76400 137193
rect 76560 137193 76583 138170
rect 79567 139170 79590 140177
rect 79750 140177 82780 140200
rect 79750 139170 79773 140177
rect 79567 138170 79773 139170
rect 79567 137193 79590 138170
rect 76560 137170 79590 137193
rect 79750 137193 79773 138170
rect 82757 139170 82780 140177
rect 82940 140177 85970 140200
rect 82940 139170 82963 140177
rect 82757 138170 82963 139170
rect 82757 137193 82780 138170
rect 79750 137170 82780 137193
rect 82940 137193 82963 138170
rect 85947 139170 85970 140177
rect 86130 140177 89160 140200
rect 86130 139170 86153 140177
rect 85947 138170 86153 139170
rect 85947 137193 85970 138170
rect 82940 137170 85970 137193
rect 86130 137193 86153 138170
rect 89137 139170 89160 140177
rect 89320 140177 92350 140200
rect 89320 139170 89343 140177
rect 89137 138170 89343 139170
rect 89137 137193 89160 138170
rect 86130 137170 89160 137193
rect 89320 137193 89343 138170
rect 92327 139170 92350 140177
rect 92510 140177 95540 140200
rect 92510 139170 92533 140177
rect 92327 138170 92533 139170
rect 92327 137193 92350 138170
rect 89320 137170 92350 137193
rect 92510 137193 92533 138170
rect 95517 139170 95540 140177
rect 95700 140177 98730 140200
rect 95700 139170 95723 140177
rect 95517 138170 95723 139170
rect 95517 137193 95540 138170
rect 92510 137170 95540 137193
rect 95700 137193 95723 138170
rect 98707 139170 98730 140177
rect 98890 140177 101920 140200
rect 98890 139170 98913 140177
rect 98707 138170 98913 139170
rect 98707 137193 98730 138170
rect 95700 137170 98730 137193
rect 98890 137193 98913 138170
rect 101897 139170 101920 140177
rect 102080 140177 105110 140200
rect 102080 139170 102103 140177
rect 101897 138170 102103 139170
rect 101897 137193 101920 138170
rect 98890 137170 101920 137193
rect 102080 137193 102103 138170
rect 105087 139170 105110 140177
rect 105270 140177 108300 140200
rect 105270 139170 105293 140177
rect 105087 138170 105293 139170
rect 105087 137193 105110 138170
rect 102080 137170 105110 137193
rect 105270 137193 105293 138170
rect 108277 139170 108300 140177
rect 108460 140177 111490 140200
rect 108460 139170 108483 140177
rect 108277 138170 108483 139170
rect 108277 137193 108300 138170
rect 105270 137170 108300 137193
rect 108460 137193 108483 138170
rect 111467 139170 111490 140177
rect 111650 140177 114680 140200
rect 111650 139170 111673 140177
rect 111467 138170 111673 139170
rect 111467 137193 111490 138170
rect 108460 137170 111490 137193
rect 111650 137193 111673 138170
rect 114657 139170 114680 140177
rect 114840 140177 117870 140200
rect 114840 139170 114863 140177
rect 114657 138170 114863 139170
rect 114657 137193 114680 138170
rect 111650 137170 114680 137193
rect 114840 137193 114863 138170
rect 117847 139170 117870 140177
rect 118030 140177 121060 140200
rect 118030 139170 118053 140177
rect 117847 138170 118053 139170
rect 117847 137193 117870 138170
rect 114840 137170 117870 137193
rect 118030 137193 118053 138170
rect 121037 139170 121060 140177
rect 121220 140177 124250 140200
rect 121220 139170 121243 140177
rect 121037 138170 121243 139170
rect 121037 137193 121060 138170
rect 118030 137170 121060 137193
rect 121220 137193 121243 138170
rect 124227 139170 124250 140177
rect 124410 140177 127440 140200
rect 124410 139170 124433 140177
rect 124227 138170 124433 139170
rect 124227 137193 124250 138170
rect 121220 137170 124250 137193
rect 124410 137193 124433 138170
rect 127417 139170 127440 140177
rect 127600 140177 130630 140200
rect 127600 139170 127623 140177
rect 127417 138170 127623 139170
rect 127417 137193 127440 138170
rect 124410 137170 127440 137193
rect 127600 137193 127623 138170
rect 130607 139170 130630 140177
rect 130790 140177 133820 140200
rect 130790 139170 130813 140177
rect 130607 138170 130813 139170
rect 130607 137193 130630 138170
rect 127600 137170 130630 137193
rect 130790 137193 130813 138170
rect 133797 139170 133820 140177
rect 133980 140177 137010 140200
rect 133980 139170 134003 140177
rect 133797 138170 134003 139170
rect 133797 137193 133820 138170
rect 130790 137170 133820 137193
rect 133980 137193 134003 138170
rect 136987 139170 137010 140177
rect 136987 138170 137170 139170
rect 136987 137193 137010 138170
rect 133980 137170 137010 137193
rect 10570 137010 11570 137170
rect 13760 137010 14760 137170
rect 16950 137010 17950 137170
rect 20140 137010 21140 137170
rect 23330 137010 24330 137170
rect 26520 137010 27520 137170
rect 29710 137010 30710 137170
rect 32900 137010 33900 137170
rect 36090 137010 37090 137170
rect 39280 137010 40280 137170
rect 42470 137010 43470 137170
rect 45660 137010 46660 137170
rect 48850 137010 49850 137170
rect 52040 137010 53040 137170
rect 55230 137010 56230 137170
rect 58420 137010 59420 137170
rect 61610 137010 62610 137170
rect 64800 137010 65800 137170
rect 67990 137010 68990 137170
rect 71180 137010 72180 137170
rect 74370 137010 75370 137170
rect 77560 137010 78560 137170
rect 80750 137010 81750 137170
rect 83940 137010 84940 137170
rect 87130 137010 88130 137170
rect 90320 137010 91320 137170
rect 93510 137010 94510 137170
rect 96700 137010 97700 137170
rect 99890 137010 100890 137170
rect 103080 137010 104080 137170
rect 106270 137010 107270 137170
rect 109460 137010 110460 137170
rect 112650 137010 113650 137170
rect 115840 137010 116840 137170
rect 119030 137010 120030 137170
rect 122220 137010 123220 137170
rect 125410 137010 126410 137170
rect 128600 137010 129600 137170
rect 131790 137010 132790 137170
rect 134980 137010 135980 137170
rect 9570 136987 12600 137010
rect 9570 134003 9593 136987
rect 12577 135980 12600 136987
rect 12760 136987 15790 137010
rect 12760 135980 12783 136987
rect 12577 134980 12783 135980
rect 12577 134003 12600 134980
rect 9570 133980 12600 134003
rect 12760 134003 12783 134980
rect 15767 135980 15790 136987
rect 15950 136987 18980 137010
rect 15950 135980 15973 136987
rect 15767 134980 15973 135980
rect 15767 134003 15790 134980
rect 12760 133980 15790 134003
rect 15950 134003 15973 134980
rect 18957 135980 18980 136987
rect 19140 136987 22170 137010
rect 19140 135980 19163 136987
rect 18957 134980 19163 135980
rect 18957 134003 18980 134980
rect 15950 133980 18980 134003
rect 19140 134003 19163 134980
rect 22147 135980 22170 136987
rect 22330 136987 25360 137010
rect 22330 135980 22353 136987
rect 22147 134980 22353 135980
rect 22147 134003 22170 134980
rect 19140 133980 22170 134003
rect 22330 134003 22353 134980
rect 25337 135980 25360 136987
rect 25520 136987 28550 137010
rect 25520 135980 25543 136987
rect 25337 134980 25543 135980
rect 25337 134003 25360 134980
rect 22330 133980 25360 134003
rect 25520 134003 25543 134980
rect 28527 135980 28550 136987
rect 28710 136987 31740 137010
rect 28710 135980 28733 136987
rect 28527 134980 28733 135980
rect 28527 134003 28550 134980
rect 25520 133980 28550 134003
rect 28710 134003 28733 134980
rect 31717 135980 31740 136987
rect 31900 136987 34930 137010
rect 31900 135980 31923 136987
rect 31717 134980 31923 135980
rect 31717 134003 31740 134980
rect 28710 133980 31740 134003
rect 31900 134003 31923 134980
rect 34907 135980 34930 136987
rect 35090 136987 38120 137010
rect 35090 135980 35113 136987
rect 34907 134980 35113 135980
rect 34907 134003 34930 134980
rect 31900 133980 34930 134003
rect 35090 134003 35113 134980
rect 38097 135980 38120 136987
rect 38280 136987 41310 137010
rect 38280 135980 38303 136987
rect 38097 134980 38303 135980
rect 38097 134003 38120 134980
rect 35090 133980 38120 134003
rect 38280 134003 38303 134980
rect 41287 135980 41310 136987
rect 41470 136987 44500 137010
rect 41470 135980 41493 136987
rect 41287 134980 41493 135980
rect 41287 134003 41310 134980
rect 38280 133980 41310 134003
rect 41470 134003 41493 134980
rect 44477 135980 44500 136987
rect 44660 136987 47690 137010
rect 44660 135980 44683 136987
rect 44477 134980 44683 135980
rect 44477 134003 44500 134980
rect 41470 133980 44500 134003
rect 44660 134003 44683 134980
rect 47667 135980 47690 136987
rect 47850 136987 50880 137010
rect 47850 135980 47873 136987
rect 47667 134980 47873 135980
rect 47667 134003 47690 134980
rect 44660 133980 47690 134003
rect 47850 134003 47873 134980
rect 50857 135980 50880 136987
rect 51040 136987 54070 137010
rect 51040 135980 51063 136987
rect 50857 134980 51063 135980
rect 50857 134003 50880 134980
rect 47850 133980 50880 134003
rect 51040 134003 51063 134980
rect 54047 135980 54070 136987
rect 54230 136987 57260 137010
rect 54230 135980 54253 136987
rect 54047 134980 54253 135980
rect 54047 134003 54070 134980
rect 51040 133980 54070 134003
rect 54230 134003 54253 134980
rect 57237 135980 57260 136987
rect 57420 136987 60450 137010
rect 57420 135980 57443 136987
rect 57237 134980 57443 135980
rect 57237 134003 57260 134980
rect 54230 133980 57260 134003
rect 57420 134003 57443 134980
rect 60427 135980 60450 136987
rect 60610 136987 63640 137010
rect 60610 135980 60633 136987
rect 60427 134980 60633 135980
rect 60427 134003 60450 134980
rect 57420 133980 60450 134003
rect 60610 134003 60633 134980
rect 63617 135980 63640 136987
rect 63800 136987 66830 137010
rect 63800 135980 63823 136987
rect 63617 134980 63823 135980
rect 63617 134003 63640 134980
rect 60610 133980 63640 134003
rect 63800 134003 63823 134980
rect 66807 135980 66830 136987
rect 66990 136987 70020 137010
rect 66990 135980 67013 136987
rect 66807 134980 67013 135980
rect 66807 134003 66830 134980
rect 63800 133980 66830 134003
rect 66990 134003 67013 134980
rect 69997 135980 70020 136987
rect 70180 136987 73210 137010
rect 70180 135980 70203 136987
rect 69997 134980 70203 135980
rect 69997 134003 70020 134980
rect 66990 133980 70020 134003
rect 70180 134003 70203 134980
rect 73187 135980 73210 136987
rect 73370 136987 76400 137010
rect 73370 135980 73393 136987
rect 73187 134980 73393 135980
rect 73187 134003 73210 134980
rect 70180 133980 73210 134003
rect 73370 134003 73393 134980
rect 76377 135980 76400 136987
rect 76560 136987 79590 137010
rect 76560 135980 76583 136987
rect 76377 134980 76583 135980
rect 76377 134003 76400 134980
rect 73370 133980 76400 134003
rect 76560 134003 76583 134980
rect 79567 135980 79590 136987
rect 79750 136987 82780 137010
rect 79750 135980 79773 136987
rect 79567 134980 79773 135980
rect 79567 134003 79590 134980
rect 76560 133980 79590 134003
rect 79750 134003 79773 134980
rect 82757 135980 82780 136987
rect 82940 136987 85970 137010
rect 82940 135980 82963 136987
rect 82757 134980 82963 135980
rect 82757 134003 82780 134980
rect 79750 133980 82780 134003
rect 82940 134003 82963 134980
rect 85947 135980 85970 136987
rect 86130 136987 89160 137010
rect 86130 135980 86153 136987
rect 85947 134980 86153 135980
rect 85947 134003 85970 134980
rect 82940 133980 85970 134003
rect 86130 134003 86153 134980
rect 89137 135980 89160 136987
rect 89320 136987 92350 137010
rect 89320 135980 89343 136987
rect 89137 134980 89343 135980
rect 89137 134003 89160 134980
rect 86130 133980 89160 134003
rect 89320 134003 89343 134980
rect 92327 135980 92350 136987
rect 92510 136987 95540 137010
rect 92510 135980 92533 136987
rect 92327 134980 92533 135980
rect 92327 134003 92350 134980
rect 89320 133980 92350 134003
rect 92510 134003 92533 134980
rect 95517 135980 95540 136987
rect 95700 136987 98730 137010
rect 95700 135980 95723 136987
rect 95517 134980 95723 135980
rect 95517 134003 95540 134980
rect 92510 133980 95540 134003
rect 95700 134003 95723 134980
rect 98707 135980 98730 136987
rect 98890 136987 101920 137010
rect 98890 135980 98913 136987
rect 98707 134980 98913 135980
rect 98707 134003 98730 134980
rect 95700 133980 98730 134003
rect 98890 134003 98913 134980
rect 101897 135980 101920 136987
rect 102080 136987 105110 137010
rect 102080 135980 102103 136987
rect 101897 134980 102103 135980
rect 101897 134003 101920 134980
rect 98890 133980 101920 134003
rect 102080 134003 102103 134980
rect 105087 135980 105110 136987
rect 105270 136987 108300 137010
rect 105270 135980 105293 136987
rect 105087 134980 105293 135980
rect 105087 134003 105110 134980
rect 102080 133980 105110 134003
rect 105270 134003 105293 134980
rect 108277 135980 108300 136987
rect 108460 136987 111490 137010
rect 108460 135980 108483 136987
rect 108277 134980 108483 135980
rect 108277 134003 108300 134980
rect 105270 133980 108300 134003
rect 108460 134003 108483 134980
rect 111467 135980 111490 136987
rect 111650 136987 114680 137010
rect 111650 135980 111673 136987
rect 111467 134980 111673 135980
rect 111467 134003 111490 134980
rect 108460 133980 111490 134003
rect 111650 134003 111673 134980
rect 114657 135980 114680 136987
rect 114840 136987 117870 137010
rect 114840 135980 114863 136987
rect 114657 134980 114863 135980
rect 114657 134003 114680 134980
rect 111650 133980 114680 134003
rect 114840 134003 114863 134980
rect 117847 135980 117870 136987
rect 118030 136987 121060 137010
rect 118030 135980 118053 136987
rect 117847 134980 118053 135980
rect 117847 134003 117870 134980
rect 114840 133980 117870 134003
rect 118030 134003 118053 134980
rect 121037 135980 121060 136987
rect 121220 136987 124250 137010
rect 121220 135980 121243 136987
rect 121037 134980 121243 135980
rect 121037 134003 121060 134980
rect 118030 133980 121060 134003
rect 121220 134003 121243 134980
rect 124227 135980 124250 136987
rect 124410 136987 127440 137010
rect 124410 135980 124433 136987
rect 124227 134980 124433 135980
rect 124227 134003 124250 134980
rect 121220 133980 124250 134003
rect 124410 134003 124433 134980
rect 127417 135980 127440 136987
rect 127600 136987 130630 137010
rect 127600 135980 127623 136987
rect 127417 134980 127623 135980
rect 127417 134003 127440 134980
rect 124410 133980 127440 134003
rect 127600 134003 127623 134980
rect 130607 135980 130630 136987
rect 130790 136987 133820 137010
rect 130790 135980 130813 136987
rect 130607 134980 130813 135980
rect 130607 134003 130630 134980
rect 127600 133980 130630 134003
rect 130790 134003 130813 134980
rect 133797 135980 133820 136987
rect 133980 136987 137010 137010
rect 133980 135980 134003 136987
rect 133797 134980 134003 135980
rect 133797 134003 133820 134980
rect 130790 133980 133820 134003
rect 133980 134003 134003 134980
rect 136987 135980 137010 136987
rect 136987 134980 137170 135980
rect 136987 134003 137010 134980
rect 133980 133980 137010 134003
rect 10570 133820 11570 133980
rect 13760 133820 14760 133980
rect 16950 133820 17950 133980
rect 20140 133820 21140 133980
rect 23330 133820 24330 133980
rect 26520 133820 27520 133980
rect 29710 133820 30710 133980
rect 32900 133820 33900 133980
rect 36090 133820 37090 133980
rect 39280 133820 40280 133980
rect 42470 133820 43470 133980
rect 45660 133820 46660 133980
rect 48850 133820 49850 133980
rect 52040 133820 53040 133980
rect 55230 133820 56230 133980
rect 58420 133820 59420 133980
rect 61610 133820 62610 133980
rect 64800 133820 65800 133980
rect 67990 133820 68990 133980
rect 71180 133820 72180 133980
rect 74370 133820 75370 133980
rect 77560 133820 78560 133980
rect 80750 133820 81750 133980
rect 83940 133820 84940 133980
rect 87130 133820 88130 133980
rect 90320 133820 91320 133980
rect 93510 133820 94510 133980
rect 96700 133820 97700 133980
rect 99890 133820 100890 133980
rect 103080 133820 104080 133980
rect 106270 133820 107270 133980
rect 109460 133820 110460 133980
rect 112650 133820 113650 133980
rect 115840 133820 116840 133980
rect 119030 133820 120030 133980
rect 122220 133820 123220 133980
rect 125410 133820 126410 133980
rect 128600 133820 129600 133980
rect 131790 133820 132790 133980
rect 134980 133820 135980 133980
rect 9570 133797 12600 133820
rect 9570 130813 9593 133797
rect 12577 132790 12600 133797
rect 12760 133797 15790 133820
rect 12760 132790 12783 133797
rect 12577 131790 12783 132790
rect 12577 130813 12600 131790
rect 9570 130790 12600 130813
rect 12760 130813 12783 131790
rect 15767 132790 15790 133797
rect 15950 133797 18980 133820
rect 15950 132790 15973 133797
rect 15767 131790 15973 132790
rect 15767 130813 15790 131790
rect 12760 130790 15790 130813
rect 15950 130813 15973 131790
rect 18957 132790 18980 133797
rect 19140 133797 22170 133820
rect 19140 132790 19163 133797
rect 18957 131790 19163 132790
rect 18957 130813 18980 131790
rect 15950 130790 18980 130813
rect 19140 130813 19163 131790
rect 22147 132790 22170 133797
rect 22330 133797 25360 133820
rect 22330 132790 22353 133797
rect 22147 131790 22353 132790
rect 22147 130813 22170 131790
rect 19140 130790 22170 130813
rect 22330 130813 22353 131790
rect 25337 132790 25360 133797
rect 25520 133797 28550 133820
rect 25520 132790 25543 133797
rect 25337 131790 25543 132790
rect 25337 130813 25360 131790
rect 22330 130790 25360 130813
rect 25520 130813 25543 131790
rect 28527 132790 28550 133797
rect 28710 133797 31740 133820
rect 28710 132790 28733 133797
rect 28527 131790 28733 132790
rect 28527 130813 28550 131790
rect 25520 130790 28550 130813
rect 28710 130813 28733 131790
rect 31717 132790 31740 133797
rect 31900 133797 34930 133820
rect 31900 132790 31923 133797
rect 31717 131790 31923 132790
rect 31717 130813 31740 131790
rect 28710 130790 31740 130813
rect 31900 130813 31923 131790
rect 34907 132790 34930 133797
rect 35090 133797 38120 133820
rect 35090 132790 35113 133797
rect 34907 131790 35113 132790
rect 34907 130813 34930 131790
rect 31900 130790 34930 130813
rect 35090 130813 35113 131790
rect 38097 132790 38120 133797
rect 38280 133797 41310 133820
rect 38280 132790 38303 133797
rect 38097 131790 38303 132790
rect 38097 130813 38120 131790
rect 35090 130790 38120 130813
rect 38280 130813 38303 131790
rect 41287 132790 41310 133797
rect 41470 133797 44500 133820
rect 41470 132790 41493 133797
rect 41287 131790 41493 132790
rect 41287 130813 41310 131790
rect 38280 130790 41310 130813
rect 41470 130813 41493 131790
rect 44477 132790 44500 133797
rect 44660 133797 47690 133820
rect 44660 132790 44683 133797
rect 44477 131790 44683 132790
rect 44477 130813 44500 131790
rect 41470 130790 44500 130813
rect 44660 130813 44683 131790
rect 47667 132790 47690 133797
rect 47850 133797 50880 133820
rect 47850 132790 47873 133797
rect 47667 131790 47873 132790
rect 47667 130813 47690 131790
rect 44660 130790 47690 130813
rect 47850 130813 47873 131790
rect 50857 132790 50880 133797
rect 51040 133797 54070 133820
rect 51040 132790 51063 133797
rect 50857 131790 51063 132790
rect 50857 130813 50880 131790
rect 47850 130790 50880 130813
rect 51040 130813 51063 131790
rect 54047 132790 54070 133797
rect 54230 133797 57260 133820
rect 54230 132790 54253 133797
rect 54047 131790 54253 132790
rect 54047 130813 54070 131790
rect 51040 130790 54070 130813
rect 54230 130813 54253 131790
rect 57237 132790 57260 133797
rect 57420 133797 60450 133820
rect 57420 132790 57443 133797
rect 57237 131790 57443 132790
rect 57237 130813 57260 131790
rect 54230 130790 57260 130813
rect 57420 130813 57443 131790
rect 60427 132790 60450 133797
rect 60610 133797 63640 133820
rect 60610 132790 60633 133797
rect 60427 131790 60633 132790
rect 60427 130813 60450 131790
rect 57420 130790 60450 130813
rect 60610 130813 60633 131790
rect 63617 132790 63640 133797
rect 63800 133797 66830 133820
rect 63800 132790 63823 133797
rect 63617 131790 63823 132790
rect 63617 130813 63640 131790
rect 60610 130790 63640 130813
rect 63800 130813 63823 131790
rect 66807 132790 66830 133797
rect 66990 133797 70020 133820
rect 66990 132790 67013 133797
rect 66807 131790 67013 132790
rect 66807 130813 66830 131790
rect 63800 130790 66830 130813
rect 66990 130813 67013 131790
rect 69997 132790 70020 133797
rect 70180 133797 73210 133820
rect 70180 132790 70203 133797
rect 69997 131790 70203 132790
rect 69997 130813 70020 131790
rect 66990 130790 70020 130813
rect 70180 130813 70203 131790
rect 73187 132790 73210 133797
rect 73370 133797 76400 133820
rect 73370 132790 73393 133797
rect 73187 131790 73393 132790
rect 73187 130813 73210 131790
rect 70180 130790 73210 130813
rect 73370 130813 73393 131790
rect 76377 132790 76400 133797
rect 76560 133797 79590 133820
rect 76560 132790 76583 133797
rect 76377 131790 76583 132790
rect 76377 130813 76400 131790
rect 73370 130790 76400 130813
rect 76560 130813 76583 131790
rect 79567 132790 79590 133797
rect 79750 133797 82780 133820
rect 79750 132790 79773 133797
rect 79567 131790 79773 132790
rect 79567 130813 79590 131790
rect 76560 130790 79590 130813
rect 79750 130813 79773 131790
rect 82757 132790 82780 133797
rect 82940 133797 85970 133820
rect 82940 132790 82963 133797
rect 82757 131790 82963 132790
rect 82757 130813 82780 131790
rect 79750 130790 82780 130813
rect 82940 130813 82963 131790
rect 85947 132790 85970 133797
rect 86130 133797 89160 133820
rect 86130 132790 86153 133797
rect 85947 131790 86153 132790
rect 85947 130813 85970 131790
rect 82940 130790 85970 130813
rect 86130 130813 86153 131790
rect 89137 132790 89160 133797
rect 89320 133797 92350 133820
rect 89320 132790 89343 133797
rect 89137 131790 89343 132790
rect 89137 130813 89160 131790
rect 86130 130790 89160 130813
rect 89320 130813 89343 131790
rect 92327 132790 92350 133797
rect 92510 133797 95540 133820
rect 92510 132790 92533 133797
rect 92327 131790 92533 132790
rect 92327 130813 92350 131790
rect 89320 130790 92350 130813
rect 92510 130813 92533 131790
rect 95517 132790 95540 133797
rect 95700 133797 98730 133820
rect 95700 132790 95723 133797
rect 95517 131790 95723 132790
rect 95517 130813 95540 131790
rect 92510 130790 95540 130813
rect 95700 130813 95723 131790
rect 98707 132790 98730 133797
rect 98890 133797 101920 133820
rect 98890 132790 98913 133797
rect 98707 131790 98913 132790
rect 98707 130813 98730 131790
rect 95700 130790 98730 130813
rect 98890 130813 98913 131790
rect 101897 132790 101920 133797
rect 102080 133797 105110 133820
rect 102080 132790 102103 133797
rect 101897 131790 102103 132790
rect 101897 130813 101920 131790
rect 98890 130790 101920 130813
rect 102080 130813 102103 131790
rect 105087 132790 105110 133797
rect 105270 133797 108300 133820
rect 105270 132790 105293 133797
rect 105087 131790 105293 132790
rect 105087 130813 105110 131790
rect 102080 130790 105110 130813
rect 105270 130813 105293 131790
rect 108277 132790 108300 133797
rect 108460 133797 111490 133820
rect 108460 132790 108483 133797
rect 108277 131790 108483 132790
rect 108277 130813 108300 131790
rect 105270 130790 108300 130813
rect 108460 130813 108483 131790
rect 111467 132790 111490 133797
rect 111650 133797 114680 133820
rect 111650 132790 111673 133797
rect 111467 131790 111673 132790
rect 111467 130813 111490 131790
rect 108460 130790 111490 130813
rect 111650 130813 111673 131790
rect 114657 132790 114680 133797
rect 114840 133797 117870 133820
rect 114840 132790 114863 133797
rect 114657 131790 114863 132790
rect 114657 130813 114680 131790
rect 111650 130790 114680 130813
rect 114840 130813 114863 131790
rect 117847 132790 117870 133797
rect 118030 133797 121060 133820
rect 118030 132790 118053 133797
rect 117847 131790 118053 132790
rect 117847 130813 117870 131790
rect 114840 130790 117870 130813
rect 118030 130813 118053 131790
rect 121037 132790 121060 133797
rect 121220 133797 124250 133820
rect 121220 132790 121243 133797
rect 121037 131790 121243 132790
rect 121037 130813 121060 131790
rect 118030 130790 121060 130813
rect 121220 130813 121243 131790
rect 124227 132790 124250 133797
rect 124410 133797 127440 133820
rect 124410 132790 124433 133797
rect 124227 131790 124433 132790
rect 124227 130813 124250 131790
rect 121220 130790 124250 130813
rect 124410 130813 124433 131790
rect 127417 132790 127440 133797
rect 127600 133797 130630 133820
rect 127600 132790 127623 133797
rect 127417 131790 127623 132790
rect 127417 130813 127440 131790
rect 124410 130790 127440 130813
rect 127600 130813 127623 131790
rect 130607 132790 130630 133797
rect 130790 133797 133820 133820
rect 130790 132790 130813 133797
rect 130607 131790 130813 132790
rect 130607 130813 130630 131790
rect 127600 130790 130630 130813
rect 130790 130813 130813 131790
rect 133797 132790 133820 133797
rect 133980 133797 137010 133820
rect 133980 132790 134003 133797
rect 133797 131790 134003 132790
rect 133797 130813 133820 131790
rect 130790 130790 133820 130813
rect 133980 130813 134003 131790
rect 136987 132790 137010 133797
rect 136987 131790 137170 132790
rect 136987 130813 137010 131790
rect 133980 130790 137010 130813
rect 10570 130630 11570 130790
rect 13760 130630 14760 130790
rect 16950 130630 17950 130790
rect 20140 130630 21140 130790
rect 23330 130630 24330 130790
rect 26520 130630 27520 130790
rect 29710 130630 30710 130790
rect 32900 130630 33900 130790
rect 36090 130630 37090 130790
rect 39280 130630 40280 130790
rect 42470 130630 43470 130790
rect 45660 130630 46660 130790
rect 48850 130630 49850 130790
rect 52040 130630 53040 130790
rect 55230 130630 56230 130790
rect 58420 130630 59420 130790
rect 61610 130630 62610 130790
rect 64800 130630 65800 130790
rect 67990 130630 68990 130790
rect 71180 130630 72180 130790
rect 74370 130630 75370 130790
rect 77560 130630 78560 130790
rect 80750 130630 81750 130790
rect 83940 130630 84940 130790
rect 87130 130630 88130 130790
rect 90320 130630 91320 130790
rect 93510 130630 94510 130790
rect 96700 130630 97700 130790
rect 99890 130630 100890 130790
rect 103080 130630 104080 130790
rect 106270 130630 107270 130790
rect 109460 130630 110460 130790
rect 112650 130630 113650 130790
rect 115840 130630 116840 130790
rect 119030 130630 120030 130790
rect 122220 130630 123220 130790
rect 125410 130630 126410 130790
rect 128600 130630 129600 130790
rect 131790 130630 132790 130790
rect 134980 130630 135980 130790
rect 9570 130607 12600 130630
rect 9570 127623 9593 130607
rect 12577 129600 12600 130607
rect 12760 130607 15790 130630
rect 12760 129600 12783 130607
rect 12577 128600 12783 129600
rect 12577 127623 12600 128600
rect 9570 127600 12600 127623
rect 12760 127623 12783 128600
rect 15767 129600 15790 130607
rect 15950 130607 18980 130630
rect 15950 129600 15973 130607
rect 15767 128600 15973 129600
rect 15767 127623 15790 128600
rect 12760 127600 15790 127623
rect 15950 127623 15973 128600
rect 18957 129600 18980 130607
rect 19140 130607 22170 130630
rect 19140 129600 19163 130607
rect 18957 128600 19163 129600
rect 18957 127623 18980 128600
rect 15950 127600 18980 127623
rect 19140 127623 19163 128600
rect 22147 129600 22170 130607
rect 22330 130607 25360 130630
rect 22330 129600 22353 130607
rect 22147 128600 22353 129600
rect 22147 127623 22170 128600
rect 19140 127600 22170 127623
rect 22330 127623 22353 128600
rect 25337 129600 25360 130607
rect 25520 130607 28550 130630
rect 25520 129600 25543 130607
rect 25337 128600 25543 129600
rect 25337 127623 25360 128600
rect 22330 127600 25360 127623
rect 25520 127623 25543 128600
rect 28527 129600 28550 130607
rect 28710 130607 31740 130630
rect 28710 129600 28733 130607
rect 28527 128600 28733 129600
rect 28527 127623 28550 128600
rect 25520 127600 28550 127623
rect 28710 127623 28733 128600
rect 31717 129600 31740 130607
rect 31900 130607 34930 130630
rect 31900 129600 31923 130607
rect 31717 128600 31923 129600
rect 31717 127623 31740 128600
rect 28710 127600 31740 127623
rect 31900 127623 31923 128600
rect 34907 129600 34930 130607
rect 35090 130607 38120 130630
rect 35090 129600 35113 130607
rect 34907 128600 35113 129600
rect 34907 127623 34930 128600
rect 31900 127600 34930 127623
rect 35090 127623 35113 128600
rect 38097 129600 38120 130607
rect 38280 130607 41310 130630
rect 38280 129600 38303 130607
rect 38097 128600 38303 129600
rect 38097 127623 38120 128600
rect 35090 127600 38120 127623
rect 38280 127623 38303 128600
rect 41287 129600 41310 130607
rect 41470 130607 44500 130630
rect 41470 129600 41493 130607
rect 41287 128600 41493 129600
rect 41287 127623 41310 128600
rect 38280 127600 41310 127623
rect 41470 127623 41493 128600
rect 44477 129600 44500 130607
rect 44660 130607 47690 130630
rect 44660 129600 44683 130607
rect 44477 128600 44683 129600
rect 44477 127623 44500 128600
rect 41470 127600 44500 127623
rect 44660 127623 44683 128600
rect 47667 129600 47690 130607
rect 47850 130607 50880 130630
rect 47850 129600 47873 130607
rect 47667 128600 47873 129600
rect 47667 127623 47690 128600
rect 44660 127600 47690 127623
rect 47850 127623 47873 128600
rect 50857 129600 50880 130607
rect 51040 130607 54070 130630
rect 51040 129600 51063 130607
rect 50857 128600 51063 129600
rect 50857 127623 50880 128600
rect 47850 127600 50880 127623
rect 51040 127623 51063 128600
rect 54047 129600 54070 130607
rect 54230 130607 57260 130630
rect 54230 129600 54253 130607
rect 54047 128600 54253 129600
rect 54047 127623 54070 128600
rect 51040 127600 54070 127623
rect 54230 127623 54253 128600
rect 57237 129600 57260 130607
rect 57420 130607 60450 130630
rect 57420 129600 57443 130607
rect 57237 128600 57443 129600
rect 57237 127623 57260 128600
rect 54230 127600 57260 127623
rect 57420 127623 57443 128600
rect 60427 129600 60450 130607
rect 60610 130607 63640 130630
rect 60610 129600 60633 130607
rect 60427 128600 60633 129600
rect 60427 127623 60450 128600
rect 57420 127600 60450 127623
rect 60610 127623 60633 128600
rect 63617 129600 63640 130607
rect 63800 130607 66830 130630
rect 63800 129600 63823 130607
rect 63617 128600 63823 129600
rect 63617 127623 63640 128600
rect 60610 127600 63640 127623
rect 63800 127623 63823 128600
rect 66807 129600 66830 130607
rect 66990 130607 70020 130630
rect 66990 129600 67013 130607
rect 66807 128600 67013 129600
rect 66807 127623 66830 128600
rect 63800 127600 66830 127623
rect 66990 127623 67013 128600
rect 69997 129600 70020 130607
rect 70180 130607 73210 130630
rect 70180 129600 70203 130607
rect 69997 128600 70203 129600
rect 69997 127623 70020 128600
rect 66990 127600 70020 127623
rect 70180 127623 70203 128600
rect 73187 129600 73210 130607
rect 73370 130607 76400 130630
rect 73370 129600 73393 130607
rect 73187 128600 73393 129600
rect 73187 127623 73210 128600
rect 70180 127600 73210 127623
rect 73370 127623 73393 128600
rect 76377 129600 76400 130607
rect 76560 130607 79590 130630
rect 76560 129600 76583 130607
rect 76377 128600 76583 129600
rect 76377 127623 76400 128600
rect 73370 127600 76400 127623
rect 76560 127623 76583 128600
rect 79567 129600 79590 130607
rect 79750 130607 82780 130630
rect 79750 129600 79773 130607
rect 79567 128600 79773 129600
rect 79567 127623 79590 128600
rect 76560 127600 79590 127623
rect 79750 127623 79773 128600
rect 82757 129600 82780 130607
rect 82940 130607 85970 130630
rect 82940 129600 82963 130607
rect 82757 128600 82963 129600
rect 82757 127623 82780 128600
rect 79750 127600 82780 127623
rect 82940 127623 82963 128600
rect 85947 129600 85970 130607
rect 86130 130607 89160 130630
rect 86130 129600 86153 130607
rect 85947 128600 86153 129600
rect 85947 127623 85970 128600
rect 82940 127600 85970 127623
rect 86130 127623 86153 128600
rect 89137 129600 89160 130607
rect 89320 130607 92350 130630
rect 89320 129600 89343 130607
rect 89137 128600 89343 129600
rect 89137 127623 89160 128600
rect 86130 127600 89160 127623
rect 89320 127623 89343 128600
rect 92327 129600 92350 130607
rect 92510 130607 95540 130630
rect 92510 129600 92533 130607
rect 92327 128600 92533 129600
rect 92327 127623 92350 128600
rect 89320 127600 92350 127623
rect 92510 127623 92533 128600
rect 95517 129600 95540 130607
rect 95700 130607 98730 130630
rect 95700 129600 95723 130607
rect 95517 128600 95723 129600
rect 95517 127623 95540 128600
rect 92510 127600 95540 127623
rect 95700 127623 95723 128600
rect 98707 129600 98730 130607
rect 98890 130607 101920 130630
rect 98890 129600 98913 130607
rect 98707 128600 98913 129600
rect 98707 127623 98730 128600
rect 95700 127600 98730 127623
rect 98890 127623 98913 128600
rect 101897 129600 101920 130607
rect 102080 130607 105110 130630
rect 102080 129600 102103 130607
rect 101897 128600 102103 129600
rect 101897 127623 101920 128600
rect 98890 127600 101920 127623
rect 102080 127623 102103 128600
rect 105087 129600 105110 130607
rect 105270 130607 108300 130630
rect 105270 129600 105293 130607
rect 105087 128600 105293 129600
rect 105087 127623 105110 128600
rect 102080 127600 105110 127623
rect 105270 127623 105293 128600
rect 108277 129600 108300 130607
rect 108460 130607 111490 130630
rect 108460 129600 108483 130607
rect 108277 128600 108483 129600
rect 108277 127623 108300 128600
rect 105270 127600 108300 127623
rect 108460 127623 108483 128600
rect 111467 129600 111490 130607
rect 111650 130607 114680 130630
rect 111650 129600 111673 130607
rect 111467 128600 111673 129600
rect 111467 127623 111490 128600
rect 108460 127600 111490 127623
rect 111650 127623 111673 128600
rect 114657 129600 114680 130607
rect 114840 130607 117870 130630
rect 114840 129600 114863 130607
rect 114657 128600 114863 129600
rect 114657 127623 114680 128600
rect 111650 127600 114680 127623
rect 114840 127623 114863 128600
rect 117847 129600 117870 130607
rect 118030 130607 121060 130630
rect 118030 129600 118053 130607
rect 117847 128600 118053 129600
rect 117847 127623 117870 128600
rect 114840 127600 117870 127623
rect 118030 127623 118053 128600
rect 121037 129600 121060 130607
rect 121220 130607 124250 130630
rect 121220 129600 121243 130607
rect 121037 128600 121243 129600
rect 121037 127623 121060 128600
rect 118030 127600 121060 127623
rect 121220 127623 121243 128600
rect 124227 129600 124250 130607
rect 124410 130607 127440 130630
rect 124410 129600 124433 130607
rect 124227 128600 124433 129600
rect 124227 127623 124250 128600
rect 121220 127600 124250 127623
rect 124410 127623 124433 128600
rect 127417 129600 127440 130607
rect 127600 130607 130630 130630
rect 127600 129600 127623 130607
rect 127417 128600 127623 129600
rect 127417 127623 127440 128600
rect 124410 127600 127440 127623
rect 127600 127623 127623 128600
rect 130607 129600 130630 130607
rect 130790 130607 133820 130630
rect 130790 129600 130813 130607
rect 130607 128600 130813 129600
rect 130607 127623 130630 128600
rect 127600 127600 130630 127623
rect 130790 127623 130813 128600
rect 133797 129600 133820 130607
rect 133980 130607 137010 130630
rect 133980 129600 134003 130607
rect 133797 128600 134003 129600
rect 133797 127623 133820 128600
rect 130790 127600 133820 127623
rect 133980 127623 134003 128600
rect 136987 129600 137010 130607
rect 136987 128600 137170 129600
rect 136987 127623 137010 128600
rect 133980 127600 137010 127623
rect 10570 127440 11570 127600
rect 13760 127440 14760 127600
rect 16950 127440 17950 127600
rect 20140 127440 21140 127600
rect 23330 127440 24330 127600
rect 26520 127440 27520 127600
rect 29710 127440 30710 127600
rect 32900 127440 33900 127600
rect 36090 127440 37090 127600
rect 39280 127440 40280 127600
rect 42470 127440 43470 127600
rect 45660 127440 46660 127600
rect 48850 127440 49850 127600
rect 52040 127440 53040 127600
rect 55230 127440 56230 127600
rect 58420 127440 59420 127600
rect 61610 127440 62610 127600
rect 64800 127440 65800 127600
rect 67990 127440 68990 127600
rect 71180 127440 72180 127600
rect 74370 127440 75370 127600
rect 77560 127440 78560 127600
rect 80750 127440 81750 127600
rect 83940 127440 84940 127600
rect 87130 127440 88130 127600
rect 90320 127440 91320 127600
rect 93510 127440 94510 127600
rect 96700 127440 97700 127600
rect 99890 127440 100890 127600
rect 103080 127440 104080 127600
rect 106270 127440 107270 127600
rect 109460 127440 110460 127600
rect 112650 127440 113650 127600
rect 115840 127440 116840 127600
rect 119030 127440 120030 127600
rect 122220 127440 123220 127600
rect 125410 127440 126410 127600
rect 128600 127440 129600 127600
rect 131790 127440 132790 127600
rect 134980 127440 135980 127600
rect 9570 127417 12600 127440
rect 9570 124433 9593 127417
rect 12577 126410 12600 127417
rect 12760 127417 15790 127440
rect 12760 126410 12783 127417
rect 12577 125410 12783 126410
rect 12577 124433 12600 125410
rect 9570 124410 12600 124433
rect 12760 124433 12783 125410
rect 15767 126410 15790 127417
rect 15950 127417 18980 127440
rect 15950 126410 15973 127417
rect 15767 125410 15973 126410
rect 15767 124433 15790 125410
rect 12760 124410 15790 124433
rect 15950 124433 15973 125410
rect 18957 126410 18980 127417
rect 19140 127417 22170 127440
rect 19140 126410 19163 127417
rect 18957 125410 19163 126410
rect 18957 124433 18980 125410
rect 15950 124410 18980 124433
rect 19140 124433 19163 125410
rect 22147 126410 22170 127417
rect 22330 127417 25360 127440
rect 22330 126410 22353 127417
rect 22147 125410 22353 126410
rect 22147 124433 22170 125410
rect 19140 124410 22170 124433
rect 22330 124433 22353 125410
rect 25337 126410 25360 127417
rect 25520 127417 28550 127440
rect 25520 126410 25543 127417
rect 25337 125410 25543 126410
rect 25337 124433 25360 125410
rect 22330 124410 25360 124433
rect 25520 124433 25543 125410
rect 28527 126410 28550 127417
rect 28710 127417 31740 127440
rect 28710 126410 28733 127417
rect 28527 125410 28733 126410
rect 28527 124433 28550 125410
rect 25520 124410 28550 124433
rect 28710 124433 28733 125410
rect 31717 126410 31740 127417
rect 31900 127417 34930 127440
rect 31900 126410 31923 127417
rect 31717 125410 31923 126410
rect 31717 124433 31740 125410
rect 28710 124410 31740 124433
rect 31900 124433 31923 125410
rect 34907 126410 34930 127417
rect 35090 127417 38120 127440
rect 35090 126410 35113 127417
rect 34907 125410 35113 126410
rect 34907 124433 34930 125410
rect 31900 124410 34930 124433
rect 35090 124433 35113 125410
rect 38097 126410 38120 127417
rect 38280 127417 41310 127440
rect 38280 126410 38303 127417
rect 38097 125410 38303 126410
rect 38097 124433 38120 125410
rect 35090 124410 38120 124433
rect 38280 124433 38303 125410
rect 41287 126410 41310 127417
rect 41470 127417 44500 127440
rect 41470 126410 41493 127417
rect 41287 125410 41493 126410
rect 41287 124433 41310 125410
rect 38280 124410 41310 124433
rect 41470 124433 41493 125410
rect 44477 126410 44500 127417
rect 44660 127417 47690 127440
rect 44660 126410 44683 127417
rect 44477 125410 44683 126410
rect 44477 124433 44500 125410
rect 41470 124410 44500 124433
rect 44660 124433 44683 125410
rect 47667 126410 47690 127417
rect 47850 127417 50880 127440
rect 47850 126410 47873 127417
rect 47667 125410 47873 126410
rect 47667 124433 47690 125410
rect 44660 124410 47690 124433
rect 47850 124433 47873 125410
rect 50857 126410 50880 127417
rect 51040 127417 54070 127440
rect 51040 126410 51063 127417
rect 50857 125410 51063 126410
rect 50857 124433 50880 125410
rect 47850 124410 50880 124433
rect 51040 124433 51063 125410
rect 54047 126410 54070 127417
rect 54230 127417 57260 127440
rect 54230 126410 54253 127417
rect 54047 125410 54253 126410
rect 54047 124433 54070 125410
rect 51040 124410 54070 124433
rect 54230 124433 54253 125410
rect 57237 126410 57260 127417
rect 57420 127417 60450 127440
rect 57420 126410 57443 127417
rect 57237 125410 57443 126410
rect 57237 124433 57260 125410
rect 54230 124410 57260 124433
rect 57420 124433 57443 125410
rect 60427 126410 60450 127417
rect 60610 127417 63640 127440
rect 60610 126410 60633 127417
rect 60427 125410 60633 126410
rect 60427 124433 60450 125410
rect 57420 124410 60450 124433
rect 60610 124433 60633 125410
rect 63617 126410 63640 127417
rect 63800 127417 66830 127440
rect 63800 126410 63823 127417
rect 63617 125410 63823 126410
rect 63617 124433 63640 125410
rect 60610 124410 63640 124433
rect 63800 124433 63823 125410
rect 66807 126410 66830 127417
rect 66990 127417 70020 127440
rect 66990 126410 67013 127417
rect 66807 125410 67013 126410
rect 66807 124433 66830 125410
rect 63800 124410 66830 124433
rect 66990 124433 67013 125410
rect 69997 126410 70020 127417
rect 70180 127417 73210 127440
rect 70180 126410 70203 127417
rect 69997 125410 70203 126410
rect 69997 124433 70020 125410
rect 66990 124410 70020 124433
rect 70180 124433 70203 125410
rect 73187 126410 73210 127417
rect 73370 127417 76400 127440
rect 73370 126410 73393 127417
rect 73187 125410 73393 126410
rect 73187 124433 73210 125410
rect 70180 124410 73210 124433
rect 73370 124433 73393 125410
rect 76377 126410 76400 127417
rect 76560 127417 79590 127440
rect 76560 126410 76583 127417
rect 76377 125410 76583 126410
rect 76377 124433 76400 125410
rect 73370 124410 76400 124433
rect 76560 124433 76583 125410
rect 79567 126410 79590 127417
rect 79750 127417 82780 127440
rect 79750 126410 79773 127417
rect 79567 125410 79773 126410
rect 79567 124433 79590 125410
rect 76560 124410 79590 124433
rect 79750 124433 79773 125410
rect 82757 126410 82780 127417
rect 82940 127417 85970 127440
rect 82940 126410 82963 127417
rect 82757 125410 82963 126410
rect 82757 124433 82780 125410
rect 79750 124410 82780 124433
rect 82940 124433 82963 125410
rect 85947 126410 85970 127417
rect 86130 127417 89160 127440
rect 86130 126410 86153 127417
rect 85947 125410 86153 126410
rect 85947 124433 85970 125410
rect 82940 124410 85970 124433
rect 86130 124433 86153 125410
rect 89137 126410 89160 127417
rect 89320 127417 92350 127440
rect 89320 126410 89343 127417
rect 89137 125410 89343 126410
rect 89137 124433 89160 125410
rect 86130 124410 89160 124433
rect 89320 124433 89343 125410
rect 92327 126410 92350 127417
rect 92510 127417 95540 127440
rect 92510 126410 92533 127417
rect 92327 125410 92533 126410
rect 92327 124433 92350 125410
rect 89320 124410 92350 124433
rect 92510 124433 92533 125410
rect 95517 126410 95540 127417
rect 95700 127417 98730 127440
rect 95700 126410 95723 127417
rect 95517 125410 95723 126410
rect 95517 124433 95540 125410
rect 92510 124410 95540 124433
rect 95700 124433 95723 125410
rect 98707 126410 98730 127417
rect 98890 127417 101920 127440
rect 98890 126410 98913 127417
rect 98707 125410 98913 126410
rect 98707 124433 98730 125410
rect 95700 124410 98730 124433
rect 98890 124433 98913 125410
rect 101897 126410 101920 127417
rect 102080 127417 105110 127440
rect 102080 126410 102103 127417
rect 101897 125410 102103 126410
rect 101897 124433 101920 125410
rect 98890 124410 101920 124433
rect 102080 124433 102103 125410
rect 105087 126410 105110 127417
rect 105270 127417 108300 127440
rect 105270 126410 105293 127417
rect 105087 125410 105293 126410
rect 105087 124433 105110 125410
rect 102080 124410 105110 124433
rect 105270 124433 105293 125410
rect 108277 126410 108300 127417
rect 108460 127417 111490 127440
rect 108460 126410 108483 127417
rect 108277 125410 108483 126410
rect 108277 124433 108300 125410
rect 105270 124410 108300 124433
rect 108460 124433 108483 125410
rect 111467 126410 111490 127417
rect 111650 127417 114680 127440
rect 111650 126410 111673 127417
rect 111467 125410 111673 126410
rect 111467 124433 111490 125410
rect 108460 124410 111490 124433
rect 111650 124433 111673 125410
rect 114657 126410 114680 127417
rect 114840 127417 117870 127440
rect 114840 126410 114863 127417
rect 114657 125410 114863 126410
rect 114657 124433 114680 125410
rect 111650 124410 114680 124433
rect 114840 124433 114863 125410
rect 117847 126410 117870 127417
rect 118030 127417 121060 127440
rect 118030 126410 118053 127417
rect 117847 125410 118053 126410
rect 117847 124433 117870 125410
rect 114840 124410 117870 124433
rect 118030 124433 118053 125410
rect 121037 126410 121060 127417
rect 121220 127417 124250 127440
rect 121220 126410 121243 127417
rect 121037 125410 121243 126410
rect 121037 124433 121060 125410
rect 118030 124410 121060 124433
rect 121220 124433 121243 125410
rect 124227 126410 124250 127417
rect 124410 127417 127440 127440
rect 124410 126410 124433 127417
rect 124227 125410 124433 126410
rect 124227 124433 124250 125410
rect 121220 124410 124250 124433
rect 124410 124433 124433 125410
rect 127417 126410 127440 127417
rect 127600 127417 130630 127440
rect 127600 126410 127623 127417
rect 127417 125410 127623 126410
rect 127417 124433 127440 125410
rect 124410 124410 127440 124433
rect 127600 124433 127623 125410
rect 130607 126410 130630 127417
rect 130790 127417 133820 127440
rect 130790 126410 130813 127417
rect 130607 125410 130813 126410
rect 130607 124433 130630 125410
rect 127600 124410 130630 124433
rect 130790 124433 130813 125410
rect 133797 126410 133820 127417
rect 133980 127417 137010 127440
rect 133980 126410 134003 127417
rect 133797 125410 134003 126410
rect 133797 124433 133820 125410
rect 130790 124410 133820 124433
rect 133980 124433 134003 125410
rect 136987 126410 137010 127417
rect 136987 125410 137170 126410
rect 136987 124433 137010 125410
rect 133980 124410 137010 124433
rect 10570 124250 11570 124410
rect 13760 124250 14760 124410
rect 16950 124250 17950 124410
rect 20140 124250 21140 124410
rect 23330 124250 24330 124410
rect 26520 124250 27520 124410
rect 29710 124250 30710 124410
rect 32900 124250 33900 124410
rect 36090 124250 37090 124410
rect 39280 124250 40280 124410
rect 42470 124250 43470 124410
rect 45660 124250 46660 124410
rect 48850 124250 49850 124410
rect 52040 124250 53040 124410
rect 55230 124250 56230 124410
rect 58420 124250 59420 124410
rect 61610 124250 62610 124410
rect 64800 124250 65800 124410
rect 67990 124250 68990 124410
rect 71180 124250 72180 124410
rect 74370 124250 75370 124410
rect 77560 124250 78560 124410
rect 80750 124250 81750 124410
rect 83940 124250 84940 124410
rect 87130 124250 88130 124410
rect 90320 124250 91320 124410
rect 93510 124250 94510 124410
rect 96700 124250 97700 124410
rect 99890 124250 100890 124410
rect 103080 124250 104080 124410
rect 106270 124250 107270 124410
rect 109460 124250 110460 124410
rect 112650 124250 113650 124410
rect 115840 124250 116840 124410
rect 119030 124250 120030 124410
rect 122220 124250 123220 124410
rect 125410 124250 126410 124410
rect 128600 124250 129600 124410
rect 131790 124250 132790 124410
rect 134980 124250 135980 124410
rect 0 121260 9370 121310
rect 9570 124227 12600 124250
rect 9570 121243 9593 124227
rect 12577 123220 12600 124227
rect 12760 124227 15790 124250
rect 12760 123220 12783 124227
rect 12577 122220 12783 123220
rect 12577 121243 12600 122220
rect 9570 121220 12600 121243
rect 12760 121243 12783 122220
rect 15767 123220 15790 124227
rect 15950 124227 18980 124250
rect 15950 123220 15973 124227
rect 15767 122220 15973 123220
rect 15767 121243 15790 122220
rect 12760 121220 15790 121243
rect 15950 121243 15973 122220
rect 18957 123220 18980 124227
rect 19140 124227 22170 124250
rect 19140 123220 19163 124227
rect 18957 122220 19163 123220
rect 18957 121243 18980 122220
rect 15950 121220 18980 121243
rect 19140 121243 19163 122220
rect 22147 123220 22170 124227
rect 22330 124227 25360 124250
rect 22330 123220 22353 124227
rect 22147 122220 22353 123220
rect 22147 121243 22170 122220
rect 19140 121220 22170 121243
rect 22330 121243 22353 122220
rect 25337 123220 25360 124227
rect 25520 124227 28550 124250
rect 25520 123220 25543 124227
rect 25337 122220 25543 123220
rect 25337 121243 25360 122220
rect 22330 121220 25360 121243
rect 25520 121243 25543 122220
rect 28527 123220 28550 124227
rect 28710 124227 31740 124250
rect 28710 123220 28733 124227
rect 28527 122220 28733 123220
rect 28527 121243 28550 122220
rect 25520 121220 28550 121243
rect 28710 121243 28733 122220
rect 31717 123220 31740 124227
rect 31900 124227 34930 124250
rect 31900 123220 31923 124227
rect 31717 122220 31923 123220
rect 31717 121243 31740 122220
rect 28710 121220 31740 121243
rect 31900 121243 31923 122220
rect 34907 123220 34930 124227
rect 35090 124227 38120 124250
rect 35090 123220 35113 124227
rect 34907 122220 35113 123220
rect 34907 121243 34930 122220
rect 31900 121220 34930 121243
rect 35090 121243 35113 122220
rect 38097 123220 38120 124227
rect 38280 124227 41310 124250
rect 38280 123220 38303 124227
rect 38097 122220 38303 123220
rect 38097 121243 38120 122220
rect 35090 121220 38120 121243
rect 38280 121243 38303 122220
rect 41287 123220 41310 124227
rect 41470 124227 44500 124250
rect 41470 123220 41493 124227
rect 41287 122220 41493 123220
rect 41287 121243 41310 122220
rect 38280 121220 41310 121243
rect 41470 121243 41493 122220
rect 44477 123220 44500 124227
rect 44660 124227 47690 124250
rect 44660 123220 44683 124227
rect 44477 122220 44683 123220
rect 44477 121243 44500 122220
rect 41470 121220 44500 121243
rect 44660 121243 44683 122220
rect 47667 123220 47690 124227
rect 47850 124227 50880 124250
rect 47850 123220 47873 124227
rect 47667 122220 47873 123220
rect 47667 121243 47690 122220
rect 44660 121220 47690 121243
rect 47850 121243 47873 122220
rect 50857 123220 50880 124227
rect 51040 124227 54070 124250
rect 51040 123220 51063 124227
rect 50857 122220 51063 123220
rect 50857 121243 50880 122220
rect 47850 121220 50880 121243
rect 51040 121243 51063 122220
rect 54047 123220 54070 124227
rect 54230 124227 57260 124250
rect 54230 123220 54253 124227
rect 54047 122220 54253 123220
rect 54047 121243 54070 122220
rect 51040 121220 54070 121243
rect 54230 121243 54253 122220
rect 57237 123220 57260 124227
rect 57420 124227 60450 124250
rect 57420 123220 57443 124227
rect 57237 122220 57443 123220
rect 57237 121243 57260 122220
rect 54230 121220 57260 121243
rect 57420 121243 57443 122220
rect 60427 123220 60450 124227
rect 60610 124227 63640 124250
rect 60610 123220 60633 124227
rect 60427 122220 60633 123220
rect 60427 121243 60450 122220
rect 57420 121220 60450 121243
rect 60610 121243 60633 122220
rect 63617 123220 63640 124227
rect 63800 124227 66830 124250
rect 63800 123220 63823 124227
rect 63617 122220 63823 123220
rect 63617 121243 63640 122220
rect 60610 121220 63640 121243
rect 63800 121243 63823 122220
rect 66807 123220 66830 124227
rect 66990 124227 70020 124250
rect 66990 123220 67013 124227
rect 66807 122220 67013 123220
rect 66807 121243 66830 122220
rect 63800 121220 66830 121243
rect 66990 121243 67013 122220
rect 69997 123220 70020 124227
rect 70180 124227 73210 124250
rect 70180 123220 70203 124227
rect 69997 122220 70203 123220
rect 69997 121243 70020 122220
rect 66990 121220 70020 121243
rect 70180 121243 70203 122220
rect 73187 123220 73210 124227
rect 73370 124227 76400 124250
rect 73370 123220 73393 124227
rect 73187 122220 73393 123220
rect 73187 121243 73210 122220
rect 70180 121220 73210 121243
rect 73370 121243 73393 122220
rect 76377 123220 76400 124227
rect 76560 124227 79590 124250
rect 76560 123220 76583 124227
rect 76377 122220 76583 123220
rect 76377 121243 76400 122220
rect 73370 121220 76400 121243
rect 76560 121243 76583 122220
rect 79567 123220 79590 124227
rect 79750 124227 82780 124250
rect 79750 123220 79773 124227
rect 79567 122220 79773 123220
rect 79567 121243 79590 122220
rect 76560 121220 79590 121243
rect 79750 121243 79773 122220
rect 82757 123220 82780 124227
rect 82940 124227 85970 124250
rect 82940 123220 82963 124227
rect 82757 122220 82963 123220
rect 82757 121243 82780 122220
rect 79750 121220 82780 121243
rect 82940 121243 82963 122220
rect 85947 123220 85970 124227
rect 86130 124227 89160 124250
rect 86130 123220 86153 124227
rect 85947 122220 86153 123220
rect 85947 121243 85970 122220
rect 82940 121220 85970 121243
rect 86130 121243 86153 122220
rect 89137 123220 89160 124227
rect 89320 124227 92350 124250
rect 89320 123220 89343 124227
rect 89137 122220 89343 123220
rect 89137 121243 89160 122220
rect 86130 121220 89160 121243
rect 89320 121243 89343 122220
rect 92327 123220 92350 124227
rect 92510 124227 95540 124250
rect 92510 123220 92533 124227
rect 92327 122220 92533 123220
rect 92327 121243 92350 122220
rect 89320 121220 92350 121243
rect 92510 121243 92533 122220
rect 95517 123220 95540 124227
rect 95700 124227 98730 124250
rect 95700 123220 95723 124227
rect 95517 122220 95723 123220
rect 95517 121243 95540 122220
rect 92510 121220 95540 121243
rect 95700 121243 95723 122220
rect 98707 123220 98730 124227
rect 98890 124227 101920 124250
rect 98890 123220 98913 124227
rect 98707 122220 98913 123220
rect 98707 121243 98730 122220
rect 95700 121220 98730 121243
rect 98890 121243 98913 122220
rect 101897 123220 101920 124227
rect 102080 124227 105110 124250
rect 102080 123220 102103 124227
rect 101897 122220 102103 123220
rect 101897 121243 101920 122220
rect 98890 121220 101920 121243
rect 102080 121243 102103 122220
rect 105087 123220 105110 124227
rect 105270 124227 108300 124250
rect 105270 123220 105293 124227
rect 105087 122220 105293 123220
rect 105087 121243 105110 122220
rect 102080 121220 105110 121243
rect 105270 121243 105293 122220
rect 108277 123220 108300 124227
rect 108460 124227 111490 124250
rect 108460 123220 108483 124227
rect 108277 122220 108483 123220
rect 108277 121243 108300 122220
rect 105270 121220 108300 121243
rect 108460 121243 108483 122220
rect 111467 123220 111490 124227
rect 111650 124227 114680 124250
rect 111650 123220 111673 124227
rect 111467 122220 111673 123220
rect 111467 121243 111490 122220
rect 108460 121220 111490 121243
rect 111650 121243 111673 122220
rect 114657 123220 114680 124227
rect 114840 124227 117870 124250
rect 114840 123220 114863 124227
rect 114657 122220 114863 123220
rect 114657 121243 114680 122220
rect 111650 121220 114680 121243
rect 114840 121243 114863 122220
rect 117847 123220 117870 124227
rect 118030 124227 121060 124250
rect 118030 123220 118053 124227
rect 117847 122220 118053 123220
rect 117847 121243 117870 122220
rect 114840 121220 117870 121243
rect 118030 121243 118053 122220
rect 121037 123220 121060 124227
rect 121220 124227 124250 124250
rect 121220 123220 121243 124227
rect 121037 122220 121243 123220
rect 121037 121243 121060 122220
rect 118030 121220 121060 121243
rect 121220 121243 121243 122220
rect 124227 123220 124250 124227
rect 124410 124227 127440 124250
rect 124410 123220 124433 124227
rect 124227 122220 124433 123220
rect 124227 121243 124250 122220
rect 121220 121220 124250 121243
rect 124410 121243 124433 122220
rect 127417 123220 127440 124227
rect 127600 124227 130630 124250
rect 127600 123220 127623 124227
rect 127417 122220 127623 123220
rect 127417 121243 127440 122220
rect 124410 121220 127440 121243
rect 127600 121243 127623 122220
rect 130607 123220 130630 124227
rect 130790 124227 133820 124250
rect 130790 123220 130813 124227
rect 130607 122220 130813 123220
rect 130607 121243 130630 122220
rect 127600 121220 130630 121243
rect 130790 121243 130813 122220
rect 133797 123220 133820 124227
rect 133980 124227 137010 124250
rect 133980 123220 134003 124227
rect 133797 122220 134003 123220
rect 133797 121243 133820 122220
rect 130790 121220 133820 121243
rect 133980 121243 134003 122220
rect 136987 123220 137010 124227
rect 136987 122220 137170 123220
rect 136987 121243 137010 122220
rect 133980 121220 137010 121243
rect 10570 121060 11570 121220
rect 13760 121060 14760 121220
rect 16950 121060 17950 121220
rect 20140 121060 21140 121220
rect 23330 121060 24330 121220
rect 26520 121060 27520 121220
rect 29710 121060 30710 121220
rect 32900 121060 33900 121220
rect 36090 121060 37090 121220
rect 39280 121060 40280 121220
rect 42470 121060 43470 121220
rect 45660 121060 46660 121220
rect 48850 121060 49850 121220
rect 52040 121060 53040 121220
rect 55230 121060 56230 121220
rect 58420 121060 59420 121220
rect 61610 121060 62610 121220
rect 64800 121060 65800 121220
rect 67990 121060 68990 121220
rect 71180 121060 72180 121220
rect 74370 121060 75370 121220
rect 77560 121060 78560 121220
rect 80750 121060 81750 121220
rect 83940 121060 84940 121220
rect 87130 121060 88130 121220
rect 90320 121060 91320 121220
rect 93510 121060 94510 121220
rect 96700 121060 97700 121220
rect 99890 121060 100890 121220
rect 103080 121060 104080 121220
rect 106270 121060 107270 121220
rect 109460 121060 110460 121220
rect 112650 121060 113650 121220
rect 115840 121060 116840 121220
rect 119030 121060 120030 121220
rect 122220 121060 123220 121220
rect 125410 121060 126410 121220
rect 128600 121060 129600 121220
rect 131790 121060 132790 121220
rect 134980 121060 135980 121220
rect 0 121037 3030 121060
rect 0 118053 23 121037
rect 3007 120030 3030 121037
rect 3190 121037 6220 121060
rect 3190 120030 3213 121037
rect 3007 119030 3213 120030
rect 3007 118053 3030 119030
rect 0 118030 3030 118053
rect 3190 118053 3213 119030
rect 6197 120030 6220 121037
rect 6380 121037 9410 121060
rect 6380 120030 6403 121037
rect 6197 119030 6403 120030
rect 6197 118053 6220 119030
rect 3190 118030 6220 118053
rect 6380 118053 6403 119030
rect 9387 120030 9410 121037
rect 9570 121037 12600 121060
rect 9570 120030 9593 121037
rect 9387 119030 9593 120030
rect 9387 118053 9410 119030
rect 6380 118030 9410 118053
rect 9570 118053 9593 119030
rect 12577 120030 12600 121037
rect 12760 121037 15790 121060
rect 12760 120030 12783 121037
rect 12577 119030 12783 120030
rect 12577 118053 12600 119030
rect 9570 118030 12600 118053
rect 12760 118053 12783 119030
rect 15767 120030 15790 121037
rect 15950 121037 18980 121060
rect 15950 120030 15973 121037
rect 15767 119030 15973 120030
rect 15767 118053 15790 119030
rect 12760 118030 15790 118053
rect 15950 118053 15973 119030
rect 18957 120030 18980 121037
rect 19140 121037 22170 121060
rect 19140 120030 19163 121037
rect 18957 119030 19163 120030
rect 18957 118053 18980 119030
rect 15950 118030 18980 118053
rect 19140 118053 19163 119030
rect 22147 120030 22170 121037
rect 22330 121037 25360 121060
rect 22330 120030 22353 121037
rect 22147 119030 22353 120030
rect 22147 118053 22170 119030
rect 19140 118030 22170 118053
rect 22330 118053 22353 119030
rect 25337 120030 25360 121037
rect 25520 121037 28550 121060
rect 25520 120030 25543 121037
rect 25337 119030 25543 120030
rect 25337 118053 25360 119030
rect 22330 118030 25360 118053
rect 25520 118053 25543 119030
rect 28527 120030 28550 121037
rect 28710 121037 31740 121060
rect 28710 120030 28733 121037
rect 28527 119030 28733 120030
rect 28527 118053 28550 119030
rect 25520 118030 28550 118053
rect 28710 118053 28733 119030
rect 31717 120030 31740 121037
rect 31900 121037 34930 121060
rect 31900 120030 31923 121037
rect 31717 119030 31923 120030
rect 31717 118053 31740 119030
rect 28710 118030 31740 118053
rect 31900 118053 31923 119030
rect 34907 120030 34930 121037
rect 35090 121037 38120 121060
rect 35090 120030 35113 121037
rect 34907 119030 35113 120030
rect 34907 118053 34930 119030
rect 31900 118030 34930 118053
rect 35090 118053 35113 119030
rect 38097 120030 38120 121037
rect 38280 121037 41310 121060
rect 38280 120030 38303 121037
rect 38097 119030 38303 120030
rect 38097 118053 38120 119030
rect 35090 118030 38120 118053
rect 38280 118053 38303 119030
rect 41287 120030 41310 121037
rect 41470 121037 44500 121060
rect 41470 120030 41493 121037
rect 41287 119030 41493 120030
rect 41287 118053 41310 119030
rect 38280 118030 41310 118053
rect 41470 118053 41493 119030
rect 44477 120030 44500 121037
rect 44660 121037 47690 121060
rect 44660 120030 44683 121037
rect 44477 119030 44683 120030
rect 44477 118053 44500 119030
rect 41470 118030 44500 118053
rect 44660 118053 44683 119030
rect 47667 120030 47690 121037
rect 47850 121037 50880 121060
rect 47850 120030 47873 121037
rect 47667 119030 47873 120030
rect 47667 118053 47690 119030
rect 44660 118030 47690 118053
rect 47850 118053 47873 119030
rect 50857 120030 50880 121037
rect 51040 121037 54070 121060
rect 51040 120030 51063 121037
rect 50857 119030 51063 120030
rect 50857 118053 50880 119030
rect 47850 118030 50880 118053
rect 51040 118053 51063 119030
rect 54047 120030 54070 121037
rect 54230 121037 57260 121060
rect 54230 120030 54253 121037
rect 54047 119030 54253 120030
rect 54047 118053 54070 119030
rect 51040 118030 54070 118053
rect 54230 118053 54253 119030
rect 57237 120030 57260 121037
rect 57420 121037 60450 121060
rect 57420 120030 57443 121037
rect 57237 119030 57443 120030
rect 57237 118053 57260 119030
rect 54230 118030 57260 118053
rect 57420 118053 57443 119030
rect 60427 120030 60450 121037
rect 60610 121037 63640 121060
rect 60610 120030 60633 121037
rect 60427 119030 60633 120030
rect 60427 118053 60450 119030
rect 57420 118030 60450 118053
rect 60610 118053 60633 119030
rect 63617 120030 63640 121037
rect 63800 121037 66830 121060
rect 63800 120030 63823 121037
rect 63617 119030 63823 120030
rect 63617 118053 63640 119030
rect 60610 118030 63640 118053
rect 63800 118053 63823 119030
rect 66807 120030 66830 121037
rect 66990 121037 70020 121060
rect 66990 120030 67013 121037
rect 66807 119030 67013 120030
rect 66807 118053 66830 119030
rect 63800 118030 66830 118053
rect 66990 118053 67013 119030
rect 69997 120030 70020 121037
rect 70180 121037 73210 121060
rect 70180 120030 70203 121037
rect 69997 119030 70203 120030
rect 69997 118053 70020 119030
rect 66990 118030 70020 118053
rect 70180 118053 70203 119030
rect 73187 120030 73210 121037
rect 73370 121037 76400 121060
rect 73370 120030 73393 121037
rect 73187 119030 73393 120030
rect 73187 118053 73210 119030
rect 70180 118030 73210 118053
rect 73370 118053 73393 119030
rect 76377 120030 76400 121037
rect 76560 121037 79590 121060
rect 76560 120030 76583 121037
rect 76377 119030 76583 120030
rect 76377 118053 76400 119030
rect 73370 118030 76400 118053
rect 76560 118053 76583 119030
rect 79567 120030 79590 121037
rect 79750 121037 82780 121060
rect 79750 120030 79773 121037
rect 79567 119030 79773 120030
rect 79567 118053 79590 119030
rect 76560 118030 79590 118053
rect 79750 118053 79773 119030
rect 82757 120030 82780 121037
rect 82940 121037 85970 121060
rect 82940 120030 82963 121037
rect 82757 119030 82963 120030
rect 82757 118053 82780 119030
rect 79750 118030 82780 118053
rect 82940 118053 82963 119030
rect 85947 120030 85970 121037
rect 86130 121037 89160 121060
rect 86130 120030 86153 121037
rect 85947 119030 86153 120030
rect 85947 118053 85970 119030
rect 82940 118030 85970 118053
rect 86130 118053 86153 119030
rect 89137 120030 89160 121037
rect 89320 121037 92350 121060
rect 89320 120030 89343 121037
rect 89137 119030 89343 120030
rect 89137 118053 89160 119030
rect 86130 118030 89160 118053
rect 89320 118053 89343 119030
rect 92327 120030 92350 121037
rect 92510 121037 95540 121060
rect 92510 120030 92533 121037
rect 92327 119030 92533 120030
rect 92327 118053 92350 119030
rect 89320 118030 92350 118053
rect 92510 118053 92533 119030
rect 95517 120030 95540 121037
rect 95700 121037 98730 121060
rect 95700 120030 95723 121037
rect 95517 119030 95723 120030
rect 95517 118053 95540 119030
rect 92510 118030 95540 118053
rect 95700 118053 95723 119030
rect 98707 120030 98730 121037
rect 98890 121037 101920 121060
rect 98890 120030 98913 121037
rect 98707 119030 98913 120030
rect 98707 118053 98730 119030
rect 95700 118030 98730 118053
rect 98890 118053 98913 119030
rect 101897 120030 101920 121037
rect 102080 121037 105110 121060
rect 102080 120030 102103 121037
rect 101897 119030 102103 120030
rect 101897 118053 101920 119030
rect 98890 118030 101920 118053
rect 102080 118053 102103 119030
rect 105087 120030 105110 121037
rect 105270 121037 108300 121060
rect 105270 120030 105293 121037
rect 105087 119030 105293 120030
rect 105087 118053 105110 119030
rect 102080 118030 105110 118053
rect 105270 118053 105293 119030
rect 108277 120030 108300 121037
rect 108460 121037 111490 121060
rect 108460 120030 108483 121037
rect 108277 119030 108483 120030
rect 108277 118053 108300 119030
rect 105270 118030 108300 118053
rect 108460 118053 108483 119030
rect 111467 120030 111490 121037
rect 111650 121037 114680 121060
rect 111650 120030 111673 121037
rect 111467 119030 111673 120030
rect 111467 118053 111490 119030
rect 108460 118030 111490 118053
rect 111650 118053 111673 119030
rect 114657 120030 114680 121037
rect 114840 121037 117870 121060
rect 114840 120030 114863 121037
rect 114657 119030 114863 120030
rect 114657 118053 114680 119030
rect 111650 118030 114680 118053
rect 114840 118053 114863 119030
rect 117847 120030 117870 121037
rect 118030 121037 121060 121060
rect 118030 120030 118053 121037
rect 117847 119030 118053 120030
rect 117847 118053 117870 119030
rect 114840 118030 117870 118053
rect 118030 118053 118053 119030
rect 121037 120030 121060 121037
rect 121220 121037 124250 121060
rect 121220 120030 121243 121037
rect 121037 119030 121243 120030
rect 121037 118053 121060 119030
rect 118030 118030 121060 118053
rect 121220 118053 121243 119030
rect 124227 120030 124250 121037
rect 124410 121037 127440 121060
rect 124410 120030 124433 121037
rect 124227 119030 124433 120030
rect 124227 118053 124250 119030
rect 121220 118030 124250 118053
rect 124410 118053 124433 119030
rect 127417 120030 127440 121037
rect 127600 121037 130630 121060
rect 127600 120030 127623 121037
rect 127417 119030 127623 120030
rect 127417 118053 127440 119030
rect 124410 118030 127440 118053
rect 127600 118053 127623 119030
rect 130607 120030 130630 121037
rect 130790 121037 133820 121060
rect 130790 120030 130813 121037
rect 130607 119030 130813 120030
rect 130607 118053 130630 119030
rect 127600 118030 130630 118053
rect 130790 118053 130813 119030
rect 133797 120030 133820 121037
rect 133980 121037 137010 121060
rect 133980 120030 134003 121037
rect 133797 119030 134003 120030
rect 133797 118053 133820 119030
rect 130790 118030 133820 118053
rect 133980 118053 134003 119030
rect 136987 120030 137010 121037
rect 136987 119030 137170 120030
rect 136987 118053 137010 119030
rect 133980 118030 137010 118053
rect 1000 117870 2000 118030
rect 4190 117870 5190 118030
rect 7380 117870 8380 118030
rect 10570 117870 11570 118030
rect 13760 117870 14760 118030
rect 16950 117870 17950 118030
rect 20140 117870 21140 118030
rect 23330 117870 24330 118030
rect 26520 117870 27520 118030
rect 29710 117870 30710 118030
rect 32900 117870 33900 118030
rect 36090 117870 37090 118030
rect 39280 117870 40280 118030
rect 42470 117870 43470 118030
rect 45660 117870 46660 118030
rect 48850 117870 49850 118030
rect 52040 117870 53040 118030
rect 55230 117870 56230 118030
rect 58420 117870 59420 118030
rect 61610 117870 62610 118030
rect 64800 117870 65800 118030
rect 67990 117870 68990 118030
rect 71180 117870 72180 118030
rect 74370 117870 75370 118030
rect 77560 117870 78560 118030
rect 80750 117870 81750 118030
rect 83940 117870 84940 118030
rect 87130 117870 88130 118030
rect 90320 117870 91320 118030
rect 93510 117870 94510 118030
rect 96700 117870 97700 118030
rect 99890 117870 100890 118030
rect 103080 117870 104080 118030
rect 106270 117870 107270 118030
rect 109460 117870 110460 118030
rect 112650 117870 113650 118030
rect 115840 117870 116840 118030
rect 119030 117870 120030 118030
rect 122220 117870 123220 118030
rect 125410 117870 126410 118030
rect 128600 117870 129600 118030
rect 131790 117870 132790 118030
rect 134980 117870 135980 118030
rect 0 117847 3030 117870
rect 0 114863 23 117847
rect 3007 116840 3030 117847
rect 3190 117847 6220 117870
rect 3190 116840 3213 117847
rect 3007 115840 3213 116840
rect 3007 114863 3030 115840
rect 0 114840 3030 114863
rect 3190 114863 3213 115840
rect 6197 116840 6220 117847
rect 6380 117847 9410 117870
rect 6380 116840 6403 117847
rect 6197 115840 6403 116840
rect 6197 114863 6220 115840
rect 3190 114840 6220 114863
rect 6380 114863 6403 115840
rect 9387 116840 9410 117847
rect 9570 117847 12600 117870
rect 9570 116840 9593 117847
rect 9387 115840 9593 116840
rect 9387 114863 9410 115840
rect 6380 114840 9410 114863
rect 9570 114863 9593 115840
rect 12577 116840 12600 117847
rect 12760 117847 15790 117870
rect 12760 116840 12783 117847
rect 12577 115840 12783 116840
rect 12577 114863 12600 115840
rect 9570 114840 12600 114863
rect 12760 114863 12783 115840
rect 15767 116840 15790 117847
rect 15950 117847 18980 117870
rect 15950 116840 15973 117847
rect 15767 115840 15973 116840
rect 15767 114863 15790 115840
rect 12760 114840 15790 114863
rect 15950 114863 15973 115840
rect 18957 116840 18980 117847
rect 19140 117847 22170 117870
rect 19140 116840 19163 117847
rect 18957 115840 19163 116840
rect 18957 114863 18980 115840
rect 15950 114840 18980 114863
rect 19140 114863 19163 115840
rect 22147 116840 22170 117847
rect 22330 117847 25360 117870
rect 22330 116840 22353 117847
rect 22147 115840 22353 116840
rect 22147 114863 22170 115840
rect 19140 114840 22170 114863
rect 22330 114863 22353 115840
rect 25337 116840 25360 117847
rect 25520 117847 28550 117870
rect 25520 116840 25543 117847
rect 25337 115840 25543 116840
rect 25337 114863 25360 115840
rect 22330 114840 25360 114863
rect 25520 114863 25543 115840
rect 28527 116840 28550 117847
rect 28710 117847 31740 117870
rect 28710 116840 28733 117847
rect 28527 115840 28733 116840
rect 28527 114863 28550 115840
rect 25520 114840 28550 114863
rect 28710 114863 28733 115840
rect 31717 116840 31740 117847
rect 31900 117847 34930 117870
rect 31900 116840 31923 117847
rect 31717 115840 31923 116840
rect 31717 114863 31740 115840
rect 28710 114840 31740 114863
rect 31900 114863 31923 115840
rect 34907 116840 34930 117847
rect 35090 117847 38120 117870
rect 35090 116840 35113 117847
rect 34907 115840 35113 116840
rect 34907 114863 34930 115840
rect 31900 114840 34930 114863
rect 35090 114863 35113 115840
rect 38097 116840 38120 117847
rect 38280 117847 41310 117870
rect 38280 116840 38303 117847
rect 38097 115840 38303 116840
rect 38097 114863 38120 115840
rect 35090 114840 38120 114863
rect 38280 114863 38303 115840
rect 41287 116840 41310 117847
rect 41470 117847 44500 117870
rect 41470 116840 41493 117847
rect 41287 115840 41493 116840
rect 41287 114863 41310 115840
rect 38280 114840 41310 114863
rect 41470 114863 41493 115840
rect 44477 116840 44500 117847
rect 44660 117847 47690 117870
rect 44660 116840 44683 117847
rect 44477 115840 44683 116840
rect 44477 114863 44500 115840
rect 41470 114840 44500 114863
rect 44660 114863 44683 115840
rect 47667 116840 47690 117847
rect 47850 117847 50880 117870
rect 47850 116840 47873 117847
rect 47667 115840 47873 116840
rect 47667 114863 47690 115840
rect 44660 114840 47690 114863
rect 47850 114863 47873 115840
rect 50857 116840 50880 117847
rect 51040 117847 54070 117870
rect 51040 116840 51063 117847
rect 50857 115840 51063 116840
rect 50857 114863 50880 115840
rect 47850 114840 50880 114863
rect 51040 114863 51063 115840
rect 54047 116840 54070 117847
rect 54230 117847 57260 117870
rect 54230 116840 54253 117847
rect 54047 115840 54253 116840
rect 54047 114863 54070 115840
rect 51040 114840 54070 114863
rect 54230 114863 54253 115840
rect 57237 116840 57260 117847
rect 57420 117847 60450 117870
rect 57420 116840 57443 117847
rect 57237 115840 57443 116840
rect 57237 114863 57260 115840
rect 54230 114840 57260 114863
rect 57420 114863 57443 115840
rect 60427 116840 60450 117847
rect 60610 117847 63640 117870
rect 60610 116840 60633 117847
rect 60427 115840 60633 116840
rect 60427 114863 60450 115840
rect 57420 114840 60450 114863
rect 60610 114863 60633 115840
rect 63617 116840 63640 117847
rect 63800 117847 66830 117870
rect 63800 116840 63823 117847
rect 63617 115840 63823 116840
rect 63617 114863 63640 115840
rect 60610 114840 63640 114863
rect 63800 114863 63823 115840
rect 66807 116840 66830 117847
rect 66990 117847 70020 117870
rect 66990 116840 67013 117847
rect 66807 115840 67013 116840
rect 66807 114863 66830 115840
rect 63800 114840 66830 114863
rect 66990 114863 67013 115840
rect 69997 116840 70020 117847
rect 70180 117847 73210 117870
rect 70180 116840 70203 117847
rect 69997 115840 70203 116840
rect 69997 114863 70020 115840
rect 66990 114840 70020 114863
rect 70180 114863 70203 115840
rect 73187 116840 73210 117847
rect 73370 117847 76400 117870
rect 73370 116840 73393 117847
rect 73187 115840 73393 116840
rect 73187 114863 73210 115840
rect 70180 114840 73210 114863
rect 73370 114863 73393 115840
rect 76377 116840 76400 117847
rect 76560 117847 79590 117870
rect 76560 116840 76583 117847
rect 76377 115840 76583 116840
rect 76377 114863 76400 115840
rect 73370 114840 76400 114863
rect 76560 114863 76583 115840
rect 79567 116840 79590 117847
rect 79750 117847 82780 117870
rect 79750 116840 79773 117847
rect 79567 115840 79773 116840
rect 79567 114863 79590 115840
rect 76560 114840 79590 114863
rect 79750 114863 79773 115840
rect 82757 116840 82780 117847
rect 82940 117847 85970 117870
rect 82940 116840 82963 117847
rect 82757 115840 82963 116840
rect 82757 114863 82780 115840
rect 79750 114840 82780 114863
rect 82940 114863 82963 115840
rect 85947 116840 85970 117847
rect 86130 117847 89160 117870
rect 86130 116840 86153 117847
rect 85947 115840 86153 116840
rect 85947 114863 85970 115840
rect 82940 114840 85970 114863
rect 86130 114863 86153 115840
rect 89137 116840 89160 117847
rect 89320 117847 92350 117870
rect 89320 116840 89343 117847
rect 89137 115840 89343 116840
rect 89137 114863 89160 115840
rect 86130 114840 89160 114863
rect 89320 114863 89343 115840
rect 92327 116840 92350 117847
rect 92510 117847 95540 117870
rect 92510 116840 92533 117847
rect 92327 115840 92533 116840
rect 92327 114863 92350 115840
rect 89320 114840 92350 114863
rect 92510 114863 92533 115840
rect 95517 116840 95540 117847
rect 95700 117847 98730 117870
rect 95700 116840 95723 117847
rect 95517 115840 95723 116840
rect 95517 114863 95540 115840
rect 92510 114840 95540 114863
rect 95700 114863 95723 115840
rect 98707 116840 98730 117847
rect 98890 117847 101920 117870
rect 98890 116840 98913 117847
rect 98707 115840 98913 116840
rect 98707 114863 98730 115840
rect 95700 114840 98730 114863
rect 98890 114863 98913 115840
rect 101897 116840 101920 117847
rect 102080 117847 105110 117870
rect 102080 116840 102103 117847
rect 101897 115840 102103 116840
rect 101897 114863 101920 115840
rect 98890 114840 101920 114863
rect 102080 114863 102103 115840
rect 105087 116840 105110 117847
rect 105270 117847 108300 117870
rect 105270 116840 105293 117847
rect 105087 115840 105293 116840
rect 105087 114863 105110 115840
rect 102080 114840 105110 114863
rect 105270 114863 105293 115840
rect 108277 116840 108300 117847
rect 108460 117847 111490 117870
rect 108460 116840 108483 117847
rect 108277 115840 108483 116840
rect 108277 114863 108300 115840
rect 105270 114840 108300 114863
rect 108460 114863 108483 115840
rect 111467 116840 111490 117847
rect 111650 117847 114680 117870
rect 111650 116840 111673 117847
rect 111467 115840 111673 116840
rect 111467 114863 111490 115840
rect 108460 114840 111490 114863
rect 111650 114863 111673 115840
rect 114657 116840 114680 117847
rect 114840 117847 117870 117870
rect 114840 116840 114863 117847
rect 114657 115840 114863 116840
rect 114657 114863 114680 115840
rect 111650 114840 114680 114863
rect 114840 114863 114863 115840
rect 117847 116840 117870 117847
rect 118030 117847 121060 117870
rect 118030 116840 118053 117847
rect 117847 115840 118053 116840
rect 117847 114863 117870 115840
rect 114840 114840 117870 114863
rect 118030 114863 118053 115840
rect 121037 116840 121060 117847
rect 121220 117847 124250 117870
rect 121220 116840 121243 117847
rect 121037 115840 121243 116840
rect 121037 114863 121060 115840
rect 118030 114840 121060 114863
rect 121220 114863 121243 115840
rect 124227 116840 124250 117847
rect 124410 117847 127440 117870
rect 124410 116840 124433 117847
rect 124227 115840 124433 116840
rect 124227 114863 124250 115840
rect 121220 114840 124250 114863
rect 124410 114863 124433 115840
rect 127417 116840 127440 117847
rect 127600 117847 130630 117870
rect 127600 116840 127623 117847
rect 127417 115840 127623 116840
rect 127417 114863 127440 115840
rect 124410 114840 127440 114863
rect 127600 114863 127623 115840
rect 130607 116840 130630 117847
rect 130790 117847 133820 117870
rect 130790 116840 130813 117847
rect 130607 115840 130813 116840
rect 130607 114863 130630 115840
rect 127600 114840 130630 114863
rect 130790 114863 130813 115840
rect 133797 116840 133820 117847
rect 133980 117847 137010 117870
rect 133980 116840 134003 117847
rect 133797 115840 134003 116840
rect 133797 114863 133820 115840
rect 130790 114840 133820 114863
rect 133980 114863 134003 115840
rect 136987 116840 137010 117847
rect 136987 115840 137170 116840
rect 136987 114863 137010 115840
rect 133980 114840 137010 114863
rect 1000 114680 2000 114840
rect 4190 114680 5190 114840
rect 7380 114680 8380 114840
rect 10570 114680 11570 114840
rect 13760 114680 14760 114840
rect 16950 114680 17950 114840
rect 20140 114680 21140 114840
rect 23330 114680 24330 114840
rect 26520 114680 27520 114840
rect 29710 114680 30710 114840
rect 32900 114680 33900 114840
rect 36090 114680 37090 114840
rect 39280 114680 40280 114840
rect 42470 114680 43470 114840
rect 45660 114680 46660 114840
rect 48850 114680 49850 114840
rect 52040 114680 53040 114840
rect 55230 114680 56230 114840
rect 58420 114680 59420 114840
rect 61610 114680 62610 114840
rect 64800 114680 65800 114840
rect 67990 114680 68990 114840
rect 71180 114680 72180 114840
rect 74370 114680 75370 114840
rect 77560 114680 78560 114840
rect 80750 114680 81750 114840
rect 83940 114680 84940 114840
rect 87130 114680 88130 114840
rect 90320 114680 91320 114840
rect 93510 114680 94510 114840
rect 96700 114680 97700 114840
rect 99890 114680 100890 114840
rect 103080 114680 104080 114840
rect 106270 114680 107270 114840
rect 109460 114680 110460 114840
rect 112650 114680 113650 114840
rect 115840 114680 116840 114840
rect 119030 114680 120030 114840
rect 122220 114680 123220 114840
rect 125410 114680 126410 114840
rect 128600 114680 129600 114840
rect 131790 114680 132790 114840
rect 134980 114680 135980 114840
rect 0 114657 3030 114680
rect 0 111673 23 114657
rect 3007 113650 3030 114657
rect 3190 114657 6220 114680
rect 3190 113650 3213 114657
rect 3007 112650 3213 113650
rect 3007 111673 3030 112650
rect 0 111650 3030 111673
rect 3190 111673 3213 112650
rect 6197 113650 6220 114657
rect 6380 114657 9410 114680
rect 6380 113650 6403 114657
rect 6197 112650 6403 113650
rect 6197 111673 6220 112650
rect 3190 111650 6220 111673
rect 6380 111673 6403 112650
rect 9387 113650 9410 114657
rect 9570 114657 12600 114680
rect 9570 113650 9593 114657
rect 9387 112650 9593 113650
rect 9387 111673 9410 112650
rect 6380 111650 9410 111673
rect 9570 111673 9593 112650
rect 12577 113650 12600 114657
rect 12760 114657 15790 114680
rect 12760 113650 12783 114657
rect 12577 112650 12783 113650
rect 12577 111673 12600 112650
rect 9570 111650 12600 111673
rect 12760 111673 12783 112650
rect 15767 113650 15790 114657
rect 15950 114657 18980 114680
rect 15950 113650 15973 114657
rect 15767 112650 15973 113650
rect 15767 111673 15790 112650
rect 12760 111650 15790 111673
rect 15950 111673 15973 112650
rect 18957 113650 18980 114657
rect 19140 114657 22170 114680
rect 19140 113650 19163 114657
rect 18957 112650 19163 113650
rect 18957 111673 18980 112650
rect 15950 111650 18980 111673
rect 19140 111673 19163 112650
rect 22147 113650 22170 114657
rect 22330 114657 25360 114680
rect 22330 113650 22353 114657
rect 22147 112650 22353 113650
rect 22147 111673 22170 112650
rect 19140 111650 22170 111673
rect 22330 111673 22353 112650
rect 25337 113650 25360 114657
rect 25520 114657 28550 114680
rect 25520 113650 25543 114657
rect 25337 112650 25543 113650
rect 25337 111673 25360 112650
rect 22330 111650 25360 111673
rect 25520 111673 25543 112650
rect 28527 113650 28550 114657
rect 28710 114657 31740 114680
rect 28710 113650 28733 114657
rect 28527 112650 28733 113650
rect 28527 111673 28550 112650
rect 25520 111650 28550 111673
rect 28710 111673 28733 112650
rect 31717 113650 31740 114657
rect 31900 114657 34930 114680
rect 31900 113650 31923 114657
rect 31717 112650 31923 113650
rect 31717 111673 31740 112650
rect 28710 111650 31740 111673
rect 31900 111673 31923 112650
rect 34907 113650 34930 114657
rect 35090 114657 38120 114680
rect 35090 113650 35113 114657
rect 34907 112650 35113 113650
rect 34907 111673 34930 112650
rect 31900 111650 34930 111673
rect 35090 111673 35113 112650
rect 38097 113650 38120 114657
rect 38280 114657 41310 114680
rect 38280 113650 38303 114657
rect 38097 112650 38303 113650
rect 38097 111673 38120 112650
rect 35090 111650 38120 111673
rect 38280 111673 38303 112650
rect 41287 113650 41310 114657
rect 41470 114657 44500 114680
rect 41470 113650 41493 114657
rect 41287 112650 41493 113650
rect 41287 111673 41310 112650
rect 38280 111650 41310 111673
rect 41470 111673 41493 112650
rect 44477 113650 44500 114657
rect 44660 114657 47690 114680
rect 44660 113650 44683 114657
rect 44477 112650 44683 113650
rect 44477 111673 44500 112650
rect 41470 111650 44500 111673
rect 44660 111673 44683 112650
rect 47667 113650 47690 114657
rect 47850 114657 50880 114680
rect 47850 113650 47873 114657
rect 47667 112650 47873 113650
rect 47667 111673 47690 112650
rect 44660 111650 47690 111673
rect 47850 111673 47873 112650
rect 50857 113650 50880 114657
rect 51040 114657 54070 114680
rect 51040 113650 51063 114657
rect 50857 112650 51063 113650
rect 50857 111673 50880 112650
rect 47850 111650 50880 111673
rect 51040 111673 51063 112650
rect 54047 113650 54070 114657
rect 54230 114657 57260 114680
rect 54230 113650 54253 114657
rect 54047 112650 54253 113650
rect 54047 111673 54070 112650
rect 51040 111650 54070 111673
rect 54230 111673 54253 112650
rect 57237 113650 57260 114657
rect 57420 114657 60450 114680
rect 57420 113650 57443 114657
rect 57237 112650 57443 113650
rect 57237 111673 57260 112650
rect 54230 111650 57260 111673
rect 57420 111673 57443 112650
rect 60427 113650 60450 114657
rect 60610 114657 63640 114680
rect 60610 113650 60633 114657
rect 60427 112650 60633 113650
rect 60427 111673 60450 112650
rect 57420 111650 60450 111673
rect 60610 111673 60633 112650
rect 63617 113650 63640 114657
rect 63800 114657 66830 114680
rect 63800 113650 63823 114657
rect 63617 112650 63823 113650
rect 63617 111673 63640 112650
rect 60610 111650 63640 111673
rect 63800 111673 63823 112650
rect 66807 113650 66830 114657
rect 66990 114657 70020 114680
rect 66990 113650 67013 114657
rect 66807 112650 67013 113650
rect 66807 111673 66830 112650
rect 63800 111650 66830 111673
rect 66990 111673 67013 112650
rect 69997 113650 70020 114657
rect 70180 114657 73210 114680
rect 70180 113650 70203 114657
rect 69997 112650 70203 113650
rect 69997 111673 70020 112650
rect 66990 111650 70020 111673
rect 70180 111673 70203 112650
rect 73187 113650 73210 114657
rect 73370 114657 76400 114680
rect 73370 113650 73393 114657
rect 73187 112650 73393 113650
rect 73187 111673 73210 112650
rect 70180 111650 73210 111673
rect 73370 111673 73393 112650
rect 76377 113650 76400 114657
rect 76560 114657 79590 114680
rect 76560 113650 76583 114657
rect 76377 112650 76583 113650
rect 76377 111673 76400 112650
rect 73370 111650 76400 111673
rect 76560 111673 76583 112650
rect 79567 113650 79590 114657
rect 79750 114657 82780 114680
rect 79750 113650 79773 114657
rect 79567 112650 79773 113650
rect 79567 111673 79590 112650
rect 76560 111650 79590 111673
rect 79750 111673 79773 112650
rect 82757 113650 82780 114657
rect 82940 114657 85970 114680
rect 82940 113650 82963 114657
rect 82757 112650 82963 113650
rect 82757 111673 82780 112650
rect 79750 111650 82780 111673
rect 82940 111673 82963 112650
rect 85947 113650 85970 114657
rect 86130 114657 89160 114680
rect 86130 113650 86153 114657
rect 85947 112650 86153 113650
rect 85947 111673 85970 112650
rect 82940 111650 85970 111673
rect 86130 111673 86153 112650
rect 89137 113650 89160 114657
rect 89320 114657 92350 114680
rect 89320 113650 89343 114657
rect 89137 112650 89343 113650
rect 89137 111673 89160 112650
rect 86130 111650 89160 111673
rect 89320 111673 89343 112650
rect 92327 113650 92350 114657
rect 92510 114657 95540 114680
rect 92510 113650 92533 114657
rect 92327 112650 92533 113650
rect 92327 111673 92350 112650
rect 89320 111650 92350 111673
rect 92510 111673 92533 112650
rect 95517 113650 95540 114657
rect 95700 114657 98730 114680
rect 95700 113650 95723 114657
rect 95517 112650 95723 113650
rect 95517 111673 95540 112650
rect 92510 111650 95540 111673
rect 95700 111673 95723 112650
rect 98707 113650 98730 114657
rect 98890 114657 101920 114680
rect 98890 113650 98913 114657
rect 98707 112650 98913 113650
rect 98707 111673 98730 112650
rect 95700 111650 98730 111673
rect 98890 111673 98913 112650
rect 101897 113650 101920 114657
rect 102080 114657 105110 114680
rect 102080 113650 102103 114657
rect 101897 112650 102103 113650
rect 101897 111673 101920 112650
rect 98890 111650 101920 111673
rect 102080 111673 102103 112650
rect 105087 113650 105110 114657
rect 105270 114657 108300 114680
rect 105270 113650 105293 114657
rect 105087 112650 105293 113650
rect 105087 111673 105110 112650
rect 102080 111650 105110 111673
rect 105270 111673 105293 112650
rect 108277 113650 108300 114657
rect 108460 114657 111490 114680
rect 108460 113650 108483 114657
rect 108277 112650 108483 113650
rect 108277 111673 108300 112650
rect 105270 111650 108300 111673
rect 108460 111673 108483 112650
rect 111467 113650 111490 114657
rect 111650 114657 114680 114680
rect 111650 113650 111673 114657
rect 111467 112650 111673 113650
rect 111467 111673 111490 112650
rect 108460 111650 111490 111673
rect 111650 111673 111673 112650
rect 114657 113650 114680 114657
rect 114840 114657 117870 114680
rect 114840 113650 114863 114657
rect 114657 112650 114863 113650
rect 114657 111673 114680 112650
rect 111650 111650 114680 111673
rect 114840 111673 114863 112650
rect 117847 113650 117870 114657
rect 118030 114657 121060 114680
rect 118030 113650 118053 114657
rect 117847 112650 118053 113650
rect 117847 111673 117870 112650
rect 114840 111650 117870 111673
rect 118030 111673 118053 112650
rect 121037 113650 121060 114657
rect 121220 114657 124250 114680
rect 121220 113650 121243 114657
rect 121037 112650 121243 113650
rect 121037 111673 121060 112650
rect 118030 111650 121060 111673
rect 121220 111673 121243 112650
rect 124227 113650 124250 114657
rect 124410 114657 127440 114680
rect 124410 113650 124433 114657
rect 124227 112650 124433 113650
rect 124227 111673 124250 112650
rect 121220 111650 124250 111673
rect 124410 111673 124433 112650
rect 127417 113650 127440 114657
rect 127600 114657 130630 114680
rect 127600 113650 127623 114657
rect 127417 112650 127623 113650
rect 127417 111673 127440 112650
rect 124410 111650 127440 111673
rect 127600 111673 127623 112650
rect 130607 113650 130630 114657
rect 130790 114657 133820 114680
rect 130790 113650 130813 114657
rect 130607 112650 130813 113650
rect 130607 111673 130630 112650
rect 127600 111650 130630 111673
rect 130790 111673 130813 112650
rect 133797 113650 133820 114657
rect 133980 114657 137010 114680
rect 133980 113650 134003 114657
rect 133797 112650 134003 113650
rect 133797 111673 133820 112650
rect 130790 111650 133820 111673
rect 133980 111673 134003 112650
rect 136987 113650 137010 114657
rect 136987 112650 137170 113650
rect 136987 111673 137010 112650
rect 133980 111650 137010 111673
rect 1000 111490 2000 111650
rect 4190 111490 5190 111650
rect 7380 111490 8380 111650
rect 10570 111490 11570 111650
rect 13760 111490 14760 111650
rect 16950 111490 17950 111650
rect 20140 111490 21140 111650
rect 23330 111490 24330 111650
rect 26520 111490 27520 111650
rect 29710 111490 30710 111650
rect 32900 111490 33900 111650
rect 36090 111490 37090 111650
rect 39280 111490 40280 111650
rect 42470 111490 43470 111650
rect 45660 111490 46660 111650
rect 48850 111490 49850 111650
rect 52040 111490 53040 111650
rect 55230 111490 56230 111650
rect 58420 111490 59420 111650
rect 61610 111490 62610 111650
rect 64800 111490 65800 111650
rect 67990 111490 68990 111650
rect 71180 111490 72180 111650
rect 74370 111490 75370 111650
rect 77560 111490 78560 111650
rect 80750 111490 81750 111650
rect 83940 111490 84940 111650
rect 87130 111490 88130 111650
rect 90320 111490 91320 111650
rect 93510 111490 94510 111650
rect 96700 111490 97700 111650
rect 99890 111490 100890 111650
rect 103080 111490 104080 111650
rect 106270 111490 107270 111650
rect 109460 111490 110460 111650
rect 112650 111490 113650 111650
rect 115840 111490 116840 111650
rect 119030 111490 120030 111650
rect 122220 111490 123220 111650
rect 125410 111490 126410 111650
rect 128600 111490 129600 111650
rect 131790 111490 132790 111650
rect 134980 111490 135980 111650
rect 0 111467 3030 111490
rect 0 108483 23 111467
rect 3007 110460 3030 111467
rect 3190 111467 6220 111490
rect 3190 110460 3213 111467
rect 3007 109460 3213 110460
rect 3007 108483 3030 109460
rect 0 108460 3030 108483
rect 3190 108483 3213 109460
rect 6197 110460 6220 111467
rect 6380 111467 9410 111490
rect 6380 110460 6403 111467
rect 6197 109460 6403 110460
rect 6197 108483 6220 109460
rect 3190 108460 6220 108483
rect 6380 108483 6403 109460
rect 9387 110460 9410 111467
rect 9570 111467 12600 111490
rect 9570 110460 9593 111467
rect 9387 109460 9593 110460
rect 9387 108483 9410 109460
rect 6380 108460 9410 108483
rect 9570 108483 9593 109460
rect 12577 110460 12600 111467
rect 12760 111467 15790 111490
rect 12760 110460 12783 111467
rect 12577 109460 12783 110460
rect 12577 108483 12600 109460
rect 9570 108460 12600 108483
rect 12760 108483 12783 109460
rect 15767 110460 15790 111467
rect 15950 111467 18980 111490
rect 15950 110460 15973 111467
rect 15767 109460 15973 110460
rect 15767 108483 15790 109460
rect 12760 108460 15790 108483
rect 15950 108483 15973 109460
rect 18957 110460 18980 111467
rect 19140 111467 22170 111490
rect 19140 110460 19163 111467
rect 18957 109460 19163 110460
rect 18957 108483 18980 109460
rect 15950 108460 18980 108483
rect 19140 108483 19163 109460
rect 22147 110460 22170 111467
rect 22330 111467 25360 111490
rect 22330 110460 22353 111467
rect 22147 109460 22353 110460
rect 22147 108483 22170 109460
rect 19140 108460 22170 108483
rect 22330 108483 22353 109460
rect 25337 110460 25360 111467
rect 25520 111467 28550 111490
rect 25520 110460 25543 111467
rect 25337 109460 25543 110460
rect 25337 108483 25360 109460
rect 22330 108460 25360 108483
rect 25520 108483 25543 109460
rect 28527 110460 28550 111467
rect 28710 111467 31740 111490
rect 28710 110460 28733 111467
rect 28527 109460 28733 110460
rect 28527 108483 28550 109460
rect 25520 108460 28550 108483
rect 28710 108483 28733 109460
rect 31717 110460 31740 111467
rect 31900 111467 34930 111490
rect 31900 110460 31923 111467
rect 31717 109460 31923 110460
rect 31717 108483 31740 109460
rect 28710 108460 31740 108483
rect 31900 108483 31923 109460
rect 34907 110460 34930 111467
rect 35090 111467 38120 111490
rect 35090 110460 35113 111467
rect 34907 109460 35113 110460
rect 34907 108483 34930 109460
rect 31900 108460 34930 108483
rect 35090 108483 35113 109460
rect 38097 110460 38120 111467
rect 38280 111467 41310 111490
rect 38280 110460 38303 111467
rect 38097 109460 38303 110460
rect 38097 108483 38120 109460
rect 35090 108460 38120 108483
rect 38280 108483 38303 109460
rect 41287 110460 41310 111467
rect 41470 111467 44500 111490
rect 41470 110460 41493 111467
rect 41287 109460 41493 110460
rect 41287 108483 41310 109460
rect 38280 108460 41310 108483
rect 41470 108483 41493 109460
rect 44477 110460 44500 111467
rect 44660 111467 47690 111490
rect 44660 110460 44683 111467
rect 44477 109460 44683 110460
rect 44477 108483 44500 109460
rect 41470 108460 44500 108483
rect 44660 108483 44683 109460
rect 47667 110460 47690 111467
rect 47850 111467 50880 111490
rect 47850 110460 47873 111467
rect 47667 109460 47873 110460
rect 47667 108483 47690 109460
rect 44660 108460 47690 108483
rect 47850 108483 47873 109460
rect 50857 110460 50880 111467
rect 51040 111467 54070 111490
rect 51040 110460 51063 111467
rect 50857 109460 51063 110460
rect 50857 108483 50880 109460
rect 47850 108460 50880 108483
rect 51040 108483 51063 109460
rect 54047 110460 54070 111467
rect 54230 111467 57260 111490
rect 54230 110460 54253 111467
rect 54047 109460 54253 110460
rect 54047 108483 54070 109460
rect 51040 108460 54070 108483
rect 54230 108483 54253 109460
rect 57237 110460 57260 111467
rect 57420 111467 60450 111490
rect 57420 110460 57443 111467
rect 57237 109460 57443 110460
rect 57237 108483 57260 109460
rect 54230 108460 57260 108483
rect 57420 108483 57443 109460
rect 60427 110460 60450 111467
rect 60610 111467 63640 111490
rect 60610 110460 60633 111467
rect 60427 109460 60633 110460
rect 60427 108483 60450 109460
rect 57420 108460 60450 108483
rect 60610 108483 60633 109460
rect 63617 110460 63640 111467
rect 63800 111467 66830 111490
rect 63800 110460 63823 111467
rect 63617 109460 63823 110460
rect 63617 108483 63640 109460
rect 60610 108460 63640 108483
rect 63800 108483 63823 109460
rect 66807 110460 66830 111467
rect 66990 111467 70020 111490
rect 66990 110460 67013 111467
rect 66807 109460 67013 110460
rect 66807 108483 66830 109460
rect 63800 108460 66830 108483
rect 66990 108483 67013 109460
rect 69997 110460 70020 111467
rect 70180 111467 73210 111490
rect 70180 110460 70203 111467
rect 69997 109460 70203 110460
rect 69997 108483 70020 109460
rect 66990 108460 70020 108483
rect 70180 108483 70203 109460
rect 73187 110460 73210 111467
rect 73370 111467 76400 111490
rect 73370 110460 73393 111467
rect 73187 109460 73393 110460
rect 73187 108483 73210 109460
rect 70180 108460 73210 108483
rect 73370 108483 73393 109460
rect 76377 110460 76400 111467
rect 76560 111467 79590 111490
rect 76560 110460 76583 111467
rect 76377 109460 76583 110460
rect 76377 108483 76400 109460
rect 73370 108460 76400 108483
rect 76560 108483 76583 109460
rect 79567 110460 79590 111467
rect 79750 111467 82780 111490
rect 79750 110460 79773 111467
rect 79567 109460 79773 110460
rect 79567 108483 79590 109460
rect 76560 108460 79590 108483
rect 79750 108483 79773 109460
rect 82757 110460 82780 111467
rect 82940 111467 85970 111490
rect 82940 110460 82963 111467
rect 82757 109460 82963 110460
rect 82757 108483 82780 109460
rect 79750 108460 82780 108483
rect 82940 108483 82963 109460
rect 85947 110460 85970 111467
rect 86130 111467 89160 111490
rect 86130 110460 86153 111467
rect 85947 109460 86153 110460
rect 85947 108483 85970 109460
rect 82940 108460 85970 108483
rect 86130 108483 86153 109460
rect 89137 110460 89160 111467
rect 89320 111467 92350 111490
rect 89320 110460 89343 111467
rect 89137 109460 89343 110460
rect 89137 108483 89160 109460
rect 86130 108460 89160 108483
rect 89320 108483 89343 109460
rect 92327 110460 92350 111467
rect 92510 111467 95540 111490
rect 92510 110460 92533 111467
rect 92327 109460 92533 110460
rect 92327 108483 92350 109460
rect 89320 108460 92350 108483
rect 92510 108483 92533 109460
rect 95517 110460 95540 111467
rect 95700 111467 98730 111490
rect 95700 110460 95723 111467
rect 95517 109460 95723 110460
rect 95517 108483 95540 109460
rect 92510 108460 95540 108483
rect 95700 108483 95723 109460
rect 98707 110460 98730 111467
rect 98890 111467 101920 111490
rect 98890 110460 98913 111467
rect 98707 109460 98913 110460
rect 98707 108483 98730 109460
rect 95700 108460 98730 108483
rect 98890 108483 98913 109460
rect 101897 110460 101920 111467
rect 102080 111467 105110 111490
rect 102080 110460 102103 111467
rect 101897 109460 102103 110460
rect 101897 108483 101920 109460
rect 98890 108460 101920 108483
rect 102080 108483 102103 109460
rect 105087 110460 105110 111467
rect 105270 111467 108300 111490
rect 105270 110460 105293 111467
rect 105087 109460 105293 110460
rect 105087 108483 105110 109460
rect 102080 108460 105110 108483
rect 105270 108483 105293 109460
rect 108277 110460 108300 111467
rect 108460 111467 111490 111490
rect 108460 110460 108483 111467
rect 108277 109460 108483 110460
rect 108277 108483 108300 109460
rect 105270 108460 108300 108483
rect 108460 108483 108483 109460
rect 111467 110460 111490 111467
rect 111650 111467 114680 111490
rect 111650 110460 111673 111467
rect 111467 109460 111673 110460
rect 111467 108483 111490 109460
rect 108460 108460 111490 108483
rect 111650 108483 111673 109460
rect 114657 110460 114680 111467
rect 114840 111467 117870 111490
rect 114840 110460 114863 111467
rect 114657 109460 114863 110460
rect 114657 108483 114680 109460
rect 111650 108460 114680 108483
rect 114840 108483 114863 109460
rect 117847 110460 117870 111467
rect 118030 111467 121060 111490
rect 118030 110460 118053 111467
rect 117847 109460 118053 110460
rect 117847 108483 117870 109460
rect 114840 108460 117870 108483
rect 118030 108483 118053 109460
rect 121037 110460 121060 111467
rect 121220 111467 124250 111490
rect 121220 110460 121243 111467
rect 121037 109460 121243 110460
rect 121037 108483 121060 109460
rect 118030 108460 121060 108483
rect 121220 108483 121243 109460
rect 124227 110460 124250 111467
rect 124410 111467 127440 111490
rect 124410 110460 124433 111467
rect 124227 109460 124433 110460
rect 124227 108483 124250 109460
rect 121220 108460 124250 108483
rect 124410 108483 124433 109460
rect 127417 110460 127440 111467
rect 127600 111467 130630 111490
rect 127600 110460 127623 111467
rect 127417 109460 127623 110460
rect 127417 108483 127440 109460
rect 124410 108460 127440 108483
rect 127600 108483 127623 109460
rect 130607 110460 130630 111467
rect 130790 111467 133820 111490
rect 130790 110460 130813 111467
rect 130607 109460 130813 110460
rect 130607 108483 130630 109460
rect 127600 108460 130630 108483
rect 130790 108483 130813 109460
rect 133797 110460 133820 111467
rect 133980 111467 137010 111490
rect 133980 110460 134003 111467
rect 133797 109460 134003 110460
rect 133797 108483 133820 109460
rect 130790 108460 133820 108483
rect 133980 108483 134003 109460
rect 136987 110460 137010 111467
rect 136987 109460 137170 110460
rect 136987 108483 137010 109460
rect 133980 108460 137010 108483
rect 1000 108300 2000 108460
rect 4190 108300 5190 108460
rect 7380 108300 8380 108460
rect 10570 108300 11570 108460
rect 13760 108300 14760 108460
rect 16950 108300 17950 108460
rect 20140 108300 21140 108460
rect 23330 108300 24330 108460
rect 26520 108300 27520 108460
rect 29710 108300 30710 108460
rect 32900 108300 33900 108460
rect 36090 108300 37090 108460
rect 39280 108300 40280 108460
rect 42470 108300 43470 108460
rect 45660 108300 46660 108460
rect 48850 108300 49850 108460
rect 52040 108300 53040 108460
rect 55230 108300 56230 108460
rect 58420 108300 59420 108460
rect 61610 108300 62610 108460
rect 64800 108300 65800 108460
rect 67990 108300 68990 108460
rect 71180 108300 72180 108460
rect 74370 108300 75370 108460
rect 77560 108300 78560 108460
rect 80750 108300 81750 108460
rect 83940 108300 84940 108460
rect 87130 108300 88130 108460
rect 90320 108300 91320 108460
rect 93510 108300 94510 108460
rect 96700 108300 97700 108460
rect 99890 108300 100890 108460
rect 103080 108300 104080 108460
rect 106270 108300 107270 108460
rect 109460 108300 110460 108460
rect 112650 108300 113650 108460
rect 115840 108300 116840 108460
rect 119030 108300 120030 108460
rect 122220 108300 123220 108460
rect 125410 108300 126410 108460
rect 128600 108300 129600 108460
rect 131790 108300 132790 108460
rect 134980 108300 135980 108460
rect 0 108277 3030 108300
rect 0 105293 23 108277
rect 3007 107270 3030 108277
rect 3190 108277 6220 108300
rect 3190 107270 3213 108277
rect 3007 106270 3213 107270
rect 3007 105293 3030 106270
rect 0 105270 3030 105293
rect 3190 105293 3213 106270
rect 6197 107270 6220 108277
rect 6380 108277 9410 108300
rect 6380 107270 6403 108277
rect 6197 106270 6403 107270
rect 6197 105293 6220 106270
rect 3190 105270 6220 105293
rect 6380 105293 6403 106270
rect 9387 107270 9410 108277
rect 9570 108277 12600 108300
rect 9570 107270 9593 108277
rect 9387 106270 9593 107270
rect 9387 105293 9410 106270
rect 6380 105270 9410 105293
rect 9570 105293 9593 106270
rect 12577 107270 12600 108277
rect 12760 108277 15790 108300
rect 12760 107270 12783 108277
rect 12577 106270 12783 107270
rect 12577 105293 12600 106270
rect 9570 105270 12600 105293
rect 12760 105293 12783 106270
rect 15767 107270 15790 108277
rect 15950 108277 18980 108300
rect 15950 107270 15973 108277
rect 15767 106270 15973 107270
rect 15767 105293 15790 106270
rect 12760 105270 15790 105293
rect 15950 105293 15973 106270
rect 18957 107270 18980 108277
rect 19140 108277 22170 108300
rect 19140 107270 19163 108277
rect 18957 106270 19163 107270
rect 18957 105293 18980 106270
rect 15950 105270 18980 105293
rect 19140 105293 19163 106270
rect 22147 107270 22170 108277
rect 22330 108277 25360 108300
rect 22330 107270 22353 108277
rect 22147 106270 22353 107270
rect 22147 105293 22170 106270
rect 19140 105270 22170 105293
rect 22330 105293 22353 106270
rect 25337 107270 25360 108277
rect 25520 108277 28550 108300
rect 25520 107270 25543 108277
rect 25337 106270 25543 107270
rect 25337 105293 25360 106270
rect 22330 105270 25360 105293
rect 25520 105293 25543 106270
rect 28527 107270 28550 108277
rect 28710 108277 31740 108300
rect 28710 107270 28733 108277
rect 28527 106270 28733 107270
rect 28527 105293 28550 106270
rect 25520 105270 28550 105293
rect 28710 105293 28733 106270
rect 31717 107270 31740 108277
rect 31900 108277 34930 108300
rect 31900 107270 31923 108277
rect 31717 106270 31923 107270
rect 31717 105293 31740 106270
rect 28710 105270 31740 105293
rect 31900 105293 31923 106270
rect 34907 107270 34930 108277
rect 35090 108277 38120 108300
rect 35090 107270 35113 108277
rect 34907 106270 35113 107270
rect 34907 105293 34930 106270
rect 31900 105270 34930 105293
rect 35090 105293 35113 106270
rect 38097 107270 38120 108277
rect 38280 108277 41310 108300
rect 38280 107270 38303 108277
rect 38097 106270 38303 107270
rect 38097 105293 38120 106270
rect 35090 105270 38120 105293
rect 38280 105293 38303 106270
rect 41287 107270 41310 108277
rect 41470 108277 44500 108300
rect 41470 107270 41493 108277
rect 41287 106270 41493 107270
rect 41287 105293 41310 106270
rect 38280 105270 41310 105293
rect 41470 105293 41493 106270
rect 44477 107270 44500 108277
rect 44660 108277 47690 108300
rect 44660 107270 44683 108277
rect 44477 106270 44683 107270
rect 44477 105293 44500 106270
rect 41470 105270 44500 105293
rect 44660 105293 44683 106270
rect 47667 107270 47690 108277
rect 47850 108277 50880 108300
rect 47850 107270 47873 108277
rect 47667 106270 47873 107270
rect 47667 105293 47690 106270
rect 44660 105270 47690 105293
rect 47850 105293 47873 106270
rect 50857 107270 50880 108277
rect 51040 108277 54070 108300
rect 51040 107270 51063 108277
rect 50857 106270 51063 107270
rect 50857 105293 50880 106270
rect 47850 105270 50880 105293
rect 51040 105293 51063 106270
rect 54047 107270 54070 108277
rect 54230 108277 57260 108300
rect 54230 107270 54253 108277
rect 54047 106270 54253 107270
rect 54047 105293 54070 106270
rect 51040 105270 54070 105293
rect 54230 105293 54253 106270
rect 57237 107270 57260 108277
rect 57420 108277 60450 108300
rect 57420 107270 57443 108277
rect 57237 106270 57443 107270
rect 57237 105293 57260 106270
rect 54230 105270 57260 105293
rect 57420 105293 57443 106270
rect 60427 107270 60450 108277
rect 60610 108277 63640 108300
rect 60610 107270 60633 108277
rect 60427 106270 60633 107270
rect 60427 105293 60450 106270
rect 57420 105270 60450 105293
rect 60610 105293 60633 106270
rect 63617 107270 63640 108277
rect 63800 108277 66830 108300
rect 63800 107270 63823 108277
rect 63617 106270 63823 107270
rect 63617 105293 63640 106270
rect 60610 105270 63640 105293
rect 63800 105293 63823 106270
rect 66807 107270 66830 108277
rect 66990 108277 70020 108300
rect 66990 107270 67013 108277
rect 66807 106270 67013 107270
rect 66807 105293 66830 106270
rect 63800 105270 66830 105293
rect 66990 105293 67013 106270
rect 69997 107270 70020 108277
rect 70180 108277 73210 108300
rect 70180 107270 70203 108277
rect 69997 106270 70203 107270
rect 69997 105293 70020 106270
rect 66990 105270 70020 105293
rect 70180 105293 70203 106270
rect 73187 107270 73210 108277
rect 73370 108277 76400 108300
rect 73370 107270 73393 108277
rect 73187 106270 73393 107270
rect 73187 105293 73210 106270
rect 70180 105270 73210 105293
rect 73370 105293 73393 106270
rect 76377 107270 76400 108277
rect 76560 108277 79590 108300
rect 76560 107270 76583 108277
rect 76377 106270 76583 107270
rect 76377 105293 76400 106270
rect 73370 105270 76400 105293
rect 76560 105293 76583 106270
rect 79567 107270 79590 108277
rect 79750 108277 82780 108300
rect 79750 107270 79773 108277
rect 79567 106270 79773 107270
rect 79567 105293 79590 106270
rect 76560 105270 79590 105293
rect 79750 105293 79773 106270
rect 82757 107270 82780 108277
rect 82940 108277 85970 108300
rect 82940 107270 82963 108277
rect 82757 106270 82963 107270
rect 82757 105293 82780 106270
rect 79750 105270 82780 105293
rect 82940 105293 82963 106270
rect 85947 107270 85970 108277
rect 86130 108277 89160 108300
rect 86130 107270 86153 108277
rect 85947 106270 86153 107270
rect 85947 105293 85970 106270
rect 82940 105270 85970 105293
rect 86130 105293 86153 106270
rect 89137 107270 89160 108277
rect 89320 108277 92350 108300
rect 89320 107270 89343 108277
rect 89137 106270 89343 107270
rect 89137 105293 89160 106270
rect 86130 105270 89160 105293
rect 89320 105293 89343 106270
rect 92327 107270 92350 108277
rect 92510 108277 95540 108300
rect 92510 107270 92533 108277
rect 92327 106270 92533 107270
rect 92327 105293 92350 106270
rect 89320 105270 92350 105293
rect 92510 105293 92533 106270
rect 95517 107270 95540 108277
rect 95700 108277 98730 108300
rect 95700 107270 95723 108277
rect 95517 106270 95723 107270
rect 95517 105293 95540 106270
rect 92510 105270 95540 105293
rect 95700 105293 95723 106270
rect 98707 107270 98730 108277
rect 98890 108277 101920 108300
rect 98890 107270 98913 108277
rect 98707 106270 98913 107270
rect 98707 105293 98730 106270
rect 95700 105270 98730 105293
rect 98890 105293 98913 106270
rect 101897 107270 101920 108277
rect 102080 108277 105110 108300
rect 102080 107270 102103 108277
rect 101897 106270 102103 107270
rect 101897 105293 101920 106270
rect 98890 105270 101920 105293
rect 102080 105293 102103 106270
rect 105087 107270 105110 108277
rect 105270 108277 108300 108300
rect 105270 107270 105293 108277
rect 105087 106270 105293 107270
rect 105087 105293 105110 106270
rect 102080 105270 105110 105293
rect 105270 105293 105293 106270
rect 108277 107270 108300 108277
rect 108460 108277 111490 108300
rect 108460 107270 108483 108277
rect 108277 106270 108483 107270
rect 108277 105293 108300 106270
rect 105270 105270 108300 105293
rect 108460 105293 108483 106270
rect 111467 107270 111490 108277
rect 111650 108277 114680 108300
rect 111650 107270 111673 108277
rect 111467 106270 111673 107270
rect 111467 105293 111490 106270
rect 108460 105270 111490 105293
rect 111650 105293 111673 106270
rect 114657 107270 114680 108277
rect 114840 108277 117870 108300
rect 114840 107270 114863 108277
rect 114657 106270 114863 107270
rect 114657 105293 114680 106270
rect 111650 105270 114680 105293
rect 114840 105293 114863 106270
rect 117847 107270 117870 108277
rect 118030 108277 121060 108300
rect 118030 107270 118053 108277
rect 117847 106270 118053 107270
rect 117847 105293 117870 106270
rect 114840 105270 117870 105293
rect 118030 105293 118053 106270
rect 121037 107270 121060 108277
rect 121220 108277 124250 108300
rect 121220 107270 121243 108277
rect 121037 106270 121243 107270
rect 121037 105293 121060 106270
rect 118030 105270 121060 105293
rect 121220 105293 121243 106270
rect 124227 107270 124250 108277
rect 124410 108277 127440 108300
rect 124410 107270 124433 108277
rect 124227 106270 124433 107270
rect 124227 105293 124250 106270
rect 121220 105270 124250 105293
rect 124410 105293 124433 106270
rect 127417 107270 127440 108277
rect 127600 108277 130630 108300
rect 127600 107270 127623 108277
rect 127417 106270 127623 107270
rect 127417 105293 127440 106270
rect 124410 105270 127440 105293
rect 127600 105293 127623 106270
rect 130607 107270 130630 108277
rect 130790 108277 133820 108300
rect 130790 107270 130813 108277
rect 130607 106270 130813 107270
rect 130607 105293 130630 106270
rect 127600 105270 130630 105293
rect 130790 105293 130813 106270
rect 133797 107270 133820 108277
rect 133980 108277 137010 108300
rect 133980 107270 134003 108277
rect 133797 106270 134003 107270
rect 133797 105293 133820 106270
rect 130790 105270 133820 105293
rect 133980 105293 134003 106270
rect 136987 107270 137010 108277
rect 136987 106270 137170 107270
rect 136987 105293 137010 106270
rect 133980 105270 137010 105293
rect 1000 105110 2000 105270
rect 4190 105110 5190 105270
rect 7380 105110 8380 105270
rect 10570 105110 11570 105270
rect 13760 105110 14760 105270
rect 16950 105110 17950 105270
rect 20140 105110 21140 105270
rect 23330 105110 24330 105270
rect 26520 105110 27520 105270
rect 29710 105110 30710 105270
rect 32900 105110 33900 105270
rect 36090 105110 37090 105270
rect 39280 105110 40280 105270
rect 42470 105110 43470 105270
rect 45660 105110 46660 105270
rect 48850 105110 49850 105270
rect 52040 105110 53040 105270
rect 55230 105110 56230 105270
rect 58420 105110 59420 105270
rect 61610 105110 62610 105270
rect 64800 105110 65800 105270
rect 67990 105110 68990 105270
rect 71180 105110 72180 105270
rect 74370 105110 75370 105270
rect 77560 105110 78560 105270
rect 80750 105110 81750 105270
rect 83940 105110 84940 105270
rect 87130 105110 88130 105270
rect 90320 105110 91320 105270
rect 93510 105110 94510 105270
rect 96700 105110 97700 105270
rect 99890 105110 100890 105270
rect 103080 105110 104080 105270
rect 106270 105110 107270 105270
rect 109460 105110 110460 105270
rect 112650 105110 113650 105270
rect 115840 105110 116840 105270
rect 119030 105110 120030 105270
rect 122220 105110 123220 105270
rect 125410 105110 126410 105270
rect 128600 105110 129600 105270
rect 131790 105110 132790 105270
rect 134980 105110 135980 105270
rect 0 105087 3030 105110
rect 0 102103 23 105087
rect 3007 104080 3030 105087
rect 3190 105087 6220 105110
rect 3190 104080 3213 105087
rect 3007 103080 3213 104080
rect 3007 102103 3030 103080
rect 0 102080 3030 102103
rect 3190 102103 3213 103080
rect 6197 104080 6220 105087
rect 6380 105087 9410 105110
rect 6380 104080 6403 105087
rect 6197 103080 6403 104080
rect 6197 102103 6220 103080
rect 3190 102080 6220 102103
rect 6380 102103 6403 103080
rect 9387 104080 9410 105087
rect 9570 105087 12600 105110
rect 9570 104080 9593 105087
rect 9387 103080 9593 104080
rect 9387 102103 9410 103080
rect 6380 102080 9410 102103
rect 9570 102103 9593 103080
rect 12577 104080 12600 105087
rect 12760 105087 15790 105110
rect 12760 104080 12783 105087
rect 12577 103080 12783 104080
rect 12577 102103 12600 103080
rect 9570 102080 12600 102103
rect 12760 102103 12783 103080
rect 15767 104080 15790 105087
rect 15950 105087 18980 105110
rect 15950 104080 15973 105087
rect 15767 103080 15973 104080
rect 15767 102103 15790 103080
rect 12760 102080 15790 102103
rect 15950 102103 15973 103080
rect 18957 104080 18980 105087
rect 19140 105087 22170 105110
rect 19140 104080 19163 105087
rect 18957 103080 19163 104080
rect 18957 102103 18980 103080
rect 15950 102080 18980 102103
rect 19140 102103 19163 103080
rect 22147 104080 22170 105087
rect 22330 105087 25360 105110
rect 22330 104080 22353 105087
rect 22147 103080 22353 104080
rect 22147 102103 22170 103080
rect 19140 102080 22170 102103
rect 22330 102103 22353 103080
rect 25337 104080 25360 105087
rect 25520 105087 28550 105110
rect 25520 104080 25543 105087
rect 25337 103080 25543 104080
rect 25337 102103 25360 103080
rect 22330 102080 25360 102103
rect 25520 102103 25543 103080
rect 28527 104080 28550 105087
rect 28710 105087 31740 105110
rect 28710 104080 28733 105087
rect 28527 103080 28733 104080
rect 28527 102103 28550 103080
rect 25520 102080 28550 102103
rect 28710 102103 28733 103080
rect 31717 104080 31740 105087
rect 31900 105087 34930 105110
rect 31900 104080 31923 105087
rect 31717 103080 31923 104080
rect 31717 102103 31740 103080
rect 28710 102080 31740 102103
rect 31900 102103 31923 103080
rect 34907 104080 34930 105087
rect 35090 105087 38120 105110
rect 35090 104080 35113 105087
rect 34907 103080 35113 104080
rect 34907 102103 34930 103080
rect 31900 102080 34930 102103
rect 35090 102103 35113 103080
rect 38097 104080 38120 105087
rect 38280 105087 41310 105110
rect 38280 104080 38303 105087
rect 38097 103080 38303 104080
rect 38097 102103 38120 103080
rect 35090 102080 38120 102103
rect 38280 102103 38303 103080
rect 41287 104080 41310 105087
rect 41470 105087 44500 105110
rect 41470 104080 41493 105087
rect 41287 103080 41493 104080
rect 41287 102103 41310 103080
rect 38280 102080 41310 102103
rect 41470 102103 41493 103080
rect 44477 104080 44500 105087
rect 44660 105087 47690 105110
rect 44660 104080 44683 105087
rect 44477 103080 44683 104080
rect 44477 102103 44500 103080
rect 41470 102080 44500 102103
rect 44660 102103 44683 103080
rect 47667 104080 47690 105087
rect 47850 105087 50880 105110
rect 47850 104080 47873 105087
rect 47667 103080 47873 104080
rect 47667 102103 47690 103080
rect 44660 102080 47690 102103
rect 47850 102103 47873 103080
rect 50857 104080 50880 105087
rect 51040 105087 54070 105110
rect 51040 104080 51063 105087
rect 50857 103080 51063 104080
rect 50857 102103 50880 103080
rect 47850 102080 50880 102103
rect 51040 102103 51063 103080
rect 54047 104080 54070 105087
rect 54230 105087 57260 105110
rect 54230 104080 54253 105087
rect 54047 103080 54253 104080
rect 54047 102103 54070 103080
rect 51040 102080 54070 102103
rect 54230 102103 54253 103080
rect 57237 104080 57260 105087
rect 57420 105087 60450 105110
rect 57420 104080 57443 105087
rect 57237 103080 57443 104080
rect 57237 102103 57260 103080
rect 54230 102080 57260 102103
rect 57420 102103 57443 103080
rect 60427 104080 60450 105087
rect 60610 105087 63640 105110
rect 60610 104080 60633 105087
rect 60427 103080 60633 104080
rect 60427 102103 60450 103080
rect 57420 102080 60450 102103
rect 60610 102103 60633 103080
rect 63617 104080 63640 105087
rect 63800 105087 66830 105110
rect 63800 104080 63823 105087
rect 63617 103080 63823 104080
rect 63617 102103 63640 103080
rect 60610 102080 63640 102103
rect 63800 102103 63823 103080
rect 66807 104080 66830 105087
rect 66990 105087 70020 105110
rect 66990 104080 67013 105087
rect 66807 103080 67013 104080
rect 66807 102103 66830 103080
rect 63800 102080 66830 102103
rect 66990 102103 67013 103080
rect 69997 104080 70020 105087
rect 70180 105087 73210 105110
rect 70180 104080 70203 105087
rect 69997 103080 70203 104080
rect 69997 102103 70020 103080
rect 66990 102080 70020 102103
rect 70180 102103 70203 103080
rect 73187 104080 73210 105087
rect 73370 105087 76400 105110
rect 73370 104080 73393 105087
rect 73187 103080 73393 104080
rect 73187 102103 73210 103080
rect 70180 102080 73210 102103
rect 73370 102103 73393 103080
rect 76377 104080 76400 105087
rect 76560 105087 79590 105110
rect 76560 104080 76583 105087
rect 76377 103080 76583 104080
rect 76377 102103 76400 103080
rect 73370 102080 76400 102103
rect 76560 102103 76583 103080
rect 79567 104080 79590 105087
rect 79750 105087 82780 105110
rect 79750 104080 79773 105087
rect 79567 103080 79773 104080
rect 79567 102103 79590 103080
rect 76560 102080 79590 102103
rect 79750 102103 79773 103080
rect 82757 104080 82780 105087
rect 82940 105087 85970 105110
rect 82940 104080 82963 105087
rect 82757 103080 82963 104080
rect 82757 102103 82780 103080
rect 79750 102080 82780 102103
rect 82940 102103 82963 103080
rect 85947 104080 85970 105087
rect 86130 105087 89160 105110
rect 86130 104080 86153 105087
rect 85947 103080 86153 104080
rect 85947 102103 85970 103080
rect 82940 102080 85970 102103
rect 86130 102103 86153 103080
rect 89137 104080 89160 105087
rect 89320 105087 92350 105110
rect 89320 104080 89343 105087
rect 89137 103080 89343 104080
rect 89137 102103 89160 103080
rect 86130 102080 89160 102103
rect 89320 102103 89343 103080
rect 92327 104080 92350 105087
rect 92510 105087 95540 105110
rect 92510 104080 92533 105087
rect 92327 103080 92533 104080
rect 92327 102103 92350 103080
rect 89320 102080 92350 102103
rect 92510 102103 92533 103080
rect 95517 104080 95540 105087
rect 95700 105087 98730 105110
rect 95700 104080 95723 105087
rect 95517 103080 95723 104080
rect 95517 102103 95540 103080
rect 92510 102080 95540 102103
rect 95700 102103 95723 103080
rect 98707 104080 98730 105087
rect 98890 105087 101920 105110
rect 98890 104080 98913 105087
rect 98707 103080 98913 104080
rect 98707 102103 98730 103080
rect 95700 102080 98730 102103
rect 98890 102103 98913 103080
rect 101897 104080 101920 105087
rect 102080 105087 105110 105110
rect 102080 104080 102103 105087
rect 101897 103080 102103 104080
rect 101897 102103 101920 103080
rect 98890 102080 101920 102103
rect 102080 102103 102103 103080
rect 105087 104080 105110 105087
rect 105270 105087 108300 105110
rect 105270 104080 105293 105087
rect 105087 103080 105293 104080
rect 105087 102103 105110 103080
rect 102080 102080 105110 102103
rect 105270 102103 105293 103080
rect 108277 104080 108300 105087
rect 108460 105087 111490 105110
rect 108460 104080 108483 105087
rect 108277 103080 108483 104080
rect 108277 102103 108300 103080
rect 105270 102080 108300 102103
rect 108460 102103 108483 103080
rect 111467 104080 111490 105087
rect 111650 105087 114680 105110
rect 111650 104080 111673 105087
rect 111467 103080 111673 104080
rect 111467 102103 111490 103080
rect 108460 102080 111490 102103
rect 111650 102103 111673 103080
rect 114657 104080 114680 105087
rect 114840 105087 117870 105110
rect 114840 104080 114863 105087
rect 114657 103080 114863 104080
rect 114657 102103 114680 103080
rect 111650 102080 114680 102103
rect 114840 102103 114863 103080
rect 117847 104080 117870 105087
rect 118030 105087 121060 105110
rect 118030 104080 118053 105087
rect 117847 103080 118053 104080
rect 117847 102103 117870 103080
rect 114840 102080 117870 102103
rect 118030 102103 118053 103080
rect 121037 104080 121060 105087
rect 121220 105087 124250 105110
rect 121220 104080 121243 105087
rect 121037 103080 121243 104080
rect 121037 102103 121060 103080
rect 118030 102080 121060 102103
rect 121220 102103 121243 103080
rect 124227 104080 124250 105087
rect 124410 105087 127440 105110
rect 124410 104080 124433 105087
rect 124227 103080 124433 104080
rect 124227 102103 124250 103080
rect 121220 102080 124250 102103
rect 124410 102103 124433 103080
rect 127417 104080 127440 105087
rect 127600 105087 130630 105110
rect 127600 104080 127623 105087
rect 127417 103080 127623 104080
rect 127417 102103 127440 103080
rect 124410 102080 127440 102103
rect 127600 102103 127623 103080
rect 130607 104080 130630 105087
rect 130790 105087 133820 105110
rect 130790 104080 130813 105087
rect 130607 103080 130813 104080
rect 130607 102103 130630 103080
rect 127600 102080 130630 102103
rect 130790 102103 130813 103080
rect 133797 104080 133820 105087
rect 133980 105087 137010 105110
rect 133980 104080 134003 105087
rect 133797 103080 134003 104080
rect 133797 102103 133820 103080
rect 130790 102080 133820 102103
rect 133980 102103 134003 103080
rect 136987 104080 137010 105087
rect 136987 103080 137170 104080
rect 136987 102103 137010 103080
rect 133980 102080 137010 102103
rect 1000 101920 2000 102080
rect 4190 101920 5190 102080
rect 7380 101920 8380 102080
rect 10570 101920 11570 102080
rect 13760 101920 14760 102080
rect 16950 101920 17950 102080
rect 20140 101920 21140 102080
rect 23330 101920 24330 102080
rect 26520 101920 27520 102080
rect 29710 101920 30710 102080
rect 32900 101920 33900 102080
rect 36090 101920 37090 102080
rect 39280 101920 40280 102080
rect 42470 101920 43470 102080
rect 45660 101920 46660 102080
rect 48850 101920 49850 102080
rect 52040 101920 53040 102080
rect 55230 101920 56230 102080
rect 58420 101920 59420 102080
rect 61610 101920 62610 102080
rect 64800 101920 65800 102080
rect 67990 101920 68990 102080
rect 71180 101920 72180 102080
rect 74370 101920 75370 102080
rect 77560 101920 78560 102080
rect 80750 101920 81750 102080
rect 83940 101920 84940 102080
rect 87130 101920 88130 102080
rect 90320 101920 91320 102080
rect 93510 101920 94510 102080
rect 96700 101920 97700 102080
rect 99890 101920 100890 102080
rect 103080 101920 104080 102080
rect 106270 101920 107270 102080
rect 109460 101920 110460 102080
rect 112650 101920 113650 102080
rect 115840 101920 116840 102080
rect 119030 101920 120030 102080
rect 122220 101920 123220 102080
rect 125410 101920 126410 102080
rect 128600 101920 129600 102080
rect 131790 101920 132790 102080
rect 134980 101920 135980 102080
rect 0 101897 3030 101920
rect 0 98913 23 101897
rect 3007 100890 3030 101897
rect 3190 101897 6220 101920
rect 3190 100890 3213 101897
rect 3007 99890 3213 100890
rect 3007 98913 3030 99890
rect 0 98890 3030 98913
rect 3190 98913 3213 99890
rect 6197 100890 6220 101897
rect 6380 101897 9410 101920
rect 6380 100890 6403 101897
rect 6197 99890 6403 100890
rect 6197 98913 6220 99890
rect 3190 98890 6220 98913
rect 6380 98913 6403 99890
rect 9387 100890 9410 101897
rect 9570 101897 12600 101920
rect 9570 100890 9593 101897
rect 9387 99890 9593 100890
rect 9387 98913 9410 99890
rect 6380 98890 9410 98913
rect 9570 98913 9593 99890
rect 12577 100890 12600 101897
rect 12760 101897 15790 101920
rect 12760 100890 12783 101897
rect 12577 99890 12783 100890
rect 12577 98913 12600 99890
rect 9570 98890 12600 98913
rect 12760 98913 12783 99890
rect 15767 100890 15790 101897
rect 15950 101897 18980 101920
rect 15950 100890 15973 101897
rect 15767 99890 15973 100890
rect 15767 98913 15790 99890
rect 12760 98890 15790 98913
rect 15950 98913 15973 99890
rect 18957 100890 18980 101897
rect 19140 101897 22170 101920
rect 19140 100890 19163 101897
rect 18957 99890 19163 100890
rect 18957 98913 18980 99890
rect 15950 98890 18980 98913
rect 19140 98913 19163 99890
rect 22147 100890 22170 101897
rect 22330 101897 25360 101920
rect 22330 100890 22353 101897
rect 22147 99890 22353 100890
rect 22147 98913 22170 99890
rect 19140 98890 22170 98913
rect 22330 98913 22353 99890
rect 25337 100890 25360 101897
rect 25520 101897 28550 101920
rect 25520 100890 25543 101897
rect 25337 99890 25543 100890
rect 25337 98913 25360 99890
rect 22330 98890 25360 98913
rect 25520 98913 25543 99890
rect 28527 100890 28550 101897
rect 28710 101897 31740 101920
rect 28710 100890 28733 101897
rect 28527 99890 28733 100890
rect 28527 98913 28550 99890
rect 25520 98890 28550 98913
rect 28710 98913 28733 99890
rect 31717 100890 31740 101897
rect 31900 101897 34930 101920
rect 31900 100890 31923 101897
rect 31717 99890 31923 100890
rect 31717 98913 31740 99890
rect 28710 98890 31740 98913
rect 31900 98913 31923 99890
rect 34907 100890 34930 101897
rect 35090 101897 38120 101920
rect 35090 100890 35113 101897
rect 34907 99890 35113 100890
rect 34907 98913 34930 99890
rect 31900 98890 34930 98913
rect 35090 98913 35113 99890
rect 38097 100890 38120 101897
rect 38280 101897 41310 101920
rect 38280 100890 38303 101897
rect 38097 99890 38303 100890
rect 38097 98913 38120 99890
rect 35090 98890 38120 98913
rect 38280 98913 38303 99890
rect 41287 100890 41310 101897
rect 41470 101897 44500 101920
rect 41470 100890 41493 101897
rect 41287 99890 41493 100890
rect 41287 98913 41310 99890
rect 38280 98890 41310 98913
rect 41470 98913 41493 99890
rect 44477 100890 44500 101897
rect 44660 101897 47690 101920
rect 44660 100890 44683 101897
rect 44477 99890 44683 100890
rect 44477 98913 44500 99890
rect 41470 98890 44500 98913
rect 44660 98913 44683 99890
rect 47667 100890 47690 101897
rect 47850 101897 50880 101920
rect 47850 100890 47873 101897
rect 47667 99890 47873 100890
rect 47667 98913 47690 99890
rect 44660 98890 47690 98913
rect 47850 98913 47873 99890
rect 50857 100890 50880 101897
rect 51040 101897 54070 101920
rect 51040 100890 51063 101897
rect 50857 99890 51063 100890
rect 50857 98913 50880 99890
rect 47850 98890 50880 98913
rect 51040 98913 51063 99890
rect 54047 100890 54070 101897
rect 54230 101897 57260 101920
rect 54230 100890 54253 101897
rect 54047 99890 54253 100890
rect 54047 98913 54070 99890
rect 51040 98890 54070 98913
rect 54230 98913 54253 99890
rect 57237 100890 57260 101897
rect 57420 101897 60450 101920
rect 57420 100890 57443 101897
rect 57237 99890 57443 100890
rect 57237 98913 57260 99890
rect 54230 98890 57260 98913
rect 57420 98913 57443 99890
rect 60427 100890 60450 101897
rect 60610 101897 63640 101920
rect 60610 100890 60633 101897
rect 60427 99890 60633 100890
rect 60427 98913 60450 99890
rect 57420 98890 60450 98913
rect 60610 98913 60633 99890
rect 63617 100890 63640 101897
rect 63800 101897 66830 101920
rect 63800 100890 63823 101897
rect 63617 99890 63823 100890
rect 63617 98913 63640 99890
rect 60610 98890 63640 98913
rect 63800 98913 63823 99890
rect 66807 100890 66830 101897
rect 66990 101897 70020 101920
rect 66990 100890 67013 101897
rect 66807 99890 67013 100890
rect 66807 98913 66830 99890
rect 63800 98890 66830 98913
rect 66990 98913 67013 99890
rect 69997 100890 70020 101897
rect 70180 101897 73210 101920
rect 70180 100890 70203 101897
rect 69997 99890 70203 100890
rect 69997 98913 70020 99890
rect 66990 98890 70020 98913
rect 70180 98913 70203 99890
rect 73187 100890 73210 101897
rect 73370 101897 76400 101920
rect 73370 100890 73393 101897
rect 73187 99890 73393 100890
rect 73187 98913 73210 99890
rect 70180 98890 73210 98913
rect 73370 98913 73393 99890
rect 76377 100890 76400 101897
rect 76560 101897 79590 101920
rect 76560 100890 76583 101897
rect 76377 99890 76583 100890
rect 76377 98913 76400 99890
rect 73370 98890 76400 98913
rect 76560 98913 76583 99890
rect 79567 100890 79590 101897
rect 79750 101897 82780 101920
rect 79750 100890 79773 101897
rect 79567 99890 79773 100890
rect 79567 98913 79590 99890
rect 76560 98890 79590 98913
rect 79750 98913 79773 99890
rect 82757 100890 82780 101897
rect 82940 101897 85970 101920
rect 82940 100890 82963 101897
rect 82757 99890 82963 100890
rect 82757 98913 82780 99890
rect 79750 98890 82780 98913
rect 82940 98913 82963 99890
rect 85947 100890 85970 101897
rect 86130 101897 89160 101920
rect 86130 100890 86153 101897
rect 85947 99890 86153 100890
rect 85947 98913 85970 99890
rect 82940 98890 85970 98913
rect 86130 98913 86153 99890
rect 89137 100890 89160 101897
rect 89320 101897 92350 101920
rect 89320 100890 89343 101897
rect 89137 99890 89343 100890
rect 89137 98913 89160 99890
rect 86130 98890 89160 98913
rect 89320 98913 89343 99890
rect 92327 100890 92350 101897
rect 92510 101897 95540 101920
rect 92510 100890 92533 101897
rect 92327 99890 92533 100890
rect 92327 98913 92350 99890
rect 89320 98890 92350 98913
rect 92510 98913 92533 99890
rect 95517 100890 95540 101897
rect 95700 101897 98730 101920
rect 95700 100890 95723 101897
rect 95517 99890 95723 100890
rect 95517 98913 95540 99890
rect 92510 98890 95540 98913
rect 95700 98913 95723 99890
rect 98707 100890 98730 101897
rect 98890 101897 101920 101920
rect 98890 100890 98913 101897
rect 98707 99890 98913 100890
rect 98707 98913 98730 99890
rect 95700 98890 98730 98913
rect 98890 98913 98913 99890
rect 101897 100890 101920 101897
rect 102080 101897 105110 101920
rect 102080 100890 102103 101897
rect 101897 99890 102103 100890
rect 101897 98913 101920 99890
rect 98890 98890 101920 98913
rect 102080 98913 102103 99890
rect 105087 100890 105110 101897
rect 105270 101897 108300 101920
rect 105270 100890 105293 101897
rect 105087 99890 105293 100890
rect 105087 98913 105110 99890
rect 102080 98890 105110 98913
rect 105270 98913 105293 99890
rect 108277 100890 108300 101897
rect 108460 101897 111490 101920
rect 108460 100890 108483 101897
rect 108277 99890 108483 100890
rect 108277 98913 108300 99890
rect 105270 98890 108300 98913
rect 108460 98913 108483 99890
rect 111467 100890 111490 101897
rect 111650 101897 114680 101920
rect 111650 100890 111673 101897
rect 111467 99890 111673 100890
rect 111467 98913 111490 99890
rect 108460 98890 111490 98913
rect 111650 98913 111673 99890
rect 114657 100890 114680 101897
rect 114840 101897 117870 101920
rect 114840 100890 114863 101897
rect 114657 99890 114863 100890
rect 114657 98913 114680 99890
rect 111650 98890 114680 98913
rect 114840 98913 114863 99890
rect 117847 100890 117870 101897
rect 118030 101897 121060 101920
rect 118030 100890 118053 101897
rect 117847 99890 118053 100890
rect 117847 98913 117870 99890
rect 114840 98890 117870 98913
rect 118030 98913 118053 99890
rect 121037 100890 121060 101897
rect 121220 101897 124250 101920
rect 121220 100890 121243 101897
rect 121037 99890 121243 100890
rect 121037 98913 121060 99890
rect 118030 98890 121060 98913
rect 121220 98913 121243 99890
rect 124227 100890 124250 101897
rect 124410 101897 127440 101920
rect 124410 100890 124433 101897
rect 124227 99890 124433 100890
rect 124227 98913 124250 99890
rect 121220 98890 124250 98913
rect 124410 98913 124433 99890
rect 127417 100890 127440 101897
rect 127600 101897 130630 101920
rect 127600 100890 127623 101897
rect 127417 99890 127623 100890
rect 127417 98913 127440 99890
rect 124410 98890 127440 98913
rect 127600 98913 127623 99890
rect 130607 100890 130630 101897
rect 130790 101897 133820 101920
rect 130790 100890 130813 101897
rect 130607 99890 130813 100890
rect 130607 98913 130630 99890
rect 127600 98890 130630 98913
rect 130790 98913 130813 99890
rect 133797 100890 133820 101897
rect 133980 101897 137010 101920
rect 133980 100890 134003 101897
rect 133797 99890 134003 100890
rect 133797 98913 133820 99890
rect 130790 98890 133820 98913
rect 133980 98913 134003 99890
rect 136987 100890 137010 101897
rect 136987 99890 137170 100890
rect 136987 98913 137010 99890
rect 133980 98890 137010 98913
rect 1000 98730 2000 98890
rect 4190 98730 5190 98890
rect 7380 98730 8380 98890
rect 10570 98730 11570 98890
rect 13760 98730 14760 98890
rect 16950 98730 17950 98890
rect 20140 98730 21140 98890
rect 23330 98730 24330 98890
rect 26520 98730 27520 98890
rect 29710 98730 30710 98890
rect 32900 98730 33900 98890
rect 36090 98730 37090 98890
rect 39280 98730 40280 98890
rect 42470 98730 43470 98890
rect 45660 98730 46660 98890
rect 48850 98730 49850 98890
rect 52040 98730 53040 98890
rect 55230 98730 56230 98890
rect 58420 98730 59420 98890
rect 61610 98730 62610 98890
rect 64800 98730 65800 98890
rect 67990 98730 68990 98890
rect 71180 98730 72180 98890
rect 74370 98730 75370 98890
rect 77560 98730 78560 98890
rect 80750 98730 81750 98890
rect 83940 98730 84940 98890
rect 87130 98730 88130 98890
rect 90320 98730 91320 98890
rect 93510 98730 94510 98890
rect 96700 98730 97700 98890
rect 99890 98730 100890 98890
rect 103080 98730 104080 98890
rect 106270 98730 107270 98890
rect 109460 98730 110460 98890
rect 112650 98730 113650 98890
rect 115840 98730 116840 98890
rect 119030 98730 120030 98890
rect 122220 98730 123220 98890
rect 125410 98730 126410 98890
rect 128600 98730 129600 98890
rect 131790 98730 132790 98890
rect 134980 98730 135980 98890
rect 0 98689 3030 98730
rect 3190 98689 6220 98730
rect 6380 98689 9410 98730
rect 0 98639 9410 98689
rect 0 79839 50 98639
rect 9320 97700 9410 98639
rect 9570 98707 12600 98730
rect 9570 97700 9593 98707
rect 9320 96700 9593 97700
rect 9320 95700 9410 96700
rect 9570 95723 9593 96700
rect 12577 97700 12600 98707
rect 12760 98707 15790 98730
rect 12760 97700 12783 98707
rect 12577 96700 12783 97700
rect 12577 95723 12600 96700
rect 9570 95700 12600 95723
rect 12760 95723 12783 96700
rect 15767 97700 15790 98707
rect 15950 98707 18980 98730
rect 15950 97700 15973 98707
rect 15767 96700 15973 97700
rect 15767 95723 15790 96700
rect 12760 95700 15790 95723
rect 15950 95723 15973 96700
rect 18957 97700 18980 98707
rect 19140 98707 22170 98730
rect 19140 97700 19163 98707
rect 18957 96700 19163 97700
rect 18957 95723 18980 96700
rect 15950 95700 18980 95723
rect 19140 95723 19163 96700
rect 22147 97700 22170 98707
rect 22330 98707 25360 98730
rect 22330 97700 22353 98707
rect 22147 96700 22353 97700
rect 22147 95723 22170 96700
rect 19140 95700 22170 95723
rect 22330 95723 22353 96700
rect 25337 97700 25360 98707
rect 25520 98707 28550 98730
rect 25520 97700 25543 98707
rect 25337 96700 25543 97700
rect 25337 95723 25360 96700
rect 22330 95700 25360 95723
rect 25520 95723 25543 96700
rect 28527 97700 28550 98707
rect 28710 98707 31740 98730
rect 28710 97700 28733 98707
rect 28527 96700 28733 97700
rect 28527 95723 28550 96700
rect 25520 95700 28550 95723
rect 28710 95723 28733 96700
rect 31717 97700 31740 98707
rect 31900 98707 34930 98730
rect 31900 97700 31923 98707
rect 31717 96700 31923 97700
rect 31717 95723 31740 96700
rect 28710 95700 31740 95723
rect 31900 95723 31923 96700
rect 34907 97700 34930 98707
rect 35090 98707 38120 98730
rect 35090 97700 35113 98707
rect 34907 96700 35113 97700
rect 34907 95723 34930 96700
rect 31900 95700 34930 95723
rect 35090 95723 35113 96700
rect 38097 97700 38120 98707
rect 38280 98707 41310 98730
rect 38280 97700 38303 98707
rect 38097 96700 38303 97700
rect 38097 95723 38120 96700
rect 35090 95700 38120 95723
rect 38280 95723 38303 96700
rect 41287 97700 41310 98707
rect 41470 98707 44500 98730
rect 41470 97700 41493 98707
rect 41287 96700 41493 97700
rect 41287 95723 41310 96700
rect 38280 95700 41310 95723
rect 41470 95723 41493 96700
rect 44477 97700 44500 98707
rect 44660 98707 47690 98730
rect 44660 97700 44683 98707
rect 44477 96700 44683 97700
rect 44477 95723 44500 96700
rect 41470 95700 44500 95723
rect 44660 95723 44683 96700
rect 47667 97700 47690 98707
rect 47850 98707 50880 98730
rect 47850 97700 47873 98707
rect 47667 96700 47873 97700
rect 47667 95723 47690 96700
rect 44660 95700 47690 95723
rect 47850 95723 47873 96700
rect 50857 97700 50880 98707
rect 51040 98707 54070 98730
rect 51040 97700 51063 98707
rect 50857 96700 51063 97700
rect 50857 95723 50880 96700
rect 47850 95700 50880 95723
rect 51040 95723 51063 96700
rect 54047 97700 54070 98707
rect 54230 98707 57260 98730
rect 54230 97700 54253 98707
rect 54047 96700 54253 97700
rect 54047 95723 54070 96700
rect 51040 95700 54070 95723
rect 54230 95723 54253 96700
rect 57237 97700 57260 98707
rect 57420 98707 60450 98730
rect 57420 97700 57443 98707
rect 57237 96700 57443 97700
rect 57237 95723 57260 96700
rect 54230 95700 57260 95723
rect 57420 95723 57443 96700
rect 60427 97700 60450 98707
rect 60610 98707 63640 98730
rect 60610 97700 60633 98707
rect 60427 96700 60633 97700
rect 60427 95723 60450 96700
rect 57420 95700 60450 95723
rect 60610 95723 60633 96700
rect 63617 97700 63640 98707
rect 63800 98707 66830 98730
rect 63800 97700 63823 98707
rect 63617 96700 63823 97700
rect 63617 95723 63640 96700
rect 60610 95700 63640 95723
rect 63800 95723 63823 96700
rect 66807 97700 66830 98707
rect 66990 98707 70020 98730
rect 66990 97700 67013 98707
rect 66807 96700 67013 97700
rect 66807 95723 66830 96700
rect 63800 95700 66830 95723
rect 66990 95723 67013 96700
rect 69997 97700 70020 98707
rect 70180 98707 73210 98730
rect 70180 97700 70203 98707
rect 69997 96700 70203 97700
rect 69997 95723 70020 96700
rect 66990 95700 70020 95723
rect 70180 95723 70203 96700
rect 73187 97700 73210 98707
rect 73370 98707 76400 98730
rect 73370 97700 73393 98707
rect 73187 96700 73393 97700
rect 73187 95723 73210 96700
rect 70180 95700 73210 95723
rect 73370 95723 73393 96700
rect 76377 97700 76400 98707
rect 76560 98707 79590 98730
rect 76560 97700 76583 98707
rect 76377 96700 76583 97700
rect 76377 95723 76400 96700
rect 73370 95700 76400 95723
rect 76560 95723 76583 96700
rect 79567 97700 79590 98707
rect 79750 98707 82780 98730
rect 79750 97700 79773 98707
rect 79567 96700 79773 97700
rect 79567 95723 79590 96700
rect 76560 95700 79590 95723
rect 79750 95723 79773 96700
rect 82757 97700 82780 98707
rect 82940 98707 85970 98730
rect 82940 97700 82963 98707
rect 82757 96700 82963 97700
rect 82757 95723 82780 96700
rect 79750 95700 82780 95723
rect 82940 95723 82963 96700
rect 85947 97700 85970 98707
rect 86130 98707 89160 98730
rect 86130 97700 86153 98707
rect 85947 96700 86153 97700
rect 85947 95723 85970 96700
rect 82940 95700 85970 95723
rect 86130 95723 86153 96700
rect 89137 97700 89160 98707
rect 89320 98707 92350 98730
rect 89320 97700 89343 98707
rect 89137 96700 89343 97700
rect 89137 95723 89160 96700
rect 86130 95700 89160 95723
rect 89320 95723 89343 96700
rect 92327 97700 92350 98707
rect 92510 98707 95540 98730
rect 92510 97700 92533 98707
rect 92327 96700 92533 97700
rect 92327 95723 92350 96700
rect 89320 95700 92350 95723
rect 92510 95723 92533 96700
rect 95517 97700 95540 98707
rect 95700 98707 98730 98730
rect 95700 97700 95723 98707
rect 95517 96700 95723 97700
rect 95517 95723 95540 96700
rect 92510 95700 95540 95723
rect 95700 95723 95723 96700
rect 98707 97700 98730 98707
rect 98890 98707 101920 98730
rect 98890 97700 98913 98707
rect 98707 96700 98913 97700
rect 98707 95723 98730 96700
rect 95700 95700 98730 95723
rect 98890 95723 98913 96700
rect 101897 97700 101920 98707
rect 102080 98707 105110 98730
rect 102080 97700 102103 98707
rect 101897 96700 102103 97700
rect 101897 95723 101920 96700
rect 98890 95700 101920 95723
rect 102080 95723 102103 96700
rect 105087 97700 105110 98707
rect 105270 98707 108300 98730
rect 105270 97700 105293 98707
rect 105087 96700 105293 97700
rect 105087 95723 105110 96700
rect 102080 95700 105110 95723
rect 105270 95723 105293 96700
rect 108277 97700 108300 98707
rect 108460 98707 111490 98730
rect 108460 97700 108483 98707
rect 108277 96700 108483 97700
rect 108277 95723 108300 96700
rect 105270 95700 108300 95723
rect 108460 95723 108483 96700
rect 111467 97700 111490 98707
rect 111650 98707 114680 98730
rect 111650 97700 111673 98707
rect 111467 96700 111673 97700
rect 111467 95723 111490 96700
rect 108460 95700 111490 95723
rect 111650 95723 111673 96700
rect 114657 97700 114680 98707
rect 114840 98707 117870 98730
rect 114840 97700 114863 98707
rect 114657 96700 114863 97700
rect 114657 95723 114680 96700
rect 111650 95700 114680 95723
rect 114840 95723 114863 96700
rect 117847 97700 117870 98707
rect 118030 98707 121060 98730
rect 118030 97700 118053 98707
rect 117847 96700 118053 97700
rect 117847 95723 117870 96700
rect 114840 95700 117870 95723
rect 118030 95723 118053 96700
rect 121037 97700 121060 98707
rect 121220 98707 124250 98730
rect 121220 97700 121243 98707
rect 121037 96700 121243 97700
rect 121037 95723 121060 96700
rect 118030 95700 121060 95723
rect 121220 95723 121243 96700
rect 124227 97700 124250 98707
rect 124410 98707 127440 98730
rect 124410 97700 124433 98707
rect 124227 96700 124433 97700
rect 124227 95723 124250 96700
rect 121220 95700 124250 95723
rect 124410 95723 124433 96700
rect 127417 97700 127440 98707
rect 127600 98707 130630 98730
rect 127600 97700 127623 98707
rect 127417 96700 127623 97700
rect 127417 95723 127440 96700
rect 124410 95700 127440 95723
rect 127600 95723 127623 96700
rect 130607 97700 130630 98707
rect 130790 98707 133820 98730
rect 130790 97700 130813 98707
rect 130607 96700 130813 97700
rect 130607 95723 130630 96700
rect 127600 95700 130630 95723
rect 130790 95723 130813 96700
rect 133797 97700 133820 98707
rect 133980 98707 137010 98730
rect 133980 97700 134003 98707
rect 133797 96700 134003 97700
rect 133797 95723 133820 96700
rect 130790 95700 133820 95723
rect 133980 95723 134003 96700
rect 136987 97700 137010 98707
rect 136987 96700 137170 97700
rect 136987 95723 137010 96700
rect 133980 95700 137010 95723
rect 9320 95540 9370 95700
rect 10570 95540 11570 95700
rect 13760 95540 14760 95700
rect 16950 95540 17950 95700
rect 20140 95540 21140 95700
rect 23330 95540 24330 95700
rect 26520 95540 27520 95700
rect 29710 95540 30710 95700
rect 32900 95540 33900 95700
rect 36090 95540 37090 95700
rect 39280 95540 40280 95700
rect 42470 95540 43470 95700
rect 45660 95540 46660 95700
rect 48850 95540 49850 95700
rect 52040 95540 53040 95700
rect 55230 95540 56230 95700
rect 58420 95540 59420 95700
rect 61610 95540 62610 95700
rect 64800 95540 65800 95700
rect 67990 95540 68990 95700
rect 71180 95540 72180 95700
rect 74370 95540 75370 95700
rect 77560 95540 78560 95700
rect 80750 95540 81750 95700
rect 83940 95540 84940 95700
rect 87130 95540 88130 95700
rect 90320 95540 91320 95700
rect 93510 95540 94510 95700
rect 96700 95540 97700 95700
rect 99890 95540 100890 95700
rect 103080 95540 104080 95700
rect 106270 95540 107270 95700
rect 109460 95540 110460 95700
rect 112650 95540 113650 95700
rect 115840 95540 116840 95700
rect 119030 95540 120030 95700
rect 122220 95540 123220 95700
rect 125410 95540 126410 95700
rect 128600 95540 129600 95700
rect 131790 95540 132790 95700
rect 134980 95540 135980 95700
rect 9320 94510 9410 95540
rect 9570 95517 12600 95540
rect 9570 94510 9593 95517
rect 9320 93510 9593 94510
rect 9320 92510 9410 93510
rect 9570 92533 9593 93510
rect 12577 94510 12600 95517
rect 12760 95517 15790 95540
rect 12760 94510 12783 95517
rect 12577 93510 12783 94510
rect 12577 92533 12600 93510
rect 9570 92510 12600 92533
rect 12760 92533 12783 93510
rect 15767 94510 15790 95517
rect 15950 95517 18980 95540
rect 15950 94510 15973 95517
rect 15767 93510 15973 94510
rect 15767 92533 15790 93510
rect 12760 92510 15790 92533
rect 15950 92533 15973 93510
rect 18957 94510 18980 95517
rect 19140 95517 22170 95540
rect 19140 94510 19163 95517
rect 18957 93510 19163 94510
rect 18957 92533 18980 93510
rect 15950 92510 18980 92533
rect 19140 92533 19163 93510
rect 22147 94510 22170 95517
rect 22330 95517 25360 95540
rect 22330 94510 22353 95517
rect 22147 93510 22353 94510
rect 22147 92533 22170 93510
rect 19140 92510 22170 92533
rect 22330 92533 22353 93510
rect 25337 94510 25360 95517
rect 25520 95517 28550 95540
rect 25520 94510 25543 95517
rect 25337 93510 25543 94510
rect 25337 92533 25360 93510
rect 22330 92510 25360 92533
rect 25520 92533 25543 93510
rect 28527 94510 28550 95517
rect 28710 95517 31740 95540
rect 28710 94510 28733 95517
rect 28527 93510 28733 94510
rect 28527 92533 28550 93510
rect 25520 92510 28550 92533
rect 28710 92533 28733 93510
rect 31717 94510 31740 95517
rect 31900 95517 34930 95540
rect 31900 94510 31923 95517
rect 31717 93510 31923 94510
rect 31717 92533 31740 93510
rect 28710 92510 31740 92533
rect 31900 92533 31923 93510
rect 34907 94510 34930 95517
rect 35090 95517 38120 95540
rect 35090 94510 35113 95517
rect 34907 93510 35113 94510
rect 34907 92533 34930 93510
rect 31900 92510 34930 92533
rect 35090 92533 35113 93510
rect 38097 94510 38120 95517
rect 38280 95517 41310 95540
rect 38280 94510 38303 95517
rect 38097 93510 38303 94510
rect 38097 92533 38120 93510
rect 35090 92510 38120 92533
rect 38280 92533 38303 93510
rect 41287 94510 41310 95517
rect 41470 95517 44500 95540
rect 41470 94510 41493 95517
rect 41287 93510 41493 94510
rect 41287 92533 41310 93510
rect 38280 92510 41310 92533
rect 41470 92533 41493 93510
rect 44477 94510 44500 95517
rect 44660 95517 47690 95540
rect 44660 94510 44683 95517
rect 44477 93510 44683 94510
rect 44477 92533 44500 93510
rect 41470 92510 44500 92533
rect 44660 92533 44683 93510
rect 47667 94510 47690 95517
rect 47850 95517 50880 95540
rect 47850 94510 47873 95517
rect 47667 93510 47873 94510
rect 47667 92533 47690 93510
rect 44660 92510 47690 92533
rect 47850 92533 47873 93510
rect 50857 94510 50880 95517
rect 51040 95517 54070 95540
rect 51040 94510 51063 95517
rect 50857 93510 51063 94510
rect 50857 92533 50880 93510
rect 47850 92510 50880 92533
rect 51040 92533 51063 93510
rect 54047 94510 54070 95517
rect 54230 95517 57260 95540
rect 54230 94510 54253 95517
rect 54047 93510 54253 94510
rect 54047 92533 54070 93510
rect 51040 92510 54070 92533
rect 54230 92533 54253 93510
rect 57237 94510 57260 95517
rect 57420 95517 60450 95540
rect 57420 94510 57443 95517
rect 57237 93510 57443 94510
rect 57237 92533 57260 93510
rect 54230 92510 57260 92533
rect 57420 92533 57443 93510
rect 60427 94510 60450 95517
rect 60610 95517 63640 95540
rect 60610 94510 60633 95517
rect 60427 93510 60633 94510
rect 60427 92533 60450 93510
rect 57420 92510 60450 92533
rect 60610 92533 60633 93510
rect 63617 94510 63640 95517
rect 63800 95517 66830 95540
rect 63800 94510 63823 95517
rect 63617 93510 63823 94510
rect 63617 92533 63640 93510
rect 60610 92510 63640 92533
rect 63800 92533 63823 93510
rect 66807 94510 66830 95517
rect 66990 95517 70020 95540
rect 66990 94510 67013 95517
rect 66807 93510 67013 94510
rect 66807 92533 66830 93510
rect 63800 92510 66830 92533
rect 66990 92533 67013 93510
rect 69997 94510 70020 95517
rect 70180 95517 73210 95540
rect 70180 94510 70203 95517
rect 69997 93510 70203 94510
rect 69997 92533 70020 93510
rect 66990 92510 70020 92533
rect 70180 92533 70203 93510
rect 73187 94510 73210 95517
rect 73370 95517 76400 95540
rect 73370 94510 73393 95517
rect 73187 93510 73393 94510
rect 73187 92533 73210 93510
rect 70180 92510 73210 92533
rect 73370 92533 73393 93510
rect 76377 94510 76400 95517
rect 76560 95517 79590 95540
rect 76560 94510 76583 95517
rect 76377 93510 76583 94510
rect 76377 92533 76400 93510
rect 73370 92510 76400 92533
rect 76560 92533 76583 93510
rect 79567 94510 79590 95517
rect 79750 95517 82780 95540
rect 79750 94510 79773 95517
rect 79567 93510 79773 94510
rect 79567 92533 79590 93510
rect 76560 92510 79590 92533
rect 79750 92533 79773 93510
rect 82757 94510 82780 95517
rect 82940 95517 85970 95540
rect 82940 94510 82963 95517
rect 82757 93510 82963 94510
rect 82757 92533 82780 93510
rect 79750 92510 82780 92533
rect 82940 92533 82963 93510
rect 85947 94510 85970 95517
rect 86130 95517 89160 95540
rect 86130 94510 86153 95517
rect 85947 93510 86153 94510
rect 85947 92533 85970 93510
rect 82940 92510 85970 92533
rect 86130 92533 86153 93510
rect 89137 94510 89160 95517
rect 89320 95517 92350 95540
rect 89320 94510 89343 95517
rect 89137 93510 89343 94510
rect 89137 92533 89160 93510
rect 86130 92510 89160 92533
rect 89320 92533 89343 93510
rect 92327 94510 92350 95517
rect 92510 95517 95540 95540
rect 92510 94510 92533 95517
rect 92327 93510 92533 94510
rect 92327 92533 92350 93510
rect 89320 92510 92350 92533
rect 92510 92533 92533 93510
rect 95517 94510 95540 95517
rect 95700 95517 98730 95540
rect 95700 94510 95723 95517
rect 95517 93510 95723 94510
rect 95517 92533 95540 93510
rect 92510 92510 95540 92533
rect 95700 92533 95723 93510
rect 98707 94510 98730 95517
rect 98890 95517 101920 95540
rect 98890 94510 98913 95517
rect 98707 93510 98913 94510
rect 98707 92533 98730 93510
rect 95700 92510 98730 92533
rect 98890 92533 98913 93510
rect 101897 94510 101920 95517
rect 102080 95517 105110 95540
rect 102080 94510 102103 95517
rect 101897 93510 102103 94510
rect 101897 92533 101920 93510
rect 98890 92510 101920 92533
rect 102080 92533 102103 93510
rect 105087 94510 105110 95517
rect 105270 95517 108300 95540
rect 105270 94510 105293 95517
rect 105087 93510 105293 94510
rect 105087 92533 105110 93510
rect 102080 92510 105110 92533
rect 105270 92533 105293 93510
rect 108277 94510 108300 95517
rect 108460 95517 111490 95540
rect 108460 94510 108483 95517
rect 108277 93510 108483 94510
rect 108277 92533 108300 93510
rect 105270 92510 108300 92533
rect 108460 92533 108483 93510
rect 111467 94510 111490 95517
rect 111650 95517 114680 95540
rect 111650 94510 111673 95517
rect 111467 93510 111673 94510
rect 111467 92533 111490 93510
rect 108460 92510 111490 92533
rect 111650 92533 111673 93510
rect 114657 94510 114680 95517
rect 114840 95517 117870 95540
rect 114840 94510 114863 95517
rect 114657 93510 114863 94510
rect 114657 92533 114680 93510
rect 111650 92510 114680 92533
rect 114840 92533 114863 93510
rect 117847 94510 117870 95517
rect 118030 95517 121060 95540
rect 118030 94510 118053 95517
rect 117847 93510 118053 94510
rect 117847 92533 117870 93510
rect 114840 92510 117870 92533
rect 118030 92533 118053 93510
rect 121037 94510 121060 95517
rect 121220 95517 124250 95540
rect 121220 94510 121243 95517
rect 121037 93510 121243 94510
rect 121037 92533 121060 93510
rect 118030 92510 121060 92533
rect 121220 92533 121243 93510
rect 124227 94510 124250 95517
rect 124410 95517 127440 95540
rect 124410 94510 124433 95517
rect 124227 93510 124433 94510
rect 124227 92533 124250 93510
rect 121220 92510 124250 92533
rect 124410 92533 124433 93510
rect 127417 94510 127440 95517
rect 127600 95517 130630 95540
rect 127600 94510 127623 95517
rect 127417 93510 127623 94510
rect 127417 92533 127440 93510
rect 124410 92510 127440 92533
rect 127600 92533 127623 93510
rect 130607 94510 130630 95517
rect 130790 95517 133820 95540
rect 130790 94510 130813 95517
rect 130607 93510 130813 94510
rect 130607 92533 130630 93510
rect 127600 92510 130630 92533
rect 130790 92533 130813 93510
rect 133797 94510 133820 95517
rect 133980 95517 137010 95540
rect 133980 94510 134003 95517
rect 133797 93510 134003 94510
rect 133797 92533 133820 93510
rect 130790 92510 133820 92533
rect 133980 92533 134003 93510
rect 136987 94510 137010 95517
rect 136987 93510 137170 94510
rect 136987 92533 137010 93510
rect 133980 92510 137010 92533
rect 9320 92350 9370 92510
rect 10570 92350 11570 92510
rect 13760 92350 14760 92510
rect 16950 92350 17950 92510
rect 20140 92350 21140 92510
rect 23330 92350 24330 92510
rect 26520 92350 27520 92510
rect 29710 92350 30710 92510
rect 32900 92350 33900 92510
rect 36090 92350 37090 92510
rect 39280 92350 40280 92510
rect 42470 92350 43470 92510
rect 45660 92350 46660 92510
rect 48850 92350 49850 92510
rect 52040 92350 53040 92510
rect 55230 92350 56230 92510
rect 58420 92350 59420 92510
rect 61610 92350 62610 92510
rect 64800 92350 65800 92510
rect 67990 92350 68990 92510
rect 71180 92350 72180 92510
rect 74370 92350 75370 92510
rect 77560 92350 78560 92510
rect 80750 92350 81750 92510
rect 83940 92350 84940 92510
rect 87130 92350 88130 92510
rect 90320 92350 91320 92510
rect 93510 92350 94510 92510
rect 96700 92350 97700 92510
rect 99890 92350 100890 92510
rect 103080 92350 104080 92510
rect 106270 92350 107270 92510
rect 109460 92350 110460 92510
rect 112650 92350 113650 92510
rect 115840 92350 116840 92510
rect 119030 92350 120030 92510
rect 122220 92350 123220 92510
rect 125410 92350 126410 92510
rect 128600 92350 129600 92510
rect 131790 92350 132790 92510
rect 134980 92350 135980 92510
rect 9320 91320 9410 92350
rect 9570 92327 12600 92350
rect 9570 91320 9593 92327
rect 9320 90320 9593 91320
rect 9320 89320 9410 90320
rect 9570 89343 9593 90320
rect 12577 91320 12600 92327
rect 12760 92327 15790 92350
rect 12760 91320 12783 92327
rect 12577 90320 12783 91320
rect 12577 89343 12600 90320
rect 9570 89320 12600 89343
rect 12760 89343 12783 90320
rect 15767 91320 15790 92327
rect 15950 92327 18980 92350
rect 15950 91320 15973 92327
rect 15767 90320 15973 91320
rect 15767 89343 15790 90320
rect 12760 89320 15790 89343
rect 15950 89343 15973 90320
rect 18957 91320 18980 92327
rect 19140 92327 22170 92350
rect 19140 91320 19163 92327
rect 18957 90320 19163 91320
rect 18957 89343 18980 90320
rect 15950 89320 18980 89343
rect 19140 89343 19163 90320
rect 22147 91320 22170 92327
rect 22330 92327 25360 92350
rect 22330 91320 22353 92327
rect 22147 90320 22353 91320
rect 22147 89343 22170 90320
rect 19140 89320 22170 89343
rect 22330 89343 22353 90320
rect 25337 91320 25360 92327
rect 25520 92327 28550 92350
rect 25520 91320 25543 92327
rect 25337 90320 25543 91320
rect 25337 89343 25360 90320
rect 22330 89320 25360 89343
rect 25520 89343 25543 90320
rect 28527 91320 28550 92327
rect 28710 92327 31740 92350
rect 28710 91320 28733 92327
rect 28527 90320 28733 91320
rect 28527 89343 28550 90320
rect 25520 89320 28550 89343
rect 28710 89343 28733 90320
rect 31717 91320 31740 92327
rect 31900 92327 34930 92350
rect 31900 91320 31923 92327
rect 31717 90320 31923 91320
rect 31717 89343 31740 90320
rect 28710 89320 31740 89343
rect 31900 89343 31923 90320
rect 34907 91320 34930 92327
rect 35090 92327 38120 92350
rect 35090 91320 35113 92327
rect 34907 90320 35113 91320
rect 34907 89343 34930 90320
rect 31900 89320 34930 89343
rect 35090 89343 35113 90320
rect 38097 91320 38120 92327
rect 38280 92327 41310 92350
rect 38280 91320 38303 92327
rect 38097 90320 38303 91320
rect 38097 89343 38120 90320
rect 35090 89320 38120 89343
rect 38280 89343 38303 90320
rect 41287 91320 41310 92327
rect 41470 92327 44500 92350
rect 41470 91320 41493 92327
rect 41287 90320 41493 91320
rect 41287 89343 41310 90320
rect 38280 89320 41310 89343
rect 41470 89343 41493 90320
rect 44477 91320 44500 92327
rect 44660 92327 47690 92350
rect 44660 91320 44683 92327
rect 44477 90320 44683 91320
rect 44477 89343 44500 90320
rect 41470 89320 44500 89343
rect 44660 89343 44683 90320
rect 47667 91320 47690 92327
rect 47850 92327 50880 92350
rect 47850 91320 47873 92327
rect 47667 90320 47873 91320
rect 47667 89343 47690 90320
rect 44660 89320 47690 89343
rect 47850 89343 47873 90320
rect 50857 91320 50880 92327
rect 51040 92327 54070 92350
rect 51040 91320 51063 92327
rect 50857 90320 51063 91320
rect 50857 89343 50880 90320
rect 47850 89320 50880 89343
rect 51040 89343 51063 90320
rect 54047 91320 54070 92327
rect 54230 92327 57260 92350
rect 54230 91320 54253 92327
rect 54047 90320 54253 91320
rect 54047 89343 54070 90320
rect 51040 89320 54070 89343
rect 54230 89343 54253 90320
rect 57237 91320 57260 92327
rect 57420 92327 60450 92350
rect 57420 91320 57443 92327
rect 57237 90320 57443 91320
rect 57237 89343 57260 90320
rect 54230 89320 57260 89343
rect 57420 89343 57443 90320
rect 60427 91320 60450 92327
rect 60610 92327 63640 92350
rect 60610 91320 60633 92327
rect 60427 90320 60633 91320
rect 60427 89343 60450 90320
rect 57420 89320 60450 89343
rect 60610 89343 60633 90320
rect 63617 91320 63640 92327
rect 63800 92327 66830 92350
rect 63800 91320 63823 92327
rect 63617 90320 63823 91320
rect 63617 89343 63640 90320
rect 60610 89320 63640 89343
rect 63800 89343 63823 90320
rect 66807 91320 66830 92327
rect 66990 92327 70020 92350
rect 66990 91320 67013 92327
rect 66807 90320 67013 91320
rect 66807 89343 66830 90320
rect 63800 89320 66830 89343
rect 66990 89343 67013 90320
rect 69997 91320 70020 92327
rect 70180 92327 73210 92350
rect 70180 91320 70203 92327
rect 69997 90320 70203 91320
rect 69997 89343 70020 90320
rect 66990 89320 70020 89343
rect 70180 89343 70203 90320
rect 73187 91320 73210 92327
rect 73370 92327 76400 92350
rect 73370 91320 73393 92327
rect 73187 90320 73393 91320
rect 73187 89343 73210 90320
rect 70180 89320 73210 89343
rect 73370 89343 73393 90320
rect 76377 91320 76400 92327
rect 76560 92327 79590 92350
rect 76560 91320 76583 92327
rect 76377 90320 76583 91320
rect 76377 89343 76400 90320
rect 73370 89320 76400 89343
rect 76560 89343 76583 90320
rect 79567 91320 79590 92327
rect 79750 92327 82780 92350
rect 79750 91320 79773 92327
rect 79567 90320 79773 91320
rect 79567 89343 79590 90320
rect 76560 89320 79590 89343
rect 79750 89343 79773 90320
rect 82757 91320 82780 92327
rect 82940 92327 85970 92350
rect 82940 91320 82963 92327
rect 82757 90320 82963 91320
rect 82757 89343 82780 90320
rect 79750 89320 82780 89343
rect 82940 89343 82963 90320
rect 85947 91320 85970 92327
rect 86130 92327 89160 92350
rect 86130 91320 86153 92327
rect 85947 90320 86153 91320
rect 85947 89343 85970 90320
rect 82940 89320 85970 89343
rect 86130 89343 86153 90320
rect 89137 91320 89160 92327
rect 89320 92327 92350 92350
rect 89320 91320 89343 92327
rect 89137 90320 89343 91320
rect 89137 89343 89160 90320
rect 86130 89320 89160 89343
rect 89320 89343 89343 90320
rect 92327 91320 92350 92327
rect 92510 92327 95540 92350
rect 92510 91320 92533 92327
rect 92327 90320 92533 91320
rect 92327 89343 92350 90320
rect 89320 89320 92350 89343
rect 92510 89343 92533 90320
rect 95517 91320 95540 92327
rect 95700 92327 98730 92350
rect 95700 91320 95723 92327
rect 95517 90320 95723 91320
rect 95517 89343 95540 90320
rect 92510 89320 95540 89343
rect 95700 89343 95723 90320
rect 98707 91320 98730 92327
rect 98890 92327 101920 92350
rect 98890 91320 98913 92327
rect 98707 90320 98913 91320
rect 98707 89343 98730 90320
rect 95700 89320 98730 89343
rect 98890 89343 98913 90320
rect 101897 91320 101920 92327
rect 102080 92327 105110 92350
rect 102080 91320 102103 92327
rect 101897 90320 102103 91320
rect 101897 89343 101920 90320
rect 98890 89320 101920 89343
rect 102080 89343 102103 90320
rect 105087 91320 105110 92327
rect 105270 92327 108300 92350
rect 105270 91320 105293 92327
rect 105087 90320 105293 91320
rect 105087 89343 105110 90320
rect 102080 89320 105110 89343
rect 105270 89343 105293 90320
rect 108277 91320 108300 92327
rect 108460 92327 111490 92350
rect 108460 91320 108483 92327
rect 108277 90320 108483 91320
rect 108277 89343 108300 90320
rect 105270 89320 108300 89343
rect 108460 89343 108483 90320
rect 111467 91320 111490 92327
rect 111650 92327 114680 92350
rect 111650 91320 111673 92327
rect 111467 90320 111673 91320
rect 111467 89343 111490 90320
rect 108460 89320 111490 89343
rect 111650 89343 111673 90320
rect 114657 91320 114680 92327
rect 114840 92327 117870 92350
rect 114840 91320 114863 92327
rect 114657 90320 114863 91320
rect 114657 89343 114680 90320
rect 111650 89320 114680 89343
rect 114840 89343 114863 90320
rect 117847 91320 117870 92327
rect 118030 92327 121060 92350
rect 118030 91320 118053 92327
rect 117847 90320 118053 91320
rect 117847 89343 117870 90320
rect 114840 89320 117870 89343
rect 118030 89343 118053 90320
rect 121037 91320 121060 92327
rect 121220 92327 124250 92350
rect 121220 91320 121243 92327
rect 121037 90320 121243 91320
rect 121037 89343 121060 90320
rect 118030 89320 121060 89343
rect 121220 89343 121243 90320
rect 124227 91320 124250 92327
rect 124410 92327 127440 92350
rect 124410 91320 124433 92327
rect 124227 90320 124433 91320
rect 124227 89343 124250 90320
rect 121220 89320 124250 89343
rect 124410 89343 124433 90320
rect 127417 91320 127440 92327
rect 127600 92327 130630 92350
rect 127600 91320 127623 92327
rect 127417 90320 127623 91320
rect 127417 89343 127440 90320
rect 124410 89320 127440 89343
rect 127600 89343 127623 90320
rect 130607 91320 130630 92327
rect 130790 92327 133820 92350
rect 130790 91320 130813 92327
rect 130607 90320 130813 91320
rect 130607 89343 130630 90320
rect 127600 89320 130630 89343
rect 130790 89343 130813 90320
rect 133797 91320 133820 92327
rect 133980 92327 137010 92350
rect 133980 91320 134003 92327
rect 133797 90320 134003 91320
rect 133797 89343 133820 90320
rect 130790 89320 133820 89343
rect 133980 89343 134003 90320
rect 136987 91320 137010 92327
rect 136987 90320 137170 91320
rect 136987 89343 137010 90320
rect 133980 89320 137010 89343
rect 9320 89160 9370 89320
rect 10570 89160 11570 89320
rect 13760 89160 14760 89320
rect 16950 89160 17950 89320
rect 20140 89160 21140 89320
rect 23330 89160 24330 89320
rect 26520 89160 27520 89320
rect 29710 89160 30710 89320
rect 32900 89160 33900 89320
rect 36090 89160 37090 89320
rect 39280 89160 40280 89320
rect 42470 89160 43470 89320
rect 45660 89160 46660 89320
rect 48850 89160 49850 89320
rect 52040 89160 53040 89320
rect 55230 89160 56230 89320
rect 58420 89160 59420 89320
rect 61610 89160 62610 89320
rect 64800 89160 65800 89320
rect 67990 89160 68990 89320
rect 71180 89160 72180 89320
rect 74370 89160 75370 89320
rect 77560 89160 78560 89320
rect 80750 89160 81750 89320
rect 83940 89160 84940 89320
rect 87130 89160 88130 89320
rect 90320 89160 91320 89320
rect 93510 89160 94510 89320
rect 96700 89160 97700 89320
rect 99890 89160 100890 89320
rect 103080 89160 104080 89320
rect 106270 89160 107270 89320
rect 109460 89160 110460 89320
rect 112650 89160 113650 89320
rect 115840 89160 116840 89320
rect 119030 89160 120030 89320
rect 122220 89160 123220 89320
rect 125410 89160 126410 89320
rect 128600 89160 129600 89320
rect 131790 89160 132790 89320
rect 134980 89160 135980 89320
rect 9320 88130 9410 89160
rect 9570 89137 12600 89160
rect 9570 88130 9593 89137
rect 9320 87130 9593 88130
rect 9320 86130 9410 87130
rect 9570 86153 9593 87130
rect 12577 88130 12600 89137
rect 12760 89137 15790 89160
rect 12760 88130 12783 89137
rect 12577 87130 12783 88130
rect 12577 86153 12600 87130
rect 9570 86130 12600 86153
rect 12760 86153 12783 87130
rect 15767 88130 15790 89137
rect 15950 89137 18980 89160
rect 15950 88130 15973 89137
rect 15767 87130 15973 88130
rect 15767 86153 15790 87130
rect 12760 86130 15790 86153
rect 15950 86153 15973 87130
rect 18957 88130 18980 89137
rect 19140 89137 22170 89160
rect 19140 88130 19163 89137
rect 18957 87130 19163 88130
rect 18957 86153 18980 87130
rect 15950 86130 18980 86153
rect 19140 86153 19163 87130
rect 22147 88130 22170 89137
rect 22330 89137 25360 89160
rect 22330 88130 22353 89137
rect 22147 87130 22353 88130
rect 22147 86153 22170 87130
rect 19140 86130 22170 86153
rect 22330 86153 22353 87130
rect 25337 88130 25360 89137
rect 25520 89137 28550 89160
rect 25520 88130 25543 89137
rect 25337 87130 25543 88130
rect 25337 86153 25360 87130
rect 22330 86130 25360 86153
rect 25520 86153 25543 87130
rect 28527 88130 28550 89137
rect 28710 89137 31740 89160
rect 28710 88130 28733 89137
rect 28527 87130 28733 88130
rect 28527 86153 28550 87130
rect 25520 86130 28550 86153
rect 28710 86153 28733 87130
rect 31717 88130 31740 89137
rect 31900 89137 34930 89160
rect 31900 88130 31923 89137
rect 31717 87130 31923 88130
rect 31717 86153 31740 87130
rect 28710 86130 31740 86153
rect 31900 86153 31923 87130
rect 34907 88130 34930 89137
rect 35090 89137 38120 89160
rect 35090 88130 35113 89137
rect 34907 87130 35113 88130
rect 34907 86153 34930 87130
rect 31900 86130 34930 86153
rect 35090 86153 35113 87130
rect 38097 88130 38120 89137
rect 38280 89137 41310 89160
rect 38280 88130 38303 89137
rect 38097 87130 38303 88130
rect 38097 86153 38120 87130
rect 35090 86130 38120 86153
rect 38280 86153 38303 87130
rect 41287 88130 41310 89137
rect 41470 89137 44500 89160
rect 41470 88130 41493 89137
rect 41287 87130 41493 88130
rect 41287 86153 41310 87130
rect 38280 86130 41310 86153
rect 41470 86153 41493 87130
rect 44477 88130 44500 89137
rect 44660 89137 47690 89160
rect 44660 88130 44683 89137
rect 44477 87130 44683 88130
rect 44477 86153 44500 87130
rect 41470 86130 44500 86153
rect 44660 86153 44683 87130
rect 47667 88130 47690 89137
rect 47850 89137 50880 89160
rect 47850 88130 47873 89137
rect 47667 87130 47873 88130
rect 47667 86153 47690 87130
rect 44660 86130 47690 86153
rect 47850 86153 47873 87130
rect 50857 88130 50880 89137
rect 51040 89137 54070 89160
rect 51040 88130 51063 89137
rect 50857 87130 51063 88130
rect 50857 86153 50880 87130
rect 47850 86130 50880 86153
rect 51040 86153 51063 87130
rect 54047 88130 54070 89137
rect 54230 89137 57260 89160
rect 54230 88130 54253 89137
rect 54047 87130 54253 88130
rect 54047 86153 54070 87130
rect 51040 86130 54070 86153
rect 54230 86153 54253 87130
rect 57237 88130 57260 89137
rect 57420 89137 60450 89160
rect 57420 88130 57443 89137
rect 57237 87130 57443 88130
rect 57237 86153 57260 87130
rect 54230 86130 57260 86153
rect 57420 86153 57443 87130
rect 60427 88130 60450 89137
rect 60610 89137 63640 89160
rect 60610 88130 60633 89137
rect 60427 87130 60633 88130
rect 60427 86153 60450 87130
rect 57420 86130 60450 86153
rect 60610 86153 60633 87130
rect 63617 88130 63640 89137
rect 63800 89137 66830 89160
rect 63800 88130 63823 89137
rect 63617 87130 63823 88130
rect 63617 86153 63640 87130
rect 60610 86130 63640 86153
rect 63800 86153 63823 87130
rect 66807 88130 66830 89137
rect 66990 89137 70020 89160
rect 66990 88130 67013 89137
rect 66807 87130 67013 88130
rect 66807 86153 66830 87130
rect 63800 86130 66830 86153
rect 66990 86153 67013 87130
rect 69997 88130 70020 89137
rect 70180 89137 73210 89160
rect 70180 88130 70203 89137
rect 69997 87130 70203 88130
rect 69997 86153 70020 87130
rect 66990 86130 70020 86153
rect 70180 86153 70203 87130
rect 73187 88130 73210 89137
rect 73370 89137 76400 89160
rect 73370 88130 73393 89137
rect 73187 87130 73393 88130
rect 73187 86153 73210 87130
rect 70180 86130 73210 86153
rect 73370 86153 73393 87130
rect 76377 88130 76400 89137
rect 76560 89137 79590 89160
rect 76560 88130 76583 89137
rect 76377 87130 76583 88130
rect 76377 86153 76400 87130
rect 73370 86130 76400 86153
rect 76560 86153 76583 87130
rect 79567 88130 79590 89137
rect 79750 89137 82780 89160
rect 79750 88130 79773 89137
rect 79567 87130 79773 88130
rect 79567 86153 79590 87130
rect 76560 86130 79590 86153
rect 79750 86153 79773 87130
rect 82757 88130 82780 89137
rect 82940 89137 85970 89160
rect 82940 88130 82963 89137
rect 82757 87130 82963 88130
rect 82757 86153 82780 87130
rect 79750 86130 82780 86153
rect 82940 86153 82963 87130
rect 85947 88130 85970 89137
rect 86130 89137 89160 89160
rect 86130 88130 86153 89137
rect 85947 87130 86153 88130
rect 85947 86153 85970 87130
rect 82940 86130 85970 86153
rect 86130 86153 86153 87130
rect 89137 88130 89160 89137
rect 89320 89137 92350 89160
rect 89320 88130 89343 89137
rect 89137 87130 89343 88130
rect 89137 86153 89160 87130
rect 86130 86130 89160 86153
rect 89320 86153 89343 87130
rect 92327 88130 92350 89137
rect 92510 89137 95540 89160
rect 92510 88130 92533 89137
rect 92327 87130 92533 88130
rect 92327 86153 92350 87130
rect 89320 86130 92350 86153
rect 92510 86153 92533 87130
rect 95517 88130 95540 89137
rect 95700 89137 98730 89160
rect 95700 88130 95723 89137
rect 95517 87130 95723 88130
rect 95517 86153 95540 87130
rect 92510 86130 95540 86153
rect 95700 86153 95723 87130
rect 98707 88130 98730 89137
rect 98890 89137 101920 89160
rect 98890 88130 98913 89137
rect 98707 87130 98913 88130
rect 98707 86153 98730 87130
rect 95700 86130 98730 86153
rect 98890 86153 98913 87130
rect 101897 88130 101920 89137
rect 102080 89137 105110 89160
rect 102080 88130 102103 89137
rect 101897 87130 102103 88130
rect 101897 86153 101920 87130
rect 98890 86130 101920 86153
rect 102080 86153 102103 87130
rect 105087 88130 105110 89137
rect 105270 89137 108300 89160
rect 105270 88130 105293 89137
rect 105087 87130 105293 88130
rect 105087 86153 105110 87130
rect 102080 86130 105110 86153
rect 105270 86153 105293 87130
rect 108277 88130 108300 89137
rect 108460 89137 111490 89160
rect 108460 88130 108483 89137
rect 108277 87130 108483 88130
rect 108277 86153 108300 87130
rect 105270 86130 108300 86153
rect 108460 86153 108483 87130
rect 111467 88130 111490 89137
rect 111650 89137 114680 89160
rect 111650 88130 111673 89137
rect 111467 87130 111673 88130
rect 111467 86153 111490 87130
rect 108460 86130 111490 86153
rect 111650 86153 111673 87130
rect 114657 88130 114680 89137
rect 114840 89137 117870 89160
rect 114840 88130 114863 89137
rect 114657 87130 114863 88130
rect 114657 86153 114680 87130
rect 111650 86130 114680 86153
rect 114840 86153 114863 87130
rect 117847 88130 117870 89137
rect 118030 89137 121060 89160
rect 118030 88130 118053 89137
rect 117847 87130 118053 88130
rect 117847 86153 117870 87130
rect 114840 86130 117870 86153
rect 118030 86153 118053 87130
rect 121037 88130 121060 89137
rect 121220 89137 124250 89160
rect 121220 88130 121243 89137
rect 121037 87130 121243 88130
rect 121037 86153 121060 87130
rect 118030 86130 121060 86153
rect 121220 86153 121243 87130
rect 124227 88130 124250 89137
rect 124410 89137 127440 89160
rect 124410 88130 124433 89137
rect 124227 87130 124433 88130
rect 124227 86153 124250 87130
rect 121220 86130 124250 86153
rect 124410 86153 124433 87130
rect 127417 88130 127440 89137
rect 127600 89137 130630 89160
rect 127600 88130 127623 89137
rect 127417 87130 127623 88130
rect 127417 86153 127440 87130
rect 124410 86130 127440 86153
rect 127600 86153 127623 87130
rect 130607 88130 130630 89137
rect 130790 89137 133820 89160
rect 130790 88130 130813 89137
rect 130607 87130 130813 88130
rect 130607 86153 130630 87130
rect 127600 86130 130630 86153
rect 130790 86153 130813 87130
rect 133797 88130 133820 89137
rect 133980 89137 137010 89160
rect 133980 88130 134003 89137
rect 133797 87130 134003 88130
rect 133797 86153 133820 87130
rect 130790 86130 133820 86153
rect 133980 86153 134003 87130
rect 136987 88130 137010 89137
rect 136987 87130 137170 88130
rect 136987 86153 137010 87130
rect 133980 86130 137010 86153
rect 9320 85970 9370 86130
rect 10570 85970 11570 86130
rect 13760 85970 14760 86130
rect 16950 85970 17950 86130
rect 20140 85970 21140 86130
rect 23330 85970 24330 86130
rect 26520 85970 27520 86130
rect 29710 85970 30710 86130
rect 32900 85970 33900 86130
rect 36090 85970 37090 86130
rect 39280 85970 40280 86130
rect 42470 85970 43470 86130
rect 45660 85970 46660 86130
rect 48850 85970 49850 86130
rect 52040 85970 53040 86130
rect 55230 85970 56230 86130
rect 58420 85970 59420 86130
rect 61610 85970 62610 86130
rect 64800 85970 65800 86130
rect 67990 85970 68990 86130
rect 71180 85970 72180 86130
rect 74370 85970 75370 86130
rect 77560 85970 78560 86130
rect 80750 85970 81750 86130
rect 83940 85970 84940 86130
rect 87130 85970 88130 86130
rect 90320 85970 91320 86130
rect 93510 85970 94510 86130
rect 96700 85970 97700 86130
rect 99890 85970 100890 86130
rect 103080 85970 104080 86130
rect 106270 85970 107270 86130
rect 109460 85970 110460 86130
rect 112650 85970 113650 86130
rect 115840 85970 116840 86130
rect 119030 85970 120030 86130
rect 122220 85970 123220 86130
rect 125410 85970 126410 86130
rect 128600 85970 129600 86130
rect 131790 85970 132790 86130
rect 134980 85970 135980 86130
rect 9320 84940 9410 85970
rect 9570 85947 12600 85970
rect 9570 84940 9593 85947
rect 9320 83940 9593 84940
rect 9320 82940 9410 83940
rect 9570 82963 9593 83940
rect 12577 84940 12600 85947
rect 12760 85947 15790 85970
rect 12760 84940 12783 85947
rect 12577 83940 12783 84940
rect 12577 82963 12600 83940
rect 9570 82940 12600 82963
rect 12760 82963 12783 83940
rect 15767 84940 15790 85947
rect 15950 85947 18980 85970
rect 15950 84940 15973 85947
rect 15767 83940 15973 84940
rect 15767 82963 15790 83940
rect 12760 82940 15790 82963
rect 15950 82963 15973 83940
rect 18957 84940 18980 85947
rect 19140 85947 22170 85970
rect 19140 84940 19163 85947
rect 18957 83940 19163 84940
rect 18957 82963 18980 83940
rect 15950 82940 18980 82963
rect 19140 82963 19163 83940
rect 22147 84940 22170 85947
rect 22330 85947 25360 85970
rect 22330 84940 22353 85947
rect 22147 83940 22353 84940
rect 22147 82963 22170 83940
rect 19140 82940 22170 82963
rect 22330 82963 22353 83940
rect 25337 84940 25360 85947
rect 25520 85947 28550 85970
rect 25520 84940 25543 85947
rect 25337 83940 25543 84940
rect 25337 82963 25360 83940
rect 22330 82940 25360 82963
rect 25520 82963 25543 83940
rect 28527 84940 28550 85947
rect 28710 85947 31740 85970
rect 28710 84940 28733 85947
rect 28527 83940 28733 84940
rect 28527 82963 28550 83940
rect 25520 82940 28550 82963
rect 28710 82963 28733 83940
rect 31717 84940 31740 85947
rect 31900 85947 34930 85970
rect 31900 84940 31923 85947
rect 31717 83940 31923 84940
rect 31717 82963 31740 83940
rect 28710 82940 31740 82963
rect 31900 82963 31923 83940
rect 34907 84940 34930 85947
rect 35090 85947 38120 85970
rect 35090 84940 35113 85947
rect 34907 83940 35113 84940
rect 34907 82963 34930 83940
rect 31900 82940 34930 82963
rect 35090 82963 35113 83940
rect 38097 84940 38120 85947
rect 38280 85947 41310 85970
rect 38280 84940 38303 85947
rect 38097 83940 38303 84940
rect 38097 82963 38120 83940
rect 35090 82940 38120 82963
rect 38280 82963 38303 83940
rect 41287 84940 41310 85947
rect 41470 85947 44500 85970
rect 41470 84940 41493 85947
rect 41287 83940 41493 84940
rect 41287 82963 41310 83940
rect 38280 82940 41310 82963
rect 41470 82963 41493 83940
rect 44477 84940 44500 85947
rect 44660 85947 47690 85970
rect 44660 84940 44683 85947
rect 44477 83940 44683 84940
rect 44477 82963 44500 83940
rect 41470 82940 44500 82963
rect 44660 82963 44683 83940
rect 47667 84940 47690 85947
rect 47850 85947 50880 85970
rect 47850 84940 47873 85947
rect 47667 83940 47873 84940
rect 47667 82963 47690 83940
rect 44660 82940 47690 82963
rect 47850 82963 47873 83940
rect 50857 84940 50880 85947
rect 51040 85947 54070 85970
rect 51040 84940 51063 85947
rect 50857 83940 51063 84940
rect 50857 82963 50880 83940
rect 47850 82940 50880 82963
rect 51040 82963 51063 83940
rect 54047 84940 54070 85947
rect 54230 85947 57260 85970
rect 54230 84940 54253 85947
rect 54047 83940 54253 84940
rect 54047 82963 54070 83940
rect 51040 82940 54070 82963
rect 54230 82963 54253 83940
rect 57237 84940 57260 85947
rect 57420 85947 60450 85970
rect 57420 84940 57443 85947
rect 57237 83940 57443 84940
rect 57237 82963 57260 83940
rect 54230 82940 57260 82963
rect 57420 82963 57443 83940
rect 60427 84940 60450 85947
rect 60610 85947 63640 85970
rect 60610 84940 60633 85947
rect 60427 83940 60633 84940
rect 60427 82963 60450 83940
rect 57420 82940 60450 82963
rect 60610 82963 60633 83940
rect 63617 84940 63640 85947
rect 63800 85947 66830 85970
rect 63800 84940 63823 85947
rect 63617 83940 63823 84940
rect 63617 82963 63640 83940
rect 60610 82940 63640 82963
rect 63800 82963 63823 83940
rect 66807 84940 66830 85947
rect 66990 85947 70020 85970
rect 66990 84940 67013 85947
rect 66807 83940 67013 84940
rect 66807 82963 66830 83940
rect 63800 82940 66830 82963
rect 66990 82963 67013 83940
rect 69997 84940 70020 85947
rect 70180 85947 73210 85970
rect 70180 84940 70203 85947
rect 69997 83940 70203 84940
rect 69997 82963 70020 83940
rect 66990 82940 70020 82963
rect 70180 82963 70203 83940
rect 73187 84940 73210 85947
rect 73370 85947 76400 85970
rect 73370 84940 73393 85947
rect 73187 83940 73393 84940
rect 73187 82963 73210 83940
rect 70180 82940 73210 82963
rect 73370 82963 73393 83940
rect 76377 84940 76400 85947
rect 76560 85947 79590 85970
rect 76560 84940 76583 85947
rect 76377 83940 76583 84940
rect 76377 82963 76400 83940
rect 73370 82940 76400 82963
rect 76560 82963 76583 83940
rect 79567 84940 79590 85947
rect 79750 85947 82780 85970
rect 79750 84940 79773 85947
rect 79567 83940 79773 84940
rect 79567 82963 79590 83940
rect 76560 82940 79590 82963
rect 79750 82963 79773 83940
rect 82757 84940 82780 85947
rect 82940 85947 85970 85970
rect 82940 84940 82963 85947
rect 82757 83940 82963 84940
rect 82757 82963 82780 83940
rect 79750 82940 82780 82963
rect 82940 82963 82963 83940
rect 85947 84940 85970 85947
rect 86130 85947 89160 85970
rect 86130 84940 86153 85947
rect 85947 83940 86153 84940
rect 85947 82963 85970 83940
rect 82940 82940 85970 82963
rect 86130 82963 86153 83940
rect 89137 84940 89160 85947
rect 89320 85947 92350 85970
rect 89320 84940 89343 85947
rect 89137 83940 89343 84940
rect 89137 82963 89160 83940
rect 86130 82940 89160 82963
rect 89320 82963 89343 83940
rect 92327 84940 92350 85947
rect 92510 85947 95540 85970
rect 92510 84940 92533 85947
rect 92327 83940 92533 84940
rect 92327 82963 92350 83940
rect 89320 82940 92350 82963
rect 92510 82963 92533 83940
rect 95517 84940 95540 85947
rect 95700 85947 98730 85970
rect 95700 84940 95723 85947
rect 95517 83940 95723 84940
rect 95517 82963 95540 83940
rect 92510 82940 95540 82963
rect 95700 82963 95723 83940
rect 98707 84940 98730 85947
rect 98890 85947 101920 85970
rect 98890 84940 98913 85947
rect 98707 83940 98913 84940
rect 98707 82963 98730 83940
rect 95700 82940 98730 82963
rect 98890 82963 98913 83940
rect 101897 84940 101920 85947
rect 102080 85947 105110 85970
rect 102080 84940 102103 85947
rect 101897 83940 102103 84940
rect 101897 82963 101920 83940
rect 98890 82940 101920 82963
rect 102080 82963 102103 83940
rect 105087 84940 105110 85947
rect 105270 85947 108300 85970
rect 105270 84940 105293 85947
rect 105087 83940 105293 84940
rect 105087 82963 105110 83940
rect 102080 82940 105110 82963
rect 105270 82963 105293 83940
rect 108277 84940 108300 85947
rect 108460 85947 111490 85970
rect 108460 84940 108483 85947
rect 108277 83940 108483 84940
rect 108277 82963 108300 83940
rect 105270 82940 108300 82963
rect 108460 82963 108483 83940
rect 111467 84940 111490 85947
rect 111650 85947 114680 85970
rect 111650 84940 111673 85947
rect 111467 83940 111673 84940
rect 111467 82963 111490 83940
rect 108460 82940 111490 82963
rect 111650 82963 111673 83940
rect 114657 84940 114680 85947
rect 114840 85947 117870 85970
rect 114840 84940 114863 85947
rect 114657 83940 114863 84940
rect 114657 82963 114680 83940
rect 111650 82940 114680 82963
rect 114840 82963 114863 83940
rect 117847 84940 117870 85947
rect 118030 85947 121060 85970
rect 118030 84940 118053 85947
rect 117847 83940 118053 84940
rect 117847 82963 117870 83940
rect 114840 82940 117870 82963
rect 118030 82963 118053 83940
rect 121037 84940 121060 85947
rect 121220 85947 124250 85970
rect 121220 84940 121243 85947
rect 121037 83940 121243 84940
rect 121037 82963 121060 83940
rect 118030 82940 121060 82963
rect 121220 82963 121243 83940
rect 124227 84940 124250 85947
rect 124410 85947 127440 85970
rect 124410 84940 124433 85947
rect 124227 83940 124433 84940
rect 124227 82963 124250 83940
rect 121220 82940 124250 82963
rect 124410 82963 124433 83940
rect 127417 84940 127440 85947
rect 127600 85947 130630 85970
rect 127600 84940 127623 85947
rect 127417 83940 127623 84940
rect 127417 82963 127440 83940
rect 124410 82940 127440 82963
rect 127600 82963 127623 83940
rect 130607 84940 130630 85947
rect 130790 85947 133820 85970
rect 130790 84940 130813 85947
rect 130607 83940 130813 84940
rect 130607 82963 130630 83940
rect 127600 82940 130630 82963
rect 130790 82963 130813 83940
rect 133797 84940 133820 85947
rect 133980 85947 137010 85970
rect 133980 84940 134003 85947
rect 133797 83940 134003 84940
rect 133797 82963 133820 83940
rect 130790 82940 133820 82963
rect 133980 82963 134003 83940
rect 136987 84940 137010 85947
rect 136987 83940 137170 84940
rect 136987 82963 137010 83940
rect 133980 82940 137010 82963
rect 9320 82780 9370 82940
rect 10570 82780 11570 82940
rect 13760 82780 14760 82940
rect 16950 82780 17950 82940
rect 20140 82780 21140 82940
rect 23330 82780 24330 82940
rect 26520 82780 27520 82940
rect 29710 82780 30710 82940
rect 32900 82780 33900 82940
rect 36090 82780 37090 82940
rect 39280 82780 40280 82940
rect 42470 82780 43470 82940
rect 45660 82780 46660 82940
rect 48850 82780 49850 82940
rect 52040 82780 53040 82940
rect 55230 82780 56230 82940
rect 58420 82780 59420 82940
rect 61610 82780 62610 82940
rect 64800 82780 65800 82940
rect 67990 82780 68990 82940
rect 71180 82780 72180 82940
rect 74370 82780 75370 82940
rect 77560 82780 78560 82940
rect 80750 82780 81750 82940
rect 83940 82780 84940 82940
rect 87130 82780 88130 82940
rect 90320 82780 91320 82940
rect 93510 82780 94510 82940
rect 96700 82780 97700 82940
rect 99890 82780 100890 82940
rect 103080 82780 104080 82940
rect 106270 82780 107270 82940
rect 109460 82780 110460 82940
rect 112650 82780 113650 82940
rect 115840 82780 116840 82940
rect 119030 82780 120030 82940
rect 122220 82780 123220 82940
rect 125410 82780 126410 82940
rect 128600 82780 129600 82940
rect 131790 82780 132790 82940
rect 134980 82780 135980 82940
rect 9320 81750 9410 82780
rect 9570 82757 12600 82780
rect 9570 81750 9593 82757
rect 9320 80750 9593 81750
rect 9320 79839 9410 80750
rect 0 79789 9410 79839
rect 0 79750 3030 79789
rect 3190 79750 6220 79789
rect 6380 79750 9410 79789
rect 9570 79773 9593 80750
rect 12577 81750 12600 82757
rect 12760 82757 15790 82780
rect 12760 81750 12783 82757
rect 12577 80750 12783 81750
rect 12577 79773 12600 80750
rect 9570 79750 12600 79773
rect 12760 79773 12783 80750
rect 15767 81750 15790 82757
rect 15950 82757 18980 82780
rect 15950 81750 15973 82757
rect 15767 80750 15973 81750
rect 15767 79773 15790 80750
rect 12760 79750 15790 79773
rect 15950 79773 15973 80750
rect 18957 81750 18980 82757
rect 19140 82757 22170 82780
rect 19140 81750 19163 82757
rect 18957 80750 19163 81750
rect 18957 79773 18980 80750
rect 15950 79750 18980 79773
rect 19140 79773 19163 80750
rect 22147 81750 22170 82757
rect 22330 82757 25360 82780
rect 22330 81750 22353 82757
rect 22147 80750 22353 81750
rect 22147 79773 22170 80750
rect 19140 79750 22170 79773
rect 22330 79773 22353 80750
rect 25337 81750 25360 82757
rect 25520 82757 28550 82780
rect 25520 81750 25543 82757
rect 25337 80750 25543 81750
rect 25337 79773 25360 80750
rect 22330 79750 25360 79773
rect 25520 79773 25543 80750
rect 28527 81750 28550 82757
rect 28710 82757 31740 82780
rect 28710 81750 28733 82757
rect 28527 80750 28733 81750
rect 28527 79773 28550 80750
rect 25520 79750 28550 79773
rect 28710 79773 28733 80750
rect 31717 81750 31740 82757
rect 31900 82757 34930 82780
rect 31900 81750 31923 82757
rect 31717 80750 31923 81750
rect 31717 79773 31740 80750
rect 28710 79750 31740 79773
rect 31900 79773 31923 80750
rect 34907 81750 34930 82757
rect 35090 82757 38120 82780
rect 35090 81750 35113 82757
rect 34907 80750 35113 81750
rect 34907 79773 34930 80750
rect 31900 79750 34930 79773
rect 35090 79773 35113 80750
rect 38097 81750 38120 82757
rect 38280 82757 41310 82780
rect 38280 81750 38303 82757
rect 38097 80750 38303 81750
rect 38097 79773 38120 80750
rect 35090 79750 38120 79773
rect 38280 79773 38303 80750
rect 41287 81750 41310 82757
rect 41470 82757 44500 82780
rect 41470 81750 41493 82757
rect 41287 80750 41493 81750
rect 41287 79773 41310 80750
rect 38280 79750 41310 79773
rect 41470 79773 41493 80750
rect 44477 81750 44500 82757
rect 44660 82757 47690 82780
rect 44660 81750 44683 82757
rect 44477 80750 44683 81750
rect 44477 79773 44500 80750
rect 41470 79750 44500 79773
rect 44660 79773 44683 80750
rect 47667 81750 47690 82757
rect 47850 82757 50880 82780
rect 47850 81750 47873 82757
rect 47667 80750 47873 81750
rect 47667 79773 47690 80750
rect 44660 79750 47690 79773
rect 47850 79773 47873 80750
rect 50857 81750 50880 82757
rect 51040 82757 54070 82780
rect 51040 81750 51063 82757
rect 50857 80750 51063 81750
rect 50857 79773 50880 80750
rect 47850 79750 50880 79773
rect 51040 79773 51063 80750
rect 54047 81750 54070 82757
rect 54230 82757 57260 82780
rect 54230 81750 54253 82757
rect 54047 80750 54253 81750
rect 54047 79773 54070 80750
rect 51040 79750 54070 79773
rect 54230 79773 54253 80750
rect 57237 81750 57260 82757
rect 57420 82757 60450 82780
rect 57420 81750 57443 82757
rect 57237 80750 57443 81750
rect 57237 79773 57260 80750
rect 54230 79750 57260 79773
rect 57420 79773 57443 80750
rect 60427 81750 60450 82757
rect 60610 82757 63640 82780
rect 60610 81750 60633 82757
rect 60427 80750 60633 81750
rect 60427 79773 60450 80750
rect 57420 79750 60450 79773
rect 60610 79773 60633 80750
rect 63617 81750 63640 82757
rect 63800 82757 66830 82780
rect 63800 81750 63823 82757
rect 63617 80750 63823 81750
rect 63617 79773 63640 80750
rect 60610 79750 63640 79773
rect 63800 79773 63823 80750
rect 66807 81750 66830 82757
rect 66990 82757 70020 82780
rect 66990 81750 67013 82757
rect 66807 80750 67013 81750
rect 66807 79773 66830 80750
rect 63800 79750 66830 79773
rect 66990 79773 67013 80750
rect 69997 81750 70020 82757
rect 70180 82757 73210 82780
rect 70180 81750 70203 82757
rect 69997 80750 70203 81750
rect 69997 79773 70020 80750
rect 66990 79750 70020 79773
rect 70180 79773 70203 80750
rect 73187 81750 73210 82757
rect 73370 82757 76400 82780
rect 73370 81750 73393 82757
rect 73187 80750 73393 81750
rect 73187 79773 73210 80750
rect 70180 79750 73210 79773
rect 73370 79773 73393 80750
rect 76377 81750 76400 82757
rect 76560 82757 79590 82780
rect 76560 81750 76583 82757
rect 76377 80750 76583 81750
rect 76377 79773 76400 80750
rect 73370 79750 76400 79773
rect 76560 79773 76583 80750
rect 79567 81750 79590 82757
rect 79750 82757 82780 82780
rect 79750 81750 79773 82757
rect 79567 80750 79773 81750
rect 79567 79773 79590 80750
rect 76560 79750 79590 79773
rect 79750 79773 79773 80750
rect 82757 81750 82780 82757
rect 82940 82757 85970 82780
rect 82940 81750 82963 82757
rect 82757 80750 82963 81750
rect 82757 79773 82780 80750
rect 79750 79750 82780 79773
rect 82940 79773 82963 80750
rect 85947 81750 85970 82757
rect 86130 82757 89160 82780
rect 86130 81750 86153 82757
rect 85947 80750 86153 81750
rect 85947 79773 85970 80750
rect 82940 79750 85970 79773
rect 86130 79773 86153 80750
rect 89137 81750 89160 82757
rect 89320 82757 92350 82780
rect 89320 81750 89343 82757
rect 89137 80750 89343 81750
rect 89137 79773 89160 80750
rect 86130 79750 89160 79773
rect 89320 79773 89343 80750
rect 92327 81750 92350 82757
rect 92510 82757 95540 82780
rect 92510 81750 92533 82757
rect 92327 80750 92533 81750
rect 92327 79773 92350 80750
rect 89320 79750 92350 79773
rect 92510 79773 92533 80750
rect 95517 81750 95540 82757
rect 95700 82757 98730 82780
rect 95700 81750 95723 82757
rect 95517 80750 95723 81750
rect 95517 79773 95540 80750
rect 92510 79750 95540 79773
rect 95700 79773 95723 80750
rect 98707 81750 98730 82757
rect 98890 82757 101920 82780
rect 98890 81750 98913 82757
rect 98707 80750 98913 81750
rect 98707 79773 98730 80750
rect 95700 79750 98730 79773
rect 98890 79773 98913 80750
rect 101897 81750 101920 82757
rect 102080 82757 105110 82780
rect 102080 81750 102103 82757
rect 101897 80750 102103 81750
rect 101897 79773 101920 80750
rect 98890 79750 101920 79773
rect 102080 79773 102103 80750
rect 105087 81750 105110 82757
rect 105270 82757 108300 82780
rect 105270 81750 105293 82757
rect 105087 80750 105293 81750
rect 105087 79773 105110 80750
rect 102080 79750 105110 79773
rect 105270 79773 105293 80750
rect 108277 81750 108300 82757
rect 108460 82757 111490 82780
rect 108460 81750 108483 82757
rect 108277 80750 108483 81750
rect 108277 79773 108300 80750
rect 105270 79750 108300 79773
rect 108460 79773 108483 80750
rect 111467 81750 111490 82757
rect 111650 82757 114680 82780
rect 111650 81750 111673 82757
rect 111467 80750 111673 81750
rect 111467 79773 111490 80750
rect 108460 79750 111490 79773
rect 111650 79773 111673 80750
rect 114657 81750 114680 82757
rect 114840 82757 117870 82780
rect 114840 81750 114863 82757
rect 114657 80750 114863 81750
rect 114657 79773 114680 80750
rect 111650 79750 114680 79773
rect 114840 79773 114863 80750
rect 117847 81750 117870 82757
rect 118030 82757 121060 82780
rect 118030 81750 118053 82757
rect 117847 80750 118053 81750
rect 117847 79773 117870 80750
rect 114840 79750 117870 79773
rect 118030 79773 118053 80750
rect 121037 81750 121060 82757
rect 121220 82757 124250 82780
rect 121220 81750 121243 82757
rect 121037 80750 121243 81750
rect 121037 79773 121060 80750
rect 118030 79750 121060 79773
rect 121220 79773 121243 80750
rect 124227 81750 124250 82757
rect 124410 82757 127440 82780
rect 124410 81750 124433 82757
rect 124227 80750 124433 81750
rect 124227 79773 124250 80750
rect 121220 79750 124250 79773
rect 124410 79773 124433 80750
rect 127417 81750 127440 82757
rect 127600 82757 130630 82780
rect 127600 81750 127623 82757
rect 127417 80750 127623 81750
rect 127417 79773 127440 80750
rect 124410 79750 127440 79773
rect 127600 79773 127623 80750
rect 130607 81750 130630 82757
rect 130790 82757 133820 82780
rect 130790 81750 130813 82757
rect 130607 80750 130813 81750
rect 130607 79773 130630 80750
rect 127600 79750 130630 79773
rect 130790 79773 130813 80750
rect 133797 81750 133820 82757
rect 133980 82757 137010 82780
rect 133980 81750 134003 82757
rect 133797 80750 134003 81750
rect 133797 79773 133820 80750
rect 130790 79750 133820 79773
rect 133980 79773 134003 80750
rect 136987 81750 137010 82757
rect 136987 80750 137170 81750
rect 136987 79773 137010 80750
rect 133980 79750 137010 79773
rect 1000 79590 2000 79750
rect 4190 79590 5190 79750
rect 7380 79590 8380 79750
rect 10570 79590 11570 79750
rect 13760 79590 14760 79750
rect 16950 79590 17950 79750
rect 20140 79590 21140 79750
rect 23330 79590 24330 79750
rect 26520 79590 27520 79750
rect 29710 79590 30710 79750
rect 32900 79590 33900 79750
rect 36090 79590 37090 79750
rect 39280 79590 40280 79750
rect 42470 79590 43470 79750
rect 45660 79590 46660 79750
rect 48850 79590 49850 79750
rect 52040 79590 53040 79750
rect 55230 79590 56230 79750
rect 58420 79590 59420 79750
rect 61610 79590 62610 79750
rect 64800 79590 65800 79750
rect 67990 79590 68990 79750
rect 71180 79590 72180 79750
rect 74370 79590 75370 79750
rect 77560 79590 78560 79750
rect 80750 79590 81750 79750
rect 83940 79590 84940 79750
rect 87130 79590 88130 79750
rect 90320 79590 91320 79750
rect 93510 79590 94510 79750
rect 96700 79590 97700 79750
rect 99890 79590 100890 79750
rect 103080 79590 104080 79750
rect 106270 79590 107270 79750
rect 109460 79590 110460 79750
rect 112650 79590 113650 79750
rect 115840 79590 116840 79750
rect 119030 79590 120030 79750
rect 122220 79590 123220 79750
rect 125410 79590 126410 79750
rect 128600 79590 129600 79750
rect 131790 79590 132790 79750
rect 134980 79590 135980 79750
rect 0 79567 3030 79590
rect 0 76583 23 79567
rect 3007 78560 3030 79567
rect 3190 79567 6220 79590
rect 3190 78560 3213 79567
rect 3007 77560 3213 78560
rect 3007 76583 3030 77560
rect 0 76560 3030 76583
rect 3190 76583 3213 77560
rect 6197 78560 6220 79567
rect 6380 79567 9410 79590
rect 6380 78560 6403 79567
rect 6197 77560 6403 78560
rect 6197 76583 6220 77560
rect 3190 76560 6220 76583
rect 6380 76583 6403 77560
rect 9387 78560 9410 79567
rect 9570 79567 12600 79590
rect 9570 78560 9593 79567
rect 9387 77560 9593 78560
rect 9387 76583 9410 77560
rect 6380 76560 9410 76583
rect 9570 76583 9593 77560
rect 12577 78560 12600 79567
rect 12760 79567 15790 79590
rect 12760 78560 12783 79567
rect 12577 77560 12783 78560
rect 12577 76583 12600 77560
rect 9570 76560 12600 76583
rect 12760 76583 12783 77560
rect 15767 78560 15790 79567
rect 15950 79567 18980 79590
rect 15950 78560 15973 79567
rect 15767 77560 15973 78560
rect 15767 76583 15790 77560
rect 12760 76560 15790 76583
rect 15950 76583 15973 77560
rect 18957 78560 18980 79567
rect 19140 79567 22170 79590
rect 19140 78560 19163 79567
rect 18957 77560 19163 78560
rect 18957 76583 18980 77560
rect 15950 76560 18980 76583
rect 19140 76583 19163 77560
rect 22147 78560 22170 79567
rect 22330 79567 25360 79590
rect 22330 78560 22353 79567
rect 22147 77560 22353 78560
rect 22147 76583 22170 77560
rect 19140 76560 22170 76583
rect 22330 76583 22353 77560
rect 25337 78560 25360 79567
rect 25520 79567 28550 79590
rect 25520 78560 25543 79567
rect 25337 77560 25543 78560
rect 25337 76583 25360 77560
rect 22330 76560 25360 76583
rect 25520 76583 25543 77560
rect 28527 78560 28550 79567
rect 28710 79567 31740 79590
rect 28710 78560 28733 79567
rect 28527 77560 28733 78560
rect 28527 76583 28550 77560
rect 25520 76560 28550 76583
rect 28710 76583 28733 77560
rect 31717 78560 31740 79567
rect 31900 79567 34930 79590
rect 31900 78560 31923 79567
rect 31717 77560 31923 78560
rect 31717 76583 31740 77560
rect 28710 76560 31740 76583
rect 31900 76583 31923 77560
rect 34907 78560 34930 79567
rect 35090 79567 38120 79590
rect 35090 78560 35113 79567
rect 34907 77560 35113 78560
rect 34907 76583 34930 77560
rect 31900 76560 34930 76583
rect 35090 76583 35113 77560
rect 38097 78560 38120 79567
rect 38280 79567 41310 79590
rect 38280 78560 38303 79567
rect 38097 77560 38303 78560
rect 38097 76583 38120 77560
rect 35090 76560 38120 76583
rect 38280 76583 38303 77560
rect 41287 78560 41310 79567
rect 41470 79567 44500 79590
rect 41470 78560 41493 79567
rect 41287 77560 41493 78560
rect 41287 76583 41310 77560
rect 38280 76560 41310 76583
rect 41470 76583 41493 77560
rect 44477 78560 44500 79567
rect 44660 79567 47690 79590
rect 44660 78560 44683 79567
rect 44477 77560 44683 78560
rect 44477 76583 44500 77560
rect 41470 76560 44500 76583
rect 44660 76583 44683 77560
rect 47667 78560 47690 79567
rect 47850 79567 50880 79590
rect 47850 78560 47873 79567
rect 47667 77560 47873 78560
rect 47667 76583 47690 77560
rect 44660 76560 47690 76583
rect 47850 76583 47873 77560
rect 50857 78560 50880 79567
rect 51040 79567 54070 79590
rect 51040 78560 51063 79567
rect 50857 77560 51063 78560
rect 50857 76583 50880 77560
rect 47850 76560 50880 76583
rect 51040 76583 51063 77560
rect 54047 78560 54070 79567
rect 54230 79567 57260 79590
rect 54230 78560 54253 79567
rect 54047 77560 54253 78560
rect 54047 76583 54070 77560
rect 51040 76560 54070 76583
rect 54230 76583 54253 77560
rect 57237 78560 57260 79567
rect 57420 79567 60450 79590
rect 57420 78560 57443 79567
rect 57237 77560 57443 78560
rect 57237 76583 57260 77560
rect 54230 76560 57260 76583
rect 57420 76583 57443 77560
rect 60427 78560 60450 79567
rect 60610 79567 63640 79590
rect 60610 78560 60633 79567
rect 60427 77560 60633 78560
rect 60427 76583 60450 77560
rect 57420 76560 60450 76583
rect 60610 76583 60633 77560
rect 63617 78560 63640 79567
rect 63800 79567 66830 79590
rect 63800 78560 63823 79567
rect 63617 77560 63823 78560
rect 63617 76583 63640 77560
rect 60610 76560 63640 76583
rect 63800 76583 63823 77560
rect 66807 78560 66830 79567
rect 66990 79567 70020 79590
rect 66990 78560 67013 79567
rect 66807 77560 67013 78560
rect 66807 76583 66830 77560
rect 63800 76560 66830 76583
rect 66990 76583 67013 77560
rect 69997 78560 70020 79567
rect 70180 79567 73210 79590
rect 70180 78560 70203 79567
rect 69997 77560 70203 78560
rect 69997 76583 70020 77560
rect 66990 76560 70020 76583
rect 70180 76583 70203 77560
rect 73187 78560 73210 79567
rect 73370 79567 76400 79590
rect 73370 78560 73393 79567
rect 73187 77560 73393 78560
rect 73187 76583 73210 77560
rect 70180 76560 73210 76583
rect 73370 76583 73393 77560
rect 76377 78560 76400 79567
rect 76560 79567 79590 79590
rect 76560 78560 76583 79567
rect 76377 77560 76583 78560
rect 76377 76583 76400 77560
rect 73370 76560 76400 76583
rect 76560 76583 76583 77560
rect 79567 78560 79590 79567
rect 79750 79567 82780 79590
rect 79750 78560 79773 79567
rect 79567 77560 79773 78560
rect 79567 76583 79590 77560
rect 76560 76560 79590 76583
rect 79750 76583 79773 77560
rect 82757 78560 82780 79567
rect 82940 79567 85970 79590
rect 82940 78560 82963 79567
rect 82757 77560 82963 78560
rect 82757 76583 82780 77560
rect 79750 76560 82780 76583
rect 82940 76583 82963 77560
rect 85947 78560 85970 79567
rect 86130 79567 89160 79590
rect 86130 78560 86153 79567
rect 85947 77560 86153 78560
rect 85947 76583 85970 77560
rect 82940 76560 85970 76583
rect 86130 76583 86153 77560
rect 89137 78560 89160 79567
rect 89320 79567 92350 79590
rect 89320 78560 89343 79567
rect 89137 77560 89343 78560
rect 89137 76583 89160 77560
rect 86130 76560 89160 76583
rect 89320 76583 89343 77560
rect 92327 78560 92350 79567
rect 92510 79567 95540 79590
rect 92510 78560 92533 79567
rect 92327 77560 92533 78560
rect 92327 76583 92350 77560
rect 89320 76560 92350 76583
rect 92510 76583 92533 77560
rect 95517 78560 95540 79567
rect 95700 79567 98730 79590
rect 95700 78560 95723 79567
rect 95517 77560 95723 78560
rect 95517 76583 95540 77560
rect 92510 76560 95540 76583
rect 95700 76583 95723 77560
rect 98707 78560 98730 79567
rect 98890 79567 101920 79590
rect 98890 78560 98913 79567
rect 98707 77560 98913 78560
rect 98707 76583 98730 77560
rect 95700 76560 98730 76583
rect 98890 76583 98913 77560
rect 101897 78560 101920 79567
rect 102080 79567 105110 79590
rect 102080 78560 102103 79567
rect 101897 77560 102103 78560
rect 101897 76583 101920 77560
rect 98890 76560 101920 76583
rect 102080 76583 102103 77560
rect 105087 78560 105110 79567
rect 105270 79567 108300 79590
rect 105270 78560 105293 79567
rect 105087 77560 105293 78560
rect 105087 76583 105110 77560
rect 102080 76560 105110 76583
rect 105270 76583 105293 77560
rect 108277 78560 108300 79567
rect 108460 79567 111490 79590
rect 108460 78560 108483 79567
rect 108277 77560 108483 78560
rect 108277 76583 108300 77560
rect 105270 76560 108300 76583
rect 108460 76583 108483 77560
rect 111467 78560 111490 79567
rect 111650 79567 114680 79590
rect 111650 78560 111673 79567
rect 111467 77560 111673 78560
rect 111467 76583 111490 77560
rect 108460 76560 111490 76583
rect 111650 76583 111673 77560
rect 114657 78560 114680 79567
rect 114840 79567 117870 79590
rect 114840 78560 114863 79567
rect 114657 77560 114863 78560
rect 114657 76583 114680 77560
rect 111650 76560 114680 76583
rect 114840 76583 114863 77560
rect 117847 78560 117870 79567
rect 118030 79567 121060 79590
rect 118030 78560 118053 79567
rect 117847 77560 118053 78560
rect 117847 76583 117870 77560
rect 114840 76560 117870 76583
rect 118030 76583 118053 77560
rect 121037 78560 121060 79567
rect 121220 79567 124250 79590
rect 121220 78560 121243 79567
rect 121037 77560 121243 78560
rect 121037 76583 121060 77560
rect 118030 76560 121060 76583
rect 121220 76583 121243 77560
rect 124227 78560 124250 79567
rect 124410 79567 127440 79590
rect 124410 78560 124433 79567
rect 124227 77560 124433 78560
rect 124227 76583 124250 77560
rect 121220 76560 124250 76583
rect 124410 76583 124433 77560
rect 127417 78560 127440 79567
rect 127600 79567 130630 79590
rect 127600 78560 127623 79567
rect 127417 77560 127623 78560
rect 127417 76583 127440 77560
rect 124410 76560 127440 76583
rect 127600 76583 127623 77560
rect 130607 78560 130630 79567
rect 130790 79567 133820 79590
rect 130790 78560 130813 79567
rect 130607 77560 130813 78560
rect 130607 76583 130630 77560
rect 127600 76560 130630 76583
rect 130790 76583 130813 77560
rect 133797 78560 133820 79567
rect 133980 79567 137010 79590
rect 133980 78560 134003 79567
rect 133797 77560 134003 78560
rect 133797 76583 133820 77560
rect 130790 76560 133820 76583
rect 133980 76583 134003 77560
rect 136987 78560 137010 79567
rect 136987 77560 137170 78560
rect 136987 76583 137010 77560
rect 133980 76560 137010 76583
rect 1000 76400 2000 76560
rect 4190 76400 5190 76560
rect 7380 76400 8380 76560
rect 10570 76400 11570 76560
rect 13760 76400 14760 76560
rect 16950 76400 17950 76560
rect 20140 76400 21140 76560
rect 23330 76400 24330 76560
rect 26520 76400 27520 76560
rect 29710 76400 30710 76560
rect 32900 76400 33900 76560
rect 36090 76400 37090 76560
rect 39280 76400 40280 76560
rect 42470 76400 43470 76560
rect 45660 76400 46660 76560
rect 48850 76400 49850 76560
rect 52040 76400 53040 76560
rect 55230 76400 56230 76560
rect 58420 76400 59420 76560
rect 61610 76400 62610 76560
rect 64800 76400 65800 76560
rect 67990 76400 68990 76560
rect 71180 76400 72180 76560
rect 74370 76400 75370 76560
rect 77560 76400 78560 76560
rect 80750 76400 81750 76560
rect 83940 76400 84940 76560
rect 87130 76400 88130 76560
rect 90320 76400 91320 76560
rect 93510 76400 94510 76560
rect 96700 76400 97700 76560
rect 99890 76400 100890 76560
rect 103080 76400 104080 76560
rect 106270 76400 107270 76560
rect 109460 76400 110460 76560
rect 112650 76400 113650 76560
rect 115840 76400 116840 76560
rect 119030 76400 120030 76560
rect 122220 76400 123220 76560
rect 125410 76400 126410 76560
rect 128600 76400 129600 76560
rect 131790 76400 132790 76560
rect 134980 76400 135980 76560
rect 0 76377 3030 76400
rect 0 73393 23 76377
rect 3007 75370 3030 76377
rect 3190 76377 6220 76400
rect 3190 75370 3213 76377
rect 3007 74370 3213 75370
rect 3007 73393 3030 74370
rect 0 73370 3030 73393
rect 3190 73393 3213 74370
rect 6197 75370 6220 76377
rect 6380 76377 9410 76400
rect 6380 75370 6403 76377
rect 6197 74370 6403 75370
rect 6197 73393 6220 74370
rect 3190 73370 6220 73393
rect 6380 73393 6403 74370
rect 9387 75370 9410 76377
rect 9570 76377 12600 76400
rect 9570 75370 9593 76377
rect 9387 74370 9593 75370
rect 9387 73393 9410 74370
rect 6380 73370 9410 73393
rect 9570 73393 9593 74370
rect 12577 75370 12600 76377
rect 12760 76377 15790 76400
rect 12760 75370 12783 76377
rect 12577 74370 12783 75370
rect 12577 73393 12600 74370
rect 9570 73370 12600 73393
rect 12760 73393 12783 74370
rect 15767 75370 15790 76377
rect 15950 76377 18980 76400
rect 15950 75370 15973 76377
rect 15767 74370 15973 75370
rect 15767 73393 15790 74370
rect 12760 73370 15790 73393
rect 15950 73393 15973 74370
rect 18957 75370 18980 76377
rect 19140 76377 22170 76400
rect 19140 75370 19163 76377
rect 18957 74370 19163 75370
rect 18957 73393 18980 74370
rect 15950 73370 18980 73393
rect 19140 73393 19163 74370
rect 22147 75370 22170 76377
rect 22330 76377 25360 76400
rect 22330 75370 22353 76377
rect 22147 74370 22353 75370
rect 22147 73393 22170 74370
rect 19140 73370 22170 73393
rect 22330 73393 22353 74370
rect 25337 75370 25360 76377
rect 25520 76377 28550 76400
rect 25520 75370 25543 76377
rect 25337 74370 25543 75370
rect 25337 73393 25360 74370
rect 22330 73370 25360 73393
rect 25520 73393 25543 74370
rect 28527 75370 28550 76377
rect 28710 76377 31740 76400
rect 28710 75370 28733 76377
rect 28527 74370 28733 75370
rect 28527 73393 28550 74370
rect 25520 73370 28550 73393
rect 28710 73393 28733 74370
rect 31717 75370 31740 76377
rect 31900 76377 34930 76400
rect 31900 75370 31923 76377
rect 31717 74370 31923 75370
rect 31717 73393 31740 74370
rect 28710 73370 31740 73393
rect 31900 73393 31923 74370
rect 34907 75370 34930 76377
rect 35090 76377 38120 76400
rect 35090 75370 35113 76377
rect 34907 74370 35113 75370
rect 34907 73393 34930 74370
rect 31900 73370 34930 73393
rect 35090 73393 35113 74370
rect 38097 75370 38120 76377
rect 38280 76377 41310 76400
rect 38280 75370 38303 76377
rect 38097 74370 38303 75370
rect 38097 73393 38120 74370
rect 35090 73370 38120 73393
rect 38280 73393 38303 74370
rect 41287 75370 41310 76377
rect 41470 76377 44500 76400
rect 41470 75370 41493 76377
rect 41287 74370 41493 75370
rect 41287 73393 41310 74370
rect 38280 73370 41310 73393
rect 41470 73393 41493 74370
rect 44477 75370 44500 76377
rect 44660 76377 47690 76400
rect 44660 75370 44683 76377
rect 44477 74370 44683 75370
rect 44477 73393 44500 74370
rect 41470 73370 44500 73393
rect 44660 73393 44683 74370
rect 47667 75370 47690 76377
rect 47850 76377 50880 76400
rect 47850 75370 47873 76377
rect 47667 74370 47873 75370
rect 47667 73393 47690 74370
rect 44660 73370 47690 73393
rect 47850 73393 47873 74370
rect 50857 75370 50880 76377
rect 51040 76377 54070 76400
rect 51040 75370 51063 76377
rect 50857 74370 51063 75370
rect 50857 73393 50880 74370
rect 47850 73370 50880 73393
rect 51040 73393 51063 74370
rect 54047 75370 54070 76377
rect 54230 76377 57260 76400
rect 54230 75370 54253 76377
rect 54047 74370 54253 75370
rect 54047 73393 54070 74370
rect 51040 73370 54070 73393
rect 54230 73393 54253 74370
rect 57237 75370 57260 76377
rect 57420 76377 60450 76400
rect 57420 75370 57443 76377
rect 57237 74370 57443 75370
rect 57237 73393 57260 74370
rect 54230 73370 57260 73393
rect 57420 73393 57443 74370
rect 60427 75370 60450 76377
rect 60610 76377 63640 76400
rect 60610 75370 60633 76377
rect 60427 74370 60633 75370
rect 60427 73393 60450 74370
rect 57420 73370 60450 73393
rect 60610 73393 60633 74370
rect 63617 75370 63640 76377
rect 63800 76377 66830 76400
rect 63800 75370 63823 76377
rect 63617 74370 63823 75370
rect 63617 73393 63640 74370
rect 60610 73370 63640 73393
rect 63800 73393 63823 74370
rect 66807 75370 66830 76377
rect 66990 76377 70020 76400
rect 66990 75370 67013 76377
rect 66807 74370 67013 75370
rect 66807 73393 66830 74370
rect 63800 73370 66830 73393
rect 66990 73393 67013 74370
rect 69997 75370 70020 76377
rect 70180 76377 73210 76400
rect 70180 75370 70203 76377
rect 69997 74370 70203 75370
rect 69997 73393 70020 74370
rect 66990 73370 70020 73393
rect 70180 73393 70203 74370
rect 73187 75370 73210 76377
rect 73370 76377 76400 76400
rect 73370 75370 73393 76377
rect 73187 74370 73393 75370
rect 73187 73393 73210 74370
rect 70180 73370 73210 73393
rect 73370 73393 73393 74370
rect 76377 75370 76400 76377
rect 76560 76377 79590 76400
rect 76560 75370 76583 76377
rect 76377 74370 76583 75370
rect 76377 73393 76400 74370
rect 73370 73370 76400 73393
rect 76560 73393 76583 74370
rect 79567 75370 79590 76377
rect 79750 76377 82780 76400
rect 79750 75370 79773 76377
rect 79567 74370 79773 75370
rect 79567 73393 79590 74370
rect 76560 73370 79590 73393
rect 79750 73393 79773 74370
rect 82757 75370 82780 76377
rect 82940 76377 85970 76400
rect 82940 75370 82963 76377
rect 82757 74370 82963 75370
rect 82757 73393 82780 74370
rect 79750 73370 82780 73393
rect 82940 73393 82963 74370
rect 85947 75370 85970 76377
rect 86130 76377 89160 76400
rect 86130 75370 86153 76377
rect 85947 74370 86153 75370
rect 85947 73393 85970 74370
rect 82940 73370 85970 73393
rect 86130 73393 86153 74370
rect 89137 75370 89160 76377
rect 89320 76377 92350 76400
rect 89320 75370 89343 76377
rect 89137 74370 89343 75370
rect 89137 73393 89160 74370
rect 86130 73370 89160 73393
rect 89320 73393 89343 74370
rect 92327 75370 92350 76377
rect 92510 76377 95540 76400
rect 92510 75370 92533 76377
rect 92327 74370 92533 75370
rect 92327 73393 92350 74370
rect 89320 73370 92350 73393
rect 92510 73393 92533 74370
rect 95517 75370 95540 76377
rect 95700 76377 98730 76400
rect 95700 75370 95723 76377
rect 95517 74370 95723 75370
rect 95517 73393 95540 74370
rect 92510 73370 95540 73393
rect 95700 73393 95723 74370
rect 98707 75370 98730 76377
rect 98890 76377 101920 76400
rect 98890 75370 98913 76377
rect 98707 74370 98913 75370
rect 98707 73393 98730 74370
rect 95700 73370 98730 73393
rect 98890 73393 98913 74370
rect 101897 75370 101920 76377
rect 102080 76377 105110 76400
rect 102080 75370 102103 76377
rect 101897 74370 102103 75370
rect 101897 73393 101920 74370
rect 98890 73370 101920 73393
rect 102080 73393 102103 74370
rect 105087 75370 105110 76377
rect 105270 76377 108300 76400
rect 105270 75370 105293 76377
rect 105087 74370 105293 75370
rect 105087 73393 105110 74370
rect 102080 73370 105110 73393
rect 105270 73393 105293 74370
rect 108277 75370 108300 76377
rect 108460 76377 111490 76400
rect 108460 75370 108483 76377
rect 108277 74370 108483 75370
rect 108277 73393 108300 74370
rect 105270 73370 108300 73393
rect 108460 73393 108483 74370
rect 111467 75370 111490 76377
rect 111650 76377 114680 76400
rect 111650 75370 111673 76377
rect 111467 74370 111673 75370
rect 111467 73393 111490 74370
rect 108460 73370 111490 73393
rect 111650 73393 111673 74370
rect 114657 75370 114680 76377
rect 114840 76377 117870 76400
rect 114840 75370 114863 76377
rect 114657 74370 114863 75370
rect 114657 73393 114680 74370
rect 111650 73370 114680 73393
rect 114840 73393 114863 74370
rect 117847 75370 117870 76377
rect 118030 76377 121060 76400
rect 118030 75370 118053 76377
rect 117847 74370 118053 75370
rect 117847 73393 117870 74370
rect 114840 73370 117870 73393
rect 118030 73393 118053 74370
rect 121037 75370 121060 76377
rect 121220 76377 124250 76400
rect 121220 75370 121243 76377
rect 121037 74370 121243 75370
rect 121037 73393 121060 74370
rect 118030 73370 121060 73393
rect 121220 73393 121243 74370
rect 124227 75370 124250 76377
rect 124410 76377 127440 76400
rect 124410 75370 124433 76377
rect 124227 74370 124433 75370
rect 124227 73393 124250 74370
rect 121220 73370 124250 73393
rect 124410 73393 124433 74370
rect 127417 75370 127440 76377
rect 127600 76377 130630 76400
rect 127600 75370 127623 76377
rect 127417 74370 127623 75370
rect 127417 73393 127440 74370
rect 124410 73370 127440 73393
rect 127600 73393 127623 74370
rect 130607 75370 130630 76377
rect 130790 76377 133820 76400
rect 130790 75370 130813 76377
rect 130607 74370 130813 75370
rect 130607 73393 130630 74370
rect 127600 73370 130630 73393
rect 130790 73393 130813 74370
rect 133797 75370 133820 76377
rect 133980 76377 137010 76400
rect 133980 75370 134003 76377
rect 133797 74370 134003 75370
rect 133797 73393 133820 74370
rect 130790 73370 133820 73393
rect 133980 73393 134003 74370
rect 136987 75370 137010 76377
rect 136987 74370 137170 75370
rect 136987 73393 137010 74370
rect 133980 73370 137010 73393
rect 1000 73210 2000 73370
rect 4190 73210 5190 73370
rect 7380 73210 8380 73370
rect 10570 73210 11570 73370
rect 13760 73210 14760 73370
rect 16950 73210 17950 73370
rect 20140 73210 21140 73370
rect 23330 73210 24330 73370
rect 26520 73210 27520 73370
rect 29710 73210 30710 73370
rect 32900 73210 33900 73370
rect 36090 73210 37090 73370
rect 39280 73210 40280 73370
rect 42470 73210 43470 73370
rect 45660 73210 46660 73370
rect 48850 73210 49850 73370
rect 52040 73210 53040 73370
rect 55230 73210 56230 73370
rect 58420 73210 59420 73370
rect 61610 73210 62610 73370
rect 64800 73210 65800 73370
rect 67990 73210 68990 73370
rect 71180 73210 72180 73370
rect 74370 73210 75370 73370
rect 77560 73210 78560 73370
rect 80750 73210 81750 73370
rect 83940 73210 84940 73370
rect 87130 73210 88130 73370
rect 90320 73210 91320 73370
rect 93510 73210 94510 73370
rect 96700 73210 97700 73370
rect 99890 73210 100890 73370
rect 103080 73210 104080 73370
rect 106270 73210 107270 73370
rect 109460 73210 110460 73370
rect 112650 73210 113650 73370
rect 115840 73210 116840 73370
rect 119030 73210 120030 73370
rect 122220 73210 123220 73370
rect 125410 73210 126410 73370
rect 128600 73210 129600 73370
rect 131790 73210 132790 73370
rect 134980 73210 135980 73370
rect 0 73187 3030 73210
rect 0 70203 23 73187
rect 3007 72180 3030 73187
rect 3190 73187 6220 73210
rect 3190 72180 3213 73187
rect 3007 71180 3213 72180
rect 3007 70203 3030 71180
rect 0 70180 3030 70203
rect 3190 70203 3213 71180
rect 6197 72180 6220 73187
rect 6380 73187 9410 73210
rect 6380 72180 6403 73187
rect 6197 71180 6403 72180
rect 6197 70203 6220 71180
rect 3190 70180 6220 70203
rect 6380 70203 6403 71180
rect 9387 72180 9410 73187
rect 9570 73187 12600 73210
rect 9570 72180 9593 73187
rect 9387 71180 9593 72180
rect 9387 70203 9410 71180
rect 6380 70180 9410 70203
rect 9570 70203 9593 71180
rect 12577 72180 12600 73187
rect 12760 73187 15790 73210
rect 12760 72180 12783 73187
rect 12577 71180 12783 72180
rect 12577 70203 12600 71180
rect 9570 70180 12600 70203
rect 12760 70203 12783 71180
rect 15767 72180 15790 73187
rect 15950 73187 18980 73210
rect 15950 72180 15973 73187
rect 15767 71180 15973 72180
rect 15767 70203 15790 71180
rect 12760 70180 15790 70203
rect 15950 70203 15973 71180
rect 18957 72180 18980 73187
rect 19140 73187 22170 73210
rect 19140 72180 19163 73187
rect 18957 71180 19163 72180
rect 18957 70203 18980 71180
rect 15950 70180 18980 70203
rect 19140 70203 19163 71180
rect 22147 72180 22170 73187
rect 22330 73187 25360 73210
rect 22330 72180 22353 73187
rect 22147 71180 22353 72180
rect 22147 70203 22170 71180
rect 19140 70180 22170 70203
rect 22330 70203 22353 71180
rect 25337 72180 25360 73187
rect 25520 73187 28550 73210
rect 25520 72180 25543 73187
rect 25337 71180 25543 72180
rect 25337 70203 25360 71180
rect 22330 70180 25360 70203
rect 25520 70203 25543 71180
rect 28527 72180 28550 73187
rect 28710 73187 31740 73210
rect 28710 72180 28733 73187
rect 28527 71180 28733 72180
rect 28527 70203 28550 71180
rect 25520 70180 28550 70203
rect 28710 70203 28733 71180
rect 31717 72180 31740 73187
rect 31900 73187 34930 73210
rect 31900 72180 31923 73187
rect 31717 71180 31923 72180
rect 31717 70203 31740 71180
rect 28710 70180 31740 70203
rect 31900 70203 31923 71180
rect 34907 72180 34930 73187
rect 35090 73187 38120 73210
rect 35090 72180 35113 73187
rect 34907 71180 35113 72180
rect 34907 70203 34930 71180
rect 31900 70180 34930 70203
rect 35090 70203 35113 71180
rect 38097 72180 38120 73187
rect 38280 73187 41310 73210
rect 38280 72180 38303 73187
rect 38097 71180 38303 72180
rect 38097 70203 38120 71180
rect 35090 70180 38120 70203
rect 38280 70203 38303 71180
rect 41287 72180 41310 73187
rect 41470 73187 44500 73210
rect 41470 72180 41493 73187
rect 41287 71180 41493 72180
rect 41287 70203 41310 71180
rect 38280 70180 41310 70203
rect 41470 70203 41493 71180
rect 44477 72180 44500 73187
rect 44660 73187 47690 73210
rect 44660 72180 44683 73187
rect 44477 71180 44683 72180
rect 44477 70203 44500 71180
rect 41470 70180 44500 70203
rect 44660 70203 44683 71180
rect 47667 72180 47690 73187
rect 47850 73187 50880 73210
rect 47850 72180 47873 73187
rect 47667 71180 47873 72180
rect 47667 70203 47690 71180
rect 44660 70180 47690 70203
rect 47850 70203 47873 71180
rect 50857 72180 50880 73187
rect 51040 73187 54070 73210
rect 51040 72180 51063 73187
rect 50857 71180 51063 72180
rect 50857 70203 50880 71180
rect 47850 70180 50880 70203
rect 51040 70203 51063 71180
rect 54047 72180 54070 73187
rect 54230 73187 57260 73210
rect 54230 72180 54253 73187
rect 54047 71180 54253 72180
rect 54047 70203 54070 71180
rect 51040 70180 54070 70203
rect 54230 70203 54253 71180
rect 57237 72180 57260 73187
rect 57420 73187 60450 73210
rect 57420 72180 57443 73187
rect 57237 71180 57443 72180
rect 57237 70203 57260 71180
rect 54230 70180 57260 70203
rect 57420 70203 57443 71180
rect 60427 72180 60450 73187
rect 60610 73187 63640 73210
rect 60610 72180 60633 73187
rect 60427 71180 60633 72180
rect 60427 70203 60450 71180
rect 57420 70180 60450 70203
rect 60610 70203 60633 71180
rect 63617 72180 63640 73187
rect 63800 73187 66830 73210
rect 63800 72180 63823 73187
rect 63617 71180 63823 72180
rect 63617 70203 63640 71180
rect 60610 70180 63640 70203
rect 63800 70203 63823 71180
rect 66807 72180 66830 73187
rect 66990 73187 70020 73210
rect 66990 72180 67013 73187
rect 66807 71180 67013 72180
rect 66807 70203 66830 71180
rect 63800 70180 66830 70203
rect 66990 70203 67013 71180
rect 69997 72180 70020 73187
rect 70180 73187 73210 73210
rect 70180 72180 70203 73187
rect 69997 71180 70203 72180
rect 69997 70203 70020 71180
rect 66990 70180 70020 70203
rect 70180 70203 70203 71180
rect 73187 72180 73210 73187
rect 73370 73187 76400 73210
rect 73370 72180 73393 73187
rect 73187 71180 73393 72180
rect 73187 70203 73210 71180
rect 70180 70180 73210 70203
rect 73370 70203 73393 71180
rect 76377 72180 76400 73187
rect 76560 73187 79590 73210
rect 76560 72180 76583 73187
rect 76377 71180 76583 72180
rect 76377 70203 76400 71180
rect 73370 70180 76400 70203
rect 76560 70203 76583 71180
rect 79567 72180 79590 73187
rect 79750 73187 82780 73210
rect 79750 72180 79773 73187
rect 79567 71180 79773 72180
rect 79567 70203 79590 71180
rect 76560 70180 79590 70203
rect 79750 70203 79773 71180
rect 82757 72180 82780 73187
rect 82940 73187 85970 73210
rect 82940 72180 82963 73187
rect 82757 71180 82963 72180
rect 82757 70203 82780 71180
rect 79750 70180 82780 70203
rect 82940 70203 82963 71180
rect 85947 72180 85970 73187
rect 86130 73187 89160 73210
rect 86130 72180 86153 73187
rect 85947 71180 86153 72180
rect 85947 70203 85970 71180
rect 82940 70180 85970 70203
rect 86130 70203 86153 71180
rect 89137 72180 89160 73187
rect 89320 73187 92350 73210
rect 89320 72180 89343 73187
rect 89137 71180 89343 72180
rect 89137 70203 89160 71180
rect 86130 70180 89160 70203
rect 89320 70203 89343 71180
rect 92327 72180 92350 73187
rect 92510 73187 95540 73210
rect 92510 72180 92533 73187
rect 92327 71180 92533 72180
rect 92327 70203 92350 71180
rect 89320 70180 92350 70203
rect 92510 70203 92533 71180
rect 95517 72180 95540 73187
rect 95700 73187 98730 73210
rect 95700 72180 95723 73187
rect 95517 71180 95723 72180
rect 95517 70203 95540 71180
rect 92510 70180 95540 70203
rect 95700 70203 95723 71180
rect 98707 72180 98730 73187
rect 98890 73187 101920 73210
rect 98890 72180 98913 73187
rect 98707 71180 98913 72180
rect 98707 70203 98730 71180
rect 95700 70180 98730 70203
rect 98890 70203 98913 71180
rect 101897 72180 101920 73187
rect 102080 73187 105110 73210
rect 102080 72180 102103 73187
rect 101897 71180 102103 72180
rect 101897 70203 101920 71180
rect 98890 70180 101920 70203
rect 102080 70203 102103 71180
rect 105087 72180 105110 73187
rect 105270 73187 108300 73210
rect 105270 72180 105293 73187
rect 105087 71180 105293 72180
rect 105087 70203 105110 71180
rect 102080 70180 105110 70203
rect 105270 70203 105293 71180
rect 108277 72180 108300 73187
rect 108460 73187 111490 73210
rect 108460 72180 108483 73187
rect 108277 71180 108483 72180
rect 108277 70203 108300 71180
rect 105270 70180 108300 70203
rect 108460 70203 108483 71180
rect 111467 72180 111490 73187
rect 111650 73187 114680 73210
rect 111650 72180 111673 73187
rect 111467 71180 111673 72180
rect 111467 70203 111490 71180
rect 108460 70180 111490 70203
rect 111650 70203 111673 71180
rect 114657 72180 114680 73187
rect 114840 73187 117870 73210
rect 114840 72180 114863 73187
rect 114657 71180 114863 72180
rect 114657 70203 114680 71180
rect 111650 70180 114680 70203
rect 114840 70203 114863 71180
rect 117847 72180 117870 73187
rect 118030 73187 121060 73210
rect 118030 72180 118053 73187
rect 117847 71180 118053 72180
rect 117847 70203 117870 71180
rect 114840 70180 117870 70203
rect 118030 70203 118053 71180
rect 121037 72180 121060 73187
rect 121220 73187 124250 73210
rect 121220 72180 121243 73187
rect 121037 71180 121243 72180
rect 121037 70203 121060 71180
rect 118030 70180 121060 70203
rect 121220 70203 121243 71180
rect 124227 72180 124250 73187
rect 124410 73187 127440 73210
rect 124410 72180 124433 73187
rect 124227 71180 124433 72180
rect 124227 70203 124250 71180
rect 121220 70180 124250 70203
rect 124410 70203 124433 71180
rect 127417 72180 127440 73187
rect 127600 73187 130630 73210
rect 127600 72180 127623 73187
rect 127417 71180 127623 72180
rect 127417 70203 127440 71180
rect 124410 70180 127440 70203
rect 127600 70203 127623 71180
rect 130607 72180 130630 73187
rect 130790 73187 133820 73210
rect 130790 72180 130813 73187
rect 130607 71180 130813 72180
rect 130607 70203 130630 71180
rect 127600 70180 130630 70203
rect 130790 70203 130813 71180
rect 133797 72180 133820 73187
rect 133980 73187 137010 73210
rect 133980 72180 134003 73187
rect 133797 71180 134003 72180
rect 133797 70203 133820 71180
rect 130790 70180 133820 70203
rect 133980 70203 134003 71180
rect 136987 72180 137010 73187
rect 136987 71180 137170 72180
rect 136987 70203 137010 71180
rect 133980 70180 137010 70203
rect 1000 70020 2000 70180
rect 4190 70020 5190 70180
rect 7380 70020 8380 70180
rect 10570 70020 11570 70180
rect 13760 70020 14760 70180
rect 16950 70020 17950 70180
rect 20140 70020 21140 70180
rect 23330 70020 24330 70180
rect 26520 70020 27520 70180
rect 29710 70020 30710 70180
rect 32900 70020 33900 70180
rect 36090 70020 37090 70180
rect 39280 70020 40280 70180
rect 42470 70020 43470 70180
rect 45660 70020 46660 70180
rect 48850 70020 49850 70180
rect 52040 70020 53040 70180
rect 55230 70020 56230 70180
rect 58420 70020 59420 70180
rect 61610 70020 62610 70180
rect 64800 70020 65800 70180
rect 67990 70020 68990 70180
rect 71180 70020 72180 70180
rect 74370 70020 75370 70180
rect 77560 70020 78560 70180
rect 80750 70020 81750 70180
rect 83940 70020 84940 70180
rect 87130 70020 88130 70180
rect 90320 70020 91320 70180
rect 93510 70020 94510 70180
rect 96700 70020 97700 70180
rect 99890 70020 100890 70180
rect 103080 70020 104080 70180
rect 106270 70020 107270 70180
rect 109460 70020 110460 70180
rect 112650 70020 113650 70180
rect 115840 70020 116840 70180
rect 119030 70020 120030 70180
rect 122220 70020 123220 70180
rect 125410 70020 126410 70180
rect 128600 70020 129600 70180
rect 131790 70020 132790 70180
rect 134980 70020 135980 70180
rect 0 69997 3030 70020
rect 0 67013 23 69997
rect 3007 68990 3030 69997
rect 3190 69997 6220 70020
rect 3190 68990 3213 69997
rect 3007 67990 3213 68990
rect 3007 67013 3030 67990
rect 0 66990 3030 67013
rect 3190 67013 3213 67990
rect 6197 68990 6220 69997
rect 6380 69997 9410 70020
rect 6380 68990 6403 69997
rect 6197 67990 6403 68990
rect 6197 67013 6220 67990
rect 3190 66990 6220 67013
rect 6380 67013 6403 67990
rect 9387 68990 9410 69997
rect 9570 69997 12600 70020
rect 9570 68990 9593 69997
rect 9387 67990 9593 68990
rect 9387 67013 9410 67990
rect 6380 66990 9410 67013
rect 9570 67013 9593 67990
rect 12577 68990 12600 69997
rect 12760 69997 15790 70020
rect 12760 68990 12783 69997
rect 12577 67990 12783 68990
rect 12577 67013 12600 67990
rect 9570 66990 12600 67013
rect 12760 67013 12783 67990
rect 15767 68990 15790 69997
rect 15950 69997 18980 70020
rect 15950 68990 15973 69997
rect 15767 67990 15973 68990
rect 15767 67013 15790 67990
rect 12760 66990 15790 67013
rect 15950 67013 15973 67990
rect 18957 68990 18980 69997
rect 19140 69997 22170 70020
rect 19140 68990 19163 69997
rect 18957 67990 19163 68990
rect 18957 67013 18980 67990
rect 15950 66990 18980 67013
rect 19140 67013 19163 67990
rect 22147 68990 22170 69997
rect 22330 69997 25360 70020
rect 22330 68990 22353 69997
rect 22147 67990 22353 68990
rect 22147 67013 22170 67990
rect 19140 66990 22170 67013
rect 22330 67013 22353 67990
rect 25337 68990 25360 69997
rect 25520 69997 28550 70020
rect 25520 68990 25543 69997
rect 25337 67990 25543 68990
rect 25337 67013 25360 67990
rect 22330 66990 25360 67013
rect 25520 67013 25543 67990
rect 28527 68990 28550 69997
rect 28710 69997 31740 70020
rect 28710 68990 28733 69997
rect 28527 67990 28733 68990
rect 28527 67013 28550 67990
rect 25520 66990 28550 67013
rect 28710 67013 28733 67990
rect 31717 68990 31740 69997
rect 31900 69997 34930 70020
rect 31900 68990 31923 69997
rect 31717 67990 31923 68990
rect 31717 67013 31740 67990
rect 28710 66990 31740 67013
rect 31900 67013 31923 67990
rect 34907 68990 34930 69997
rect 35090 69997 38120 70020
rect 35090 68990 35113 69997
rect 34907 67990 35113 68990
rect 34907 67013 34930 67990
rect 31900 66990 34930 67013
rect 35090 67013 35113 67990
rect 38097 68990 38120 69997
rect 38280 69997 41310 70020
rect 38280 68990 38303 69997
rect 38097 67990 38303 68990
rect 38097 67013 38120 67990
rect 35090 66990 38120 67013
rect 38280 67013 38303 67990
rect 41287 68990 41310 69997
rect 41470 69997 44500 70020
rect 41470 68990 41493 69997
rect 41287 67990 41493 68990
rect 41287 67013 41310 67990
rect 38280 66990 41310 67013
rect 41470 67013 41493 67990
rect 44477 68990 44500 69997
rect 44660 69997 47690 70020
rect 44660 68990 44683 69997
rect 44477 67990 44683 68990
rect 44477 67013 44500 67990
rect 41470 66990 44500 67013
rect 44660 67013 44683 67990
rect 47667 68990 47690 69997
rect 47850 69997 50880 70020
rect 47850 68990 47873 69997
rect 47667 67990 47873 68990
rect 47667 67013 47690 67990
rect 44660 66990 47690 67013
rect 47850 67013 47873 67990
rect 50857 68990 50880 69997
rect 51040 69997 54070 70020
rect 51040 68990 51063 69997
rect 50857 67990 51063 68990
rect 50857 67013 50880 67990
rect 47850 66990 50880 67013
rect 51040 67013 51063 67990
rect 54047 68990 54070 69997
rect 54230 69997 57260 70020
rect 54230 68990 54253 69997
rect 54047 67990 54253 68990
rect 54047 67013 54070 67990
rect 51040 66990 54070 67013
rect 54230 67013 54253 67990
rect 57237 68990 57260 69997
rect 57420 69997 60450 70020
rect 57420 68990 57443 69997
rect 57237 67990 57443 68990
rect 57237 67013 57260 67990
rect 54230 66990 57260 67013
rect 57420 67013 57443 67990
rect 60427 68990 60450 69997
rect 60610 69997 63640 70020
rect 60610 68990 60633 69997
rect 60427 67990 60633 68990
rect 60427 67013 60450 67990
rect 57420 66990 60450 67013
rect 60610 67013 60633 67990
rect 63617 68990 63640 69997
rect 63800 69997 66830 70020
rect 63800 68990 63823 69997
rect 63617 67990 63823 68990
rect 63617 67013 63640 67990
rect 60610 66990 63640 67013
rect 63800 67013 63823 67990
rect 66807 68990 66830 69997
rect 66990 69997 70020 70020
rect 66990 68990 67013 69997
rect 66807 67990 67013 68990
rect 66807 67013 66830 67990
rect 63800 66990 66830 67013
rect 66990 67013 67013 67990
rect 69997 68990 70020 69997
rect 70180 69997 73210 70020
rect 70180 68990 70203 69997
rect 69997 67990 70203 68990
rect 69997 67013 70020 67990
rect 66990 66990 70020 67013
rect 70180 67013 70203 67990
rect 73187 68990 73210 69997
rect 73370 69997 76400 70020
rect 73370 68990 73393 69997
rect 73187 67990 73393 68990
rect 73187 67013 73210 67990
rect 70180 66990 73210 67013
rect 73370 67013 73393 67990
rect 76377 68990 76400 69997
rect 76560 69997 79590 70020
rect 76560 68990 76583 69997
rect 76377 67990 76583 68990
rect 76377 67013 76400 67990
rect 73370 66990 76400 67013
rect 76560 67013 76583 67990
rect 79567 68990 79590 69997
rect 79750 69997 82780 70020
rect 79750 68990 79773 69997
rect 79567 67990 79773 68990
rect 79567 67013 79590 67990
rect 76560 66990 79590 67013
rect 79750 67013 79773 67990
rect 82757 68990 82780 69997
rect 82940 69997 85970 70020
rect 82940 68990 82963 69997
rect 82757 67990 82963 68990
rect 82757 67013 82780 67990
rect 79750 66990 82780 67013
rect 82940 67013 82963 67990
rect 85947 68990 85970 69997
rect 86130 69997 89160 70020
rect 86130 68990 86153 69997
rect 85947 67990 86153 68990
rect 85947 67013 85970 67990
rect 82940 66990 85970 67013
rect 86130 67013 86153 67990
rect 89137 68990 89160 69997
rect 89320 69997 92350 70020
rect 89320 68990 89343 69997
rect 89137 67990 89343 68990
rect 89137 67013 89160 67990
rect 86130 66990 89160 67013
rect 89320 67013 89343 67990
rect 92327 68990 92350 69997
rect 92510 69997 95540 70020
rect 92510 68990 92533 69997
rect 92327 67990 92533 68990
rect 92327 67013 92350 67990
rect 89320 66990 92350 67013
rect 92510 67013 92533 67990
rect 95517 68990 95540 69997
rect 95700 69997 98730 70020
rect 95700 68990 95723 69997
rect 95517 67990 95723 68990
rect 95517 67013 95540 67990
rect 92510 66990 95540 67013
rect 95700 67013 95723 67990
rect 98707 68990 98730 69997
rect 98890 69997 101920 70020
rect 98890 68990 98913 69997
rect 98707 67990 98913 68990
rect 98707 67013 98730 67990
rect 95700 66990 98730 67013
rect 98890 67013 98913 67990
rect 101897 68990 101920 69997
rect 102080 69997 105110 70020
rect 102080 68990 102103 69997
rect 101897 67990 102103 68990
rect 101897 67013 101920 67990
rect 98890 66990 101920 67013
rect 102080 67013 102103 67990
rect 105087 68990 105110 69997
rect 105270 69997 108300 70020
rect 105270 68990 105293 69997
rect 105087 67990 105293 68990
rect 105087 67013 105110 67990
rect 102080 66990 105110 67013
rect 105270 67013 105293 67990
rect 108277 68990 108300 69997
rect 108460 69997 111490 70020
rect 108460 68990 108483 69997
rect 108277 67990 108483 68990
rect 108277 67013 108300 67990
rect 105270 66990 108300 67013
rect 108460 67013 108483 67990
rect 111467 68990 111490 69997
rect 111650 69997 114680 70020
rect 111650 68990 111673 69997
rect 111467 67990 111673 68990
rect 111467 67013 111490 67990
rect 108460 66990 111490 67013
rect 111650 67013 111673 67990
rect 114657 68990 114680 69997
rect 114840 69997 117870 70020
rect 114840 68990 114863 69997
rect 114657 67990 114863 68990
rect 114657 67013 114680 67990
rect 111650 66990 114680 67013
rect 114840 67013 114863 67990
rect 117847 68990 117870 69997
rect 118030 69997 121060 70020
rect 118030 68990 118053 69997
rect 117847 67990 118053 68990
rect 117847 67013 117870 67990
rect 114840 66990 117870 67013
rect 118030 67013 118053 67990
rect 121037 68990 121060 69997
rect 121220 69997 124250 70020
rect 121220 68990 121243 69997
rect 121037 67990 121243 68990
rect 121037 67013 121060 67990
rect 118030 66990 121060 67013
rect 121220 67013 121243 67990
rect 124227 68990 124250 69997
rect 124410 69997 127440 70020
rect 124410 68990 124433 69997
rect 124227 67990 124433 68990
rect 124227 67013 124250 67990
rect 121220 66990 124250 67013
rect 124410 67013 124433 67990
rect 127417 68990 127440 69997
rect 127600 69997 130630 70020
rect 127600 68990 127623 69997
rect 127417 67990 127623 68990
rect 127417 67013 127440 67990
rect 124410 66990 127440 67013
rect 127600 67013 127623 67990
rect 130607 68990 130630 69997
rect 130790 69997 133820 70020
rect 130790 68990 130813 69997
rect 130607 67990 130813 68990
rect 130607 67013 130630 67990
rect 127600 66990 130630 67013
rect 130790 67013 130813 67990
rect 133797 68990 133820 69997
rect 133980 69997 137010 70020
rect 133980 68990 134003 69997
rect 133797 67990 134003 68990
rect 133797 67013 133820 67990
rect 130790 66990 133820 67013
rect 133980 67013 134003 67990
rect 136987 68990 137010 69997
rect 136987 67990 137170 68990
rect 136987 67013 137010 67990
rect 133980 66990 137010 67013
rect 1000 66830 2000 66990
rect 4190 66830 5190 66990
rect 7380 66830 8380 66990
rect 10570 66830 11570 66990
rect 13760 66830 14760 66990
rect 16950 66830 17950 66990
rect 20140 66830 21140 66990
rect 23330 66830 24330 66990
rect 26520 66830 27520 66990
rect 29710 66830 30710 66990
rect 32900 66830 33900 66990
rect 36090 66830 37090 66990
rect 39280 66830 40280 66990
rect 42470 66830 43470 66990
rect 45660 66830 46660 66990
rect 48850 66830 49850 66990
rect 52040 66830 53040 66990
rect 55230 66830 56230 66990
rect 58420 66830 59420 66990
rect 61610 66830 62610 66990
rect 64800 66830 65800 66990
rect 67990 66830 68990 66990
rect 71180 66830 72180 66990
rect 74370 66830 75370 66990
rect 77560 66830 78560 66990
rect 80750 66830 81750 66990
rect 83940 66830 84940 66990
rect 87130 66830 88130 66990
rect 90320 66830 91320 66990
rect 93510 66830 94510 66990
rect 96700 66830 97700 66990
rect 99890 66830 100890 66990
rect 103080 66830 104080 66990
rect 106270 66830 107270 66990
rect 109460 66830 110460 66990
rect 112650 66830 113650 66990
rect 115840 66830 116840 66990
rect 119030 66830 120030 66990
rect 122220 66830 123220 66990
rect 125410 66830 126410 66990
rect 128600 66830 129600 66990
rect 131790 66830 132790 66990
rect 134980 66830 135980 66990
rect 0 66807 3030 66830
rect 0 63823 23 66807
rect 3007 65800 3030 66807
rect 3190 66807 6220 66830
rect 3190 65800 3213 66807
rect 3007 64800 3213 65800
rect 3007 63823 3030 64800
rect 0 63800 3030 63823
rect 3190 63823 3213 64800
rect 6197 65800 6220 66807
rect 6380 66807 9410 66830
rect 6380 65800 6403 66807
rect 6197 64800 6403 65800
rect 6197 63823 6220 64800
rect 3190 63800 6220 63823
rect 6380 63823 6403 64800
rect 9387 65800 9410 66807
rect 9570 66807 12600 66830
rect 9570 65800 9593 66807
rect 9387 64800 9593 65800
rect 9387 63823 9410 64800
rect 6380 63800 9410 63823
rect 9570 63823 9593 64800
rect 12577 65800 12600 66807
rect 12760 66807 15790 66830
rect 12760 65800 12783 66807
rect 12577 64800 12783 65800
rect 12577 63823 12600 64800
rect 9570 63800 12600 63823
rect 12760 63823 12783 64800
rect 15767 65800 15790 66807
rect 15950 66807 18980 66830
rect 15950 65800 15973 66807
rect 15767 64800 15973 65800
rect 15767 63823 15790 64800
rect 12760 63800 15790 63823
rect 15950 63823 15973 64800
rect 18957 65800 18980 66807
rect 19140 66807 22170 66830
rect 19140 65800 19163 66807
rect 18957 64800 19163 65800
rect 18957 63823 18980 64800
rect 15950 63800 18980 63823
rect 19140 63823 19163 64800
rect 22147 65800 22170 66807
rect 22330 66807 25360 66830
rect 22330 65800 22353 66807
rect 22147 64800 22353 65800
rect 22147 63823 22170 64800
rect 19140 63800 22170 63823
rect 22330 63823 22353 64800
rect 25337 65800 25360 66807
rect 25520 66807 28550 66830
rect 25520 65800 25543 66807
rect 25337 64800 25543 65800
rect 25337 63823 25360 64800
rect 22330 63800 25360 63823
rect 25520 63823 25543 64800
rect 28527 65800 28550 66807
rect 28710 66807 31740 66830
rect 28710 65800 28733 66807
rect 28527 64800 28733 65800
rect 28527 63823 28550 64800
rect 25520 63800 28550 63823
rect 28710 63823 28733 64800
rect 31717 65800 31740 66807
rect 31900 66807 34930 66830
rect 31900 65800 31923 66807
rect 31717 64800 31923 65800
rect 31717 63823 31740 64800
rect 28710 63800 31740 63823
rect 31900 63823 31923 64800
rect 34907 65800 34930 66807
rect 35090 66807 38120 66830
rect 35090 65800 35113 66807
rect 34907 64800 35113 65800
rect 34907 63823 34930 64800
rect 31900 63800 34930 63823
rect 35090 63823 35113 64800
rect 38097 65800 38120 66807
rect 38280 66807 41310 66830
rect 38280 65800 38303 66807
rect 38097 64800 38303 65800
rect 38097 63823 38120 64800
rect 35090 63800 38120 63823
rect 38280 63823 38303 64800
rect 41287 65800 41310 66807
rect 41470 66807 44500 66830
rect 41470 65800 41493 66807
rect 41287 64800 41493 65800
rect 41287 63823 41310 64800
rect 38280 63800 41310 63823
rect 41470 63823 41493 64800
rect 44477 65800 44500 66807
rect 44660 66807 47690 66830
rect 44660 65800 44683 66807
rect 44477 64800 44683 65800
rect 44477 63823 44500 64800
rect 41470 63800 44500 63823
rect 44660 63823 44683 64800
rect 47667 65800 47690 66807
rect 47850 66807 50880 66830
rect 47850 65800 47873 66807
rect 47667 64800 47873 65800
rect 47667 63823 47690 64800
rect 44660 63800 47690 63823
rect 47850 63823 47873 64800
rect 50857 65800 50880 66807
rect 51040 66807 54070 66830
rect 51040 65800 51063 66807
rect 50857 64800 51063 65800
rect 50857 63823 50880 64800
rect 47850 63800 50880 63823
rect 51040 63823 51063 64800
rect 54047 65800 54070 66807
rect 54230 66807 57260 66830
rect 54230 65800 54253 66807
rect 54047 64800 54253 65800
rect 54047 63823 54070 64800
rect 51040 63800 54070 63823
rect 54230 63823 54253 64800
rect 57237 65800 57260 66807
rect 57420 66807 60450 66830
rect 57420 65800 57443 66807
rect 57237 64800 57443 65800
rect 57237 63823 57260 64800
rect 54230 63800 57260 63823
rect 57420 63823 57443 64800
rect 60427 65800 60450 66807
rect 60610 66807 63640 66830
rect 60610 65800 60633 66807
rect 60427 64800 60633 65800
rect 60427 63823 60450 64800
rect 57420 63800 60450 63823
rect 60610 63823 60633 64800
rect 63617 65800 63640 66807
rect 63800 66807 66830 66830
rect 63800 65800 63823 66807
rect 63617 64800 63823 65800
rect 63617 63823 63640 64800
rect 60610 63800 63640 63823
rect 63800 63823 63823 64800
rect 66807 65800 66830 66807
rect 66990 66807 70020 66830
rect 66990 65800 67013 66807
rect 66807 64800 67013 65800
rect 66807 63823 66830 64800
rect 63800 63800 66830 63823
rect 66990 63823 67013 64800
rect 69997 65800 70020 66807
rect 70180 66807 73210 66830
rect 70180 65800 70203 66807
rect 69997 64800 70203 65800
rect 69997 63823 70020 64800
rect 66990 63800 70020 63823
rect 70180 63823 70203 64800
rect 73187 65800 73210 66807
rect 73370 66807 76400 66830
rect 73370 65800 73393 66807
rect 73187 64800 73393 65800
rect 73187 63823 73210 64800
rect 70180 63800 73210 63823
rect 73370 63823 73393 64800
rect 76377 65800 76400 66807
rect 76560 66807 79590 66830
rect 76560 65800 76583 66807
rect 76377 64800 76583 65800
rect 76377 63823 76400 64800
rect 73370 63800 76400 63823
rect 76560 63823 76583 64800
rect 79567 65800 79590 66807
rect 79750 66807 82780 66830
rect 79750 65800 79773 66807
rect 79567 64800 79773 65800
rect 79567 63823 79590 64800
rect 76560 63800 79590 63823
rect 79750 63823 79773 64800
rect 82757 65800 82780 66807
rect 82940 66807 85970 66830
rect 82940 65800 82963 66807
rect 82757 64800 82963 65800
rect 82757 63823 82780 64800
rect 79750 63800 82780 63823
rect 82940 63823 82963 64800
rect 85947 65800 85970 66807
rect 86130 66807 89160 66830
rect 86130 65800 86153 66807
rect 85947 64800 86153 65800
rect 85947 63823 85970 64800
rect 82940 63800 85970 63823
rect 86130 63823 86153 64800
rect 89137 65800 89160 66807
rect 89320 66807 92350 66830
rect 89320 65800 89343 66807
rect 89137 64800 89343 65800
rect 89137 63823 89160 64800
rect 86130 63800 89160 63823
rect 89320 63823 89343 64800
rect 92327 65800 92350 66807
rect 92510 66807 95540 66830
rect 92510 65800 92533 66807
rect 92327 64800 92533 65800
rect 92327 63823 92350 64800
rect 89320 63800 92350 63823
rect 92510 63823 92533 64800
rect 95517 65800 95540 66807
rect 95700 66807 98730 66830
rect 95700 65800 95723 66807
rect 95517 64800 95723 65800
rect 95517 63823 95540 64800
rect 92510 63800 95540 63823
rect 95700 63823 95723 64800
rect 98707 65800 98730 66807
rect 98890 66807 101920 66830
rect 98890 65800 98913 66807
rect 98707 64800 98913 65800
rect 98707 63823 98730 64800
rect 95700 63800 98730 63823
rect 98890 63823 98913 64800
rect 101897 65800 101920 66807
rect 102080 66807 105110 66830
rect 102080 65800 102103 66807
rect 101897 64800 102103 65800
rect 101897 63823 101920 64800
rect 98890 63800 101920 63823
rect 102080 63823 102103 64800
rect 105087 65800 105110 66807
rect 105270 66807 108300 66830
rect 105270 65800 105293 66807
rect 105087 64800 105293 65800
rect 105087 63823 105110 64800
rect 102080 63800 105110 63823
rect 105270 63823 105293 64800
rect 108277 65800 108300 66807
rect 108460 66807 111490 66830
rect 108460 65800 108483 66807
rect 108277 64800 108483 65800
rect 108277 63823 108300 64800
rect 105270 63800 108300 63823
rect 108460 63823 108483 64800
rect 111467 65800 111490 66807
rect 111650 66807 114680 66830
rect 111650 65800 111673 66807
rect 111467 64800 111673 65800
rect 111467 63823 111490 64800
rect 108460 63800 111490 63823
rect 111650 63823 111673 64800
rect 114657 65800 114680 66807
rect 114840 66807 117870 66830
rect 114840 65800 114863 66807
rect 114657 64800 114863 65800
rect 114657 63823 114680 64800
rect 111650 63800 114680 63823
rect 114840 63823 114863 64800
rect 117847 65800 117870 66807
rect 118030 66807 121060 66830
rect 118030 65800 118053 66807
rect 117847 64800 118053 65800
rect 117847 63823 117870 64800
rect 114840 63800 117870 63823
rect 118030 63823 118053 64800
rect 121037 65800 121060 66807
rect 121220 66807 124250 66830
rect 121220 65800 121243 66807
rect 121037 64800 121243 65800
rect 121037 63823 121060 64800
rect 118030 63800 121060 63823
rect 121220 63823 121243 64800
rect 124227 65800 124250 66807
rect 124410 66807 127440 66830
rect 124410 65800 124433 66807
rect 124227 64800 124433 65800
rect 124227 63823 124250 64800
rect 121220 63800 124250 63823
rect 124410 63823 124433 64800
rect 127417 65800 127440 66807
rect 127600 66807 130630 66830
rect 127600 65800 127623 66807
rect 127417 64800 127623 65800
rect 127417 63823 127440 64800
rect 124410 63800 127440 63823
rect 127600 63823 127623 64800
rect 130607 65800 130630 66807
rect 130790 66807 133820 66830
rect 130790 65800 130813 66807
rect 130607 64800 130813 65800
rect 130607 63823 130630 64800
rect 127600 63800 130630 63823
rect 130790 63823 130813 64800
rect 133797 65800 133820 66807
rect 133980 66807 137010 66830
rect 133980 65800 134003 66807
rect 133797 64800 134003 65800
rect 133797 63823 133820 64800
rect 130790 63800 133820 63823
rect 133980 63823 134003 64800
rect 136987 65800 137010 66807
rect 136987 64800 137170 65800
rect 136987 63823 137010 64800
rect 133980 63800 137010 63823
rect 1000 63640 2000 63800
rect 4190 63640 5190 63800
rect 7380 63640 8380 63800
rect 10570 63640 11570 63800
rect 13760 63640 14760 63800
rect 16950 63640 17950 63800
rect 20140 63640 21140 63800
rect 23330 63640 24330 63800
rect 26520 63640 27520 63800
rect 29710 63640 30710 63800
rect 32900 63640 33900 63800
rect 36090 63640 37090 63800
rect 39280 63640 40280 63800
rect 42470 63640 43470 63800
rect 45660 63640 46660 63800
rect 48850 63640 49850 63800
rect 52040 63640 53040 63800
rect 55230 63640 56230 63800
rect 58420 63640 59420 63800
rect 61610 63640 62610 63800
rect 64800 63640 65800 63800
rect 67990 63640 68990 63800
rect 71180 63640 72180 63800
rect 74370 63640 75370 63800
rect 77560 63640 78560 63800
rect 80750 63640 81750 63800
rect 83940 63640 84940 63800
rect 87130 63640 88130 63800
rect 90320 63640 91320 63800
rect 93510 63640 94510 63800
rect 96700 63640 97700 63800
rect 99890 63640 100890 63800
rect 103080 63640 104080 63800
rect 106270 63640 107270 63800
rect 109460 63640 110460 63800
rect 112650 63640 113650 63800
rect 115840 63640 116840 63800
rect 119030 63640 120030 63800
rect 122220 63640 123220 63800
rect 125410 63640 126410 63800
rect 128600 63640 129600 63800
rect 131790 63640 132790 63800
rect 134980 63640 135980 63800
rect 0 63617 3030 63640
rect 0 60633 23 63617
rect 3007 62610 3030 63617
rect 3190 63617 6220 63640
rect 3190 62610 3213 63617
rect 3007 61610 3213 62610
rect 3007 60633 3030 61610
rect 0 60610 3030 60633
rect 3190 60633 3213 61610
rect 6197 62610 6220 63617
rect 6380 63617 9410 63640
rect 6380 62610 6403 63617
rect 6197 61610 6403 62610
rect 6197 60633 6220 61610
rect 3190 60610 6220 60633
rect 6380 60633 6403 61610
rect 9387 62610 9410 63617
rect 9570 63617 12600 63640
rect 9570 62610 9593 63617
rect 9387 61610 9593 62610
rect 9387 60633 9410 61610
rect 6380 60610 9410 60633
rect 9570 60633 9593 61610
rect 12577 62610 12600 63617
rect 12760 63617 15790 63640
rect 12760 62610 12783 63617
rect 12577 61610 12783 62610
rect 12577 60633 12600 61610
rect 9570 60610 12600 60633
rect 12760 60633 12783 61610
rect 15767 62610 15790 63617
rect 15950 63617 18980 63640
rect 15950 62610 15973 63617
rect 15767 61610 15973 62610
rect 15767 60633 15790 61610
rect 12760 60610 15790 60633
rect 15950 60633 15973 61610
rect 18957 62610 18980 63617
rect 19140 63617 22170 63640
rect 19140 62610 19163 63617
rect 18957 61610 19163 62610
rect 18957 60633 18980 61610
rect 15950 60610 18980 60633
rect 19140 60633 19163 61610
rect 22147 62610 22170 63617
rect 22330 63617 25360 63640
rect 22330 62610 22353 63617
rect 22147 61610 22353 62610
rect 22147 60633 22170 61610
rect 19140 60610 22170 60633
rect 22330 60633 22353 61610
rect 25337 62610 25360 63617
rect 25520 63617 28550 63640
rect 25520 62610 25543 63617
rect 25337 61610 25543 62610
rect 25337 60633 25360 61610
rect 22330 60610 25360 60633
rect 25520 60633 25543 61610
rect 28527 62610 28550 63617
rect 28710 63617 31740 63640
rect 28710 62610 28733 63617
rect 28527 61610 28733 62610
rect 28527 60633 28550 61610
rect 25520 60610 28550 60633
rect 28710 60633 28733 61610
rect 31717 62610 31740 63617
rect 31900 63617 34930 63640
rect 31900 62610 31923 63617
rect 31717 61610 31923 62610
rect 31717 60633 31740 61610
rect 28710 60610 31740 60633
rect 31900 60633 31923 61610
rect 34907 62610 34930 63617
rect 35090 63617 38120 63640
rect 35090 62610 35113 63617
rect 34907 61610 35113 62610
rect 34907 60633 34930 61610
rect 31900 60610 34930 60633
rect 35090 60633 35113 61610
rect 38097 62610 38120 63617
rect 38280 63617 41310 63640
rect 38280 62610 38303 63617
rect 38097 61610 38303 62610
rect 38097 60633 38120 61610
rect 35090 60610 38120 60633
rect 38280 60633 38303 61610
rect 41287 62610 41310 63617
rect 41470 63617 44500 63640
rect 41470 62610 41493 63617
rect 41287 61610 41493 62610
rect 41287 60633 41310 61610
rect 38280 60610 41310 60633
rect 41470 60633 41493 61610
rect 44477 62610 44500 63617
rect 44660 63617 47690 63640
rect 44660 62610 44683 63617
rect 44477 61610 44683 62610
rect 44477 60633 44500 61610
rect 41470 60610 44500 60633
rect 44660 60633 44683 61610
rect 47667 62610 47690 63617
rect 47850 63617 50880 63640
rect 47850 62610 47873 63617
rect 47667 61610 47873 62610
rect 47667 60633 47690 61610
rect 44660 60610 47690 60633
rect 47850 60633 47873 61610
rect 50857 62610 50880 63617
rect 51040 63617 54070 63640
rect 51040 62610 51063 63617
rect 50857 61610 51063 62610
rect 50857 60633 50880 61610
rect 47850 60610 50880 60633
rect 51040 60633 51063 61610
rect 54047 62610 54070 63617
rect 54230 63617 57260 63640
rect 54230 62610 54253 63617
rect 54047 61610 54253 62610
rect 54047 60633 54070 61610
rect 51040 60610 54070 60633
rect 54230 60633 54253 61610
rect 57237 62610 57260 63617
rect 57420 63617 60450 63640
rect 57420 62610 57443 63617
rect 57237 61610 57443 62610
rect 57237 60633 57260 61610
rect 54230 60610 57260 60633
rect 57420 60633 57443 61610
rect 60427 62610 60450 63617
rect 60610 63617 63640 63640
rect 60610 62610 60633 63617
rect 60427 61610 60633 62610
rect 60427 60633 60450 61610
rect 57420 60610 60450 60633
rect 60610 60633 60633 61610
rect 63617 62610 63640 63617
rect 63800 63617 66830 63640
rect 63800 62610 63823 63617
rect 63617 61610 63823 62610
rect 63617 60633 63640 61610
rect 60610 60610 63640 60633
rect 63800 60633 63823 61610
rect 66807 62610 66830 63617
rect 66990 63617 70020 63640
rect 66990 62610 67013 63617
rect 66807 61610 67013 62610
rect 66807 60633 66830 61610
rect 63800 60610 66830 60633
rect 66990 60633 67013 61610
rect 69997 62610 70020 63617
rect 70180 63617 73210 63640
rect 70180 62610 70203 63617
rect 69997 61610 70203 62610
rect 69997 60633 70020 61610
rect 66990 60610 70020 60633
rect 70180 60633 70203 61610
rect 73187 62610 73210 63617
rect 73370 63617 76400 63640
rect 73370 62610 73393 63617
rect 73187 61610 73393 62610
rect 73187 60633 73210 61610
rect 70180 60610 73210 60633
rect 73370 60633 73393 61610
rect 76377 62610 76400 63617
rect 76560 63617 79590 63640
rect 76560 62610 76583 63617
rect 76377 61610 76583 62610
rect 76377 60633 76400 61610
rect 73370 60610 76400 60633
rect 76560 60633 76583 61610
rect 79567 62610 79590 63617
rect 79750 63617 82780 63640
rect 79750 62610 79773 63617
rect 79567 61610 79773 62610
rect 79567 60633 79590 61610
rect 76560 60610 79590 60633
rect 79750 60633 79773 61610
rect 82757 62610 82780 63617
rect 82940 63617 85970 63640
rect 82940 62610 82963 63617
rect 82757 61610 82963 62610
rect 82757 60633 82780 61610
rect 79750 60610 82780 60633
rect 82940 60633 82963 61610
rect 85947 62610 85970 63617
rect 86130 63617 89160 63640
rect 86130 62610 86153 63617
rect 85947 61610 86153 62610
rect 85947 60633 85970 61610
rect 82940 60610 85970 60633
rect 86130 60633 86153 61610
rect 89137 62610 89160 63617
rect 89320 63617 92350 63640
rect 89320 62610 89343 63617
rect 89137 61610 89343 62610
rect 89137 60633 89160 61610
rect 86130 60610 89160 60633
rect 89320 60633 89343 61610
rect 92327 62610 92350 63617
rect 92510 63617 95540 63640
rect 92510 62610 92533 63617
rect 92327 61610 92533 62610
rect 92327 60633 92350 61610
rect 89320 60610 92350 60633
rect 92510 60633 92533 61610
rect 95517 62610 95540 63617
rect 95700 63617 98730 63640
rect 95700 62610 95723 63617
rect 95517 61610 95723 62610
rect 95517 60633 95540 61610
rect 92510 60610 95540 60633
rect 95700 60633 95723 61610
rect 98707 62610 98730 63617
rect 98890 63617 101920 63640
rect 98890 62610 98913 63617
rect 98707 61610 98913 62610
rect 98707 60633 98730 61610
rect 95700 60610 98730 60633
rect 98890 60633 98913 61610
rect 101897 62610 101920 63617
rect 102080 63617 105110 63640
rect 102080 62610 102103 63617
rect 101897 61610 102103 62610
rect 101897 60633 101920 61610
rect 98890 60610 101920 60633
rect 102080 60633 102103 61610
rect 105087 62610 105110 63617
rect 105270 63617 108300 63640
rect 105270 62610 105293 63617
rect 105087 61610 105293 62610
rect 105087 60633 105110 61610
rect 102080 60610 105110 60633
rect 105270 60633 105293 61610
rect 108277 62610 108300 63617
rect 108460 63617 111490 63640
rect 108460 62610 108483 63617
rect 108277 61610 108483 62610
rect 108277 60633 108300 61610
rect 105270 60610 108300 60633
rect 108460 60633 108483 61610
rect 111467 62610 111490 63617
rect 111650 63617 114680 63640
rect 111650 62610 111673 63617
rect 111467 61610 111673 62610
rect 111467 60633 111490 61610
rect 108460 60610 111490 60633
rect 111650 60633 111673 61610
rect 114657 62610 114680 63617
rect 114840 63617 117870 63640
rect 114840 62610 114863 63617
rect 114657 61610 114863 62610
rect 114657 60633 114680 61610
rect 111650 60610 114680 60633
rect 114840 60633 114863 61610
rect 117847 62610 117870 63617
rect 118030 63617 121060 63640
rect 118030 62610 118053 63617
rect 117847 61610 118053 62610
rect 117847 60633 117870 61610
rect 114840 60610 117870 60633
rect 118030 60633 118053 61610
rect 121037 62610 121060 63617
rect 121220 63617 124250 63640
rect 121220 62610 121243 63617
rect 121037 61610 121243 62610
rect 121037 60633 121060 61610
rect 118030 60610 121060 60633
rect 121220 60633 121243 61610
rect 124227 62610 124250 63617
rect 124410 63617 127440 63640
rect 124410 62610 124433 63617
rect 124227 61610 124433 62610
rect 124227 60633 124250 61610
rect 121220 60610 124250 60633
rect 124410 60633 124433 61610
rect 127417 62610 127440 63617
rect 127600 63617 130630 63640
rect 127600 62610 127623 63617
rect 127417 61610 127623 62610
rect 127417 60633 127440 61610
rect 124410 60610 127440 60633
rect 127600 60633 127623 61610
rect 130607 62610 130630 63617
rect 130790 63617 133820 63640
rect 130790 62610 130813 63617
rect 130607 61610 130813 62610
rect 130607 60633 130630 61610
rect 127600 60610 130630 60633
rect 130790 60633 130813 61610
rect 133797 62610 133820 63617
rect 133980 63617 137010 63640
rect 133980 62610 134003 63617
rect 133797 61610 134003 62610
rect 133797 60633 133820 61610
rect 130790 60610 133820 60633
rect 133980 60633 134003 61610
rect 136987 62610 137010 63617
rect 136987 61610 137170 62610
rect 136987 60633 137010 61610
rect 133980 60610 137010 60633
rect 1000 60450 2000 60610
rect 4190 60450 5190 60610
rect 7380 60450 8380 60610
rect 10570 60450 11570 60610
rect 13760 60450 14760 60610
rect 16950 60450 17950 60610
rect 20140 60450 21140 60610
rect 23330 60450 24330 60610
rect 26520 60450 27520 60610
rect 29710 60450 30710 60610
rect 32900 60450 33900 60610
rect 36090 60450 37090 60610
rect 39280 60450 40280 60610
rect 42470 60450 43470 60610
rect 45660 60450 46660 60610
rect 48850 60450 49850 60610
rect 52040 60450 53040 60610
rect 55230 60450 56230 60610
rect 58420 60450 59420 60610
rect 61610 60450 62610 60610
rect 64800 60450 65800 60610
rect 67990 60450 68990 60610
rect 71180 60450 72180 60610
rect 74370 60450 75370 60610
rect 77560 60450 78560 60610
rect 80750 60450 81750 60610
rect 83940 60450 84940 60610
rect 87130 60450 88130 60610
rect 90320 60450 91320 60610
rect 93510 60450 94510 60610
rect 96700 60450 97700 60610
rect 99890 60450 100890 60610
rect 103080 60450 104080 60610
rect 106270 60450 107270 60610
rect 109460 60450 110460 60610
rect 112650 60450 113650 60610
rect 115840 60450 116840 60610
rect 119030 60450 120030 60610
rect 122220 60450 123220 60610
rect 125410 60450 126410 60610
rect 128600 60450 129600 60610
rect 131790 60450 132790 60610
rect 134980 60450 135980 60610
rect 0 60427 3030 60450
rect 0 57443 23 60427
rect 3007 59420 3030 60427
rect 3190 60427 6220 60450
rect 3190 59420 3213 60427
rect 3007 58420 3213 59420
rect 3007 57443 3030 58420
rect 0 57420 3030 57443
rect 3190 57443 3213 58420
rect 6197 59420 6220 60427
rect 6380 60427 9410 60450
rect 6380 59420 6403 60427
rect 6197 58420 6403 59420
rect 6197 57443 6220 58420
rect 3190 57420 6220 57443
rect 6380 57443 6403 58420
rect 9387 59420 9410 60427
rect 9570 60427 12600 60450
rect 9570 59420 9593 60427
rect 9387 58420 9593 59420
rect 9387 57443 9410 58420
rect 6380 57420 9410 57443
rect 9570 57443 9593 58420
rect 12577 59420 12600 60427
rect 12760 60427 15790 60450
rect 12760 59420 12783 60427
rect 12577 58420 12783 59420
rect 12577 57443 12600 58420
rect 9570 57420 12600 57443
rect 12760 57443 12783 58420
rect 15767 59420 15790 60427
rect 15950 60427 18980 60450
rect 15950 59420 15973 60427
rect 15767 58420 15973 59420
rect 15767 57443 15790 58420
rect 12760 57420 15790 57443
rect 15950 57443 15973 58420
rect 18957 59420 18980 60427
rect 19140 60427 22170 60450
rect 19140 59420 19163 60427
rect 18957 58420 19163 59420
rect 18957 57443 18980 58420
rect 15950 57420 18980 57443
rect 19140 57443 19163 58420
rect 22147 59420 22170 60427
rect 22330 60427 25360 60450
rect 22330 59420 22353 60427
rect 22147 58420 22353 59420
rect 22147 57443 22170 58420
rect 19140 57420 22170 57443
rect 22330 57443 22353 58420
rect 25337 59420 25360 60427
rect 25520 60427 28550 60450
rect 25520 59420 25543 60427
rect 25337 58420 25543 59420
rect 25337 57443 25360 58420
rect 22330 57420 25360 57443
rect 25520 57443 25543 58420
rect 28527 59420 28550 60427
rect 28710 60427 31740 60450
rect 28710 59420 28733 60427
rect 28527 58420 28733 59420
rect 28527 57443 28550 58420
rect 25520 57420 28550 57443
rect 28710 57443 28733 58420
rect 31717 59420 31740 60427
rect 31900 60427 34930 60450
rect 31900 59420 31923 60427
rect 31717 58420 31923 59420
rect 31717 57443 31740 58420
rect 28710 57420 31740 57443
rect 31900 57443 31923 58420
rect 34907 59420 34930 60427
rect 35090 60427 38120 60450
rect 35090 59420 35113 60427
rect 34907 58420 35113 59420
rect 34907 57443 34930 58420
rect 31900 57420 34930 57443
rect 35090 57443 35113 58420
rect 38097 59420 38120 60427
rect 38280 60427 41310 60450
rect 38280 59420 38303 60427
rect 38097 58420 38303 59420
rect 38097 57443 38120 58420
rect 35090 57420 38120 57443
rect 38280 57443 38303 58420
rect 41287 59420 41310 60427
rect 41470 60427 44500 60450
rect 41470 59420 41493 60427
rect 41287 58420 41493 59420
rect 41287 57443 41310 58420
rect 38280 57420 41310 57443
rect 41470 57443 41493 58420
rect 44477 59420 44500 60427
rect 44660 60427 47690 60450
rect 44660 59420 44683 60427
rect 44477 58420 44683 59420
rect 44477 57443 44500 58420
rect 41470 57420 44500 57443
rect 44660 57443 44683 58420
rect 47667 59420 47690 60427
rect 47850 60427 50880 60450
rect 47850 59420 47873 60427
rect 47667 58420 47873 59420
rect 47667 57443 47690 58420
rect 44660 57420 47690 57443
rect 47850 57443 47873 58420
rect 50857 59420 50880 60427
rect 51040 60427 54070 60450
rect 51040 59420 51063 60427
rect 50857 58420 51063 59420
rect 50857 57443 50880 58420
rect 47850 57420 50880 57443
rect 51040 57443 51063 58420
rect 54047 59420 54070 60427
rect 54230 60427 57260 60450
rect 54230 59420 54253 60427
rect 54047 58420 54253 59420
rect 54047 57443 54070 58420
rect 51040 57420 54070 57443
rect 54230 57443 54253 58420
rect 57237 59420 57260 60427
rect 57420 60427 60450 60450
rect 57420 59420 57443 60427
rect 57237 58420 57443 59420
rect 57237 57443 57260 58420
rect 54230 57420 57260 57443
rect 57420 57443 57443 58420
rect 60427 59420 60450 60427
rect 60610 60427 63640 60450
rect 60610 59420 60633 60427
rect 60427 58420 60633 59420
rect 60427 57443 60450 58420
rect 57420 57420 60450 57443
rect 60610 57443 60633 58420
rect 63617 59420 63640 60427
rect 63800 60427 66830 60450
rect 63800 59420 63823 60427
rect 63617 58420 63823 59420
rect 63617 57443 63640 58420
rect 60610 57420 63640 57443
rect 63800 57443 63823 58420
rect 66807 59420 66830 60427
rect 66990 60427 70020 60450
rect 66990 59420 67013 60427
rect 66807 58420 67013 59420
rect 66807 57443 66830 58420
rect 63800 57420 66830 57443
rect 66990 57443 67013 58420
rect 69997 59420 70020 60427
rect 70180 60427 73210 60450
rect 70180 59420 70203 60427
rect 69997 58420 70203 59420
rect 69997 57443 70020 58420
rect 66990 57420 70020 57443
rect 70180 57443 70203 58420
rect 73187 59420 73210 60427
rect 73370 60427 76400 60450
rect 73370 59420 73393 60427
rect 73187 58420 73393 59420
rect 73187 57443 73210 58420
rect 70180 57420 73210 57443
rect 73370 57443 73393 58420
rect 76377 59420 76400 60427
rect 76560 60427 79590 60450
rect 76560 59420 76583 60427
rect 76377 58420 76583 59420
rect 76377 57443 76400 58420
rect 73370 57420 76400 57443
rect 76560 57443 76583 58420
rect 79567 59420 79590 60427
rect 79750 60427 82780 60450
rect 79750 59420 79773 60427
rect 79567 58420 79773 59420
rect 79567 57443 79590 58420
rect 76560 57420 79590 57443
rect 79750 57443 79773 58420
rect 82757 59420 82780 60427
rect 82940 60427 85970 60450
rect 82940 59420 82963 60427
rect 82757 58420 82963 59420
rect 82757 57443 82780 58420
rect 79750 57420 82780 57443
rect 82940 57443 82963 58420
rect 85947 59420 85970 60427
rect 86130 60427 89160 60450
rect 86130 59420 86153 60427
rect 85947 58420 86153 59420
rect 85947 57443 85970 58420
rect 82940 57420 85970 57443
rect 86130 57443 86153 58420
rect 89137 59420 89160 60427
rect 89320 60427 92350 60450
rect 89320 59420 89343 60427
rect 89137 58420 89343 59420
rect 89137 57443 89160 58420
rect 86130 57420 89160 57443
rect 89320 57443 89343 58420
rect 92327 59420 92350 60427
rect 92510 60427 95540 60450
rect 92510 59420 92533 60427
rect 92327 58420 92533 59420
rect 92327 57443 92350 58420
rect 89320 57420 92350 57443
rect 92510 57443 92533 58420
rect 95517 59420 95540 60427
rect 95700 60427 98730 60450
rect 95700 59420 95723 60427
rect 95517 58420 95723 59420
rect 95517 57443 95540 58420
rect 92510 57420 95540 57443
rect 95700 57443 95723 58420
rect 98707 59420 98730 60427
rect 98890 60427 101920 60450
rect 98890 59420 98913 60427
rect 98707 58420 98913 59420
rect 98707 57443 98730 58420
rect 95700 57420 98730 57443
rect 98890 57443 98913 58420
rect 101897 59420 101920 60427
rect 102080 60427 105110 60450
rect 102080 59420 102103 60427
rect 101897 58420 102103 59420
rect 101897 57443 101920 58420
rect 98890 57420 101920 57443
rect 102080 57443 102103 58420
rect 105087 59420 105110 60427
rect 105270 60427 108300 60450
rect 105270 59420 105293 60427
rect 105087 58420 105293 59420
rect 105087 57443 105110 58420
rect 102080 57420 105110 57443
rect 105270 57443 105293 58420
rect 108277 59420 108300 60427
rect 108460 60427 111490 60450
rect 108460 59420 108483 60427
rect 108277 58420 108483 59420
rect 108277 57443 108300 58420
rect 105270 57420 108300 57443
rect 108460 57443 108483 58420
rect 111467 59420 111490 60427
rect 111650 60427 114680 60450
rect 111650 59420 111673 60427
rect 111467 58420 111673 59420
rect 111467 57443 111490 58420
rect 108460 57420 111490 57443
rect 111650 57443 111673 58420
rect 114657 59420 114680 60427
rect 114840 60427 117870 60450
rect 114840 59420 114863 60427
rect 114657 58420 114863 59420
rect 114657 57443 114680 58420
rect 111650 57420 114680 57443
rect 114840 57443 114863 58420
rect 117847 59420 117870 60427
rect 118030 60427 121060 60450
rect 118030 59420 118053 60427
rect 117847 58420 118053 59420
rect 117847 57443 117870 58420
rect 114840 57420 117870 57443
rect 118030 57443 118053 58420
rect 121037 59420 121060 60427
rect 121220 60427 124250 60450
rect 121220 59420 121243 60427
rect 121037 58420 121243 59420
rect 121037 57443 121060 58420
rect 118030 57420 121060 57443
rect 121220 57443 121243 58420
rect 124227 59420 124250 60427
rect 124410 60427 127440 60450
rect 124410 59420 124433 60427
rect 124227 58420 124433 59420
rect 124227 57443 124250 58420
rect 121220 57420 124250 57443
rect 124410 57443 124433 58420
rect 127417 59420 127440 60427
rect 127600 60427 130630 60450
rect 127600 59420 127623 60427
rect 127417 58420 127623 59420
rect 127417 57443 127440 58420
rect 124410 57420 127440 57443
rect 127600 57443 127623 58420
rect 130607 59420 130630 60427
rect 130790 60427 133820 60450
rect 130790 59420 130813 60427
rect 130607 58420 130813 59420
rect 130607 57443 130630 58420
rect 127600 57420 130630 57443
rect 130790 57443 130813 58420
rect 133797 59420 133820 60427
rect 133980 60427 137010 60450
rect 133980 59420 134003 60427
rect 133797 58420 134003 59420
rect 133797 57443 133820 58420
rect 130790 57420 133820 57443
rect 133980 57443 134003 58420
rect 136987 59420 137010 60427
rect 136987 58420 137170 59420
rect 136987 57443 137010 58420
rect 133980 57420 137010 57443
rect 1000 57260 2000 57420
rect 4190 57260 5190 57420
rect 7380 57260 8380 57420
rect 10570 57260 11570 57420
rect 13760 57260 14760 57420
rect 16950 57260 17950 57420
rect 20140 57260 21140 57420
rect 23330 57260 24330 57420
rect 26520 57260 27520 57420
rect 29710 57260 30710 57420
rect 32900 57260 33900 57420
rect 36090 57260 37090 57420
rect 39280 57260 40280 57420
rect 42470 57260 43470 57420
rect 45660 57260 46660 57420
rect 48850 57260 49850 57420
rect 52040 57260 53040 57420
rect 55230 57260 56230 57420
rect 58420 57260 59420 57420
rect 61610 57260 62610 57420
rect 64800 57260 65800 57420
rect 67990 57260 68990 57420
rect 71180 57260 72180 57420
rect 74370 57260 75370 57420
rect 77560 57260 78560 57420
rect 80750 57260 81750 57420
rect 83940 57260 84940 57420
rect 87130 57260 88130 57420
rect 90320 57260 91320 57420
rect 93510 57260 94510 57420
rect 96700 57260 97700 57420
rect 99890 57260 100890 57420
rect 103080 57260 104080 57420
rect 106270 57260 107270 57420
rect 109460 57260 110460 57420
rect 112650 57260 113650 57420
rect 115840 57260 116840 57420
rect 119030 57260 120030 57420
rect 122220 57260 123220 57420
rect 125410 57260 126410 57420
rect 128600 57260 129600 57420
rect 131790 57260 132790 57420
rect 134980 57260 135980 57420
rect 0 57237 3030 57260
rect 0 54253 23 57237
rect 3007 56230 3030 57237
rect 3190 57237 6220 57260
rect 3190 56230 3213 57237
rect 3007 55230 3213 56230
rect 3007 54253 3030 55230
rect 0 54230 3030 54253
rect 3190 54253 3213 55230
rect 6197 56230 6220 57237
rect 6380 57237 9410 57260
rect 6380 56230 6403 57237
rect 6197 55230 6403 56230
rect 6197 54253 6220 55230
rect 3190 54230 6220 54253
rect 6380 54253 6403 55230
rect 9387 56230 9410 57237
rect 9570 57237 12600 57260
rect 9570 56230 9593 57237
rect 9387 55230 9593 56230
rect 9387 54253 9410 55230
rect 6380 54230 9410 54253
rect 9570 54253 9593 55230
rect 12577 56230 12600 57237
rect 12760 57237 15790 57260
rect 12760 56230 12783 57237
rect 12577 55230 12783 56230
rect 12577 54253 12600 55230
rect 9570 54230 12600 54253
rect 12760 54253 12783 55230
rect 15767 56230 15790 57237
rect 15950 57237 18980 57260
rect 15950 56230 15973 57237
rect 15767 55230 15973 56230
rect 15767 54253 15790 55230
rect 12760 54230 15790 54253
rect 15950 54253 15973 55230
rect 18957 56230 18980 57237
rect 19140 57237 22170 57260
rect 19140 56230 19163 57237
rect 18957 55230 19163 56230
rect 18957 54253 18980 55230
rect 15950 54230 18980 54253
rect 19140 54253 19163 55230
rect 22147 56230 22170 57237
rect 22330 57237 25360 57260
rect 22330 56230 22353 57237
rect 22147 55230 22353 56230
rect 22147 54253 22170 55230
rect 19140 54230 22170 54253
rect 22330 54253 22353 55230
rect 25337 56230 25360 57237
rect 25520 57237 28550 57260
rect 25520 56230 25543 57237
rect 25337 55230 25543 56230
rect 25337 54253 25360 55230
rect 22330 54230 25360 54253
rect 25520 54253 25543 55230
rect 28527 56230 28550 57237
rect 28710 57237 31740 57260
rect 28710 56230 28733 57237
rect 28527 55230 28733 56230
rect 28527 54253 28550 55230
rect 25520 54230 28550 54253
rect 28710 54253 28733 55230
rect 31717 56230 31740 57237
rect 31900 57237 34930 57260
rect 31900 56230 31923 57237
rect 31717 55230 31923 56230
rect 31717 54253 31740 55230
rect 28710 54230 31740 54253
rect 31900 54253 31923 55230
rect 34907 56230 34930 57237
rect 35090 57237 38120 57260
rect 35090 56230 35113 57237
rect 34907 55230 35113 56230
rect 34907 54253 34930 55230
rect 31900 54230 34930 54253
rect 35090 54253 35113 55230
rect 38097 56230 38120 57237
rect 38280 57237 41310 57260
rect 38280 56230 38303 57237
rect 38097 55230 38303 56230
rect 38097 54253 38120 55230
rect 35090 54230 38120 54253
rect 38280 54253 38303 55230
rect 41287 56230 41310 57237
rect 41470 57237 44500 57260
rect 41470 56230 41493 57237
rect 41287 55230 41493 56230
rect 41287 54253 41310 55230
rect 38280 54230 41310 54253
rect 41470 54253 41493 55230
rect 44477 56230 44500 57237
rect 44660 57237 47690 57260
rect 44660 56230 44683 57237
rect 44477 55230 44683 56230
rect 44477 54253 44500 55230
rect 41470 54230 44500 54253
rect 44660 54253 44683 55230
rect 47667 56230 47690 57237
rect 47850 57237 50880 57260
rect 47850 56230 47873 57237
rect 47667 55230 47873 56230
rect 47667 54253 47690 55230
rect 44660 54230 47690 54253
rect 47850 54253 47873 55230
rect 50857 56230 50880 57237
rect 51040 57237 54070 57260
rect 51040 56230 51063 57237
rect 50857 55230 51063 56230
rect 50857 54253 50880 55230
rect 47850 54230 50880 54253
rect 51040 54253 51063 55230
rect 54047 56230 54070 57237
rect 54230 57237 57260 57260
rect 54230 56230 54253 57237
rect 54047 55230 54253 56230
rect 54047 54253 54070 55230
rect 51040 54230 54070 54253
rect 54230 54253 54253 55230
rect 57237 56230 57260 57237
rect 57420 57237 60450 57260
rect 57420 56230 57443 57237
rect 57237 55230 57443 56230
rect 57237 54253 57260 55230
rect 54230 54230 57260 54253
rect 57420 54253 57443 55230
rect 60427 56230 60450 57237
rect 60610 57237 63640 57260
rect 60610 56230 60633 57237
rect 60427 55230 60633 56230
rect 60427 54253 60450 55230
rect 57420 54230 60450 54253
rect 60610 54253 60633 55230
rect 63617 56230 63640 57237
rect 63800 57237 66830 57260
rect 63800 56230 63823 57237
rect 63617 55230 63823 56230
rect 63617 54253 63640 55230
rect 60610 54230 63640 54253
rect 63800 54253 63823 55230
rect 66807 56230 66830 57237
rect 66990 57237 70020 57260
rect 66990 56230 67013 57237
rect 66807 55230 67013 56230
rect 66807 54253 66830 55230
rect 63800 54230 66830 54253
rect 66990 54253 67013 55230
rect 69997 56230 70020 57237
rect 70180 57237 73210 57260
rect 70180 56230 70203 57237
rect 69997 55230 70203 56230
rect 69997 54253 70020 55230
rect 66990 54230 70020 54253
rect 70180 54253 70203 55230
rect 73187 56230 73210 57237
rect 73370 57237 76400 57260
rect 73370 56230 73393 57237
rect 73187 55230 73393 56230
rect 73187 54253 73210 55230
rect 70180 54230 73210 54253
rect 73370 54253 73393 55230
rect 76377 56230 76400 57237
rect 76560 57237 79590 57260
rect 76560 56230 76583 57237
rect 76377 55230 76583 56230
rect 76377 54253 76400 55230
rect 73370 54230 76400 54253
rect 76560 54253 76583 55230
rect 79567 56230 79590 57237
rect 79750 57237 82780 57260
rect 79750 56230 79773 57237
rect 79567 55230 79773 56230
rect 79567 54253 79590 55230
rect 76560 54230 79590 54253
rect 79750 54253 79773 55230
rect 82757 56230 82780 57237
rect 82940 57237 85970 57260
rect 82940 56230 82963 57237
rect 82757 55230 82963 56230
rect 82757 54253 82780 55230
rect 79750 54230 82780 54253
rect 82940 54253 82963 55230
rect 85947 56230 85970 57237
rect 86130 57237 89160 57260
rect 86130 56230 86153 57237
rect 85947 55230 86153 56230
rect 85947 54253 85970 55230
rect 82940 54230 85970 54253
rect 86130 54253 86153 55230
rect 89137 56230 89160 57237
rect 89320 57237 92350 57260
rect 89320 56230 89343 57237
rect 89137 55230 89343 56230
rect 89137 54253 89160 55230
rect 86130 54230 89160 54253
rect 89320 54253 89343 55230
rect 92327 56230 92350 57237
rect 92510 57237 95540 57260
rect 92510 56230 92533 57237
rect 92327 55230 92533 56230
rect 92327 54253 92350 55230
rect 89320 54230 92350 54253
rect 92510 54253 92533 55230
rect 95517 56230 95540 57237
rect 95700 57237 98730 57260
rect 95700 56230 95723 57237
rect 95517 55230 95723 56230
rect 95517 54253 95540 55230
rect 92510 54230 95540 54253
rect 95700 54253 95723 55230
rect 98707 56230 98730 57237
rect 98890 57237 101920 57260
rect 98890 56230 98913 57237
rect 98707 55230 98913 56230
rect 98707 54253 98730 55230
rect 95700 54230 98730 54253
rect 98890 54253 98913 55230
rect 101897 56230 101920 57237
rect 102080 57237 105110 57260
rect 102080 56230 102103 57237
rect 101897 55230 102103 56230
rect 101897 54253 101920 55230
rect 98890 54230 101920 54253
rect 102080 54253 102103 55230
rect 105087 56230 105110 57237
rect 105270 57237 108300 57260
rect 105270 56230 105293 57237
rect 105087 55230 105293 56230
rect 105087 54253 105110 55230
rect 102080 54230 105110 54253
rect 105270 54253 105293 55230
rect 108277 56230 108300 57237
rect 108460 57237 111490 57260
rect 108460 56230 108483 57237
rect 108277 55230 108483 56230
rect 108277 54253 108300 55230
rect 105270 54230 108300 54253
rect 108460 54253 108483 55230
rect 111467 56230 111490 57237
rect 111650 57237 114680 57260
rect 111650 56230 111673 57237
rect 111467 55230 111673 56230
rect 111467 54253 111490 55230
rect 108460 54230 111490 54253
rect 111650 54253 111673 55230
rect 114657 56230 114680 57237
rect 114840 57237 117870 57260
rect 114840 56230 114863 57237
rect 114657 55230 114863 56230
rect 114657 54253 114680 55230
rect 111650 54230 114680 54253
rect 114840 54253 114863 55230
rect 117847 56230 117870 57237
rect 118030 57237 121060 57260
rect 118030 56230 118053 57237
rect 117847 55230 118053 56230
rect 117847 54253 117870 55230
rect 114840 54230 117870 54253
rect 118030 54253 118053 55230
rect 121037 56230 121060 57237
rect 121220 57237 124250 57260
rect 121220 56230 121243 57237
rect 121037 55230 121243 56230
rect 121037 54253 121060 55230
rect 118030 54230 121060 54253
rect 121220 54253 121243 55230
rect 124227 56230 124250 57237
rect 124410 57237 127440 57260
rect 124410 56230 124433 57237
rect 124227 55230 124433 56230
rect 124227 54253 124250 55230
rect 121220 54230 124250 54253
rect 124410 54253 124433 55230
rect 127417 56230 127440 57237
rect 127600 57237 130630 57260
rect 127600 56230 127623 57237
rect 127417 55230 127623 56230
rect 127417 54253 127440 55230
rect 124410 54230 127440 54253
rect 127600 54253 127623 55230
rect 130607 56230 130630 57237
rect 130790 57237 133820 57260
rect 130790 56230 130813 57237
rect 130607 55230 130813 56230
rect 130607 54253 130630 55230
rect 127600 54230 130630 54253
rect 130790 54253 130813 55230
rect 133797 56230 133820 57237
rect 133980 57237 137010 57260
rect 133980 56230 134003 57237
rect 133797 55230 134003 56230
rect 133797 54253 133820 55230
rect 130790 54230 133820 54253
rect 133980 54253 134003 55230
rect 136987 56230 137010 57237
rect 136987 55230 137170 56230
rect 136987 54253 137010 55230
rect 133980 54230 137010 54253
rect 1000 54070 2000 54230
rect 4190 54070 5190 54230
rect 7380 54070 8380 54230
rect 10570 54070 11570 54230
rect 13760 54070 14760 54230
rect 16950 54070 17950 54230
rect 20140 54070 21140 54230
rect 23330 54070 24330 54230
rect 26520 54070 27520 54230
rect 29710 54070 30710 54230
rect 32900 54070 33900 54230
rect 36090 54070 37090 54230
rect 39280 54070 40280 54230
rect 42470 54070 43470 54230
rect 45660 54070 46660 54230
rect 48850 54070 49850 54230
rect 52040 54070 53040 54230
rect 55230 54070 56230 54230
rect 58420 54070 59420 54230
rect 61610 54070 62610 54230
rect 64800 54070 65800 54230
rect 67990 54070 68990 54230
rect 71180 54070 72180 54230
rect 74370 54070 75370 54230
rect 77560 54070 78560 54230
rect 80750 54070 81750 54230
rect 83940 54070 84940 54230
rect 87130 54070 88130 54230
rect 90320 54070 91320 54230
rect 93510 54070 94510 54230
rect 96700 54070 97700 54230
rect 99890 54070 100890 54230
rect 103080 54070 104080 54230
rect 106270 54070 107270 54230
rect 109460 54070 110460 54230
rect 112650 54070 113650 54230
rect 115840 54070 116840 54230
rect 119030 54070 120030 54230
rect 122220 54070 123220 54230
rect 125410 54070 126410 54230
rect 128600 54070 129600 54230
rect 131790 54070 132790 54230
rect 134980 54070 135980 54230
rect 0 54047 3030 54070
rect 0 51063 23 54047
rect 3007 53040 3030 54047
rect 3190 54047 6220 54070
rect 3190 53040 3213 54047
rect 3007 52040 3213 53040
rect 3007 51063 3030 52040
rect 0 51040 3030 51063
rect 3190 51063 3213 52040
rect 6197 53040 6220 54047
rect 6380 54047 9410 54070
rect 6380 53040 6403 54047
rect 6197 52040 6403 53040
rect 6197 51063 6220 52040
rect 3190 51040 6220 51063
rect 6380 51063 6403 52040
rect 9387 53040 9410 54047
rect 9570 54047 12600 54070
rect 9570 53040 9593 54047
rect 9387 52040 9593 53040
rect 9387 51063 9410 52040
rect 6380 51040 9410 51063
rect 9570 51063 9593 52040
rect 12577 53040 12600 54047
rect 12760 54047 15790 54070
rect 12760 53040 12783 54047
rect 12577 52040 12783 53040
rect 12577 51063 12600 52040
rect 9570 51040 12600 51063
rect 12760 51063 12783 52040
rect 15767 53040 15790 54047
rect 15950 54047 18980 54070
rect 15950 53040 15973 54047
rect 15767 52040 15973 53040
rect 15767 51063 15790 52040
rect 12760 51040 15790 51063
rect 15950 51063 15973 52040
rect 18957 53040 18980 54047
rect 19140 54047 22170 54070
rect 19140 53040 19163 54047
rect 18957 52040 19163 53040
rect 18957 51063 18980 52040
rect 15950 51040 18980 51063
rect 19140 51063 19163 52040
rect 22147 53040 22170 54047
rect 22330 54047 25360 54070
rect 22330 53040 22353 54047
rect 22147 52040 22353 53040
rect 22147 51063 22170 52040
rect 19140 51040 22170 51063
rect 22330 51063 22353 52040
rect 25337 53040 25360 54047
rect 25520 54047 28550 54070
rect 25520 53040 25543 54047
rect 25337 52040 25543 53040
rect 25337 51063 25360 52040
rect 22330 51040 25360 51063
rect 25520 51063 25543 52040
rect 28527 53040 28550 54047
rect 28710 54047 31740 54070
rect 28710 53040 28733 54047
rect 28527 52040 28733 53040
rect 28527 51063 28550 52040
rect 25520 51040 28550 51063
rect 28710 51063 28733 52040
rect 31717 53040 31740 54047
rect 31900 54047 34930 54070
rect 31900 53040 31923 54047
rect 31717 52040 31923 53040
rect 31717 51063 31740 52040
rect 28710 51040 31740 51063
rect 31900 51063 31923 52040
rect 34907 53040 34930 54047
rect 35090 54047 38120 54070
rect 35090 53040 35113 54047
rect 34907 52040 35113 53040
rect 34907 51063 34930 52040
rect 31900 51040 34930 51063
rect 35090 51063 35113 52040
rect 38097 53040 38120 54047
rect 38280 54047 41310 54070
rect 38280 53040 38303 54047
rect 38097 52040 38303 53040
rect 38097 51063 38120 52040
rect 35090 51040 38120 51063
rect 38280 51063 38303 52040
rect 41287 53040 41310 54047
rect 41470 54047 44500 54070
rect 41470 53040 41493 54047
rect 41287 52040 41493 53040
rect 41287 51063 41310 52040
rect 38280 51040 41310 51063
rect 41470 51063 41493 52040
rect 44477 53040 44500 54047
rect 44660 54047 47690 54070
rect 44660 53040 44683 54047
rect 44477 52040 44683 53040
rect 44477 51063 44500 52040
rect 41470 51040 44500 51063
rect 44660 51063 44683 52040
rect 47667 53040 47690 54047
rect 47850 54047 50880 54070
rect 47850 53040 47873 54047
rect 47667 52040 47873 53040
rect 47667 51063 47690 52040
rect 44660 51040 47690 51063
rect 47850 51063 47873 52040
rect 50857 53040 50880 54047
rect 51040 54047 54070 54070
rect 51040 53040 51063 54047
rect 50857 52040 51063 53040
rect 50857 51063 50880 52040
rect 47850 51040 50880 51063
rect 51040 51063 51063 52040
rect 54047 53040 54070 54047
rect 54230 54047 57260 54070
rect 54230 53040 54253 54047
rect 54047 52040 54253 53040
rect 54047 51063 54070 52040
rect 51040 51040 54070 51063
rect 54230 51063 54253 52040
rect 57237 53040 57260 54047
rect 57420 54047 60450 54070
rect 57420 53040 57443 54047
rect 57237 52040 57443 53040
rect 57237 51063 57260 52040
rect 54230 51040 57260 51063
rect 57420 51063 57443 52040
rect 60427 53040 60450 54047
rect 60610 54047 63640 54070
rect 60610 53040 60633 54047
rect 60427 52040 60633 53040
rect 60427 51063 60450 52040
rect 57420 51040 60450 51063
rect 60610 51063 60633 52040
rect 63617 53040 63640 54047
rect 63800 54047 66830 54070
rect 63800 53040 63823 54047
rect 63617 52040 63823 53040
rect 63617 51063 63640 52040
rect 60610 51040 63640 51063
rect 63800 51063 63823 52040
rect 66807 53040 66830 54047
rect 66990 54047 70020 54070
rect 66990 53040 67013 54047
rect 66807 52040 67013 53040
rect 66807 51063 66830 52040
rect 63800 51040 66830 51063
rect 66990 51063 67013 52040
rect 69997 53040 70020 54047
rect 70180 54047 73210 54070
rect 70180 53040 70203 54047
rect 69997 52040 70203 53040
rect 69997 51063 70020 52040
rect 66990 51040 70020 51063
rect 70180 51063 70203 52040
rect 73187 53040 73210 54047
rect 73370 54047 76400 54070
rect 73370 53040 73393 54047
rect 73187 52040 73393 53040
rect 73187 51063 73210 52040
rect 70180 51040 73210 51063
rect 73370 51063 73393 52040
rect 76377 53040 76400 54047
rect 76560 54047 79590 54070
rect 76560 53040 76583 54047
rect 76377 52040 76583 53040
rect 76377 51063 76400 52040
rect 73370 51040 76400 51063
rect 76560 51063 76583 52040
rect 79567 53040 79590 54047
rect 79750 54047 82780 54070
rect 79750 53040 79773 54047
rect 79567 52040 79773 53040
rect 79567 51063 79590 52040
rect 76560 51040 79590 51063
rect 79750 51063 79773 52040
rect 82757 53040 82780 54047
rect 82940 54047 85970 54070
rect 82940 53040 82963 54047
rect 82757 52040 82963 53040
rect 82757 51063 82780 52040
rect 79750 51040 82780 51063
rect 82940 51063 82963 52040
rect 85947 53040 85970 54047
rect 86130 54047 89160 54070
rect 86130 53040 86153 54047
rect 85947 52040 86153 53040
rect 85947 51063 85970 52040
rect 82940 51040 85970 51063
rect 86130 51063 86153 52040
rect 89137 53040 89160 54047
rect 89320 54047 92350 54070
rect 89320 53040 89343 54047
rect 89137 52040 89343 53040
rect 89137 51063 89160 52040
rect 86130 51040 89160 51063
rect 89320 51063 89343 52040
rect 92327 53040 92350 54047
rect 92510 54047 95540 54070
rect 92510 53040 92533 54047
rect 92327 52040 92533 53040
rect 92327 51063 92350 52040
rect 89320 51040 92350 51063
rect 92510 51063 92533 52040
rect 95517 53040 95540 54047
rect 95700 54047 98730 54070
rect 95700 53040 95723 54047
rect 95517 52040 95723 53040
rect 95517 51063 95540 52040
rect 92510 51040 95540 51063
rect 95700 51063 95723 52040
rect 98707 53040 98730 54047
rect 98890 54047 101920 54070
rect 98890 53040 98913 54047
rect 98707 52040 98913 53040
rect 98707 51063 98730 52040
rect 95700 51040 98730 51063
rect 98890 51063 98913 52040
rect 101897 53040 101920 54047
rect 102080 54047 105110 54070
rect 102080 53040 102103 54047
rect 101897 52040 102103 53040
rect 101897 51063 101920 52040
rect 98890 51040 101920 51063
rect 102080 51063 102103 52040
rect 105087 53040 105110 54047
rect 105270 54047 108300 54070
rect 105270 53040 105293 54047
rect 105087 52040 105293 53040
rect 105087 51063 105110 52040
rect 102080 51040 105110 51063
rect 105270 51063 105293 52040
rect 108277 53040 108300 54047
rect 108460 54047 111490 54070
rect 108460 53040 108483 54047
rect 108277 52040 108483 53040
rect 108277 51063 108300 52040
rect 105270 51040 108300 51063
rect 108460 51063 108483 52040
rect 111467 53040 111490 54047
rect 111650 54047 114680 54070
rect 111650 53040 111673 54047
rect 111467 52040 111673 53040
rect 111467 51063 111490 52040
rect 108460 51040 111490 51063
rect 111650 51063 111673 52040
rect 114657 53040 114680 54047
rect 114840 54047 117870 54070
rect 114840 53040 114863 54047
rect 114657 52040 114863 53040
rect 114657 51063 114680 52040
rect 111650 51040 114680 51063
rect 114840 51063 114863 52040
rect 117847 53040 117870 54047
rect 118030 54047 121060 54070
rect 118030 53040 118053 54047
rect 117847 52040 118053 53040
rect 117847 51063 117870 52040
rect 114840 51040 117870 51063
rect 118030 51063 118053 52040
rect 121037 53040 121060 54047
rect 121220 54047 124250 54070
rect 121220 53040 121243 54047
rect 121037 52040 121243 53040
rect 121037 51063 121060 52040
rect 118030 51040 121060 51063
rect 121220 51063 121243 52040
rect 124227 53040 124250 54047
rect 124410 54047 127440 54070
rect 124410 53040 124433 54047
rect 124227 52040 124433 53040
rect 124227 51063 124250 52040
rect 121220 51040 124250 51063
rect 124410 51063 124433 52040
rect 127417 53040 127440 54047
rect 127600 54047 130630 54070
rect 127600 53040 127623 54047
rect 127417 52040 127623 53040
rect 127417 51063 127440 52040
rect 124410 51040 127440 51063
rect 127600 51063 127623 52040
rect 130607 53040 130630 54047
rect 130790 54047 133820 54070
rect 130790 53040 130813 54047
rect 130607 52040 130813 53040
rect 130607 51063 130630 52040
rect 127600 51040 130630 51063
rect 130790 51063 130813 52040
rect 133797 53040 133820 54047
rect 133980 54047 137010 54070
rect 133980 53040 134003 54047
rect 133797 52040 134003 53040
rect 133797 51063 133820 52040
rect 130790 51040 133820 51063
rect 133980 51063 134003 52040
rect 136987 53040 137010 54047
rect 136987 52040 137170 53040
rect 136987 51063 137010 52040
rect 133980 51040 137010 51063
rect 1000 50880 2000 51040
rect 4190 50880 5190 51040
rect 7380 50880 8380 51040
rect 10570 50880 11570 51040
rect 13760 50880 14760 51040
rect 16950 50880 17950 51040
rect 20140 50880 21140 51040
rect 23330 50880 24330 51040
rect 26520 50880 27520 51040
rect 29710 50880 30710 51040
rect 32900 50880 33900 51040
rect 36090 50880 37090 51040
rect 39280 50880 40280 51040
rect 42470 50880 43470 51040
rect 45660 50880 46660 51040
rect 48850 50880 49850 51040
rect 52040 50880 53040 51040
rect 55230 50880 56230 51040
rect 58420 50880 59420 51040
rect 61610 50880 62610 51040
rect 64800 50880 65800 51040
rect 67990 50880 68990 51040
rect 71180 50880 72180 51040
rect 74370 50880 75370 51040
rect 77560 50880 78560 51040
rect 80750 50880 81750 51040
rect 83940 50880 84940 51040
rect 87130 50880 88130 51040
rect 90320 50880 91320 51040
rect 93510 50880 94510 51040
rect 96700 50880 97700 51040
rect 99890 50880 100890 51040
rect 103080 50880 104080 51040
rect 106270 50880 107270 51040
rect 109460 50880 110460 51040
rect 112650 50880 113650 51040
rect 115840 50880 116840 51040
rect 119030 50880 120030 51040
rect 122220 50880 123220 51040
rect 125410 50880 126410 51040
rect 128600 50880 129600 51040
rect 131790 50880 132790 51040
rect 134980 50880 135980 51040
rect 0 50857 3030 50880
rect 0 47873 23 50857
rect 3007 49850 3030 50857
rect 3190 50857 6220 50880
rect 3190 49850 3213 50857
rect 3007 48850 3213 49850
rect 3007 47873 3030 48850
rect 0 47850 3030 47873
rect 3190 47873 3213 48850
rect 6197 49850 6220 50857
rect 6380 50857 9410 50880
rect 6380 49850 6403 50857
rect 6197 48850 6403 49850
rect 6197 47873 6220 48850
rect 3190 47850 6220 47873
rect 6380 47873 6403 48850
rect 9387 49850 9410 50857
rect 9570 50857 12600 50880
rect 9570 49850 9593 50857
rect 9387 48850 9593 49850
rect 9387 47873 9410 48850
rect 6380 47850 9410 47873
rect 9570 47873 9593 48850
rect 12577 49850 12600 50857
rect 12760 50857 15790 50880
rect 12760 49850 12783 50857
rect 12577 48850 12783 49850
rect 12577 47873 12600 48850
rect 9570 47850 12600 47873
rect 12760 47873 12783 48850
rect 15767 49850 15790 50857
rect 15950 50857 18980 50880
rect 15950 49850 15973 50857
rect 15767 48850 15973 49850
rect 15767 47873 15790 48850
rect 12760 47850 15790 47873
rect 15950 47873 15973 48850
rect 18957 49850 18980 50857
rect 19140 50857 22170 50880
rect 19140 49850 19163 50857
rect 18957 48850 19163 49850
rect 18957 47873 18980 48850
rect 15950 47850 18980 47873
rect 19140 47873 19163 48850
rect 22147 49850 22170 50857
rect 22330 50857 25360 50880
rect 22330 49850 22353 50857
rect 22147 48850 22353 49850
rect 22147 47873 22170 48850
rect 19140 47850 22170 47873
rect 22330 47873 22353 48850
rect 25337 49850 25360 50857
rect 25520 50857 28550 50880
rect 25520 49850 25543 50857
rect 25337 48850 25543 49850
rect 25337 47873 25360 48850
rect 22330 47850 25360 47873
rect 25520 47873 25543 48850
rect 28527 49850 28550 50857
rect 28710 50857 31740 50880
rect 28710 49850 28733 50857
rect 28527 48850 28733 49850
rect 28527 47873 28550 48850
rect 25520 47850 28550 47873
rect 28710 47873 28733 48850
rect 31717 49850 31740 50857
rect 31900 50857 34930 50880
rect 31900 49850 31923 50857
rect 31717 48850 31923 49850
rect 31717 47873 31740 48850
rect 28710 47850 31740 47873
rect 31900 47873 31923 48850
rect 34907 49850 34930 50857
rect 35090 50857 38120 50880
rect 35090 49850 35113 50857
rect 34907 48850 35113 49850
rect 34907 47873 34930 48850
rect 31900 47850 34930 47873
rect 35090 47873 35113 48850
rect 38097 49850 38120 50857
rect 38280 50857 41310 50880
rect 38280 49850 38303 50857
rect 38097 48850 38303 49850
rect 38097 47873 38120 48850
rect 35090 47850 38120 47873
rect 38280 47873 38303 48850
rect 41287 49850 41310 50857
rect 41470 50857 44500 50880
rect 41470 49850 41493 50857
rect 41287 48850 41493 49850
rect 41287 47873 41310 48850
rect 38280 47850 41310 47873
rect 41470 47873 41493 48850
rect 44477 49850 44500 50857
rect 44660 50857 47690 50880
rect 44660 49850 44683 50857
rect 44477 48850 44683 49850
rect 44477 47873 44500 48850
rect 41470 47850 44500 47873
rect 44660 47873 44683 48850
rect 47667 49850 47690 50857
rect 47850 50857 50880 50880
rect 47850 49850 47873 50857
rect 47667 48850 47873 49850
rect 47667 47873 47690 48850
rect 44660 47850 47690 47873
rect 47850 47873 47873 48850
rect 50857 49850 50880 50857
rect 51040 50857 54070 50880
rect 51040 49850 51063 50857
rect 50857 48850 51063 49850
rect 50857 47873 50880 48850
rect 47850 47850 50880 47873
rect 51040 47873 51063 48850
rect 54047 49850 54070 50857
rect 54230 50857 57260 50880
rect 54230 49850 54253 50857
rect 54047 48850 54253 49850
rect 54047 47873 54070 48850
rect 51040 47850 54070 47873
rect 54230 47873 54253 48850
rect 57237 49850 57260 50857
rect 57420 50857 60450 50880
rect 57420 49850 57443 50857
rect 57237 48850 57443 49850
rect 57237 47873 57260 48850
rect 54230 47850 57260 47873
rect 57420 47873 57443 48850
rect 60427 49850 60450 50857
rect 60610 50857 63640 50880
rect 60610 49850 60633 50857
rect 60427 48850 60633 49850
rect 60427 47873 60450 48850
rect 57420 47850 60450 47873
rect 60610 47873 60633 48850
rect 63617 49850 63640 50857
rect 63800 50857 66830 50880
rect 63800 49850 63823 50857
rect 63617 48850 63823 49850
rect 63617 47873 63640 48850
rect 60610 47850 63640 47873
rect 63800 47873 63823 48850
rect 66807 49850 66830 50857
rect 66990 50857 70020 50880
rect 66990 49850 67013 50857
rect 66807 48850 67013 49850
rect 66807 47873 66830 48850
rect 63800 47850 66830 47873
rect 66990 47873 67013 48850
rect 69997 49850 70020 50857
rect 70180 50857 73210 50880
rect 70180 49850 70203 50857
rect 69997 48850 70203 49850
rect 69997 47873 70020 48850
rect 66990 47850 70020 47873
rect 70180 47873 70203 48850
rect 73187 49850 73210 50857
rect 73370 50857 76400 50880
rect 73370 49850 73393 50857
rect 73187 48850 73393 49850
rect 73187 47873 73210 48850
rect 70180 47850 73210 47873
rect 73370 47873 73393 48850
rect 76377 49850 76400 50857
rect 76560 50857 79590 50880
rect 76560 49850 76583 50857
rect 76377 48850 76583 49850
rect 76377 47873 76400 48850
rect 73370 47850 76400 47873
rect 76560 47873 76583 48850
rect 79567 49850 79590 50857
rect 79750 50857 82780 50880
rect 79750 49850 79773 50857
rect 79567 48850 79773 49850
rect 79567 47873 79590 48850
rect 76560 47850 79590 47873
rect 79750 47873 79773 48850
rect 82757 49850 82780 50857
rect 82940 50857 85970 50880
rect 82940 49850 82963 50857
rect 82757 48850 82963 49850
rect 82757 47873 82780 48850
rect 79750 47850 82780 47873
rect 82940 47873 82963 48850
rect 85947 49850 85970 50857
rect 86130 50857 89160 50880
rect 86130 49850 86153 50857
rect 85947 48850 86153 49850
rect 85947 47873 85970 48850
rect 82940 47850 85970 47873
rect 86130 47873 86153 48850
rect 89137 49850 89160 50857
rect 89320 50857 92350 50880
rect 89320 49850 89343 50857
rect 89137 48850 89343 49850
rect 89137 47873 89160 48850
rect 86130 47850 89160 47873
rect 89320 47873 89343 48850
rect 92327 49850 92350 50857
rect 92510 50857 95540 50880
rect 92510 49850 92533 50857
rect 92327 48850 92533 49850
rect 92327 47873 92350 48850
rect 89320 47850 92350 47873
rect 92510 47873 92533 48850
rect 95517 49850 95540 50857
rect 95700 50857 98730 50880
rect 95700 49850 95723 50857
rect 95517 48850 95723 49850
rect 95517 47873 95540 48850
rect 92510 47850 95540 47873
rect 95700 47873 95723 48850
rect 98707 49850 98730 50857
rect 98890 50857 101920 50880
rect 98890 49850 98913 50857
rect 98707 48850 98913 49850
rect 98707 47873 98730 48850
rect 95700 47850 98730 47873
rect 98890 47873 98913 48850
rect 101897 49850 101920 50857
rect 102080 50857 105110 50880
rect 102080 49850 102103 50857
rect 101897 48850 102103 49850
rect 101897 47873 101920 48850
rect 98890 47850 101920 47873
rect 102080 47873 102103 48850
rect 105087 49850 105110 50857
rect 105270 50857 108300 50880
rect 105270 49850 105293 50857
rect 105087 48850 105293 49850
rect 105087 47873 105110 48850
rect 102080 47850 105110 47873
rect 105270 47873 105293 48850
rect 108277 49850 108300 50857
rect 108460 50857 111490 50880
rect 108460 49850 108483 50857
rect 108277 48850 108483 49850
rect 108277 47873 108300 48850
rect 105270 47850 108300 47873
rect 108460 47873 108483 48850
rect 111467 49850 111490 50857
rect 111650 50857 114680 50880
rect 111650 49850 111673 50857
rect 111467 48850 111673 49850
rect 111467 47873 111490 48850
rect 108460 47850 111490 47873
rect 111650 47873 111673 48850
rect 114657 49850 114680 50857
rect 114840 50857 117870 50880
rect 114840 49850 114863 50857
rect 114657 48850 114863 49850
rect 114657 47873 114680 48850
rect 111650 47850 114680 47873
rect 114840 47873 114863 48850
rect 117847 49850 117870 50857
rect 118030 50857 121060 50880
rect 118030 49850 118053 50857
rect 117847 48850 118053 49850
rect 117847 47873 117870 48850
rect 114840 47850 117870 47873
rect 118030 47873 118053 48850
rect 121037 49850 121060 50857
rect 121220 50857 124250 50880
rect 121220 49850 121243 50857
rect 121037 48850 121243 49850
rect 121037 47873 121060 48850
rect 118030 47850 121060 47873
rect 121220 47873 121243 48850
rect 124227 49850 124250 50857
rect 124410 50857 127440 50880
rect 124410 49850 124433 50857
rect 124227 48850 124433 49850
rect 124227 47873 124250 48850
rect 121220 47850 124250 47873
rect 124410 47873 124433 48850
rect 127417 49850 127440 50857
rect 127600 50857 130630 50880
rect 127600 49850 127623 50857
rect 127417 48850 127623 49850
rect 127417 47873 127440 48850
rect 124410 47850 127440 47873
rect 127600 47873 127623 48850
rect 130607 49850 130630 50857
rect 130790 50857 133820 50880
rect 130790 49850 130813 50857
rect 130607 48850 130813 49850
rect 130607 47873 130630 48850
rect 127600 47850 130630 47873
rect 130790 47873 130813 48850
rect 133797 49850 133820 50857
rect 133980 50857 137010 50880
rect 133980 49850 134003 50857
rect 133797 48850 134003 49850
rect 133797 47873 133820 48850
rect 130790 47850 133820 47873
rect 133980 47873 134003 48850
rect 136987 49850 137010 50857
rect 136987 48850 137170 49850
rect 136987 47873 137010 48850
rect 133980 47850 137010 47873
rect 1000 47690 2000 47850
rect 4190 47690 5190 47850
rect 7380 47690 8380 47850
rect 10570 47690 11570 47850
rect 13760 47690 14760 47850
rect 16950 47690 17950 47850
rect 20140 47690 21140 47850
rect 23330 47690 24330 47850
rect 26520 47690 27520 47850
rect 29710 47690 30710 47850
rect 32900 47690 33900 47850
rect 36090 47690 37090 47850
rect 39280 47690 40280 47850
rect 42470 47690 43470 47850
rect 45660 47690 46660 47850
rect 48850 47690 49850 47850
rect 52040 47690 53040 47850
rect 55230 47690 56230 47850
rect 58420 47690 59420 47850
rect 61610 47690 62610 47850
rect 64800 47690 65800 47850
rect 67990 47690 68990 47850
rect 71180 47690 72180 47850
rect 74370 47690 75370 47850
rect 77560 47690 78560 47850
rect 80750 47690 81750 47850
rect 83940 47690 84940 47850
rect 87130 47690 88130 47850
rect 90320 47690 91320 47850
rect 93510 47690 94510 47850
rect 96700 47690 97700 47850
rect 99890 47690 100890 47850
rect 103080 47690 104080 47850
rect 106270 47690 107270 47850
rect 109460 47690 110460 47850
rect 112650 47690 113650 47850
rect 115840 47690 116840 47850
rect 119030 47690 120030 47850
rect 122220 47690 123220 47850
rect 125410 47690 126410 47850
rect 128600 47690 129600 47850
rect 131790 47690 132790 47850
rect 134980 47690 135980 47850
rect 0 47667 3030 47690
rect 0 44683 23 47667
rect 3007 46660 3030 47667
rect 3190 47667 6220 47690
rect 3190 46660 3213 47667
rect 3007 45660 3213 46660
rect 3007 44683 3030 45660
rect 0 44660 3030 44683
rect 3190 44683 3213 45660
rect 6197 46660 6220 47667
rect 6380 47667 9410 47690
rect 6380 46660 6403 47667
rect 6197 45660 6403 46660
rect 6197 44683 6220 45660
rect 3190 44660 6220 44683
rect 6380 44683 6403 45660
rect 9387 46660 9410 47667
rect 9570 47667 12600 47690
rect 9570 46660 9593 47667
rect 9387 45660 9593 46660
rect 9387 44683 9410 45660
rect 6380 44660 9410 44683
rect 9570 44683 9593 45660
rect 12577 46660 12600 47667
rect 12760 47667 15790 47690
rect 12760 46660 12783 47667
rect 12577 45660 12783 46660
rect 12577 44683 12600 45660
rect 9570 44660 12600 44683
rect 12760 44683 12783 45660
rect 15767 46660 15790 47667
rect 15950 47667 18980 47690
rect 15950 46660 15973 47667
rect 15767 45660 15973 46660
rect 15767 44683 15790 45660
rect 12760 44660 15790 44683
rect 15950 44683 15973 45660
rect 18957 46660 18980 47667
rect 19140 47667 22170 47690
rect 19140 46660 19163 47667
rect 18957 45660 19163 46660
rect 18957 44683 18980 45660
rect 15950 44660 18980 44683
rect 19140 44683 19163 45660
rect 22147 46660 22170 47667
rect 22330 47667 25360 47690
rect 22330 46660 22353 47667
rect 22147 45660 22353 46660
rect 22147 44683 22170 45660
rect 19140 44660 22170 44683
rect 22330 44683 22353 45660
rect 25337 46660 25360 47667
rect 25520 47667 28550 47690
rect 25520 46660 25543 47667
rect 25337 45660 25543 46660
rect 25337 44683 25360 45660
rect 22330 44660 25360 44683
rect 25520 44683 25543 45660
rect 28527 46660 28550 47667
rect 28710 47667 31740 47690
rect 28710 46660 28733 47667
rect 28527 45660 28733 46660
rect 28527 44683 28550 45660
rect 25520 44660 28550 44683
rect 28710 44683 28733 45660
rect 31717 46660 31740 47667
rect 31900 47667 34930 47690
rect 31900 46660 31923 47667
rect 31717 45660 31923 46660
rect 31717 44683 31740 45660
rect 28710 44660 31740 44683
rect 31900 44683 31923 45660
rect 34907 46660 34930 47667
rect 35090 47667 38120 47690
rect 35090 46660 35113 47667
rect 34907 45660 35113 46660
rect 34907 44683 34930 45660
rect 31900 44660 34930 44683
rect 35090 44683 35113 45660
rect 38097 46660 38120 47667
rect 38280 47667 41310 47690
rect 38280 46660 38303 47667
rect 38097 45660 38303 46660
rect 38097 44683 38120 45660
rect 35090 44660 38120 44683
rect 38280 44683 38303 45660
rect 41287 46660 41310 47667
rect 41470 47667 44500 47690
rect 41470 46660 41493 47667
rect 41287 45660 41493 46660
rect 41287 44683 41310 45660
rect 38280 44660 41310 44683
rect 41470 44683 41493 45660
rect 44477 46660 44500 47667
rect 44660 47667 47690 47690
rect 44660 46660 44683 47667
rect 44477 45660 44683 46660
rect 44477 44683 44500 45660
rect 41470 44660 44500 44683
rect 44660 44683 44683 45660
rect 47667 46660 47690 47667
rect 47850 47667 50880 47690
rect 47850 46660 47873 47667
rect 47667 45660 47873 46660
rect 47667 44683 47690 45660
rect 44660 44660 47690 44683
rect 47850 44683 47873 45660
rect 50857 46660 50880 47667
rect 51040 47667 54070 47690
rect 51040 46660 51063 47667
rect 50857 45660 51063 46660
rect 50857 44683 50880 45660
rect 47850 44660 50880 44683
rect 51040 44683 51063 45660
rect 54047 46660 54070 47667
rect 54230 47667 57260 47690
rect 54230 46660 54253 47667
rect 54047 45660 54253 46660
rect 54047 44683 54070 45660
rect 51040 44660 54070 44683
rect 54230 44683 54253 45660
rect 57237 46660 57260 47667
rect 57420 47667 60450 47690
rect 57420 46660 57443 47667
rect 57237 45660 57443 46660
rect 57237 44683 57260 45660
rect 54230 44660 57260 44683
rect 57420 44683 57443 45660
rect 60427 46660 60450 47667
rect 60610 47667 63640 47690
rect 60610 46660 60633 47667
rect 60427 45660 60633 46660
rect 60427 44683 60450 45660
rect 57420 44660 60450 44683
rect 60610 44683 60633 45660
rect 63617 46660 63640 47667
rect 63800 47667 66830 47690
rect 63800 46660 63823 47667
rect 63617 45660 63823 46660
rect 63617 44683 63640 45660
rect 60610 44660 63640 44683
rect 63800 44683 63823 45660
rect 66807 46660 66830 47667
rect 66990 47667 70020 47690
rect 66990 46660 67013 47667
rect 66807 45660 67013 46660
rect 66807 44683 66830 45660
rect 63800 44660 66830 44683
rect 66990 44683 67013 45660
rect 69997 46660 70020 47667
rect 70180 47667 73210 47690
rect 70180 46660 70203 47667
rect 69997 45660 70203 46660
rect 69997 44683 70020 45660
rect 66990 44660 70020 44683
rect 70180 44683 70203 45660
rect 73187 46660 73210 47667
rect 73370 47667 76400 47690
rect 73370 46660 73393 47667
rect 73187 45660 73393 46660
rect 73187 44683 73210 45660
rect 70180 44660 73210 44683
rect 73370 44683 73393 45660
rect 76377 46660 76400 47667
rect 76560 47667 79590 47690
rect 76560 46660 76583 47667
rect 76377 45660 76583 46660
rect 76377 44683 76400 45660
rect 73370 44660 76400 44683
rect 76560 44683 76583 45660
rect 79567 46660 79590 47667
rect 79750 47667 82780 47690
rect 79750 46660 79773 47667
rect 79567 45660 79773 46660
rect 79567 44683 79590 45660
rect 76560 44660 79590 44683
rect 79750 44683 79773 45660
rect 82757 46660 82780 47667
rect 82940 47667 85970 47690
rect 82940 46660 82963 47667
rect 82757 45660 82963 46660
rect 82757 44683 82780 45660
rect 79750 44660 82780 44683
rect 82940 44683 82963 45660
rect 85947 46660 85970 47667
rect 86130 47667 89160 47690
rect 86130 46660 86153 47667
rect 85947 45660 86153 46660
rect 85947 44683 85970 45660
rect 82940 44660 85970 44683
rect 86130 44683 86153 45660
rect 89137 46660 89160 47667
rect 89320 47667 92350 47690
rect 89320 46660 89343 47667
rect 89137 45660 89343 46660
rect 89137 44683 89160 45660
rect 86130 44660 89160 44683
rect 89320 44683 89343 45660
rect 92327 46660 92350 47667
rect 92510 47667 95540 47690
rect 92510 46660 92533 47667
rect 92327 45660 92533 46660
rect 92327 44683 92350 45660
rect 89320 44660 92350 44683
rect 92510 44683 92533 45660
rect 95517 46660 95540 47667
rect 95700 47667 98730 47690
rect 95700 46660 95723 47667
rect 95517 45660 95723 46660
rect 95517 44683 95540 45660
rect 92510 44660 95540 44683
rect 95700 44683 95723 45660
rect 98707 46660 98730 47667
rect 98890 47667 101920 47690
rect 98890 46660 98913 47667
rect 98707 45660 98913 46660
rect 98707 44683 98730 45660
rect 95700 44660 98730 44683
rect 98890 44683 98913 45660
rect 101897 46660 101920 47667
rect 102080 47667 105110 47690
rect 102080 46660 102103 47667
rect 101897 45660 102103 46660
rect 101897 44683 101920 45660
rect 98890 44660 101920 44683
rect 102080 44683 102103 45660
rect 105087 46660 105110 47667
rect 105270 47667 108300 47690
rect 105270 46660 105293 47667
rect 105087 45660 105293 46660
rect 105087 44683 105110 45660
rect 102080 44660 105110 44683
rect 105270 44683 105293 45660
rect 108277 46660 108300 47667
rect 108460 47667 111490 47690
rect 108460 46660 108483 47667
rect 108277 45660 108483 46660
rect 108277 44683 108300 45660
rect 105270 44660 108300 44683
rect 108460 44683 108483 45660
rect 111467 46660 111490 47667
rect 111650 47667 114680 47690
rect 111650 46660 111673 47667
rect 111467 45660 111673 46660
rect 111467 44683 111490 45660
rect 108460 44660 111490 44683
rect 111650 44683 111673 45660
rect 114657 46660 114680 47667
rect 114840 47667 117870 47690
rect 114840 46660 114863 47667
rect 114657 45660 114863 46660
rect 114657 44683 114680 45660
rect 111650 44660 114680 44683
rect 114840 44683 114863 45660
rect 117847 46660 117870 47667
rect 118030 47667 121060 47690
rect 118030 46660 118053 47667
rect 117847 45660 118053 46660
rect 117847 44683 117870 45660
rect 114840 44660 117870 44683
rect 118030 44683 118053 45660
rect 121037 46660 121060 47667
rect 121220 47667 124250 47690
rect 121220 46660 121243 47667
rect 121037 45660 121243 46660
rect 121037 44683 121060 45660
rect 118030 44660 121060 44683
rect 121220 44683 121243 45660
rect 124227 46660 124250 47667
rect 124410 47667 127440 47690
rect 124410 46660 124433 47667
rect 124227 45660 124433 46660
rect 124227 44683 124250 45660
rect 121220 44660 124250 44683
rect 124410 44683 124433 45660
rect 127417 46660 127440 47667
rect 127600 47667 130630 47690
rect 127600 46660 127623 47667
rect 127417 45660 127623 46660
rect 127417 44683 127440 45660
rect 124410 44660 127440 44683
rect 127600 44683 127623 45660
rect 130607 46660 130630 47667
rect 130790 47667 133820 47690
rect 130790 46660 130813 47667
rect 130607 45660 130813 46660
rect 130607 44683 130630 45660
rect 127600 44660 130630 44683
rect 130790 44683 130813 45660
rect 133797 46660 133820 47667
rect 133980 47667 137010 47690
rect 133980 46660 134003 47667
rect 133797 45660 134003 46660
rect 133797 44683 133820 45660
rect 130790 44660 133820 44683
rect 133980 44683 134003 45660
rect 136987 46660 137010 47667
rect 136987 45660 137170 46660
rect 136987 44683 137010 45660
rect 133980 44660 137010 44683
rect 1000 44500 2000 44660
rect 4190 44500 5190 44660
rect 7380 44500 8380 44660
rect 10570 44500 11570 44660
rect 13760 44500 14760 44660
rect 16950 44500 17950 44660
rect 20140 44500 21140 44660
rect 23330 44500 24330 44660
rect 26520 44500 27520 44660
rect 29710 44500 30710 44660
rect 32900 44500 33900 44660
rect 36090 44500 37090 44660
rect 39280 44500 40280 44660
rect 42470 44500 43470 44660
rect 45660 44500 46660 44660
rect 48850 44500 49850 44660
rect 52040 44500 53040 44660
rect 55230 44500 56230 44660
rect 58420 44500 59420 44660
rect 61610 44500 62610 44660
rect 64800 44500 65800 44660
rect 67990 44500 68990 44660
rect 71180 44500 72180 44660
rect 74370 44500 75370 44660
rect 77560 44500 78560 44660
rect 80750 44500 81750 44660
rect 83940 44500 84940 44660
rect 87130 44500 88130 44660
rect 90320 44500 91320 44660
rect 93510 44500 94510 44660
rect 96700 44500 97700 44660
rect 99890 44500 100890 44660
rect 103080 44500 104080 44660
rect 106270 44500 107270 44660
rect 109460 44500 110460 44660
rect 112650 44500 113650 44660
rect 115840 44500 116840 44660
rect 119030 44500 120030 44660
rect 122220 44500 123220 44660
rect 125410 44500 126410 44660
rect 128600 44500 129600 44660
rect 131790 44500 132790 44660
rect 134980 44500 135980 44660
rect 0 44477 3030 44500
rect 0 41493 23 44477
rect 3007 43470 3030 44477
rect 3190 44477 6220 44500
rect 3190 43470 3213 44477
rect 3007 42470 3213 43470
rect 3007 41493 3030 42470
rect 0 41470 3030 41493
rect 3190 41493 3213 42470
rect 6197 43470 6220 44477
rect 6380 44477 9410 44500
rect 6380 43470 6403 44477
rect 6197 42470 6403 43470
rect 6197 41493 6220 42470
rect 3190 41470 6220 41493
rect 6380 41493 6403 42470
rect 9387 43470 9410 44477
rect 9570 44477 12600 44500
rect 9570 43470 9593 44477
rect 9387 42470 9593 43470
rect 9387 41493 9410 42470
rect 6380 41470 9410 41493
rect 9570 41493 9593 42470
rect 12577 43470 12600 44477
rect 12760 44477 15790 44500
rect 12760 43470 12783 44477
rect 12577 42470 12783 43470
rect 12577 41493 12600 42470
rect 9570 41470 12600 41493
rect 12760 41493 12783 42470
rect 15767 43470 15790 44477
rect 15950 44477 18980 44500
rect 15950 43470 15973 44477
rect 15767 42470 15973 43470
rect 15767 41493 15790 42470
rect 12760 41470 15790 41493
rect 15950 41493 15973 42470
rect 18957 43470 18980 44477
rect 19140 44477 22170 44500
rect 19140 43470 19163 44477
rect 18957 42470 19163 43470
rect 18957 41493 18980 42470
rect 15950 41470 18980 41493
rect 19140 41493 19163 42470
rect 22147 43470 22170 44477
rect 22330 44477 25360 44500
rect 22330 43470 22353 44477
rect 22147 42470 22353 43470
rect 22147 41493 22170 42470
rect 19140 41470 22170 41493
rect 22330 41493 22353 42470
rect 25337 43470 25360 44477
rect 25520 44477 28550 44500
rect 25520 43470 25543 44477
rect 25337 42470 25543 43470
rect 25337 41493 25360 42470
rect 22330 41470 25360 41493
rect 25520 41493 25543 42470
rect 28527 43470 28550 44477
rect 28710 44477 31740 44500
rect 28710 43470 28733 44477
rect 28527 42470 28733 43470
rect 28527 41493 28550 42470
rect 25520 41470 28550 41493
rect 28710 41493 28733 42470
rect 31717 43470 31740 44477
rect 31900 44477 34930 44500
rect 31900 43470 31923 44477
rect 31717 42470 31923 43470
rect 31717 41493 31740 42470
rect 28710 41470 31740 41493
rect 31900 41493 31923 42470
rect 34907 43470 34930 44477
rect 35090 44477 38120 44500
rect 35090 43470 35113 44477
rect 34907 42470 35113 43470
rect 34907 41493 34930 42470
rect 31900 41470 34930 41493
rect 35090 41493 35113 42470
rect 38097 43470 38120 44477
rect 38280 44477 41310 44500
rect 38280 43470 38303 44477
rect 38097 42470 38303 43470
rect 38097 41493 38120 42470
rect 35090 41470 38120 41493
rect 38280 41493 38303 42470
rect 41287 43470 41310 44477
rect 41470 44477 44500 44500
rect 41470 43470 41493 44477
rect 41287 42470 41493 43470
rect 41287 41493 41310 42470
rect 38280 41470 41310 41493
rect 41470 41493 41493 42470
rect 44477 43470 44500 44477
rect 44660 44477 47690 44500
rect 44660 43470 44683 44477
rect 44477 42470 44683 43470
rect 44477 41493 44500 42470
rect 41470 41470 44500 41493
rect 44660 41493 44683 42470
rect 47667 43470 47690 44477
rect 47850 44477 50880 44500
rect 47850 43470 47873 44477
rect 47667 42470 47873 43470
rect 47667 41493 47690 42470
rect 44660 41470 47690 41493
rect 47850 41493 47873 42470
rect 50857 43470 50880 44477
rect 51040 44477 54070 44500
rect 51040 43470 51063 44477
rect 50857 42470 51063 43470
rect 50857 41493 50880 42470
rect 47850 41470 50880 41493
rect 51040 41493 51063 42470
rect 54047 43470 54070 44477
rect 54230 44477 57260 44500
rect 54230 43470 54253 44477
rect 54047 42470 54253 43470
rect 54047 41493 54070 42470
rect 51040 41470 54070 41493
rect 54230 41493 54253 42470
rect 57237 43470 57260 44477
rect 57420 44477 60450 44500
rect 57420 43470 57443 44477
rect 57237 42470 57443 43470
rect 57237 41493 57260 42470
rect 54230 41470 57260 41493
rect 57420 41493 57443 42470
rect 60427 43470 60450 44477
rect 60610 44477 63640 44500
rect 60610 43470 60633 44477
rect 60427 42470 60633 43470
rect 60427 41493 60450 42470
rect 57420 41470 60450 41493
rect 60610 41493 60633 42470
rect 63617 43470 63640 44477
rect 63800 44477 66830 44500
rect 63800 43470 63823 44477
rect 63617 42470 63823 43470
rect 63617 41493 63640 42470
rect 60610 41470 63640 41493
rect 63800 41493 63823 42470
rect 66807 43470 66830 44477
rect 66990 44477 70020 44500
rect 66990 43470 67013 44477
rect 66807 42470 67013 43470
rect 66807 41493 66830 42470
rect 63800 41470 66830 41493
rect 66990 41493 67013 42470
rect 69997 43470 70020 44477
rect 70180 44477 73210 44500
rect 70180 43470 70203 44477
rect 69997 42470 70203 43470
rect 69997 41493 70020 42470
rect 66990 41470 70020 41493
rect 70180 41493 70203 42470
rect 73187 43470 73210 44477
rect 73370 44477 76400 44500
rect 73370 43470 73393 44477
rect 73187 42470 73393 43470
rect 73187 41493 73210 42470
rect 70180 41470 73210 41493
rect 73370 41493 73393 42470
rect 76377 43470 76400 44477
rect 76560 44477 79590 44500
rect 76560 43470 76583 44477
rect 76377 42470 76583 43470
rect 76377 41493 76400 42470
rect 73370 41470 76400 41493
rect 76560 41493 76583 42470
rect 79567 43470 79590 44477
rect 79750 44477 82780 44500
rect 79750 43470 79773 44477
rect 79567 42470 79773 43470
rect 79567 41493 79590 42470
rect 76560 41470 79590 41493
rect 79750 41493 79773 42470
rect 82757 43470 82780 44477
rect 82940 44477 85970 44500
rect 82940 43470 82963 44477
rect 82757 42470 82963 43470
rect 82757 41493 82780 42470
rect 79750 41470 82780 41493
rect 82940 41493 82963 42470
rect 85947 43470 85970 44477
rect 86130 44477 89160 44500
rect 86130 43470 86153 44477
rect 85947 42470 86153 43470
rect 85947 41493 85970 42470
rect 82940 41470 85970 41493
rect 86130 41493 86153 42470
rect 89137 43470 89160 44477
rect 89320 44477 92350 44500
rect 89320 43470 89343 44477
rect 89137 42470 89343 43470
rect 89137 41493 89160 42470
rect 86130 41470 89160 41493
rect 89320 41493 89343 42470
rect 92327 43470 92350 44477
rect 92510 44477 95540 44500
rect 92510 43470 92533 44477
rect 92327 42470 92533 43470
rect 92327 41493 92350 42470
rect 89320 41470 92350 41493
rect 92510 41493 92533 42470
rect 95517 43470 95540 44477
rect 95700 44477 98730 44500
rect 95700 43470 95723 44477
rect 95517 42470 95723 43470
rect 95517 41493 95540 42470
rect 92510 41470 95540 41493
rect 95700 41493 95723 42470
rect 98707 43470 98730 44477
rect 98890 44477 101920 44500
rect 98890 43470 98913 44477
rect 98707 42470 98913 43470
rect 98707 41493 98730 42470
rect 95700 41470 98730 41493
rect 98890 41493 98913 42470
rect 101897 43470 101920 44477
rect 102080 44477 105110 44500
rect 102080 43470 102103 44477
rect 101897 42470 102103 43470
rect 101897 41493 101920 42470
rect 98890 41470 101920 41493
rect 102080 41493 102103 42470
rect 105087 43470 105110 44477
rect 105270 44477 108300 44500
rect 105270 43470 105293 44477
rect 105087 42470 105293 43470
rect 105087 41493 105110 42470
rect 102080 41470 105110 41493
rect 105270 41493 105293 42470
rect 108277 43470 108300 44477
rect 108460 44477 111490 44500
rect 108460 43470 108483 44477
rect 108277 42470 108483 43470
rect 108277 41493 108300 42470
rect 105270 41470 108300 41493
rect 108460 41493 108483 42470
rect 111467 43470 111490 44477
rect 111650 44477 114680 44500
rect 111650 43470 111673 44477
rect 111467 42470 111673 43470
rect 111467 41493 111490 42470
rect 108460 41470 111490 41493
rect 111650 41493 111673 42470
rect 114657 43470 114680 44477
rect 114840 44477 117870 44500
rect 114840 43470 114863 44477
rect 114657 42470 114863 43470
rect 114657 41493 114680 42470
rect 111650 41470 114680 41493
rect 114840 41493 114863 42470
rect 117847 43470 117870 44477
rect 118030 44477 121060 44500
rect 118030 43470 118053 44477
rect 117847 42470 118053 43470
rect 117847 41493 117870 42470
rect 114840 41470 117870 41493
rect 118030 41493 118053 42470
rect 121037 43470 121060 44477
rect 121220 44477 124250 44500
rect 121220 43470 121243 44477
rect 121037 42470 121243 43470
rect 121037 41493 121060 42470
rect 118030 41470 121060 41493
rect 121220 41493 121243 42470
rect 124227 43470 124250 44477
rect 124410 44477 127440 44500
rect 124410 43470 124433 44477
rect 124227 42470 124433 43470
rect 124227 41493 124250 42470
rect 121220 41470 124250 41493
rect 124410 41493 124433 42470
rect 127417 43470 127440 44477
rect 127600 44477 130630 44500
rect 127600 43470 127623 44477
rect 127417 42470 127623 43470
rect 127417 41493 127440 42470
rect 124410 41470 127440 41493
rect 127600 41493 127623 42470
rect 130607 43470 130630 44477
rect 130790 44477 133820 44500
rect 130790 43470 130813 44477
rect 130607 42470 130813 43470
rect 130607 41493 130630 42470
rect 127600 41470 130630 41493
rect 130790 41493 130813 42470
rect 133797 43470 133820 44477
rect 133980 44477 137010 44500
rect 133980 43470 134003 44477
rect 133797 42470 134003 43470
rect 133797 41493 133820 42470
rect 130790 41470 133820 41493
rect 133980 41493 134003 42470
rect 136987 43470 137010 44477
rect 136987 42470 137170 43470
rect 136987 41493 137010 42470
rect 133980 41470 137010 41493
rect 1000 41310 2000 41470
rect 4190 41310 5190 41470
rect 7380 41310 8380 41470
rect 10570 41310 11570 41470
rect 13760 41310 14760 41470
rect 16950 41310 17950 41470
rect 20140 41310 21140 41470
rect 23330 41310 24330 41470
rect 26520 41310 27520 41470
rect 29710 41310 30710 41470
rect 32900 41310 33900 41470
rect 36090 41310 37090 41470
rect 39280 41310 40280 41470
rect 42470 41310 43470 41470
rect 45660 41310 46660 41470
rect 48850 41310 49850 41470
rect 52040 41310 53040 41470
rect 55230 41310 56230 41470
rect 58420 41310 59420 41470
rect 61610 41310 62610 41470
rect 64800 41310 65800 41470
rect 67990 41310 68990 41470
rect 71180 41310 72180 41470
rect 74370 41310 75370 41470
rect 77560 41310 78560 41470
rect 80750 41310 81750 41470
rect 83940 41310 84940 41470
rect 87130 41310 88130 41470
rect 90320 41310 91320 41470
rect 93510 41310 94510 41470
rect 96700 41310 97700 41470
rect 99890 41310 100890 41470
rect 103080 41310 104080 41470
rect 106270 41310 107270 41470
rect 109460 41310 110460 41470
rect 112650 41310 113650 41470
rect 115840 41310 116840 41470
rect 119030 41310 120030 41470
rect 122220 41310 123220 41470
rect 125410 41310 126410 41470
rect 128600 41310 129600 41470
rect 131790 41310 132790 41470
rect 134980 41310 135980 41470
rect 0 41287 3030 41310
rect 0 38303 23 41287
rect 3007 40280 3030 41287
rect 3190 41287 6220 41310
rect 3190 40280 3213 41287
rect 3007 39280 3213 40280
rect 3007 38303 3030 39280
rect 0 38280 3030 38303
rect 3190 38303 3213 39280
rect 6197 40280 6220 41287
rect 6380 41287 9410 41310
rect 6380 40280 6403 41287
rect 6197 39280 6403 40280
rect 6197 38303 6220 39280
rect 3190 38280 6220 38303
rect 6380 38303 6403 39280
rect 9387 40280 9410 41287
rect 9570 41287 12600 41310
rect 9570 40280 9593 41287
rect 9387 39280 9593 40280
rect 9387 38303 9410 39280
rect 6380 38280 9410 38303
rect 9570 38303 9593 39280
rect 12577 40280 12600 41287
rect 12760 41287 15790 41310
rect 12760 40280 12783 41287
rect 12577 39280 12783 40280
rect 12577 38303 12600 39280
rect 9570 38280 12600 38303
rect 12760 38303 12783 39280
rect 15767 40280 15790 41287
rect 15950 41287 18980 41310
rect 15950 40280 15973 41287
rect 15767 39280 15973 40280
rect 15767 38303 15790 39280
rect 12760 38280 15790 38303
rect 15950 38303 15973 39280
rect 18957 40280 18980 41287
rect 19140 41287 22170 41310
rect 19140 40280 19163 41287
rect 18957 39280 19163 40280
rect 18957 38303 18980 39280
rect 15950 38280 18980 38303
rect 19140 38303 19163 39280
rect 22147 40280 22170 41287
rect 22330 41287 25360 41310
rect 22330 40280 22353 41287
rect 22147 39280 22353 40280
rect 22147 38303 22170 39280
rect 19140 38280 22170 38303
rect 22330 38303 22353 39280
rect 25337 40280 25360 41287
rect 25520 41287 28550 41310
rect 25520 40280 25543 41287
rect 25337 39280 25543 40280
rect 25337 38303 25360 39280
rect 22330 38280 25360 38303
rect 25520 38303 25543 39280
rect 28527 40280 28550 41287
rect 28710 41287 31740 41310
rect 28710 40280 28733 41287
rect 28527 39280 28733 40280
rect 28527 38303 28550 39280
rect 25520 38280 28550 38303
rect 28710 38303 28733 39280
rect 31717 40280 31740 41287
rect 31900 41287 34930 41310
rect 31900 40280 31923 41287
rect 31717 39280 31923 40280
rect 31717 38303 31740 39280
rect 28710 38280 31740 38303
rect 31900 38303 31923 39280
rect 34907 40280 34930 41287
rect 35090 41287 38120 41310
rect 35090 40280 35113 41287
rect 34907 39280 35113 40280
rect 34907 38303 34930 39280
rect 31900 38280 34930 38303
rect 35090 38303 35113 39280
rect 38097 40280 38120 41287
rect 38280 41287 41310 41310
rect 38280 40280 38303 41287
rect 38097 39280 38303 40280
rect 38097 38303 38120 39280
rect 35090 38280 38120 38303
rect 38280 38303 38303 39280
rect 41287 40280 41310 41287
rect 41470 41287 44500 41310
rect 41470 40280 41493 41287
rect 41287 39280 41493 40280
rect 41287 38303 41310 39280
rect 38280 38280 41310 38303
rect 41470 38303 41493 39280
rect 44477 40280 44500 41287
rect 44660 41287 47690 41310
rect 44660 40280 44683 41287
rect 44477 39280 44683 40280
rect 44477 38303 44500 39280
rect 41470 38280 44500 38303
rect 44660 38303 44683 39280
rect 47667 40280 47690 41287
rect 47850 41287 50880 41310
rect 47850 40280 47873 41287
rect 47667 39280 47873 40280
rect 47667 38303 47690 39280
rect 44660 38280 47690 38303
rect 47850 38303 47873 39280
rect 50857 40280 50880 41287
rect 51040 41287 54070 41310
rect 51040 40280 51063 41287
rect 50857 39280 51063 40280
rect 50857 38303 50880 39280
rect 47850 38280 50880 38303
rect 51040 38303 51063 39280
rect 54047 40280 54070 41287
rect 54230 41287 57260 41310
rect 54230 40280 54253 41287
rect 54047 39280 54253 40280
rect 54047 38303 54070 39280
rect 51040 38280 54070 38303
rect 54230 38303 54253 39280
rect 57237 40280 57260 41287
rect 57420 41287 60450 41310
rect 57420 40280 57443 41287
rect 57237 39280 57443 40280
rect 57237 38303 57260 39280
rect 54230 38280 57260 38303
rect 57420 38303 57443 39280
rect 60427 40280 60450 41287
rect 60610 41287 63640 41310
rect 60610 40280 60633 41287
rect 60427 39280 60633 40280
rect 60427 38303 60450 39280
rect 57420 38280 60450 38303
rect 60610 38303 60633 39280
rect 63617 40280 63640 41287
rect 63800 41287 66830 41310
rect 63800 40280 63823 41287
rect 63617 39280 63823 40280
rect 63617 38303 63640 39280
rect 60610 38280 63640 38303
rect 63800 38303 63823 39280
rect 66807 40280 66830 41287
rect 66990 41287 70020 41310
rect 66990 40280 67013 41287
rect 66807 39280 67013 40280
rect 66807 38303 66830 39280
rect 63800 38280 66830 38303
rect 66990 38303 67013 39280
rect 69997 40280 70020 41287
rect 70180 41287 73210 41310
rect 70180 40280 70203 41287
rect 69997 39280 70203 40280
rect 69997 38303 70020 39280
rect 66990 38280 70020 38303
rect 70180 38303 70203 39280
rect 73187 40280 73210 41287
rect 73370 41287 76400 41310
rect 73370 40280 73393 41287
rect 73187 39280 73393 40280
rect 73187 38303 73210 39280
rect 70180 38280 73210 38303
rect 73370 38303 73393 39280
rect 76377 40280 76400 41287
rect 76560 41287 79590 41310
rect 76560 40280 76583 41287
rect 76377 39280 76583 40280
rect 76377 38303 76400 39280
rect 73370 38280 76400 38303
rect 76560 38303 76583 39280
rect 79567 40280 79590 41287
rect 79750 41287 82780 41310
rect 79750 40280 79773 41287
rect 79567 39280 79773 40280
rect 79567 38303 79590 39280
rect 76560 38280 79590 38303
rect 79750 38303 79773 39280
rect 82757 40280 82780 41287
rect 82940 41287 85970 41310
rect 82940 40280 82963 41287
rect 82757 39280 82963 40280
rect 82757 38303 82780 39280
rect 79750 38280 82780 38303
rect 82940 38303 82963 39280
rect 85947 40280 85970 41287
rect 86130 41287 89160 41310
rect 86130 40280 86153 41287
rect 85947 39280 86153 40280
rect 85947 38303 85970 39280
rect 82940 38280 85970 38303
rect 86130 38303 86153 39280
rect 89137 40280 89160 41287
rect 89320 41287 92350 41310
rect 89320 40280 89343 41287
rect 89137 39280 89343 40280
rect 89137 38303 89160 39280
rect 86130 38280 89160 38303
rect 89320 38303 89343 39280
rect 92327 40280 92350 41287
rect 92510 41287 95540 41310
rect 92510 40280 92533 41287
rect 92327 39280 92533 40280
rect 92327 38303 92350 39280
rect 89320 38280 92350 38303
rect 92510 38303 92533 39280
rect 95517 40280 95540 41287
rect 95700 41287 98730 41310
rect 95700 40280 95723 41287
rect 95517 39280 95723 40280
rect 95517 38303 95540 39280
rect 92510 38280 95540 38303
rect 95700 38303 95723 39280
rect 98707 40280 98730 41287
rect 98890 41287 101920 41310
rect 98890 40280 98913 41287
rect 98707 39280 98913 40280
rect 98707 38303 98730 39280
rect 95700 38280 98730 38303
rect 98890 38303 98913 39280
rect 101897 40280 101920 41287
rect 102080 41287 105110 41310
rect 102080 40280 102103 41287
rect 101897 39280 102103 40280
rect 101897 38303 101920 39280
rect 98890 38280 101920 38303
rect 102080 38303 102103 39280
rect 105087 40280 105110 41287
rect 105270 41287 108300 41310
rect 105270 40280 105293 41287
rect 105087 39280 105293 40280
rect 105087 38303 105110 39280
rect 102080 38280 105110 38303
rect 105270 38303 105293 39280
rect 108277 40280 108300 41287
rect 108460 41287 111490 41310
rect 108460 40280 108483 41287
rect 108277 39280 108483 40280
rect 108277 38303 108300 39280
rect 105270 38280 108300 38303
rect 108460 38303 108483 39280
rect 111467 40280 111490 41287
rect 111650 41287 114680 41310
rect 111650 40280 111673 41287
rect 111467 39280 111673 40280
rect 111467 38303 111490 39280
rect 108460 38280 111490 38303
rect 111650 38303 111673 39280
rect 114657 40280 114680 41287
rect 114840 41287 117870 41310
rect 114840 40280 114863 41287
rect 114657 39280 114863 40280
rect 114657 38303 114680 39280
rect 111650 38280 114680 38303
rect 114840 38303 114863 39280
rect 117847 40280 117870 41287
rect 118030 41287 121060 41310
rect 118030 40280 118053 41287
rect 117847 39280 118053 40280
rect 117847 38303 117870 39280
rect 114840 38280 117870 38303
rect 118030 38303 118053 39280
rect 121037 40280 121060 41287
rect 121220 41287 124250 41310
rect 121220 40280 121243 41287
rect 121037 39280 121243 40280
rect 121037 38303 121060 39280
rect 118030 38280 121060 38303
rect 121220 38303 121243 39280
rect 124227 40280 124250 41287
rect 124410 41287 127440 41310
rect 124410 40280 124433 41287
rect 124227 39280 124433 40280
rect 124227 38303 124250 39280
rect 121220 38280 124250 38303
rect 124410 38303 124433 39280
rect 127417 40280 127440 41287
rect 127600 41287 130630 41310
rect 127600 40280 127623 41287
rect 127417 39280 127623 40280
rect 127417 38303 127440 39280
rect 124410 38280 127440 38303
rect 127600 38303 127623 39280
rect 130607 40280 130630 41287
rect 130790 41287 133820 41310
rect 130790 40280 130813 41287
rect 130607 39280 130813 40280
rect 130607 38303 130630 39280
rect 127600 38280 130630 38303
rect 130790 38303 130813 39280
rect 133797 40280 133820 41287
rect 133980 41287 137010 41310
rect 133980 40280 134003 41287
rect 133797 39280 134003 40280
rect 133797 38303 133820 39280
rect 130790 38280 133820 38303
rect 133980 38303 134003 39280
rect 136987 40280 137010 41287
rect 136987 39280 137170 40280
rect 136987 38303 137010 39280
rect 133980 38280 137010 38303
rect 1000 38120 2000 38280
rect 4190 38120 5190 38280
rect 7380 38120 8380 38280
rect 10570 38120 11570 38280
rect 13760 38120 14760 38280
rect 16950 38120 17950 38280
rect 20140 38120 21140 38280
rect 23330 38120 24330 38280
rect 26520 38120 27520 38280
rect 29710 38120 30710 38280
rect 32900 38120 33900 38280
rect 36090 38120 37090 38280
rect 39280 38120 40280 38280
rect 42470 38120 43470 38280
rect 45660 38120 46660 38280
rect 48850 38120 49850 38280
rect 52040 38120 53040 38280
rect 55230 38120 56230 38280
rect 58420 38120 59420 38280
rect 61610 38120 62610 38280
rect 64800 38120 65800 38280
rect 67990 38120 68990 38280
rect 71180 38120 72180 38280
rect 74370 38120 75370 38280
rect 77560 38120 78560 38280
rect 80750 38120 81750 38280
rect 83940 38120 84940 38280
rect 87130 38120 88130 38280
rect 90320 38120 91320 38280
rect 93510 38120 94510 38280
rect 96700 38120 97700 38280
rect 99890 38120 100890 38280
rect 103080 38120 104080 38280
rect 106270 38120 107270 38280
rect 109460 38120 110460 38280
rect 112650 38120 113650 38280
rect 115840 38120 116840 38280
rect 119030 38120 120030 38280
rect 122220 38120 123220 38280
rect 125410 38120 126410 38280
rect 128600 38120 129600 38280
rect 131790 38120 132790 38280
rect 134980 38120 135980 38280
rect 0 38097 3030 38120
rect 0 35113 23 38097
rect 3007 37090 3030 38097
rect 3190 38097 6220 38120
rect 3190 37090 3213 38097
rect 3007 36090 3213 37090
rect 3007 35113 3030 36090
rect 0 35090 3030 35113
rect 3190 35113 3213 36090
rect 6197 37090 6220 38097
rect 6380 38097 9410 38120
rect 6380 37090 6403 38097
rect 6197 36090 6403 37090
rect 6197 35113 6220 36090
rect 3190 35090 6220 35113
rect 6380 35113 6403 36090
rect 9387 37090 9410 38097
rect 9570 38097 12600 38120
rect 9570 37090 9593 38097
rect 9387 36090 9593 37090
rect 9387 35113 9410 36090
rect 6380 35090 9410 35113
rect 9570 35113 9593 36090
rect 12577 37090 12600 38097
rect 12760 38097 15790 38120
rect 12760 37090 12783 38097
rect 12577 36090 12783 37090
rect 12577 35113 12600 36090
rect 9570 35090 12600 35113
rect 12760 35113 12783 36090
rect 15767 37090 15790 38097
rect 15950 38097 18980 38120
rect 15950 37090 15973 38097
rect 15767 36090 15973 37090
rect 15767 35113 15790 36090
rect 12760 35090 15790 35113
rect 15950 35113 15973 36090
rect 18957 37090 18980 38097
rect 19140 38097 22170 38120
rect 19140 37090 19163 38097
rect 18957 36090 19163 37090
rect 18957 35113 18980 36090
rect 15950 35090 18980 35113
rect 19140 35113 19163 36090
rect 22147 37090 22170 38097
rect 22330 38097 25360 38120
rect 22330 37090 22353 38097
rect 22147 36090 22353 37090
rect 22147 35113 22170 36090
rect 19140 35090 22170 35113
rect 22330 35113 22353 36090
rect 25337 37090 25360 38097
rect 25520 38097 28550 38120
rect 25520 37090 25543 38097
rect 25337 36090 25543 37090
rect 25337 35113 25360 36090
rect 22330 35090 25360 35113
rect 25520 35113 25543 36090
rect 28527 37090 28550 38097
rect 28710 38097 31740 38120
rect 28710 37090 28733 38097
rect 28527 36090 28733 37090
rect 28527 35113 28550 36090
rect 25520 35090 28550 35113
rect 28710 35113 28733 36090
rect 31717 37090 31740 38097
rect 31900 38097 34930 38120
rect 31900 37090 31923 38097
rect 31717 36090 31923 37090
rect 31717 35113 31740 36090
rect 28710 35090 31740 35113
rect 31900 35113 31923 36090
rect 34907 37090 34930 38097
rect 35090 38097 38120 38120
rect 35090 37090 35113 38097
rect 34907 36090 35113 37090
rect 34907 35113 34930 36090
rect 31900 35090 34930 35113
rect 35090 35113 35113 36090
rect 38097 37090 38120 38097
rect 38280 38097 41310 38120
rect 38280 37090 38303 38097
rect 38097 36090 38303 37090
rect 38097 35113 38120 36090
rect 35090 35090 38120 35113
rect 38280 35113 38303 36090
rect 41287 37090 41310 38097
rect 41470 38097 44500 38120
rect 41470 37090 41493 38097
rect 41287 36090 41493 37090
rect 41287 35113 41310 36090
rect 38280 35090 41310 35113
rect 41470 35113 41493 36090
rect 44477 37090 44500 38097
rect 44660 38097 47690 38120
rect 44660 37090 44683 38097
rect 44477 36090 44683 37090
rect 44477 35113 44500 36090
rect 41470 35090 44500 35113
rect 44660 35113 44683 36090
rect 47667 37090 47690 38097
rect 47850 38097 50880 38120
rect 47850 37090 47873 38097
rect 47667 36090 47873 37090
rect 47667 35113 47690 36090
rect 44660 35090 47690 35113
rect 47850 35113 47873 36090
rect 50857 37090 50880 38097
rect 51040 38097 54070 38120
rect 51040 37090 51063 38097
rect 50857 36090 51063 37090
rect 50857 35113 50880 36090
rect 47850 35090 50880 35113
rect 51040 35113 51063 36090
rect 54047 37090 54070 38097
rect 54230 38097 57260 38120
rect 54230 37090 54253 38097
rect 54047 36090 54253 37090
rect 54047 35113 54070 36090
rect 51040 35090 54070 35113
rect 54230 35113 54253 36090
rect 57237 37090 57260 38097
rect 57420 38097 60450 38120
rect 57420 37090 57443 38097
rect 57237 36090 57443 37090
rect 57237 35113 57260 36090
rect 54230 35090 57260 35113
rect 57420 35113 57443 36090
rect 60427 37090 60450 38097
rect 60610 38097 63640 38120
rect 60610 37090 60633 38097
rect 60427 36090 60633 37090
rect 60427 35113 60450 36090
rect 57420 35090 60450 35113
rect 60610 35113 60633 36090
rect 63617 37090 63640 38097
rect 63800 38097 66830 38120
rect 63800 37090 63823 38097
rect 63617 36090 63823 37090
rect 63617 35113 63640 36090
rect 60610 35090 63640 35113
rect 63800 35113 63823 36090
rect 66807 37090 66830 38097
rect 66990 38097 70020 38120
rect 66990 37090 67013 38097
rect 66807 36090 67013 37090
rect 66807 35113 66830 36090
rect 63800 35090 66830 35113
rect 66990 35113 67013 36090
rect 69997 37090 70020 38097
rect 70180 38097 73210 38120
rect 70180 37090 70203 38097
rect 69997 36090 70203 37090
rect 69997 35113 70020 36090
rect 66990 35090 70020 35113
rect 70180 35113 70203 36090
rect 73187 37090 73210 38097
rect 73370 38097 76400 38120
rect 73370 37090 73393 38097
rect 73187 36090 73393 37090
rect 73187 35113 73210 36090
rect 70180 35090 73210 35113
rect 73370 35113 73393 36090
rect 76377 37090 76400 38097
rect 76560 38097 79590 38120
rect 76560 37090 76583 38097
rect 76377 36090 76583 37090
rect 76377 35113 76400 36090
rect 73370 35090 76400 35113
rect 76560 35113 76583 36090
rect 79567 37090 79590 38097
rect 79750 38097 82780 38120
rect 79750 37090 79773 38097
rect 79567 36090 79773 37090
rect 79567 35113 79590 36090
rect 76560 35090 79590 35113
rect 79750 35113 79773 36090
rect 82757 37090 82780 38097
rect 82940 38097 85970 38120
rect 82940 37090 82963 38097
rect 82757 36090 82963 37090
rect 82757 35113 82780 36090
rect 79750 35090 82780 35113
rect 82940 35113 82963 36090
rect 85947 37090 85970 38097
rect 86130 38097 89160 38120
rect 86130 37090 86153 38097
rect 85947 36090 86153 37090
rect 85947 35113 85970 36090
rect 82940 35090 85970 35113
rect 86130 35113 86153 36090
rect 89137 37090 89160 38097
rect 89320 38097 92350 38120
rect 89320 37090 89343 38097
rect 89137 36090 89343 37090
rect 89137 35113 89160 36090
rect 86130 35090 89160 35113
rect 89320 35113 89343 36090
rect 92327 37090 92350 38097
rect 92510 38097 95540 38120
rect 92510 37090 92533 38097
rect 92327 36090 92533 37090
rect 92327 35113 92350 36090
rect 89320 35090 92350 35113
rect 92510 35113 92533 36090
rect 95517 37090 95540 38097
rect 95700 38097 98730 38120
rect 95700 37090 95723 38097
rect 95517 36090 95723 37090
rect 95517 35113 95540 36090
rect 92510 35090 95540 35113
rect 95700 35113 95723 36090
rect 98707 37090 98730 38097
rect 98890 38097 101920 38120
rect 98890 37090 98913 38097
rect 98707 36090 98913 37090
rect 98707 35113 98730 36090
rect 95700 35090 98730 35113
rect 98890 35113 98913 36090
rect 101897 37090 101920 38097
rect 102080 38097 105110 38120
rect 102080 37090 102103 38097
rect 101897 36090 102103 37090
rect 101897 35113 101920 36090
rect 98890 35090 101920 35113
rect 102080 35113 102103 36090
rect 105087 37090 105110 38097
rect 105270 38097 108300 38120
rect 105270 37090 105293 38097
rect 105087 36090 105293 37090
rect 105087 35113 105110 36090
rect 102080 35090 105110 35113
rect 105270 35113 105293 36090
rect 108277 37090 108300 38097
rect 108460 38097 111490 38120
rect 108460 37090 108483 38097
rect 108277 36090 108483 37090
rect 108277 35113 108300 36090
rect 105270 35090 108300 35113
rect 108460 35113 108483 36090
rect 111467 37090 111490 38097
rect 111650 38097 114680 38120
rect 111650 37090 111673 38097
rect 111467 36090 111673 37090
rect 111467 35113 111490 36090
rect 108460 35090 111490 35113
rect 111650 35113 111673 36090
rect 114657 37090 114680 38097
rect 114840 38097 117870 38120
rect 114840 37090 114863 38097
rect 114657 36090 114863 37090
rect 114657 35113 114680 36090
rect 111650 35090 114680 35113
rect 114840 35113 114863 36090
rect 117847 37090 117870 38097
rect 118030 38097 121060 38120
rect 118030 37090 118053 38097
rect 117847 36090 118053 37090
rect 117847 35113 117870 36090
rect 114840 35090 117870 35113
rect 118030 35113 118053 36090
rect 121037 37090 121060 38097
rect 121220 38097 124250 38120
rect 121220 37090 121243 38097
rect 121037 36090 121243 37090
rect 121037 35113 121060 36090
rect 118030 35090 121060 35113
rect 121220 35113 121243 36090
rect 124227 37090 124250 38097
rect 124410 38097 127440 38120
rect 124410 37090 124433 38097
rect 124227 36090 124433 37090
rect 124227 35113 124250 36090
rect 121220 35090 124250 35113
rect 124410 35113 124433 36090
rect 127417 37090 127440 38097
rect 127600 38097 130630 38120
rect 127600 37090 127623 38097
rect 127417 36090 127623 37090
rect 127417 35113 127440 36090
rect 124410 35090 127440 35113
rect 127600 35113 127623 36090
rect 130607 37090 130630 38097
rect 130790 38097 133820 38120
rect 130790 37090 130813 38097
rect 130607 36090 130813 37090
rect 130607 35113 130630 36090
rect 127600 35090 130630 35113
rect 130790 35113 130813 36090
rect 133797 37090 133820 38097
rect 133980 38097 137010 38120
rect 133980 37090 134003 38097
rect 133797 36090 134003 37090
rect 133797 35113 133820 36090
rect 130790 35090 133820 35113
rect 133980 35113 134003 36090
rect 136987 37090 137010 38097
rect 136987 36090 137170 37090
rect 136987 35113 137010 36090
rect 133980 35090 137010 35113
rect 1000 34930 2000 35090
rect 4190 34930 5190 35090
rect 7380 34930 8380 35090
rect 10570 34930 11570 35090
rect 13760 34930 14760 35090
rect 16950 34930 17950 35090
rect 20140 34930 21140 35090
rect 23330 34930 24330 35090
rect 26520 34930 27520 35090
rect 29710 34930 30710 35090
rect 32900 34930 33900 35090
rect 36090 34930 37090 35090
rect 39280 34930 40280 35090
rect 42470 34930 43470 35090
rect 45660 34930 46660 35090
rect 48850 34930 49850 35090
rect 52040 34930 53040 35090
rect 55230 34930 56230 35090
rect 58420 34930 59420 35090
rect 61610 34930 62610 35090
rect 64800 34930 65800 35090
rect 67990 34930 68990 35090
rect 71180 34930 72180 35090
rect 74370 34930 75370 35090
rect 77560 34930 78560 35090
rect 80750 34930 81750 35090
rect 83940 34930 84940 35090
rect 87130 34930 88130 35090
rect 90320 34930 91320 35090
rect 93510 34930 94510 35090
rect 96700 34930 97700 35090
rect 99890 34930 100890 35090
rect 103080 34930 104080 35090
rect 106270 34930 107270 35090
rect 109460 34930 110460 35090
rect 112650 34930 113650 35090
rect 115840 34930 116840 35090
rect 119030 34930 120030 35090
rect 122220 34930 123220 35090
rect 125410 34930 126410 35090
rect 128600 34930 129600 35090
rect 131790 34930 132790 35090
rect 134980 34930 135980 35090
rect 0 34907 3030 34930
rect 0 31923 23 34907
rect 3007 33900 3030 34907
rect 3190 34907 6220 34930
rect 3190 33900 3213 34907
rect 3007 32900 3213 33900
rect 3007 31923 3030 32900
rect 0 31900 3030 31923
rect 3190 31923 3213 32900
rect 6197 33900 6220 34907
rect 6380 34907 9410 34930
rect 6380 33900 6403 34907
rect 6197 32900 6403 33900
rect 6197 31923 6220 32900
rect 3190 31900 6220 31923
rect 6380 31923 6403 32900
rect 9387 33900 9410 34907
rect 9570 34907 12600 34930
rect 9570 33900 9593 34907
rect 9387 32900 9593 33900
rect 9387 31923 9410 32900
rect 6380 31900 9410 31923
rect 9570 31923 9593 32900
rect 12577 33900 12600 34907
rect 12760 34907 15790 34930
rect 12760 33900 12783 34907
rect 12577 32900 12783 33900
rect 12577 31923 12600 32900
rect 9570 31900 12600 31923
rect 12760 31923 12783 32900
rect 15767 33900 15790 34907
rect 15950 34907 18980 34930
rect 15950 33900 15973 34907
rect 15767 32900 15973 33900
rect 15767 31923 15790 32900
rect 12760 31900 15790 31923
rect 15950 31923 15973 32900
rect 18957 33900 18980 34907
rect 19140 34907 22170 34930
rect 19140 33900 19163 34907
rect 18957 32900 19163 33900
rect 18957 31923 18980 32900
rect 15950 31900 18980 31923
rect 19140 31923 19163 32900
rect 22147 33900 22170 34907
rect 22330 34907 25360 34930
rect 22330 33900 22353 34907
rect 22147 32900 22353 33900
rect 22147 31923 22170 32900
rect 19140 31900 22170 31923
rect 22330 31923 22353 32900
rect 25337 33900 25360 34907
rect 25520 34907 28550 34930
rect 25520 33900 25543 34907
rect 25337 32900 25543 33900
rect 25337 31923 25360 32900
rect 22330 31900 25360 31923
rect 25520 31923 25543 32900
rect 28527 33900 28550 34907
rect 28710 34907 31740 34930
rect 28710 33900 28733 34907
rect 28527 32900 28733 33900
rect 28527 31923 28550 32900
rect 25520 31900 28550 31923
rect 28710 31923 28733 32900
rect 31717 33900 31740 34907
rect 31900 34907 34930 34930
rect 31900 33900 31923 34907
rect 31717 32900 31923 33900
rect 31717 31923 31740 32900
rect 28710 31900 31740 31923
rect 31900 31923 31923 32900
rect 34907 33900 34930 34907
rect 35090 34907 38120 34930
rect 35090 33900 35113 34907
rect 34907 32900 35113 33900
rect 34907 31923 34930 32900
rect 31900 31900 34930 31923
rect 35090 31923 35113 32900
rect 38097 33900 38120 34907
rect 38280 34907 41310 34930
rect 38280 33900 38303 34907
rect 38097 32900 38303 33900
rect 38097 31923 38120 32900
rect 35090 31900 38120 31923
rect 38280 31923 38303 32900
rect 41287 33900 41310 34907
rect 41470 34907 44500 34930
rect 41470 33900 41493 34907
rect 41287 32900 41493 33900
rect 41287 31923 41310 32900
rect 38280 31900 41310 31923
rect 41470 31923 41493 32900
rect 44477 33900 44500 34907
rect 44660 34907 47690 34930
rect 44660 33900 44683 34907
rect 44477 32900 44683 33900
rect 44477 31923 44500 32900
rect 41470 31900 44500 31923
rect 44660 31923 44683 32900
rect 47667 33900 47690 34907
rect 47850 34907 50880 34930
rect 47850 33900 47873 34907
rect 47667 32900 47873 33900
rect 47667 31923 47690 32900
rect 44660 31900 47690 31923
rect 47850 31923 47873 32900
rect 50857 33900 50880 34907
rect 51040 34907 54070 34930
rect 51040 33900 51063 34907
rect 50857 32900 51063 33900
rect 50857 31923 50880 32900
rect 47850 31900 50880 31923
rect 51040 31923 51063 32900
rect 54047 33900 54070 34907
rect 54230 34907 57260 34930
rect 54230 33900 54253 34907
rect 54047 32900 54253 33900
rect 54047 31923 54070 32900
rect 51040 31900 54070 31923
rect 54230 31923 54253 32900
rect 57237 33900 57260 34907
rect 57420 34907 60450 34930
rect 57420 33900 57443 34907
rect 57237 32900 57443 33900
rect 57237 31923 57260 32900
rect 54230 31900 57260 31923
rect 57420 31923 57443 32900
rect 60427 33900 60450 34907
rect 60610 34907 63640 34930
rect 60610 33900 60633 34907
rect 60427 32900 60633 33900
rect 60427 31923 60450 32900
rect 57420 31900 60450 31923
rect 60610 31923 60633 32900
rect 63617 33900 63640 34907
rect 63800 34907 66830 34930
rect 63800 33900 63823 34907
rect 63617 32900 63823 33900
rect 63617 31923 63640 32900
rect 60610 31900 63640 31923
rect 63800 31923 63823 32900
rect 66807 33900 66830 34907
rect 66990 34907 70020 34930
rect 66990 33900 67013 34907
rect 66807 32900 67013 33900
rect 66807 31923 66830 32900
rect 63800 31900 66830 31923
rect 66990 31923 67013 32900
rect 69997 33900 70020 34907
rect 70180 34907 73210 34930
rect 70180 33900 70203 34907
rect 69997 32900 70203 33900
rect 69997 31923 70020 32900
rect 66990 31900 70020 31923
rect 70180 31923 70203 32900
rect 73187 33900 73210 34907
rect 73370 34907 76400 34930
rect 73370 33900 73393 34907
rect 73187 32900 73393 33900
rect 73187 31923 73210 32900
rect 70180 31900 73210 31923
rect 73370 31923 73393 32900
rect 76377 33900 76400 34907
rect 76560 34907 79590 34930
rect 76560 33900 76583 34907
rect 76377 32900 76583 33900
rect 76377 31923 76400 32900
rect 73370 31900 76400 31923
rect 76560 31923 76583 32900
rect 79567 33900 79590 34907
rect 79750 34907 82780 34930
rect 79750 33900 79773 34907
rect 79567 32900 79773 33900
rect 79567 31923 79590 32900
rect 76560 31900 79590 31923
rect 79750 31923 79773 32900
rect 82757 33900 82780 34907
rect 82940 34907 85970 34930
rect 82940 33900 82963 34907
rect 82757 32900 82963 33900
rect 82757 31923 82780 32900
rect 79750 31900 82780 31923
rect 82940 31923 82963 32900
rect 85947 33900 85970 34907
rect 86130 34907 89160 34930
rect 86130 33900 86153 34907
rect 85947 32900 86153 33900
rect 85947 31923 85970 32900
rect 82940 31900 85970 31923
rect 86130 31923 86153 32900
rect 89137 33900 89160 34907
rect 89320 34907 92350 34930
rect 89320 33900 89343 34907
rect 89137 32900 89343 33900
rect 89137 31923 89160 32900
rect 86130 31900 89160 31923
rect 89320 31923 89343 32900
rect 92327 33900 92350 34907
rect 92510 34907 95540 34930
rect 92510 33900 92533 34907
rect 92327 32900 92533 33900
rect 92327 31923 92350 32900
rect 89320 31900 92350 31923
rect 92510 31923 92533 32900
rect 95517 33900 95540 34907
rect 95700 34907 98730 34930
rect 95700 33900 95723 34907
rect 95517 32900 95723 33900
rect 95517 31923 95540 32900
rect 92510 31900 95540 31923
rect 95700 31923 95723 32900
rect 98707 33900 98730 34907
rect 98890 34907 101920 34930
rect 98890 33900 98913 34907
rect 98707 32900 98913 33900
rect 98707 31923 98730 32900
rect 95700 31900 98730 31923
rect 98890 31923 98913 32900
rect 101897 33900 101920 34907
rect 102080 34907 105110 34930
rect 102080 33900 102103 34907
rect 101897 32900 102103 33900
rect 101897 31923 101920 32900
rect 98890 31900 101920 31923
rect 102080 31923 102103 32900
rect 105087 33900 105110 34907
rect 105270 34907 108300 34930
rect 105270 33900 105293 34907
rect 105087 32900 105293 33900
rect 105087 31923 105110 32900
rect 102080 31900 105110 31923
rect 105270 31923 105293 32900
rect 108277 33900 108300 34907
rect 108460 34907 111490 34930
rect 108460 33900 108483 34907
rect 108277 32900 108483 33900
rect 108277 31923 108300 32900
rect 105270 31900 108300 31923
rect 108460 31923 108483 32900
rect 111467 33900 111490 34907
rect 111650 34907 114680 34930
rect 111650 33900 111673 34907
rect 111467 32900 111673 33900
rect 111467 31923 111490 32900
rect 108460 31900 111490 31923
rect 111650 31923 111673 32900
rect 114657 33900 114680 34907
rect 114840 34907 117870 34930
rect 114840 33900 114863 34907
rect 114657 32900 114863 33900
rect 114657 31923 114680 32900
rect 111650 31900 114680 31923
rect 114840 31923 114863 32900
rect 117847 33900 117870 34907
rect 118030 34907 121060 34930
rect 118030 33900 118053 34907
rect 117847 32900 118053 33900
rect 117847 31923 117870 32900
rect 114840 31900 117870 31923
rect 118030 31923 118053 32900
rect 121037 33900 121060 34907
rect 121220 34907 124250 34930
rect 121220 33900 121243 34907
rect 121037 32900 121243 33900
rect 121037 31923 121060 32900
rect 118030 31900 121060 31923
rect 121220 31923 121243 32900
rect 124227 33900 124250 34907
rect 124410 34907 127440 34930
rect 124410 33900 124433 34907
rect 124227 32900 124433 33900
rect 124227 31923 124250 32900
rect 121220 31900 124250 31923
rect 124410 31923 124433 32900
rect 127417 33900 127440 34907
rect 127600 34907 130630 34930
rect 127600 33900 127623 34907
rect 127417 32900 127623 33900
rect 127417 31923 127440 32900
rect 124410 31900 127440 31923
rect 127600 31923 127623 32900
rect 130607 33900 130630 34907
rect 130790 34907 133820 34930
rect 130790 33900 130813 34907
rect 130607 32900 130813 33900
rect 130607 31923 130630 32900
rect 127600 31900 130630 31923
rect 130790 31923 130813 32900
rect 133797 33900 133820 34907
rect 133980 34907 137010 34930
rect 133980 33900 134003 34907
rect 133797 32900 134003 33900
rect 133797 31923 133820 32900
rect 130790 31900 133820 31923
rect 133980 31923 134003 32900
rect 136987 33900 137010 34907
rect 136987 32900 137170 33900
rect 136987 31923 137010 32900
rect 133980 31900 137010 31923
rect 1000 31740 2000 31900
rect 4190 31740 5190 31900
rect 7380 31740 8380 31900
rect 10570 31740 11570 31900
rect 13760 31740 14760 31900
rect 16950 31740 17950 31900
rect 20140 31740 21140 31900
rect 23330 31740 24330 31900
rect 26520 31740 27520 31900
rect 29710 31740 30710 31900
rect 32900 31740 33900 31900
rect 36090 31740 37090 31900
rect 39280 31740 40280 31900
rect 42470 31740 43470 31900
rect 45660 31740 46660 31900
rect 48850 31740 49850 31900
rect 52040 31740 53040 31900
rect 55230 31740 56230 31900
rect 58420 31740 59420 31900
rect 61610 31740 62610 31900
rect 64800 31740 65800 31900
rect 67990 31740 68990 31900
rect 71180 31740 72180 31900
rect 74370 31740 75370 31900
rect 77560 31740 78560 31900
rect 80750 31740 81750 31900
rect 83940 31740 84940 31900
rect 87130 31740 88130 31900
rect 90320 31740 91320 31900
rect 93510 31740 94510 31900
rect 96700 31740 97700 31900
rect 99890 31740 100890 31900
rect 103080 31740 104080 31900
rect 106270 31740 107270 31900
rect 109460 31740 110460 31900
rect 112650 31740 113650 31900
rect 115840 31740 116840 31900
rect 119030 31740 120030 31900
rect 122220 31740 123220 31900
rect 125410 31740 126410 31900
rect 128600 31740 129600 31900
rect 131790 31740 132790 31900
rect 134980 31740 135980 31900
rect 0 31717 3030 31740
rect 0 28733 23 31717
rect 3007 30710 3030 31717
rect 3190 31717 6220 31740
rect 3190 30710 3213 31717
rect 3007 29710 3213 30710
rect 3007 28733 3030 29710
rect 0 28710 3030 28733
rect 3190 28733 3213 29710
rect 6197 30710 6220 31717
rect 6380 31717 9410 31740
rect 6380 30710 6403 31717
rect 6197 29710 6403 30710
rect 6197 28733 6220 29710
rect 3190 28710 6220 28733
rect 6380 28733 6403 29710
rect 9387 30710 9410 31717
rect 9570 31717 12600 31740
rect 9570 30710 9593 31717
rect 9387 29710 9593 30710
rect 9387 28733 9410 29710
rect 6380 28710 9410 28733
rect 9570 28733 9593 29710
rect 12577 30710 12600 31717
rect 12760 31717 15790 31740
rect 12760 30710 12783 31717
rect 12577 29710 12783 30710
rect 12577 28733 12600 29710
rect 9570 28710 12600 28733
rect 12760 28733 12783 29710
rect 15767 30710 15790 31717
rect 15950 31717 18980 31740
rect 15950 30710 15973 31717
rect 15767 29710 15973 30710
rect 15767 28733 15790 29710
rect 12760 28710 15790 28733
rect 15950 28733 15973 29710
rect 18957 30710 18980 31717
rect 19140 31717 22170 31740
rect 19140 30710 19163 31717
rect 18957 29710 19163 30710
rect 18957 28733 18980 29710
rect 15950 28710 18980 28733
rect 19140 28733 19163 29710
rect 22147 30710 22170 31717
rect 22330 31717 25360 31740
rect 22330 30710 22353 31717
rect 22147 29710 22353 30710
rect 22147 28733 22170 29710
rect 19140 28710 22170 28733
rect 22330 28733 22353 29710
rect 25337 30710 25360 31717
rect 25520 31717 28550 31740
rect 25520 30710 25543 31717
rect 25337 29710 25543 30710
rect 25337 28733 25360 29710
rect 22330 28710 25360 28733
rect 25520 28733 25543 29710
rect 28527 30710 28550 31717
rect 28710 31717 31740 31740
rect 28710 30710 28733 31717
rect 28527 29710 28733 30710
rect 28527 28733 28550 29710
rect 25520 28710 28550 28733
rect 28710 28733 28733 29710
rect 31717 30710 31740 31717
rect 31900 31717 34930 31740
rect 31900 30710 31923 31717
rect 31717 29710 31923 30710
rect 31717 28733 31740 29710
rect 28710 28710 31740 28733
rect 31900 28733 31923 29710
rect 34907 30710 34930 31717
rect 35090 31717 38120 31740
rect 35090 30710 35113 31717
rect 34907 29710 35113 30710
rect 34907 28733 34930 29710
rect 31900 28710 34930 28733
rect 35090 28733 35113 29710
rect 38097 30710 38120 31717
rect 38280 31717 41310 31740
rect 38280 30710 38303 31717
rect 38097 29710 38303 30710
rect 38097 28733 38120 29710
rect 35090 28710 38120 28733
rect 38280 28733 38303 29710
rect 41287 30710 41310 31717
rect 41470 31717 44500 31740
rect 41470 30710 41493 31717
rect 41287 29710 41493 30710
rect 41287 28733 41310 29710
rect 38280 28710 41310 28733
rect 41470 28733 41493 29710
rect 44477 30710 44500 31717
rect 44660 31717 47690 31740
rect 44660 30710 44683 31717
rect 44477 29710 44683 30710
rect 44477 28733 44500 29710
rect 41470 28710 44500 28733
rect 44660 28733 44683 29710
rect 47667 30710 47690 31717
rect 47850 31717 50880 31740
rect 47850 30710 47873 31717
rect 47667 29710 47873 30710
rect 47667 28733 47690 29710
rect 44660 28710 47690 28733
rect 47850 28733 47873 29710
rect 50857 30710 50880 31717
rect 51040 31717 54070 31740
rect 51040 30710 51063 31717
rect 50857 29710 51063 30710
rect 50857 28733 50880 29710
rect 47850 28710 50880 28733
rect 51040 28733 51063 29710
rect 54047 30710 54070 31717
rect 54230 31717 57260 31740
rect 54230 30710 54253 31717
rect 54047 29710 54253 30710
rect 54047 28733 54070 29710
rect 51040 28710 54070 28733
rect 54230 28733 54253 29710
rect 57237 30710 57260 31717
rect 57420 31717 60450 31740
rect 57420 30710 57443 31717
rect 57237 29710 57443 30710
rect 57237 28733 57260 29710
rect 54230 28710 57260 28733
rect 57420 28733 57443 29710
rect 60427 30710 60450 31717
rect 60610 31717 63640 31740
rect 60610 30710 60633 31717
rect 60427 29710 60633 30710
rect 60427 28733 60450 29710
rect 57420 28710 60450 28733
rect 60610 28733 60633 29710
rect 63617 30710 63640 31717
rect 63800 31717 66830 31740
rect 63800 30710 63823 31717
rect 63617 29710 63823 30710
rect 63617 28733 63640 29710
rect 60610 28710 63640 28733
rect 63800 28733 63823 29710
rect 66807 30710 66830 31717
rect 66990 31717 70020 31740
rect 66990 30710 67013 31717
rect 66807 29710 67013 30710
rect 66807 28733 66830 29710
rect 63800 28710 66830 28733
rect 66990 28733 67013 29710
rect 69997 30710 70020 31717
rect 70180 31717 73210 31740
rect 70180 30710 70203 31717
rect 69997 29710 70203 30710
rect 69997 28733 70020 29710
rect 66990 28710 70020 28733
rect 70180 28733 70203 29710
rect 73187 30710 73210 31717
rect 73370 31717 76400 31740
rect 73370 30710 73393 31717
rect 73187 29710 73393 30710
rect 73187 28733 73210 29710
rect 70180 28710 73210 28733
rect 73370 28733 73393 29710
rect 76377 30710 76400 31717
rect 76560 31717 79590 31740
rect 76560 30710 76583 31717
rect 76377 29710 76583 30710
rect 76377 28733 76400 29710
rect 73370 28710 76400 28733
rect 76560 28733 76583 29710
rect 79567 30710 79590 31717
rect 79750 31717 82780 31740
rect 79750 30710 79773 31717
rect 79567 29710 79773 30710
rect 79567 28733 79590 29710
rect 76560 28710 79590 28733
rect 79750 28733 79773 29710
rect 82757 30710 82780 31717
rect 82940 31717 85970 31740
rect 82940 30710 82963 31717
rect 82757 29710 82963 30710
rect 82757 28733 82780 29710
rect 79750 28710 82780 28733
rect 82940 28733 82963 29710
rect 85947 30710 85970 31717
rect 86130 31717 89160 31740
rect 86130 30710 86153 31717
rect 85947 29710 86153 30710
rect 85947 28733 85970 29710
rect 82940 28710 85970 28733
rect 86130 28733 86153 29710
rect 89137 30710 89160 31717
rect 89320 31717 92350 31740
rect 89320 30710 89343 31717
rect 89137 29710 89343 30710
rect 89137 28733 89160 29710
rect 86130 28710 89160 28733
rect 89320 28733 89343 29710
rect 92327 30710 92350 31717
rect 92510 31717 95540 31740
rect 92510 30710 92533 31717
rect 92327 29710 92533 30710
rect 92327 28733 92350 29710
rect 89320 28710 92350 28733
rect 92510 28733 92533 29710
rect 95517 30710 95540 31717
rect 95700 31717 98730 31740
rect 95700 30710 95723 31717
rect 95517 29710 95723 30710
rect 95517 28733 95540 29710
rect 92510 28710 95540 28733
rect 95700 28733 95723 29710
rect 98707 30710 98730 31717
rect 98890 31717 101920 31740
rect 98890 30710 98913 31717
rect 98707 29710 98913 30710
rect 98707 28733 98730 29710
rect 95700 28710 98730 28733
rect 98890 28733 98913 29710
rect 101897 30710 101920 31717
rect 102080 31717 105110 31740
rect 102080 30710 102103 31717
rect 101897 29710 102103 30710
rect 101897 28733 101920 29710
rect 98890 28710 101920 28733
rect 102080 28733 102103 29710
rect 105087 30710 105110 31717
rect 105270 31717 108300 31740
rect 105270 30710 105293 31717
rect 105087 29710 105293 30710
rect 105087 28733 105110 29710
rect 102080 28710 105110 28733
rect 105270 28733 105293 29710
rect 108277 30710 108300 31717
rect 108460 31717 111490 31740
rect 108460 30710 108483 31717
rect 108277 29710 108483 30710
rect 108277 28733 108300 29710
rect 105270 28710 108300 28733
rect 108460 28733 108483 29710
rect 111467 30710 111490 31717
rect 111650 31717 114680 31740
rect 111650 30710 111673 31717
rect 111467 29710 111673 30710
rect 111467 28733 111490 29710
rect 108460 28710 111490 28733
rect 111650 28733 111673 29710
rect 114657 30710 114680 31717
rect 114840 31717 117870 31740
rect 114840 30710 114863 31717
rect 114657 29710 114863 30710
rect 114657 28733 114680 29710
rect 111650 28710 114680 28733
rect 114840 28733 114863 29710
rect 117847 30710 117870 31717
rect 118030 31717 121060 31740
rect 118030 30710 118053 31717
rect 117847 29710 118053 30710
rect 117847 28733 117870 29710
rect 114840 28710 117870 28733
rect 118030 28733 118053 29710
rect 121037 30710 121060 31717
rect 121220 31717 124250 31740
rect 121220 30710 121243 31717
rect 121037 29710 121243 30710
rect 121037 28733 121060 29710
rect 118030 28710 121060 28733
rect 121220 28733 121243 29710
rect 124227 30710 124250 31717
rect 124410 31717 127440 31740
rect 124410 30710 124433 31717
rect 124227 29710 124433 30710
rect 124227 28733 124250 29710
rect 121220 28710 124250 28733
rect 124410 28733 124433 29710
rect 127417 30710 127440 31717
rect 127600 31717 130630 31740
rect 127600 30710 127623 31717
rect 127417 29710 127623 30710
rect 127417 28733 127440 29710
rect 124410 28710 127440 28733
rect 127600 28733 127623 29710
rect 130607 30710 130630 31717
rect 130790 31717 133820 31740
rect 130790 30710 130813 31717
rect 130607 29710 130813 30710
rect 130607 28733 130630 29710
rect 127600 28710 130630 28733
rect 130790 28733 130813 29710
rect 133797 30710 133820 31717
rect 133980 31717 137010 31740
rect 133980 30710 134003 31717
rect 133797 29710 134003 30710
rect 133797 28733 133820 29710
rect 130790 28710 133820 28733
rect 133980 28733 134003 29710
rect 136987 30710 137010 31717
rect 136987 29710 137170 30710
rect 136987 28733 137010 29710
rect 133980 28710 137010 28733
rect 1000 28550 2000 28710
rect 4190 28550 5190 28710
rect 7380 28550 8380 28710
rect 10570 28550 11570 28710
rect 13760 28550 14760 28710
rect 16950 28550 17950 28710
rect 20140 28550 21140 28710
rect 23330 28550 24330 28710
rect 26520 28550 27520 28710
rect 29710 28550 30710 28710
rect 32900 28550 33900 28710
rect 36090 28550 37090 28710
rect 39280 28550 40280 28710
rect 42470 28550 43470 28710
rect 45660 28550 46660 28710
rect 48850 28550 49850 28710
rect 52040 28550 53040 28710
rect 55230 28550 56230 28710
rect 58420 28550 59420 28710
rect 61610 28550 62610 28710
rect 64800 28550 65800 28710
rect 67990 28550 68990 28710
rect 71180 28550 72180 28710
rect 74370 28550 75370 28710
rect 77560 28550 78560 28710
rect 80750 28550 81750 28710
rect 83940 28550 84940 28710
rect 87130 28550 88130 28710
rect 90320 28550 91320 28710
rect 93510 28550 94510 28710
rect 96700 28550 97700 28710
rect 99890 28550 100890 28710
rect 103080 28550 104080 28710
rect 106270 28550 107270 28710
rect 109460 28550 110460 28710
rect 112650 28550 113650 28710
rect 115840 28550 116840 28710
rect 119030 28550 120030 28710
rect 122220 28550 123220 28710
rect 125410 28550 126410 28710
rect 128600 28550 129600 28710
rect 131790 28550 132790 28710
rect 134980 28550 135980 28710
rect 0 28527 3030 28550
rect 0 25543 23 28527
rect 3007 27520 3030 28527
rect 3190 28527 6220 28550
rect 3190 27520 3213 28527
rect 3007 26520 3213 27520
rect 3007 25543 3030 26520
rect 0 25520 3030 25543
rect 3190 25543 3213 26520
rect 6197 27520 6220 28527
rect 6380 28527 9410 28550
rect 6380 27520 6403 28527
rect 6197 26520 6403 27520
rect 6197 25543 6220 26520
rect 3190 25520 6220 25543
rect 6380 25543 6403 26520
rect 9387 27520 9410 28527
rect 9570 28527 12600 28550
rect 9570 27520 9593 28527
rect 9387 26520 9593 27520
rect 9387 25543 9410 26520
rect 6380 25520 9410 25543
rect 9570 25543 9593 26520
rect 12577 27520 12600 28527
rect 12760 28527 15790 28550
rect 12760 27520 12783 28527
rect 12577 26520 12783 27520
rect 12577 25543 12600 26520
rect 9570 25520 12600 25543
rect 12760 25543 12783 26520
rect 15767 27520 15790 28527
rect 15950 28527 18980 28550
rect 15950 27520 15973 28527
rect 15767 26520 15973 27520
rect 15767 25543 15790 26520
rect 12760 25520 15790 25543
rect 15950 25543 15973 26520
rect 18957 27520 18980 28527
rect 19140 28527 22170 28550
rect 19140 27520 19163 28527
rect 18957 26520 19163 27520
rect 18957 25543 18980 26520
rect 15950 25520 18980 25543
rect 19140 25543 19163 26520
rect 22147 27520 22170 28527
rect 22330 28527 25360 28550
rect 22330 27520 22353 28527
rect 22147 26520 22353 27520
rect 22147 25543 22170 26520
rect 19140 25520 22170 25543
rect 22330 25543 22353 26520
rect 25337 27520 25360 28527
rect 25520 28527 28550 28550
rect 25520 27520 25543 28527
rect 25337 26520 25543 27520
rect 25337 25543 25360 26520
rect 22330 25520 25360 25543
rect 25520 25543 25543 26520
rect 28527 27520 28550 28527
rect 28710 28527 31740 28550
rect 28710 27520 28733 28527
rect 28527 26520 28733 27520
rect 28527 25543 28550 26520
rect 25520 25520 28550 25543
rect 28710 25543 28733 26520
rect 31717 27520 31740 28527
rect 31900 28527 34930 28550
rect 31900 27520 31923 28527
rect 31717 26520 31923 27520
rect 31717 25543 31740 26520
rect 28710 25520 31740 25543
rect 31900 25543 31923 26520
rect 34907 27520 34930 28527
rect 35090 28527 38120 28550
rect 35090 27520 35113 28527
rect 34907 26520 35113 27520
rect 34907 25543 34930 26520
rect 31900 25520 34930 25543
rect 35090 25543 35113 26520
rect 38097 27520 38120 28527
rect 38280 28527 41310 28550
rect 38280 27520 38303 28527
rect 38097 26520 38303 27520
rect 38097 25543 38120 26520
rect 35090 25520 38120 25543
rect 38280 25543 38303 26520
rect 41287 27520 41310 28527
rect 41470 28527 44500 28550
rect 41470 27520 41493 28527
rect 41287 26520 41493 27520
rect 41287 25543 41310 26520
rect 38280 25520 41310 25543
rect 41470 25543 41493 26520
rect 44477 27520 44500 28527
rect 44660 28527 47690 28550
rect 44660 27520 44683 28527
rect 44477 26520 44683 27520
rect 44477 25543 44500 26520
rect 41470 25520 44500 25543
rect 44660 25543 44683 26520
rect 47667 27520 47690 28527
rect 47850 28527 50880 28550
rect 47850 27520 47873 28527
rect 47667 26520 47873 27520
rect 47667 25543 47690 26520
rect 44660 25520 47690 25543
rect 47850 25543 47873 26520
rect 50857 27520 50880 28527
rect 51040 28527 54070 28550
rect 51040 27520 51063 28527
rect 50857 26520 51063 27520
rect 50857 25543 50880 26520
rect 47850 25520 50880 25543
rect 51040 25543 51063 26520
rect 54047 27520 54070 28527
rect 54230 28527 57260 28550
rect 54230 27520 54253 28527
rect 54047 26520 54253 27520
rect 54047 25543 54070 26520
rect 51040 25520 54070 25543
rect 54230 25543 54253 26520
rect 57237 27520 57260 28527
rect 57420 28527 60450 28550
rect 57420 27520 57443 28527
rect 57237 26520 57443 27520
rect 57237 25543 57260 26520
rect 54230 25520 57260 25543
rect 57420 25543 57443 26520
rect 60427 27520 60450 28527
rect 60610 28527 63640 28550
rect 60610 27520 60633 28527
rect 60427 26520 60633 27520
rect 60427 25543 60450 26520
rect 57420 25520 60450 25543
rect 60610 25543 60633 26520
rect 63617 27520 63640 28527
rect 63800 28527 66830 28550
rect 63800 27520 63823 28527
rect 63617 26520 63823 27520
rect 63617 25543 63640 26520
rect 60610 25520 63640 25543
rect 63800 25543 63823 26520
rect 66807 27520 66830 28527
rect 66990 28527 70020 28550
rect 66990 27520 67013 28527
rect 66807 26520 67013 27520
rect 66807 25543 66830 26520
rect 63800 25520 66830 25543
rect 66990 25543 67013 26520
rect 69997 27520 70020 28527
rect 70180 28527 73210 28550
rect 70180 27520 70203 28527
rect 69997 26520 70203 27520
rect 69997 25543 70020 26520
rect 66990 25520 70020 25543
rect 70180 25543 70203 26520
rect 73187 27520 73210 28527
rect 73370 28527 76400 28550
rect 73370 27520 73393 28527
rect 73187 26520 73393 27520
rect 73187 25543 73210 26520
rect 70180 25520 73210 25543
rect 73370 25543 73393 26520
rect 76377 27520 76400 28527
rect 76560 28527 79590 28550
rect 76560 27520 76583 28527
rect 76377 26520 76583 27520
rect 76377 25543 76400 26520
rect 73370 25520 76400 25543
rect 76560 25543 76583 26520
rect 79567 27520 79590 28527
rect 79750 28527 82780 28550
rect 79750 27520 79773 28527
rect 79567 26520 79773 27520
rect 79567 25543 79590 26520
rect 76560 25520 79590 25543
rect 79750 25543 79773 26520
rect 82757 27520 82780 28527
rect 82940 28527 85970 28550
rect 82940 27520 82963 28527
rect 82757 26520 82963 27520
rect 82757 25543 82780 26520
rect 79750 25520 82780 25543
rect 82940 25543 82963 26520
rect 85947 27520 85970 28527
rect 86130 28527 89160 28550
rect 86130 27520 86153 28527
rect 85947 26520 86153 27520
rect 85947 25543 85970 26520
rect 82940 25520 85970 25543
rect 86130 25543 86153 26520
rect 89137 27520 89160 28527
rect 89320 28527 92350 28550
rect 89320 27520 89343 28527
rect 89137 26520 89343 27520
rect 89137 25543 89160 26520
rect 86130 25520 89160 25543
rect 89320 25543 89343 26520
rect 92327 27520 92350 28527
rect 92510 28527 95540 28550
rect 92510 27520 92533 28527
rect 92327 26520 92533 27520
rect 92327 25543 92350 26520
rect 89320 25520 92350 25543
rect 92510 25543 92533 26520
rect 95517 27520 95540 28527
rect 95700 28527 98730 28550
rect 95700 27520 95723 28527
rect 95517 26520 95723 27520
rect 95517 25543 95540 26520
rect 92510 25520 95540 25543
rect 95700 25543 95723 26520
rect 98707 27520 98730 28527
rect 98890 28527 101920 28550
rect 98890 27520 98913 28527
rect 98707 26520 98913 27520
rect 98707 25543 98730 26520
rect 95700 25520 98730 25543
rect 98890 25543 98913 26520
rect 101897 27520 101920 28527
rect 102080 28527 105110 28550
rect 102080 27520 102103 28527
rect 101897 26520 102103 27520
rect 101897 25543 101920 26520
rect 98890 25520 101920 25543
rect 102080 25543 102103 26520
rect 105087 27520 105110 28527
rect 105270 28527 108300 28550
rect 105270 27520 105293 28527
rect 105087 26520 105293 27520
rect 105087 25543 105110 26520
rect 102080 25520 105110 25543
rect 105270 25543 105293 26520
rect 108277 27520 108300 28527
rect 108460 28527 111490 28550
rect 108460 27520 108483 28527
rect 108277 26520 108483 27520
rect 108277 25543 108300 26520
rect 105270 25520 108300 25543
rect 108460 25543 108483 26520
rect 111467 27520 111490 28527
rect 111650 28527 114680 28550
rect 111650 27520 111673 28527
rect 111467 26520 111673 27520
rect 111467 25543 111490 26520
rect 108460 25520 111490 25543
rect 111650 25543 111673 26520
rect 114657 27520 114680 28527
rect 114840 28527 117870 28550
rect 114840 27520 114863 28527
rect 114657 26520 114863 27520
rect 114657 25543 114680 26520
rect 111650 25520 114680 25543
rect 114840 25543 114863 26520
rect 117847 27520 117870 28527
rect 118030 28527 121060 28550
rect 118030 27520 118053 28527
rect 117847 26520 118053 27520
rect 117847 25543 117870 26520
rect 114840 25520 117870 25543
rect 118030 25543 118053 26520
rect 121037 27520 121060 28527
rect 121220 28527 124250 28550
rect 121220 27520 121243 28527
rect 121037 26520 121243 27520
rect 121037 25543 121060 26520
rect 118030 25520 121060 25543
rect 121220 25543 121243 26520
rect 124227 27520 124250 28527
rect 124410 28527 127440 28550
rect 124410 27520 124433 28527
rect 124227 26520 124433 27520
rect 124227 25543 124250 26520
rect 121220 25520 124250 25543
rect 124410 25543 124433 26520
rect 127417 27520 127440 28527
rect 127600 28527 130630 28550
rect 127600 27520 127623 28527
rect 127417 26520 127623 27520
rect 127417 25543 127440 26520
rect 124410 25520 127440 25543
rect 127600 25543 127623 26520
rect 130607 27520 130630 28527
rect 130790 28527 133820 28550
rect 130790 27520 130813 28527
rect 130607 26520 130813 27520
rect 130607 25543 130630 26520
rect 127600 25520 130630 25543
rect 130790 25543 130813 26520
rect 133797 27520 133820 28527
rect 133980 28527 137010 28550
rect 133980 27520 134003 28527
rect 133797 26520 134003 27520
rect 133797 25543 133820 26520
rect 130790 25520 133820 25543
rect 133980 25543 134003 26520
rect 136987 27520 137010 28527
rect 136987 26520 137170 27520
rect 136987 25543 137010 26520
rect 133980 25520 137010 25543
rect 1000 25360 2000 25520
rect 4190 25360 5190 25520
rect 7380 25360 8380 25520
rect 10570 25360 11570 25520
rect 13760 25360 14760 25520
rect 16950 25360 17950 25520
rect 20140 25360 21140 25520
rect 23330 25360 24330 25520
rect 26520 25360 27520 25520
rect 29710 25360 30710 25520
rect 32900 25360 33900 25520
rect 36090 25360 37090 25520
rect 39280 25360 40280 25520
rect 42470 25360 43470 25520
rect 45660 25360 46660 25520
rect 48850 25360 49850 25520
rect 52040 25360 53040 25520
rect 55230 25360 56230 25520
rect 58420 25360 59420 25520
rect 61610 25360 62610 25520
rect 64800 25360 65800 25520
rect 67990 25360 68990 25520
rect 71180 25360 72180 25520
rect 74370 25360 75370 25520
rect 77560 25360 78560 25520
rect 80750 25360 81750 25520
rect 83940 25360 84940 25520
rect 87130 25360 88130 25520
rect 90320 25360 91320 25520
rect 93510 25360 94510 25520
rect 96700 25360 97700 25520
rect 99890 25360 100890 25520
rect 103080 25360 104080 25520
rect 106270 25360 107270 25520
rect 109460 25360 110460 25520
rect 112650 25360 113650 25520
rect 115840 25360 116840 25520
rect 119030 25360 120030 25520
rect 122220 25360 123220 25520
rect 125410 25360 126410 25520
rect 128600 25360 129600 25520
rect 131790 25360 132790 25520
rect 134980 25360 135980 25520
rect 0 25337 3030 25360
rect 0 22353 23 25337
rect 3007 24330 3030 25337
rect 3190 25337 6220 25360
rect 3190 24330 3213 25337
rect 3007 23330 3213 24330
rect 3007 22353 3030 23330
rect 0 22330 3030 22353
rect 3190 22353 3213 23330
rect 6197 24330 6220 25337
rect 6380 25337 9410 25360
rect 6380 24330 6403 25337
rect 6197 23330 6403 24330
rect 6197 22353 6220 23330
rect 3190 22330 6220 22353
rect 6380 22353 6403 23330
rect 9387 24330 9410 25337
rect 9570 25337 12600 25360
rect 9570 24330 9593 25337
rect 9387 23330 9593 24330
rect 9387 22353 9410 23330
rect 6380 22330 9410 22353
rect 9570 22353 9593 23330
rect 12577 24330 12600 25337
rect 12760 25337 15790 25360
rect 12760 24330 12783 25337
rect 12577 23330 12783 24330
rect 12577 22353 12600 23330
rect 9570 22330 12600 22353
rect 12760 22353 12783 23330
rect 15767 24330 15790 25337
rect 15950 25337 18980 25360
rect 15950 24330 15973 25337
rect 15767 23330 15973 24330
rect 15767 22353 15790 23330
rect 12760 22330 15790 22353
rect 15950 22353 15973 23330
rect 18957 24330 18980 25337
rect 19140 25337 22170 25360
rect 19140 24330 19163 25337
rect 18957 23330 19163 24330
rect 18957 22353 18980 23330
rect 15950 22330 18980 22353
rect 19140 22353 19163 23330
rect 22147 24330 22170 25337
rect 22330 25337 25360 25360
rect 22330 24330 22353 25337
rect 22147 23330 22353 24330
rect 22147 22353 22170 23330
rect 19140 22330 22170 22353
rect 22330 22353 22353 23330
rect 25337 24330 25360 25337
rect 25520 25337 28550 25360
rect 25520 24330 25543 25337
rect 25337 23330 25543 24330
rect 25337 22353 25360 23330
rect 22330 22330 25360 22353
rect 25520 22353 25543 23330
rect 28527 24330 28550 25337
rect 28710 25337 31740 25360
rect 28710 24330 28733 25337
rect 28527 23330 28733 24330
rect 28527 22353 28550 23330
rect 25520 22330 28550 22353
rect 28710 22353 28733 23330
rect 31717 24330 31740 25337
rect 31900 25337 34930 25360
rect 31900 24330 31923 25337
rect 31717 23330 31923 24330
rect 31717 22353 31740 23330
rect 28710 22330 31740 22353
rect 31900 22353 31923 23330
rect 34907 24330 34930 25337
rect 35090 25337 38120 25360
rect 35090 24330 35113 25337
rect 34907 23330 35113 24330
rect 34907 22353 34930 23330
rect 31900 22330 34930 22353
rect 35090 22353 35113 23330
rect 38097 24330 38120 25337
rect 38280 25337 41310 25360
rect 38280 24330 38303 25337
rect 38097 23330 38303 24330
rect 38097 22353 38120 23330
rect 35090 22330 38120 22353
rect 38280 22353 38303 23330
rect 41287 24330 41310 25337
rect 41470 25337 44500 25360
rect 41470 24330 41493 25337
rect 41287 23330 41493 24330
rect 41287 22353 41310 23330
rect 38280 22330 41310 22353
rect 41470 22353 41493 23330
rect 44477 24330 44500 25337
rect 44660 25337 47690 25360
rect 44660 24330 44683 25337
rect 44477 23330 44683 24330
rect 44477 22353 44500 23330
rect 41470 22330 44500 22353
rect 44660 22353 44683 23330
rect 47667 24330 47690 25337
rect 47850 25337 50880 25360
rect 47850 24330 47873 25337
rect 47667 23330 47873 24330
rect 47667 22353 47690 23330
rect 44660 22330 47690 22353
rect 47850 22353 47873 23330
rect 50857 24330 50880 25337
rect 51040 25337 54070 25360
rect 51040 24330 51063 25337
rect 50857 23330 51063 24330
rect 50857 22353 50880 23330
rect 47850 22330 50880 22353
rect 51040 22353 51063 23330
rect 54047 24330 54070 25337
rect 54230 25337 57260 25360
rect 54230 24330 54253 25337
rect 54047 23330 54253 24330
rect 54047 22353 54070 23330
rect 51040 22330 54070 22353
rect 54230 22353 54253 23330
rect 57237 24330 57260 25337
rect 57420 25337 60450 25360
rect 57420 24330 57443 25337
rect 57237 23330 57443 24330
rect 57237 22353 57260 23330
rect 54230 22330 57260 22353
rect 57420 22353 57443 23330
rect 60427 24330 60450 25337
rect 60610 25337 63640 25360
rect 60610 24330 60633 25337
rect 60427 23330 60633 24330
rect 60427 22353 60450 23330
rect 57420 22330 60450 22353
rect 60610 22353 60633 23330
rect 63617 24330 63640 25337
rect 63800 25337 66830 25360
rect 63800 24330 63823 25337
rect 63617 23330 63823 24330
rect 63617 22353 63640 23330
rect 60610 22330 63640 22353
rect 63800 22353 63823 23330
rect 66807 24330 66830 25337
rect 66990 25337 70020 25360
rect 66990 24330 67013 25337
rect 66807 23330 67013 24330
rect 66807 22353 66830 23330
rect 63800 22330 66830 22353
rect 66990 22353 67013 23330
rect 69997 24330 70020 25337
rect 70180 25337 73210 25360
rect 70180 24330 70203 25337
rect 69997 23330 70203 24330
rect 69997 22353 70020 23330
rect 66990 22330 70020 22353
rect 70180 22353 70203 23330
rect 73187 24330 73210 25337
rect 73370 25337 76400 25360
rect 73370 24330 73393 25337
rect 73187 23330 73393 24330
rect 73187 22353 73210 23330
rect 70180 22330 73210 22353
rect 73370 22353 73393 23330
rect 76377 24330 76400 25337
rect 76560 25337 79590 25360
rect 76560 24330 76583 25337
rect 76377 23330 76583 24330
rect 76377 22353 76400 23330
rect 73370 22330 76400 22353
rect 76560 22353 76583 23330
rect 79567 24330 79590 25337
rect 79750 25337 82780 25360
rect 79750 24330 79773 25337
rect 79567 23330 79773 24330
rect 79567 22353 79590 23330
rect 76560 22330 79590 22353
rect 79750 22353 79773 23330
rect 82757 24330 82780 25337
rect 82940 25337 85970 25360
rect 82940 24330 82963 25337
rect 82757 23330 82963 24330
rect 82757 22353 82780 23330
rect 79750 22330 82780 22353
rect 82940 22353 82963 23330
rect 85947 24330 85970 25337
rect 86130 25337 89160 25360
rect 86130 24330 86153 25337
rect 85947 23330 86153 24330
rect 85947 22353 85970 23330
rect 82940 22330 85970 22353
rect 86130 22353 86153 23330
rect 89137 24330 89160 25337
rect 89320 25337 92350 25360
rect 89320 24330 89343 25337
rect 89137 23330 89343 24330
rect 89137 22353 89160 23330
rect 86130 22330 89160 22353
rect 89320 22353 89343 23330
rect 92327 24330 92350 25337
rect 92510 25337 95540 25360
rect 92510 24330 92533 25337
rect 92327 23330 92533 24330
rect 92327 22353 92350 23330
rect 89320 22330 92350 22353
rect 92510 22353 92533 23330
rect 95517 24330 95540 25337
rect 95700 25337 98730 25360
rect 95700 24330 95723 25337
rect 95517 23330 95723 24330
rect 95517 22353 95540 23330
rect 92510 22330 95540 22353
rect 95700 22353 95723 23330
rect 98707 24330 98730 25337
rect 98890 25337 101920 25360
rect 98890 24330 98913 25337
rect 98707 23330 98913 24330
rect 98707 22353 98730 23330
rect 95700 22330 98730 22353
rect 98890 22353 98913 23330
rect 101897 24330 101920 25337
rect 102080 25337 105110 25360
rect 102080 24330 102103 25337
rect 101897 23330 102103 24330
rect 101897 22353 101920 23330
rect 98890 22330 101920 22353
rect 102080 22353 102103 23330
rect 105087 24330 105110 25337
rect 105270 25337 108300 25360
rect 105270 24330 105293 25337
rect 105087 23330 105293 24330
rect 105087 22353 105110 23330
rect 102080 22330 105110 22353
rect 105270 22353 105293 23330
rect 108277 24330 108300 25337
rect 108460 25337 111490 25360
rect 108460 24330 108483 25337
rect 108277 23330 108483 24330
rect 108277 22353 108300 23330
rect 105270 22330 108300 22353
rect 108460 22353 108483 23330
rect 111467 24330 111490 25337
rect 111650 25337 114680 25360
rect 111650 24330 111673 25337
rect 111467 23330 111673 24330
rect 111467 22353 111490 23330
rect 108460 22330 111490 22353
rect 111650 22353 111673 23330
rect 114657 24330 114680 25337
rect 114840 25337 117870 25360
rect 114840 24330 114863 25337
rect 114657 23330 114863 24330
rect 114657 22353 114680 23330
rect 111650 22330 114680 22353
rect 114840 22353 114863 23330
rect 117847 24330 117870 25337
rect 118030 25337 121060 25360
rect 118030 24330 118053 25337
rect 117847 23330 118053 24330
rect 117847 22353 117870 23330
rect 114840 22330 117870 22353
rect 118030 22353 118053 23330
rect 121037 24330 121060 25337
rect 121220 25337 124250 25360
rect 121220 24330 121243 25337
rect 121037 23330 121243 24330
rect 121037 22353 121060 23330
rect 118030 22330 121060 22353
rect 121220 22353 121243 23330
rect 124227 24330 124250 25337
rect 124410 25337 127440 25360
rect 124410 24330 124433 25337
rect 124227 23330 124433 24330
rect 124227 22353 124250 23330
rect 121220 22330 124250 22353
rect 124410 22353 124433 23330
rect 127417 24330 127440 25337
rect 127600 25337 130630 25360
rect 127600 24330 127623 25337
rect 127417 23330 127623 24330
rect 127417 22353 127440 23330
rect 124410 22330 127440 22353
rect 127600 22353 127623 23330
rect 130607 24330 130630 25337
rect 130790 25337 133820 25360
rect 130790 24330 130813 25337
rect 130607 23330 130813 24330
rect 130607 22353 130630 23330
rect 127600 22330 130630 22353
rect 130790 22353 130813 23330
rect 133797 24330 133820 25337
rect 133980 25337 137010 25360
rect 133980 24330 134003 25337
rect 133797 23330 134003 24330
rect 133797 22353 133820 23330
rect 130790 22330 133820 22353
rect 133980 22353 134003 23330
rect 136987 24330 137010 25337
rect 136987 23330 137170 24330
rect 136987 22353 137010 23330
rect 133980 22330 137010 22353
rect 1000 22170 2000 22330
rect 4190 22170 5190 22330
rect 7380 22170 8380 22330
rect 10570 22170 11570 22330
rect 13760 22170 14760 22330
rect 16950 22170 17950 22330
rect 20140 22170 21140 22330
rect 23330 22170 24330 22330
rect 26520 22170 27520 22330
rect 29710 22170 30710 22330
rect 32900 22170 33900 22330
rect 36090 22170 37090 22330
rect 39280 22170 40280 22330
rect 42470 22170 43470 22330
rect 45660 22170 46660 22330
rect 48850 22170 49850 22330
rect 52040 22170 53040 22330
rect 55230 22170 56230 22330
rect 58420 22170 59420 22330
rect 61610 22170 62610 22330
rect 64800 22170 65800 22330
rect 67990 22170 68990 22330
rect 71180 22170 72180 22330
rect 74370 22170 75370 22330
rect 77560 22170 78560 22330
rect 80750 22170 81750 22330
rect 83940 22170 84940 22330
rect 87130 22170 88130 22330
rect 90320 22170 91320 22330
rect 93510 22170 94510 22330
rect 96700 22170 97700 22330
rect 99890 22170 100890 22330
rect 103080 22170 104080 22330
rect 106270 22170 107270 22330
rect 109460 22170 110460 22330
rect 112650 22170 113650 22330
rect 115840 22170 116840 22330
rect 119030 22170 120030 22330
rect 122220 22170 123220 22330
rect 125410 22170 126410 22330
rect 128600 22170 129600 22330
rect 131790 22170 132790 22330
rect 134980 22170 135980 22330
rect 0 22147 3030 22170
rect 0 19163 23 22147
rect 3007 21140 3030 22147
rect 3190 22147 6220 22170
rect 3190 21140 3213 22147
rect 3007 20140 3213 21140
rect 3007 19163 3030 20140
rect 0 19140 3030 19163
rect 3190 19163 3213 20140
rect 6197 21140 6220 22147
rect 6380 22147 9410 22170
rect 6380 21140 6403 22147
rect 6197 20140 6403 21140
rect 6197 19163 6220 20140
rect 3190 19140 6220 19163
rect 6380 19163 6403 20140
rect 9387 21140 9410 22147
rect 9570 22147 12600 22170
rect 9570 21140 9593 22147
rect 9387 20140 9593 21140
rect 9387 19163 9410 20140
rect 6380 19140 9410 19163
rect 9570 19163 9593 20140
rect 12577 21140 12600 22147
rect 12760 22147 15790 22170
rect 12760 21140 12783 22147
rect 12577 20140 12783 21140
rect 12577 19163 12600 20140
rect 9570 19140 12600 19163
rect 12760 19163 12783 20140
rect 15767 21140 15790 22147
rect 15950 22147 18980 22170
rect 15950 21140 15973 22147
rect 15767 20140 15973 21140
rect 15767 19163 15790 20140
rect 12760 19140 15790 19163
rect 15950 19163 15973 20140
rect 18957 21140 18980 22147
rect 19140 22147 22170 22170
rect 19140 21140 19163 22147
rect 18957 20140 19163 21140
rect 18957 19163 18980 20140
rect 15950 19140 18980 19163
rect 19140 19163 19163 20140
rect 22147 21140 22170 22147
rect 22330 22147 25360 22170
rect 22330 21140 22353 22147
rect 22147 20140 22353 21140
rect 22147 19163 22170 20140
rect 19140 19140 22170 19163
rect 22330 19163 22353 20140
rect 25337 21140 25360 22147
rect 25520 22147 28550 22170
rect 25520 21140 25543 22147
rect 25337 20140 25543 21140
rect 25337 19163 25360 20140
rect 22330 19140 25360 19163
rect 25520 19163 25543 20140
rect 28527 21140 28550 22147
rect 28710 22147 31740 22170
rect 28710 21140 28733 22147
rect 28527 20140 28733 21140
rect 28527 19163 28550 20140
rect 25520 19140 28550 19163
rect 28710 19163 28733 20140
rect 31717 21140 31740 22147
rect 31900 22147 34930 22170
rect 31900 21140 31923 22147
rect 31717 20140 31923 21140
rect 31717 19163 31740 20140
rect 28710 19140 31740 19163
rect 31900 19163 31923 20140
rect 34907 21140 34930 22147
rect 35090 22147 38120 22170
rect 35090 21140 35113 22147
rect 34907 20140 35113 21140
rect 34907 19163 34930 20140
rect 31900 19140 34930 19163
rect 35090 19163 35113 20140
rect 38097 21140 38120 22147
rect 38280 22147 41310 22170
rect 38280 21140 38303 22147
rect 38097 20140 38303 21140
rect 38097 19163 38120 20140
rect 35090 19140 38120 19163
rect 38280 19163 38303 20140
rect 41287 21140 41310 22147
rect 41470 22147 44500 22170
rect 41470 21140 41493 22147
rect 41287 20140 41493 21140
rect 41287 19163 41310 20140
rect 38280 19140 41310 19163
rect 41470 19163 41493 20140
rect 44477 21140 44500 22147
rect 44660 22147 47690 22170
rect 44660 21140 44683 22147
rect 44477 20140 44683 21140
rect 44477 19163 44500 20140
rect 41470 19140 44500 19163
rect 44660 19163 44683 20140
rect 47667 21140 47690 22147
rect 47850 22147 50880 22170
rect 47850 21140 47873 22147
rect 47667 20140 47873 21140
rect 47667 19163 47690 20140
rect 44660 19140 47690 19163
rect 47850 19163 47873 20140
rect 50857 21140 50880 22147
rect 51040 22147 54070 22170
rect 51040 21140 51063 22147
rect 50857 20140 51063 21140
rect 50857 19163 50880 20140
rect 47850 19140 50880 19163
rect 51040 19163 51063 20140
rect 54047 21140 54070 22147
rect 54230 22147 57260 22170
rect 54230 21140 54253 22147
rect 54047 20140 54253 21140
rect 54047 19163 54070 20140
rect 51040 19140 54070 19163
rect 54230 19163 54253 20140
rect 57237 21140 57260 22147
rect 57420 22147 60450 22170
rect 57420 21140 57443 22147
rect 57237 20140 57443 21140
rect 57237 19163 57260 20140
rect 54230 19140 57260 19163
rect 57420 19163 57443 20140
rect 60427 21140 60450 22147
rect 60610 22147 63640 22170
rect 60610 21140 60633 22147
rect 60427 20140 60633 21140
rect 60427 19163 60450 20140
rect 57420 19140 60450 19163
rect 60610 19163 60633 20140
rect 63617 21140 63640 22147
rect 63800 22147 66830 22170
rect 63800 21140 63823 22147
rect 63617 20140 63823 21140
rect 63617 19163 63640 20140
rect 60610 19140 63640 19163
rect 63800 19163 63823 20140
rect 66807 21140 66830 22147
rect 66990 22147 70020 22170
rect 66990 21140 67013 22147
rect 66807 20140 67013 21140
rect 66807 19163 66830 20140
rect 63800 19140 66830 19163
rect 66990 19163 67013 20140
rect 69997 21140 70020 22147
rect 70180 22147 73210 22170
rect 70180 21140 70203 22147
rect 69997 20140 70203 21140
rect 69997 19163 70020 20140
rect 66990 19140 70020 19163
rect 70180 19163 70203 20140
rect 73187 21140 73210 22147
rect 73370 22147 76400 22170
rect 73370 21140 73393 22147
rect 73187 20140 73393 21140
rect 73187 19163 73210 20140
rect 70180 19140 73210 19163
rect 73370 19163 73393 20140
rect 76377 21140 76400 22147
rect 76560 22147 79590 22170
rect 76560 21140 76583 22147
rect 76377 20140 76583 21140
rect 76377 19163 76400 20140
rect 73370 19140 76400 19163
rect 76560 19163 76583 20140
rect 79567 21140 79590 22147
rect 79750 22147 82780 22170
rect 79750 21140 79773 22147
rect 79567 20140 79773 21140
rect 79567 19163 79590 20140
rect 76560 19140 79590 19163
rect 79750 19163 79773 20140
rect 82757 21140 82780 22147
rect 82940 22147 85970 22170
rect 82940 21140 82963 22147
rect 82757 20140 82963 21140
rect 82757 19163 82780 20140
rect 79750 19140 82780 19163
rect 82940 19163 82963 20140
rect 85947 21140 85970 22147
rect 86130 22147 89160 22170
rect 86130 21140 86153 22147
rect 85947 20140 86153 21140
rect 85947 19163 85970 20140
rect 82940 19140 85970 19163
rect 86130 19163 86153 20140
rect 89137 21140 89160 22147
rect 89320 22147 92350 22170
rect 89320 21140 89343 22147
rect 89137 20140 89343 21140
rect 89137 19163 89160 20140
rect 86130 19140 89160 19163
rect 89320 19163 89343 20140
rect 92327 21140 92350 22147
rect 92510 22147 95540 22170
rect 92510 21140 92533 22147
rect 92327 20140 92533 21140
rect 92327 19163 92350 20140
rect 89320 19140 92350 19163
rect 92510 19163 92533 20140
rect 95517 21140 95540 22147
rect 95700 22147 98730 22170
rect 95700 21140 95723 22147
rect 95517 20140 95723 21140
rect 95517 19163 95540 20140
rect 92510 19140 95540 19163
rect 95700 19163 95723 20140
rect 98707 21140 98730 22147
rect 98890 22147 101920 22170
rect 98890 21140 98913 22147
rect 98707 20140 98913 21140
rect 98707 19163 98730 20140
rect 95700 19140 98730 19163
rect 98890 19163 98913 20140
rect 101897 21140 101920 22147
rect 102080 22147 105110 22170
rect 102080 21140 102103 22147
rect 101897 20140 102103 21140
rect 101897 19163 101920 20140
rect 98890 19140 101920 19163
rect 102080 19163 102103 20140
rect 105087 21140 105110 22147
rect 105270 22147 108300 22170
rect 105270 21140 105293 22147
rect 105087 20140 105293 21140
rect 105087 19163 105110 20140
rect 102080 19140 105110 19163
rect 105270 19163 105293 20140
rect 108277 21140 108300 22147
rect 108460 22147 111490 22170
rect 108460 21140 108483 22147
rect 108277 20140 108483 21140
rect 108277 19163 108300 20140
rect 105270 19140 108300 19163
rect 108460 19163 108483 20140
rect 111467 21140 111490 22147
rect 111650 22147 114680 22170
rect 111650 21140 111673 22147
rect 111467 20140 111673 21140
rect 111467 19163 111490 20140
rect 108460 19140 111490 19163
rect 111650 19163 111673 20140
rect 114657 21140 114680 22147
rect 114840 22147 117870 22170
rect 114840 21140 114863 22147
rect 114657 20140 114863 21140
rect 114657 19163 114680 20140
rect 111650 19140 114680 19163
rect 114840 19163 114863 20140
rect 117847 21140 117870 22147
rect 118030 22147 121060 22170
rect 118030 21140 118053 22147
rect 117847 20140 118053 21140
rect 117847 19163 117870 20140
rect 114840 19140 117870 19163
rect 118030 19163 118053 20140
rect 121037 21140 121060 22147
rect 121220 22147 124250 22170
rect 121220 21140 121243 22147
rect 121037 20140 121243 21140
rect 121037 19163 121060 20140
rect 118030 19140 121060 19163
rect 121220 19163 121243 20140
rect 124227 21140 124250 22147
rect 124410 22147 127440 22170
rect 124410 21140 124433 22147
rect 124227 20140 124433 21140
rect 124227 19163 124250 20140
rect 121220 19140 124250 19163
rect 124410 19163 124433 20140
rect 127417 21140 127440 22147
rect 127600 22147 130630 22170
rect 127600 21140 127623 22147
rect 127417 20140 127623 21140
rect 127417 19163 127440 20140
rect 124410 19140 127440 19163
rect 127600 19163 127623 20140
rect 130607 21140 130630 22147
rect 130790 22147 133820 22170
rect 130790 21140 130813 22147
rect 130607 20140 130813 21140
rect 130607 19163 130630 20140
rect 127600 19140 130630 19163
rect 130790 19163 130813 20140
rect 133797 21140 133820 22147
rect 133980 22147 137010 22170
rect 133980 21140 134003 22147
rect 133797 20140 134003 21140
rect 133797 19163 133820 20140
rect 130790 19140 133820 19163
rect 133980 19163 134003 20140
rect 136987 21140 137010 22147
rect 136987 20140 137170 21140
rect 136987 19163 137010 20140
rect 133980 19140 137010 19163
rect 1000 18980 2000 19140
rect 4190 18980 5190 19140
rect 7380 18980 8380 19140
rect 10570 18980 11570 19140
rect 13760 18980 14760 19140
rect 16950 18980 17950 19140
rect 20140 18980 21140 19140
rect 23330 18980 24330 19140
rect 26520 18980 27520 19140
rect 29710 18980 30710 19140
rect 32900 18980 33900 19140
rect 36090 18980 37090 19140
rect 39280 18980 40280 19140
rect 42470 18980 43470 19140
rect 45660 18980 46660 19140
rect 48850 18980 49850 19140
rect 52040 18980 53040 19140
rect 55230 18980 56230 19140
rect 58420 18980 59420 19140
rect 61610 18980 62610 19140
rect 64800 18980 65800 19140
rect 67990 18980 68990 19140
rect 71180 18980 72180 19140
rect 74370 18980 75370 19140
rect 77560 18980 78560 19140
rect 80750 18980 81750 19140
rect 83940 18980 84940 19140
rect 87130 18980 88130 19140
rect 90320 18980 91320 19140
rect 93510 18980 94510 19140
rect 96700 18980 97700 19140
rect 99890 18980 100890 19140
rect 103080 18980 104080 19140
rect 106270 18980 107270 19140
rect 109460 18980 110460 19140
rect 112650 18980 113650 19140
rect 115840 18980 116840 19140
rect 119030 18980 120030 19140
rect 122220 18980 123220 19140
rect 125410 18980 126410 19140
rect 128600 18980 129600 19140
rect 131790 18980 132790 19140
rect 134980 18980 135980 19140
rect 0 18957 3030 18980
rect 0 15973 23 18957
rect 3007 17950 3030 18957
rect 3190 18957 6220 18980
rect 3190 17950 3213 18957
rect 3007 16950 3213 17950
rect 3007 15973 3030 16950
rect 0 15950 3030 15973
rect 3190 15973 3213 16950
rect 6197 17950 6220 18957
rect 6380 18957 9410 18980
rect 6380 17950 6403 18957
rect 6197 16950 6403 17950
rect 6197 15973 6220 16950
rect 3190 15950 6220 15973
rect 6380 15973 6403 16950
rect 9387 17950 9410 18957
rect 9570 18957 12600 18980
rect 9570 17950 9593 18957
rect 9387 16950 9593 17950
rect 9387 15973 9410 16950
rect 6380 15950 9410 15973
rect 9570 15973 9593 16950
rect 12577 17950 12600 18957
rect 12760 18957 15790 18980
rect 12760 17950 12783 18957
rect 12577 16950 12783 17950
rect 12577 15973 12600 16950
rect 9570 15950 12600 15973
rect 12760 15973 12783 16950
rect 15767 17950 15790 18957
rect 15950 18957 18980 18980
rect 15950 17950 15973 18957
rect 15767 16950 15973 17950
rect 15767 15973 15790 16950
rect 12760 15950 15790 15973
rect 15950 15973 15973 16950
rect 18957 17950 18980 18957
rect 19140 18957 22170 18980
rect 19140 17950 19163 18957
rect 18957 16950 19163 17950
rect 18957 15973 18980 16950
rect 15950 15950 18980 15973
rect 19140 15973 19163 16950
rect 22147 17950 22170 18957
rect 22330 18957 25360 18980
rect 22330 17950 22353 18957
rect 22147 16950 22353 17950
rect 22147 15973 22170 16950
rect 19140 15950 22170 15973
rect 22330 15973 22353 16950
rect 25337 17950 25360 18957
rect 25520 18957 28550 18980
rect 25520 17950 25543 18957
rect 25337 16950 25543 17950
rect 25337 15973 25360 16950
rect 22330 15950 25360 15973
rect 25520 15973 25543 16950
rect 28527 17950 28550 18957
rect 28710 18957 31740 18980
rect 28710 17950 28733 18957
rect 28527 16950 28733 17950
rect 28527 15973 28550 16950
rect 25520 15950 28550 15973
rect 28710 15973 28733 16950
rect 31717 17950 31740 18957
rect 31900 18957 34930 18980
rect 31900 17950 31923 18957
rect 31717 16950 31923 17950
rect 31717 15973 31740 16950
rect 28710 15950 31740 15973
rect 31900 15973 31923 16950
rect 34907 17950 34930 18957
rect 35090 18957 38120 18980
rect 35090 17950 35113 18957
rect 34907 16950 35113 17950
rect 34907 15973 34930 16950
rect 31900 15950 34930 15973
rect 35090 15973 35113 16950
rect 38097 17950 38120 18957
rect 38280 18957 41310 18980
rect 38280 17950 38303 18957
rect 38097 16950 38303 17950
rect 38097 15973 38120 16950
rect 35090 15950 38120 15973
rect 38280 15973 38303 16950
rect 41287 17950 41310 18957
rect 41470 18957 44500 18980
rect 41470 17950 41493 18957
rect 41287 16950 41493 17950
rect 41287 15973 41310 16950
rect 38280 15950 41310 15973
rect 41470 15973 41493 16950
rect 44477 17950 44500 18957
rect 44660 18957 47690 18980
rect 44660 17950 44683 18957
rect 44477 16950 44683 17950
rect 44477 15973 44500 16950
rect 41470 15950 44500 15973
rect 44660 15973 44683 16950
rect 47667 17950 47690 18957
rect 47850 18957 50880 18980
rect 47850 17950 47873 18957
rect 47667 16950 47873 17950
rect 47667 15973 47690 16950
rect 44660 15950 47690 15973
rect 47850 15973 47873 16950
rect 50857 17950 50880 18957
rect 51040 18957 54070 18980
rect 51040 17950 51063 18957
rect 50857 16950 51063 17950
rect 50857 15973 50880 16950
rect 47850 15950 50880 15973
rect 51040 15973 51063 16950
rect 54047 17950 54070 18957
rect 54230 18957 57260 18980
rect 54230 17950 54253 18957
rect 54047 16950 54253 17950
rect 54047 15973 54070 16950
rect 51040 15950 54070 15973
rect 54230 15973 54253 16950
rect 57237 17950 57260 18957
rect 57420 18957 60450 18980
rect 57420 17950 57443 18957
rect 57237 16950 57443 17950
rect 57237 15973 57260 16950
rect 54230 15950 57260 15973
rect 57420 15973 57443 16950
rect 60427 17950 60450 18957
rect 60610 18957 63640 18980
rect 60610 17950 60633 18957
rect 60427 16950 60633 17950
rect 60427 15973 60450 16950
rect 57420 15950 60450 15973
rect 60610 15973 60633 16950
rect 63617 17950 63640 18957
rect 63800 18957 66830 18980
rect 63800 17950 63823 18957
rect 63617 16950 63823 17950
rect 63617 15973 63640 16950
rect 60610 15950 63640 15973
rect 63800 15973 63823 16950
rect 66807 17950 66830 18957
rect 66990 18957 70020 18980
rect 66990 17950 67013 18957
rect 66807 16950 67013 17950
rect 66807 15973 66830 16950
rect 63800 15950 66830 15973
rect 66990 15973 67013 16950
rect 69997 17950 70020 18957
rect 70180 18957 73210 18980
rect 70180 17950 70203 18957
rect 69997 16950 70203 17950
rect 69997 15973 70020 16950
rect 66990 15950 70020 15973
rect 70180 15973 70203 16950
rect 73187 17950 73210 18957
rect 73370 18957 76400 18980
rect 73370 17950 73393 18957
rect 73187 16950 73393 17950
rect 73187 15973 73210 16950
rect 70180 15950 73210 15973
rect 73370 15973 73393 16950
rect 76377 17950 76400 18957
rect 76560 18957 79590 18980
rect 76560 17950 76583 18957
rect 76377 16950 76583 17950
rect 76377 15973 76400 16950
rect 73370 15950 76400 15973
rect 76560 15973 76583 16950
rect 79567 17950 79590 18957
rect 79750 18957 82780 18980
rect 79750 17950 79773 18957
rect 79567 16950 79773 17950
rect 79567 15973 79590 16950
rect 76560 15950 79590 15973
rect 79750 15973 79773 16950
rect 82757 17950 82780 18957
rect 82940 18957 85970 18980
rect 82940 17950 82963 18957
rect 82757 16950 82963 17950
rect 82757 15973 82780 16950
rect 79750 15950 82780 15973
rect 82940 15973 82963 16950
rect 85947 17950 85970 18957
rect 86130 18957 89160 18980
rect 86130 17950 86153 18957
rect 85947 16950 86153 17950
rect 85947 15973 85970 16950
rect 82940 15950 85970 15973
rect 86130 15973 86153 16950
rect 89137 17950 89160 18957
rect 89320 18957 92350 18980
rect 89320 17950 89343 18957
rect 89137 16950 89343 17950
rect 89137 15973 89160 16950
rect 86130 15950 89160 15973
rect 89320 15973 89343 16950
rect 92327 17950 92350 18957
rect 92510 18957 95540 18980
rect 92510 17950 92533 18957
rect 92327 16950 92533 17950
rect 92327 15973 92350 16950
rect 89320 15950 92350 15973
rect 92510 15973 92533 16950
rect 95517 17950 95540 18957
rect 95700 18957 98730 18980
rect 95700 17950 95723 18957
rect 95517 16950 95723 17950
rect 95517 15973 95540 16950
rect 92510 15950 95540 15973
rect 95700 15973 95723 16950
rect 98707 17950 98730 18957
rect 98890 18957 101920 18980
rect 98890 17950 98913 18957
rect 98707 16950 98913 17950
rect 98707 15973 98730 16950
rect 95700 15950 98730 15973
rect 98890 15973 98913 16950
rect 101897 17950 101920 18957
rect 102080 18957 105110 18980
rect 102080 17950 102103 18957
rect 101897 16950 102103 17950
rect 101897 15973 101920 16950
rect 98890 15950 101920 15973
rect 102080 15973 102103 16950
rect 105087 17950 105110 18957
rect 105270 18957 108300 18980
rect 105270 17950 105293 18957
rect 105087 16950 105293 17950
rect 105087 15973 105110 16950
rect 102080 15950 105110 15973
rect 105270 15973 105293 16950
rect 108277 17950 108300 18957
rect 108460 18957 111490 18980
rect 108460 17950 108483 18957
rect 108277 16950 108483 17950
rect 108277 15973 108300 16950
rect 105270 15950 108300 15973
rect 108460 15973 108483 16950
rect 111467 17950 111490 18957
rect 111650 18957 114680 18980
rect 111650 17950 111673 18957
rect 111467 16950 111673 17950
rect 111467 15973 111490 16950
rect 108460 15950 111490 15973
rect 111650 15973 111673 16950
rect 114657 17950 114680 18957
rect 114840 18957 117870 18980
rect 114840 17950 114863 18957
rect 114657 16950 114863 17950
rect 114657 15973 114680 16950
rect 111650 15950 114680 15973
rect 114840 15973 114863 16950
rect 117847 17950 117870 18957
rect 118030 18957 121060 18980
rect 118030 17950 118053 18957
rect 117847 16950 118053 17950
rect 117847 15973 117870 16950
rect 114840 15950 117870 15973
rect 118030 15973 118053 16950
rect 121037 17950 121060 18957
rect 121220 18957 124250 18980
rect 121220 17950 121243 18957
rect 121037 16950 121243 17950
rect 121037 15973 121060 16950
rect 118030 15950 121060 15973
rect 121220 15973 121243 16950
rect 124227 17950 124250 18957
rect 124410 18957 127440 18980
rect 124410 17950 124433 18957
rect 124227 16950 124433 17950
rect 124227 15973 124250 16950
rect 121220 15950 124250 15973
rect 124410 15973 124433 16950
rect 127417 17950 127440 18957
rect 127600 18957 130630 18980
rect 127600 17950 127623 18957
rect 127417 16950 127623 17950
rect 127417 15973 127440 16950
rect 124410 15950 127440 15973
rect 127600 15973 127623 16950
rect 130607 17950 130630 18957
rect 130790 18957 133820 18980
rect 130790 17950 130813 18957
rect 130607 16950 130813 17950
rect 130607 15973 130630 16950
rect 127600 15950 130630 15973
rect 130790 15973 130813 16950
rect 133797 17950 133820 18957
rect 133980 18957 137010 18980
rect 133980 17950 134003 18957
rect 133797 16950 134003 17950
rect 133797 15973 133820 16950
rect 130790 15950 133820 15973
rect 133980 15973 134003 16950
rect 136987 17950 137010 18957
rect 136987 16950 137170 17950
rect 136987 15973 137010 16950
rect 133980 15950 137010 15973
rect 1000 15790 2000 15950
rect 4190 15790 5190 15950
rect 7380 15790 8380 15950
rect 10570 15790 11570 15950
rect 13760 15790 14760 15950
rect 16950 15790 17950 15950
rect 20140 15790 21140 15950
rect 23330 15790 24330 15950
rect 26520 15790 27520 15950
rect 29710 15790 30710 15950
rect 32900 15790 33900 15950
rect 36090 15790 37090 15950
rect 39280 15790 40280 15950
rect 42470 15790 43470 15950
rect 45660 15790 46660 15950
rect 48850 15790 49850 15950
rect 52040 15790 53040 15950
rect 55230 15790 56230 15950
rect 58420 15790 59420 15950
rect 61610 15790 62610 15950
rect 64800 15790 65800 15950
rect 67990 15790 68990 15950
rect 71180 15790 72180 15950
rect 74370 15790 75370 15950
rect 77560 15790 78560 15950
rect 80750 15790 81750 15950
rect 83940 15790 84940 15950
rect 87130 15790 88130 15950
rect 90320 15790 91320 15950
rect 93510 15790 94510 15950
rect 96700 15790 97700 15950
rect 99890 15790 100890 15950
rect 103080 15790 104080 15950
rect 106270 15790 107270 15950
rect 109460 15790 110460 15950
rect 112650 15790 113650 15950
rect 115840 15790 116840 15950
rect 119030 15790 120030 15950
rect 122220 15790 123220 15950
rect 125410 15790 126410 15950
rect 128600 15790 129600 15950
rect 131790 15790 132790 15950
rect 134980 15790 135980 15950
rect 0 15767 3030 15790
rect 0 12783 23 15767
rect 3007 14760 3030 15767
rect 3190 15767 6220 15790
rect 3190 14760 3213 15767
rect 3007 13760 3213 14760
rect 3007 12783 3030 13760
rect 0 12760 3030 12783
rect 3190 12783 3213 13760
rect 6197 14760 6220 15767
rect 6380 15767 9410 15790
rect 6380 14760 6403 15767
rect 6197 13760 6403 14760
rect 6197 12783 6220 13760
rect 3190 12760 6220 12783
rect 6380 12783 6403 13760
rect 9387 14760 9410 15767
rect 9570 15767 12600 15790
rect 9570 14760 9593 15767
rect 9387 13760 9593 14760
rect 9387 12783 9410 13760
rect 6380 12760 9410 12783
rect 9570 12783 9593 13760
rect 12577 14760 12600 15767
rect 12760 15767 15790 15790
rect 12760 14760 12783 15767
rect 12577 13760 12783 14760
rect 12577 12783 12600 13760
rect 9570 12760 12600 12783
rect 12760 12783 12783 13760
rect 15767 14760 15790 15767
rect 15950 15767 18980 15790
rect 15950 14760 15973 15767
rect 15767 13760 15973 14760
rect 15767 12783 15790 13760
rect 12760 12760 15790 12783
rect 15950 12783 15973 13760
rect 18957 14760 18980 15767
rect 19140 15767 22170 15790
rect 19140 14760 19163 15767
rect 18957 13760 19163 14760
rect 18957 12783 18980 13760
rect 15950 12760 18980 12783
rect 19140 12783 19163 13760
rect 22147 14760 22170 15767
rect 22330 15767 25360 15790
rect 22330 14760 22353 15767
rect 22147 13760 22353 14760
rect 22147 12783 22170 13760
rect 19140 12760 22170 12783
rect 22330 12783 22353 13760
rect 25337 14760 25360 15767
rect 25520 15767 28550 15790
rect 25520 14760 25543 15767
rect 25337 13760 25543 14760
rect 25337 12783 25360 13760
rect 22330 12760 25360 12783
rect 25520 12783 25543 13760
rect 28527 14760 28550 15767
rect 28710 15767 31740 15790
rect 28710 14760 28733 15767
rect 28527 13760 28733 14760
rect 28527 12783 28550 13760
rect 25520 12760 28550 12783
rect 28710 12783 28733 13760
rect 31717 14760 31740 15767
rect 31900 15767 34930 15790
rect 31900 14760 31923 15767
rect 31717 13760 31923 14760
rect 31717 12783 31740 13760
rect 28710 12760 31740 12783
rect 31900 12783 31923 13760
rect 34907 14760 34930 15767
rect 35090 15767 38120 15790
rect 35090 14760 35113 15767
rect 34907 13760 35113 14760
rect 34907 12783 34930 13760
rect 31900 12760 34930 12783
rect 35090 12783 35113 13760
rect 38097 14760 38120 15767
rect 38280 15767 41310 15790
rect 38280 14760 38303 15767
rect 38097 13760 38303 14760
rect 38097 12783 38120 13760
rect 35090 12760 38120 12783
rect 38280 12783 38303 13760
rect 41287 14760 41310 15767
rect 41470 15767 44500 15790
rect 41470 14760 41493 15767
rect 41287 13760 41493 14760
rect 41287 12783 41310 13760
rect 38280 12760 41310 12783
rect 41470 12783 41493 13760
rect 44477 14760 44500 15767
rect 44660 15767 47690 15790
rect 44660 14760 44683 15767
rect 44477 13760 44683 14760
rect 44477 12783 44500 13760
rect 41470 12760 44500 12783
rect 44660 12783 44683 13760
rect 47667 14760 47690 15767
rect 47850 15767 50880 15790
rect 47850 14760 47873 15767
rect 47667 13760 47873 14760
rect 47667 12783 47690 13760
rect 44660 12760 47690 12783
rect 47850 12783 47873 13760
rect 50857 14760 50880 15767
rect 51040 15767 54070 15790
rect 51040 14760 51063 15767
rect 50857 13760 51063 14760
rect 50857 12783 50880 13760
rect 47850 12760 50880 12783
rect 51040 12783 51063 13760
rect 54047 14760 54070 15767
rect 54230 15767 57260 15790
rect 54230 14760 54253 15767
rect 54047 13760 54253 14760
rect 54047 12783 54070 13760
rect 51040 12760 54070 12783
rect 54230 12783 54253 13760
rect 57237 14760 57260 15767
rect 57420 15767 60450 15790
rect 57420 14760 57443 15767
rect 57237 13760 57443 14760
rect 57237 12783 57260 13760
rect 54230 12760 57260 12783
rect 57420 12783 57443 13760
rect 60427 14760 60450 15767
rect 60610 15767 63640 15790
rect 60610 14760 60633 15767
rect 60427 13760 60633 14760
rect 60427 12783 60450 13760
rect 57420 12760 60450 12783
rect 60610 12783 60633 13760
rect 63617 14760 63640 15767
rect 63800 15767 66830 15790
rect 63800 14760 63823 15767
rect 63617 13760 63823 14760
rect 63617 12783 63640 13760
rect 60610 12760 63640 12783
rect 63800 12783 63823 13760
rect 66807 14760 66830 15767
rect 66990 15767 70020 15790
rect 66990 14760 67013 15767
rect 66807 13760 67013 14760
rect 66807 12783 66830 13760
rect 63800 12760 66830 12783
rect 66990 12783 67013 13760
rect 69997 14760 70020 15767
rect 70180 15767 73210 15790
rect 70180 14760 70203 15767
rect 69997 13760 70203 14760
rect 69997 12783 70020 13760
rect 66990 12760 70020 12783
rect 70180 12783 70203 13760
rect 73187 14760 73210 15767
rect 73370 15767 76400 15790
rect 73370 14760 73393 15767
rect 73187 13760 73393 14760
rect 73187 12783 73210 13760
rect 70180 12760 73210 12783
rect 73370 12783 73393 13760
rect 76377 14760 76400 15767
rect 76560 15767 79590 15790
rect 76560 14760 76583 15767
rect 76377 13760 76583 14760
rect 76377 12783 76400 13760
rect 73370 12760 76400 12783
rect 76560 12783 76583 13760
rect 79567 14760 79590 15767
rect 79750 15767 82780 15790
rect 79750 14760 79773 15767
rect 79567 13760 79773 14760
rect 79567 12783 79590 13760
rect 76560 12760 79590 12783
rect 79750 12783 79773 13760
rect 82757 14760 82780 15767
rect 82940 15767 85970 15790
rect 82940 14760 82963 15767
rect 82757 13760 82963 14760
rect 82757 12783 82780 13760
rect 79750 12760 82780 12783
rect 82940 12783 82963 13760
rect 85947 14760 85970 15767
rect 86130 15767 89160 15790
rect 86130 14760 86153 15767
rect 85947 13760 86153 14760
rect 85947 12783 85970 13760
rect 82940 12760 85970 12783
rect 86130 12783 86153 13760
rect 89137 14760 89160 15767
rect 89320 15767 92350 15790
rect 89320 14760 89343 15767
rect 89137 13760 89343 14760
rect 89137 12783 89160 13760
rect 86130 12760 89160 12783
rect 89320 12783 89343 13760
rect 92327 14760 92350 15767
rect 92510 15767 95540 15790
rect 92510 14760 92533 15767
rect 92327 13760 92533 14760
rect 92327 12783 92350 13760
rect 89320 12760 92350 12783
rect 92510 12783 92533 13760
rect 95517 14760 95540 15767
rect 95700 15767 98730 15790
rect 95700 14760 95723 15767
rect 95517 13760 95723 14760
rect 95517 12783 95540 13760
rect 92510 12760 95540 12783
rect 95700 12783 95723 13760
rect 98707 14760 98730 15767
rect 98890 15767 101920 15790
rect 98890 14760 98913 15767
rect 98707 13760 98913 14760
rect 98707 12783 98730 13760
rect 95700 12760 98730 12783
rect 98890 12783 98913 13760
rect 101897 14760 101920 15767
rect 102080 15767 105110 15790
rect 102080 14760 102103 15767
rect 101897 13760 102103 14760
rect 101897 12783 101920 13760
rect 98890 12760 101920 12783
rect 102080 12783 102103 13760
rect 105087 14760 105110 15767
rect 105270 15767 108300 15790
rect 105270 14760 105293 15767
rect 105087 13760 105293 14760
rect 105087 12783 105110 13760
rect 102080 12760 105110 12783
rect 105270 12783 105293 13760
rect 108277 14760 108300 15767
rect 108460 15767 111490 15790
rect 108460 14760 108483 15767
rect 108277 13760 108483 14760
rect 108277 12783 108300 13760
rect 105270 12760 108300 12783
rect 108460 12783 108483 13760
rect 111467 14760 111490 15767
rect 111650 15767 114680 15790
rect 111650 14760 111673 15767
rect 111467 13760 111673 14760
rect 111467 12783 111490 13760
rect 108460 12760 111490 12783
rect 111650 12783 111673 13760
rect 114657 14760 114680 15767
rect 114840 15767 117870 15790
rect 114840 14760 114863 15767
rect 114657 13760 114863 14760
rect 114657 12783 114680 13760
rect 111650 12760 114680 12783
rect 114840 12783 114863 13760
rect 117847 14760 117870 15767
rect 118030 15767 121060 15790
rect 118030 14760 118053 15767
rect 117847 13760 118053 14760
rect 117847 12783 117870 13760
rect 114840 12760 117870 12783
rect 118030 12783 118053 13760
rect 121037 14760 121060 15767
rect 121220 15767 124250 15790
rect 121220 14760 121243 15767
rect 121037 13760 121243 14760
rect 121037 12783 121060 13760
rect 118030 12760 121060 12783
rect 121220 12783 121243 13760
rect 124227 14760 124250 15767
rect 124410 15767 127440 15790
rect 124410 14760 124433 15767
rect 124227 13760 124433 14760
rect 124227 12783 124250 13760
rect 121220 12760 124250 12783
rect 124410 12783 124433 13760
rect 127417 14760 127440 15767
rect 127600 15767 130630 15790
rect 127600 14760 127623 15767
rect 127417 13760 127623 14760
rect 127417 12783 127440 13760
rect 124410 12760 127440 12783
rect 127600 12783 127623 13760
rect 130607 14760 130630 15767
rect 130790 15767 133820 15790
rect 130790 14760 130813 15767
rect 130607 13760 130813 14760
rect 130607 12783 130630 13760
rect 127600 12760 130630 12783
rect 130790 12783 130813 13760
rect 133797 14760 133820 15767
rect 133980 15767 137010 15790
rect 133980 14760 134003 15767
rect 133797 13760 134003 14760
rect 133797 12783 133820 13760
rect 130790 12760 133820 12783
rect 133980 12783 134003 13760
rect 136987 14760 137010 15767
rect 136987 13760 137170 14760
rect 136987 12783 137010 13760
rect 133980 12760 137010 12783
rect 1000 12600 2000 12760
rect 4190 12600 5190 12760
rect 7380 12600 8380 12760
rect 10570 12600 11570 12760
rect 13760 12600 14760 12760
rect 16950 12600 17950 12760
rect 20140 12600 21140 12760
rect 23330 12600 24330 12760
rect 26520 12600 27520 12760
rect 29710 12600 30710 12760
rect 32900 12600 33900 12760
rect 36090 12600 37090 12760
rect 39280 12600 40280 12760
rect 42470 12600 43470 12760
rect 45660 12600 46660 12760
rect 48850 12600 49850 12760
rect 52040 12600 53040 12760
rect 55230 12600 56230 12760
rect 58420 12600 59420 12760
rect 61610 12600 62610 12760
rect 64800 12600 65800 12760
rect 67990 12600 68990 12760
rect 71180 12600 72180 12760
rect 74370 12600 75370 12760
rect 77560 12600 78560 12760
rect 80750 12600 81750 12760
rect 83940 12600 84940 12760
rect 87130 12600 88130 12760
rect 90320 12600 91320 12760
rect 93510 12600 94510 12760
rect 96700 12600 97700 12760
rect 99890 12600 100890 12760
rect 103080 12600 104080 12760
rect 106270 12600 107270 12760
rect 109460 12600 110460 12760
rect 112650 12600 113650 12760
rect 115840 12600 116840 12760
rect 119030 12600 120030 12760
rect 122220 12600 123220 12760
rect 125410 12600 126410 12760
rect 128600 12600 129600 12760
rect 131790 12600 132790 12760
rect 134980 12600 135980 12760
rect 0 12577 3030 12600
rect 0 9593 23 12577
rect 3007 11570 3030 12577
rect 3190 12577 6220 12600
rect 3190 11570 3213 12577
rect 3007 10570 3213 11570
rect 3007 9593 3030 10570
rect 0 9570 3030 9593
rect 3190 9593 3213 10570
rect 6197 11570 6220 12577
rect 6380 12577 9410 12600
rect 6380 11570 6403 12577
rect 6197 10570 6403 11570
rect 6197 9593 6220 10570
rect 3190 9570 6220 9593
rect 6380 9593 6403 10570
rect 9387 11570 9410 12577
rect 9570 12577 12600 12600
rect 9570 11570 9593 12577
rect 9387 10570 9593 11570
rect 9387 9593 9410 10570
rect 6380 9570 9410 9593
rect 9570 9593 9593 10570
rect 12577 11570 12600 12577
rect 12760 12577 15790 12600
rect 12760 11570 12783 12577
rect 12577 10570 12783 11570
rect 12577 9593 12600 10570
rect 9570 9570 12600 9593
rect 12760 9593 12783 10570
rect 15767 11570 15790 12577
rect 15950 12577 18980 12600
rect 15950 11570 15973 12577
rect 15767 10570 15973 11570
rect 15767 9593 15790 10570
rect 12760 9570 15790 9593
rect 15950 9593 15973 10570
rect 18957 11570 18980 12577
rect 19140 12577 22170 12600
rect 19140 11570 19163 12577
rect 18957 10570 19163 11570
rect 18957 9593 18980 10570
rect 15950 9570 18980 9593
rect 19140 9593 19163 10570
rect 22147 11570 22170 12577
rect 22330 12577 25360 12600
rect 22330 11570 22353 12577
rect 22147 10570 22353 11570
rect 22147 9593 22170 10570
rect 19140 9570 22170 9593
rect 22330 9593 22353 10570
rect 25337 11570 25360 12577
rect 25520 12577 28550 12600
rect 25520 11570 25543 12577
rect 25337 10570 25543 11570
rect 25337 9593 25360 10570
rect 22330 9570 25360 9593
rect 25520 9593 25543 10570
rect 28527 11570 28550 12577
rect 28710 12577 31740 12600
rect 28710 11570 28733 12577
rect 28527 10570 28733 11570
rect 28527 9593 28550 10570
rect 25520 9570 28550 9593
rect 28710 9593 28733 10570
rect 31717 11570 31740 12577
rect 31900 12577 34930 12600
rect 31900 11570 31923 12577
rect 31717 10570 31923 11570
rect 31717 9593 31740 10570
rect 28710 9570 31740 9593
rect 31900 9593 31923 10570
rect 34907 11570 34930 12577
rect 35090 12577 38120 12600
rect 35090 11570 35113 12577
rect 34907 10570 35113 11570
rect 34907 9593 34930 10570
rect 31900 9570 34930 9593
rect 35090 9593 35113 10570
rect 38097 11570 38120 12577
rect 38280 12577 41310 12600
rect 38280 11570 38303 12577
rect 38097 10570 38303 11570
rect 38097 9593 38120 10570
rect 35090 9570 38120 9593
rect 38280 9593 38303 10570
rect 41287 11570 41310 12577
rect 41470 12577 44500 12600
rect 41470 11570 41493 12577
rect 41287 10570 41493 11570
rect 41287 9593 41310 10570
rect 38280 9570 41310 9593
rect 41470 9593 41493 10570
rect 44477 11570 44500 12577
rect 44660 12577 47690 12600
rect 44660 11570 44683 12577
rect 44477 10570 44683 11570
rect 44477 9593 44500 10570
rect 41470 9570 44500 9593
rect 44660 9593 44683 10570
rect 47667 11570 47690 12577
rect 47850 12577 50880 12600
rect 47850 11570 47873 12577
rect 47667 10570 47873 11570
rect 47667 9593 47690 10570
rect 44660 9570 47690 9593
rect 47850 9593 47873 10570
rect 50857 11570 50880 12577
rect 51040 12577 54070 12600
rect 51040 11570 51063 12577
rect 50857 10570 51063 11570
rect 50857 9593 50880 10570
rect 47850 9570 50880 9593
rect 51040 9593 51063 10570
rect 54047 11570 54070 12577
rect 54230 12577 57260 12600
rect 54230 11570 54253 12577
rect 54047 10570 54253 11570
rect 54047 9593 54070 10570
rect 51040 9570 54070 9593
rect 54230 9593 54253 10570
rect 57237 11570 57260 12577
rect 57420 12577 60450 12600
rect 57420 11570 57443 12577
rect 57237 10570 57443 11570
rect 57237 9593 57260 10570
rect 54230 9570 57260 9593
rect 57420 9593 57443 10570
rect 60427 11570 60450 12577
rect 60610 12577 63640 12600
rect 60610 11570 60633 12577
rect 60427 10570 60633 11570
rect 60427 9593 60450 10570
rect 57420 9570 60450 9593
rect 60610 9593 60633 10570
rect 63617 11570 63640 12577
rect 63800 12577 66830 12600
rect 63800 11570 63823 12577
rect 63617 10570 63823 11570
rect 63617 9593 63640 10570
rect 60610 9570 63640 9593
rect 63800 9593 63823 10570
rect 66807 11570 66830 12577
rect 66990 12577 70020 12600
rect 66990 11570 67013 12577
rect 66807 10570 67013 11570
rect 66807 9593 66830 10570
rect 63800 9570 66830 9593
rect 66990 9593 67013 10570
rect 69997 11570 70020 12577
rect 70180 12577 73210 12600
rect 70180 11570 70203 12577
rect 69997 10570 70203 11570
rect 69997 9593 70020 10570
rect 66990 9570 70020 9593
rect 70180 9593 70203 10570
rect 73187 11570 73210 12577
rect 73370 12577 76400 12600
rect 73370 11570 73393 12577
rect 73187 10570 73393 11570
rect 73187 9593 73210 10570
rect 70180 9570 73210 9593
rect 73370 9593 73393 10570
rect 76377 11570 76400 12577
rect 76560 12577 79590 12600
rect 76560 11570 76583 12577
rect 76377 10570 76583 11570
rect 76377 9593 76400 10570
rect 73370 9570 76400 9593
rect 76560 9593 76583 10570
rect 79567 11570 79590 12577
rect 79750 12577 82780 12600
rect 79750 11570 79773 12577
rect 79567 10570 79773 11570
rect 79567 9593 79590 10570
rect 76560 9570 79590 9593
rect 79750 9593 79773 10570
rect 82757 11570 82780 12577
rect 82940 12577 85970 12600
rect 82940 11570 82963 12577
rect 82757 10570 82963 11570
rect 82757 9593 82780 10570
rect 79750 9570 82780 9593
rect 82940 9593 82963 10570
rect 85947 11570 85970 12577
rect 86130 12577 89160 12600
rect 86130 11570 86153 12577
rect 85947 10570 86153 11570
rect 85947 9593 85970 10570
rect 82940 9570 85970 9593
rect 86130 9593 86153 10570
rect 89137 11570 89160 12577
rect 89320 12577 92350 12600
rect 89320 11570 89343 12577
rect 89137 10570 89343 11570
rect 89137 9593 89160 10570
rect 86130 9570 89160 9593
rect 89320 9593 89343 10570
rect 92327 11570 92350 12577
rect 92510 12577 95540 12600
rect 92510 11570 92533 12577
rect 92327 10570 92533 11570
rect 92327 9593 92350 10570
rect 89320 9570 92350 9593
rect 92510 9593 92533 10570
rect 95517 11570 95540 12577
rect 95700 12577 98730 12600
rect 95700 11570 95723 12577
rect 95517 10570 95723 11570
rect 95517 9593 95540 10570
rect 92510 9570 95540 9593
rect 95700 9593 95723 10570
rect 98707 11570 98730 12577
rect 98890 12577 101920 12600
rect 98890 11570 98913 12577
rect 98707 10570 98913 11570
rect 98707 9593 98730 10570
rect 95700 9570 98730 9593
rect 98890 9593 98913 10570
rect 101897 11570 101920 12577
rect 102080 12577 105110 12600
rect 102080 11570 102103 12577
rect 101897 10570 102103 11570
rect 101897 9593 101920 10570
rect 98890 9570 101920 9593
rect 102080 9593 102103 10570
rect 105087 11570 105110 12577
rect 105270 12577 108300 12600
rect 105270 11570 105293 12577
rect 105087 10570 105293 11570
rect 105087 9593 105110 10570
rect 102080 9570 105110 9593
rect 105270 9593 105293 10570
rect 108277 11570 108300 12577
rect 108460 12577 111490 12600
rect 108460 11570 108483 12577
rect 108277 10570 108483 11570
rect 108277 9593 108300 10570
rect 105270 9570 108300 9593
rect 108460 9593 108483 10570
rect 111467 11570 111490 12577
rect 111650 12577 114680 12600
rect 111650 11570 111673 12577
rect 111467 10570 111673 11570
rect 111467 9593 111490 10570
rect 108460 9570 111490 9593
rect 111650 9593 111673 10570
rect 114657 11570 114680 12577
rect 114840 12577 117870 12600
rect 114840 11570 114863 12577
rect 114657 10570 114863 11570
rect 114657 9593 114680 10570
rect 111650 9570 114680 9593
rect 114840 9593 114863 10570
rect 117847 11570 117870 12577
rect 118030 12577 121060 12600
rect 118030 11570 118053 12577
rect 117847 10570 118053 11570
rect 117847 9593 117870 10570
rect 114840 9570 117870 9593
rect 118030 9593 118053 10570
rect 121037 11570 121060 12577
rect 121220 12577 124250 12600
rect 121220 11570 121243 12577
rect 121037 10570 121243 11570
rect 121037 9593 121060 10570
rect 118030 9570 121060 9593
rect 121220 9593 121243 10570
rect 124227 11570 124250 12577
rect 124410 12577 127440 12600
rect 124410 11570 124433 12577
rect 124227 10570 124433 11570
rect 124227 9593 124250 10570
rect 121220 9570 124250 9593
rect 124410 9593 124433 10570
rect 127417 11570 127440 12577
rect 127600 12577 130630 12600
rect 127600 11570 127623 12577
rect 127417 10570 127623 11570
rect 127417 9593 127440 10570
rect 124410 9570 127440 9593
rect 127600 9593 127623 10570
rect 130607 11570 130630 12577
rect 130790 12577 133820 12600
rect 130790 11570 130813 12577
rect 130607 10570 130813 11570
rect 130607 9593 130630 10570
rect 127600 9570 130630 9593
rect 130790 9593 130813 10570
rect 133797 11570 133820 12577
rect 133980 12577 137010 12600
rect 133980 11570 134003 12577
rect 133797 10570 134003 11570
rect 133797 9593 133820 10570
rect 130790 9570 133820 9593
rect 133980 9593 134003 10570
rect 136987 11570 137010 12577
rect 136987 10570 137170 11570
rect 136987 9593 137010 10570
rect 133980 9570 137010 9593
rect 1000 9410 2000 9570
rect 4190 9410 5190 9570
rect 7380 9410 8380 9570
rect 10570 9410 11570 9570
rect 13760 9410 14760 9570
rect 16950 9410 17950 9570
rect 20140 9410 21140 9570
rect 23330 9410 24330 9570
rect 26520 9410 27520 9570
rect 29710 9410 30710 9570
rect 32900 9410 33900 9570
rect 36090 9410 37090 9570
rect 39280 9410 40280 9570
rect 42470 9410 43470 9570
rect 45660 9410 46660 9570
rect 48850 9410 49850 9570
rect 52040 9410 53040 9570
rect 55230 9410 56230 9570
rect 58420 9410 59420 9570
rect 61610 9410 62610 9570
rect 64800 9410 65800 9570
rect 67990 9410 68990 9570
rect 71180 9410 72180 9570
rect 74370 9410 75370 9570
rect 77560 9410 78560 9570
rect 80750 9410 81750 9570
rect 83940 9410 84940 9570
rect 87130 9410 88130 9570
rect 90320 9410 91320 9570
rect 93510 9410 94510 9570
rect 96700 9410 97700 9570
rect 99890 9410 100890 9570
rect 103080 9410 104080 9570
rect 106270 9410 107270 9570
rect 109460 9410 110460 9570
rect 112650 9410 113650 9570
rect 115840 9410 116840 9570
rect 119030 9410 120030 9570
rect 122220 9410 123220 9570
rect 125410 9410 126410 9570
rect 128600 9410 129600 9570
rect 131790 9410 132790 9570
rect 134980 9410 135980 9570
rect 0 9387 3030 9410
rect 0 6403 23 9387
rect 3007 8380 3030 9387
rect 3190 9387 6220 9410
rect 3190 8380 3213 9387
rect 3007 7380 3213 8380
rect 3007 6403 3030 7380
rect 0 6380 3030 6403
rect 3190 6403 3213 7380
rect 6197 8380 6220 9387
rect 6380 9387 9410 9410
rect 6380 8380 6403 9387
rect 6197 7380 6403 8380
rect 6197 6403 6220 7380
rect 3190 6380 6220 6403
rect 6380 6403 6403 7380
rect 9387 8380 9410 9387
rect 9570 9387 12600 9410
rect 9570 8380 9593 9387
rect 9387 7380 9593 8380
rect 9387 6403 9410 7380
rect 6380 6380 9410 6403
rect 9570 6403 9593 7380
rect 12577 8380 12600 9387
rect 12760 9387 15790 9410
rect 12760 8380 12783 9387
rect 12577 7380 12783 8380
rect 12577 6403 12600 7380
rect 9570 6380 12600 6403
rect 12760 6403 12783 7380
rect 15767 8380 15790 9387
rect 15950 9387 18980 9410
rect 15950 8380 15973 9387
rect 15767 7380 15973 8380
rect 15767 6403 15790 7380
rect 12760 6380 15790 6403
rect 15950 6403 15973 7380
rect 18957 8380 18980 9387
rect 19140 9387 22170 9410
rect 19140 8380 19163 9387
rect 18957 7380 19163 8380
rect 18957 6403 18980 7380
rect 15950 6380 18980 6403
rect 19140 6403 19163 7380
rect 22147 8380 22170 9387
rect 22330 9387 25360 9410
rect 22330 8380 22353 9387
rect 22147 7380 22353 8380
rect 22147 6403 22170 7380
rect 19140 6380 22170 6403
rect 22330 6403 22353 7380
rect 25337 8380 25360 9387
rect 25520 9387 28550 9410
rect 25520 8380 25543 9387
rect 25337 7380 25543 8380
rect 25337 6403 25360 7380
rect 22330 6380 25360 6403
rect 25520 6403 25543 7380
rect 28527 8380 28550 9387
rect 28710 9387 31740 9410
rect 28710 8380 28733 9387
rect 28527 7380 28733 8380
rect 28527 6403 28550 7380
rect 25520 6380 28550 6403
rect 28710 6403 28733 7380
rect 31717 8380 31740 9387
rect 31900 9387 34930 9410
rect 31900 8380 31923 9387
rect 31717 7380 31923 8380
rect 31717 6403 31740 7380
rect 28710 6380 31740 6403
rect 31900 6403 31923 7380
rect 34907 8380 34930 9387
rect 35090 9387 38120 9410
rect 35090 8380 35113 9387
rect 34907 7380 35113 8380
rect 34907 6403 34930 7380
rect 31900 6380 34930 6403
rect 35090 6403 35113 7380
rect 38097 8380 38120 9387
rect 38280 9387 41310 9410
rect 38280 8380 38303 9387
rect 38097 7380 38303 8380
rect 38097 6403 38120 7380
rect 35090 6380 38120 6403
rect 38280 6403 38303 7380
rect 41287 8380 41310 9387
rect 41470 9387 44500 9410
rect 41470 8380 41493 9387
rect 41287 7380 41493 8380
rect 41287 6403 41310 7380
rect 38280 6380 41310 6403
rect 41470 6403 41493 7380
rect 44477 8380 44500 9387
rect 44660 9387 47690 9410
rect 44660 8380 44683 9387
rect 44477 7380 44683 8380
rect 44477 6403 44500 7380
rect 41470 6380 44500 6403
rect 44660 6403 44683 7380
rect 47667 8380 47690 9387
rect 47850 9387 50880 9410
rect 47850 8380 47873 9387
rect 47667 7380 47873 8380
rect 47667 6403 47690 7380
rect 44660 6380 47690 6403
rect 47850 6403 47873 7380
rect 50857 8380 50880 9387
rect 51040 9387 54070 9410
rect 51040 8380 51063 9387
rect 50857 7380 51063 8380
rect 50857 6403 50880 7380
rect 47850 6380 50880 6403
rect 51040 6403 51063 7380
rect 54047 8380 54070 9387
rect 54230 9387 57260 9410
rect 54230 8380 54253 9387
rect 54047 7380 54253 8380
rect 54047 6403 54070 7380
rect 51040 6380 54070 6403
rect 54230 6403 54253 7380
rect 57237 8380 57260 9387
rect 57420 9387 60450 9410
rect 57420 8380 57443 9387
rect 57237 7380 57443 8380
rect 57237 6403 57260 7380
rect 54230 6380 57260 6403
rect 57420 6403 57443 7380
rect 60427 8380 60450 9387
rect 60610 9387 63640 9410
rect 60610 8380 60633 9387
rect 60427 7380 60633 8380
rect 60427 6403 60450 7380
rect 57420 6380 60450 6403
rect 60610 6403 60633 7380
rect 63617 8380 63640 9387
rect 63800 9387 66830 9410
rect 63800 8380 63823 9387
rect 63617 7380 63823 8380
rect 63617 6403 63640 7380
rect 60610 6380 63640 6403
rect 63800 6403 63823 7380
rect 66807 8380 66830 9387
rect 66990 9387 70020 9410
rect 66990 8380 67013 9387
rect 66807 7380 67013 8380
rect 66807 6403 66830 7380
rect 63800 6380 66830 6403
rect 66990 6403 67013 7380
rect 69997 8380 70020 9387
rect 70180 9387 73210 9410
rect 70180 8380 70203 9387
rect 69997 7380 70203 8380
rect 69997 6403 70020 7380
rect 66990 6380 70020 6403
rect 70180 6403 70203 7380
rect 73187 8380 73210 9387
rect 73370 9387 76400 9410
rect 73370 8380 73393 9387
rect 73187 7380 73393 8380
rect 73187 6403 73210 7380
rect 70180 6380 73210 6403
rect 73370 6403 73393 7380
rect 76377 8380 76400 9387
rect 76560 9387 79590 9410
rect 76560 8380 76583 9387
rect 76377 7380 76583 8380
rect 76377 6403 76400 7380
rect 73370 6380 76400 6403
rect 76560 6403 76583 7380
rect 79567 8380 79590 9387
rect 79750 9387 82780 9410
rect 79750 8380 79773 9387
rect 79567 7380 79773 8380
rect 79567 6403 79590 7380
rect 76560 6380 79590 6403
rect 79750 6403 79773 7380
rect 82757 8380 82780 9387
rect 82940 9387 85970 9410
rect 82940 8380 82963 9387
rect 82757 7380 82963 8380
rect 82757 6403 82780 7380
rect 79750 6380 82780 6403
rect 82940 6403 82963 7380
rect 85947 8380 85970 9387
rect 86130 9387 89160 9410
rect 86130 8380 86153 9387
rect 85947 7380 86153 8380
rect 85947 6403 85970 7380
rect 82940 6380 85970 6403
rect 86130 6403 86153 7380
rect 89137 8380 89160 9387
rect 89320 9387 92350 9410
rect 89320 8380 89343 9387
rect 89137 7380 89343 8380
rect 89137 6403 89160 7380
rect 86130 6380 89160 6403
rect 89320 6403 89343 7380
rect 92327 8380 92350 9387
rect 92510 9387 95540 9410
rect 92510 8380 92533 9387
rect 92327 7380 92533 8380
rect 92327 6403 92350 7380
rect 89320 6380 92350 6403
rect 92510 6403 92533 7380
rect 95517 8380 95540 9387
rect 95700 9387 98730 9410
rect 95700 8380 95723 9387
rect 95517 7380 95723 8380
rect 95517 6403 95540 7380
rect 92510 6380 95540 6403
rect 95700 6403 95723 7380
rect 98707 8380 98730 9387
rect 98890 9387 101920 9410
rect 98890 8380 98913 9387
rect 98707 7380 98913 8380
rect 98707 6403 98730 7380
rect 95700 6380 98730 6403
rect 98890 6403 98913 7380
rect 101897 8380 101920 9387
rect 102080 9387 105110 9410
rect 102080 8380 102103 9387
rect 101897 7380 102103 8380
rect 101897 6403 101920 7380
rect 98890 6380 101920 6403
rect 102080 6403 102103 7380
rect 105087 8380 105110 9387
rect 105270 9387 108300 9410
rect 105270 8380 105293 9387
rect 105087 7380 105293 8380
rect 105087 6403 105110 7380
rect 102080 6380 105110 6403
rect 105270 6403 105293 7380
rect 108277 8380 108300 9387
rect 108460 9387 111490 9410
rect 108460 8380 108483 9387
rect 108277 7380 108483 8380
rect 108277 6403 108300 7380
rect 105270 6380 108300 6403
rect 108460 6403 108483 7380
rect 111467 8380 111490 9387
rect 111650 9387 114680 9410
rect 111650 8380 111673 9387
rect 111467 7380 111673 8380
rect 111467 6403 111490 7380
rect 108460 6380 111490 6403
rect 111650 6403 111673 7380
rect 114657 8380 114680 9387
rect 114840 9387 117870 9410
rect 114840 8380 114863 9387
rect 114657 7380 114863 8380
rect 114657 6403 114680 7380
rect 111650 6380 114680 6403
rect 114840 6403 114863 7380
rect 117847 8380 117870 9387
rect 118030 9387 121060 9410
rect 118030 8380 118053 9387
rect 117847 7380 118053 8380
rect 117847 6403 117870 7380
rect 114840 6380 117870 6403
rect 118030 6403 118053 7380
rect 121037 8380 121060 9387
rect 121220 9387 124250 9410
rect 121220 8380 121243 9387
rect 121037 7380 121243 8380
rect 121037 6403 121060 7380
rect 118030 6380 121060 6403
rect 121220 6403 121243 7380
rect 124227 8380 124250 9387
rect 124410 9387 127440 9410
rect 124410 8380 124433 9387
rect 124227 7380 124433 8380
rect 124227 6403 124250 7380
rect 121220 6380 124250 6403
rect 124410 6403 124433 7380
rect 127417 8380 127440 9387
rect 127600 9387 130630 9410
rect 127600 8380 127623 9387
rect 127417 7380 127623 8380
rect 127417 6403 127440 7380
rect 124410 6380 127440 6403
rect 127600 6403 127623 7380
rect 130607 8380 130630 9387
rect 130790 9387 133820 9410
rect 130790 8380 130813 9387
rect 130607 7380 130813 8380
rect 130607 6403 130630 7380
rect 127600 6380 130630 6403
rect 130790 6403 130813 7380
rect 133797 8380 133820 9387
rect 133980 9387 137010 9410
rect 133980 8380 134003 9387
rect 133797 7380 134003 8380
rect 133797 6403 133820 7380
rect 130790 6380 133820 6403
rect 133980 6403 134003 7380
rect 136987 8380 137010 9387
rect 136987 7380 137170 8380
rect 136987 6403 137010 7380
rect 133980 6380 137010 6403
rect 1000 6220 2000 6380
rect 4190 6220 5190 6380
rect 7380 6220 8380 6380
rect 10570 6220 11570 6380
rect 13760 6220 14760 6380
rect 16950 6220 17950 6380
rect 20140 6220 21140 6380
rect 23330 6220 24330 6380
rect 26520 6220 27520 6380
rect 29710 6220 30710 6380
rect 32900 6220 33900 6380
rect 36090 6220 37090 6380
rect 39280 6220 40280 6380
rect 42470 6220 43470 6380
rect 45660 6220 46660 6380
rect 48850 6220 49850 6380
rect 52040 6220 53040 6380
rect 55230 6220 56230 6380
rect 58420 6220 59420 6380
rect 61610 6220 62610 6380
rect 64800 6220 65800 6380
rect 67990 6220 68990 6380
rect 71180 6220 72180 6380
rect 74370 6220 75370 6380
rect 77560 6220 78560 6380
rect 80750 6220 81750 6380
rect 83940 6220 84940 6380
rect 87130 6220 88130 6380
rect 90320 6220 91320 6380
rect 93510 6220 94510 6380
rect 96700 6220 97700 6380
rect 99890 6220 100890 6380
rect 103080 6220 104080 6380
rect 106270 6220 107270 6380
rect 109460 6220 110460 6380
rect 112650 6220 113650 6380
rect 115840 6220 116840 6380
rect 119030 6220 120030 6380
rect 122220 6220 123220 6380
rect 125410 6220 126410 6380
rect 128600 6220 129600 6380
rect 131790 6220 132790 6380
rect 134980 6220 135980 6380
rect 0 6197 3030 6220
rect 0 3213 23 6197
rect 3007 5190 3030 6197
rect 3190 6197 6220 6220
rect 3190 5190 3213 6197
rect 3007 4190 3213 5190
rect 3007 3213 3030 4190
rect 0 3190 3030 3213
rect 3190 3213 3213 4190
rect 6197 5190 6220 6197
rect 6380 6197 9410 6220
rect 6380 5190 6403 6197
rect 6197 4190 6403 5190
rect 6197 3213 6220 4190
rect 3190 3190 6220 3213
rect 6380 3213 6403 4190
rect 9387 5190 9410 6197
rect 9570 6197 12600 6220
rect 9570 5190 9593 6197
rect 9387 4190 9593 5190
rect 9387 3213 9410 4190
rect 6380 3190 9410 3213
rect 9570 3213 9593 4190
rect 12577 5190 12600 6197
rect 12760 6197 15790 6220
rect 12760 5190 12783 6197
rect 12577 4190 12783 5190
rect 12577 3213 12600 4190
rect 9570 3190 12600 3213
rect 12760 3213 12783 4190
rect 15767 5190 15790 6197
rect 15950 6197 18980 6220
rect 15950 5190 15973 6197
rect 15767 4190 15973 5190
rect 15767 3213 15790 4190
rect 12760 3190 15790 3213
rect 15950 3213 15973 4190
rect 18957 5190 18980 6197
rect 19140 6197 22170 6220
rect 19140 5190 19163 6197
rect 18957 4190 19163 5190
rect 18957 3213 18980 4190
rect 15950 3190 18980 3213
rect 19140 3213 19163 4190
rect 22147 5190 22170 6197
rect 22330 6197 25360 6220
rect 22330 5190 22353 6197
rect 22147 4190 22353 5190
rect 22147 3213 22170 4190
rect 19140 3190 22170 3213
rect 22330 3213 22353 4190
rect 25337 5190 25360 6197
rect 25520 6197 28550 6220
rect 25520 5190 25543 6197
rect 25337 4190 25543 5190
rect 25337 3213 25360 4190
rect 22330 3190 25360 3213
rect 25520 3213 25543 4190
rect 28527 5190 28550 6197
rect 28710 6197 31740 6220
rect 28710 5190 28733 6197
rect 28527 4190 28733 5190
rect 28527 3213 28550 4190
rect 25520 3190 28550 3213
rect 28710 3213 28733 4190
rect 31717 5190 31740 6197
rect 31900 6197 34930 6220
rect 31900 5190 31923 6197
rect 31717 4190 31923 5190
rect 31717 3213 31740 4190
rect 28710 3190 31740 3213
rect 31900 3213 31923 4190
rect 34907 5190 34930 6197
rect 35090 6197 38120 6220
rect 35090 5190 35113 6197
rect 34907 4190 35113 5190
rect 34907 3213 34930 4190
rect 31900 3190 34930 3213
rect 35090 3213 35113 4190
rect 38097 5190 38120 6197
rect 38280 6197 41310 6220
rect 38280 5190 38303 6197
rect 38097 4190 38303 5190
rect 38097 3213 38120 4190
rect 35090 3190 38120 3213
rect 38280 3213 38303 4190
rect 41287 5190 41310 6197
rect 41470 6197 44500 6220
rect 41470 5190 41493 6197
rect 41287 4190 41493 5190
rect 41287 3213 41310 4190
rect 38280 3190 41310 3213
rect 41470 3213 41493 4190
rect 44477 5190 44500 6197
rect 44660 6197 47690 6220
rect 44660 5190 44683 6197
rect 44477 4190 44683 5190
rect 44477 3213 44500 4190
rect 41470 3190 44500 3213
rect 44660 3213 44683 4190
rect 47667 5190 47690 6197
rect 47850 6197 50880 6220
rect 47850 5190 47873 6197
rect 47667 4190 47873 5190
rect 47667 3213 47690 4190
rect 44660 3190 47690 3213
rect 47850 3213 47873 4190
rect 50857 5190 50880 6197
rect 51040 6197 54070 6220
rect 51040 5190 51063 6197
rect 50857 4190 51063 5190
rect 50857 3213 50880 4190
rect 47850 3190 50880 3213
rect 51040 3213 51063 4190
rect 54047 5190 54070 6197
rect 54230 6197 57260 6220
rect 54230 5190 54253 6197
rect 54047 4190 54253 5190
rect 54047 3213 54070 4190
rect 51040 3190 54070 3213
rect 54230 3213 54253 4190
rect 57237 5190 57260 6197
rect 57420 6197 60450 6220
rect 57420 5190 57443 6197
rect 57237 4190 57443 5190
rect 57237 3213 57260 4190
rect 54230 3190 57260 3213
rect 57420 3213 57443 4190
rect 60427 5190 60450 6197
rect 60610 6197 63640 6220
rect 60610 5190 60633 6197
rect 60427 4190 60633 5190
rect 60427 3213 60450 4190
rect 57420 3190 60450 3213
rect 60610 3213 60633 4190
rect 63617 5190 63640 6197
rect 63800 6197 66830 6220
rect 63800 5190 63823 6197
rect 63617 4190 63823 5190
rect 63617 3213 63640 4190
rect 60610 3190 63640 3213
rect 63800 3213 63823 4190
rect 66807 5190 66830 6197
rect 66990 6197 70020 6220
rect 66990 5190 67013 6197
rect 66807 4190 67013 5190
rect 66807 3213 66830 4190
rect 63800 3190 66830 3213
rect 66990 3213 67013 4190
rect 69997 5190 70020 6197
rect 70180 6197 73210 6220
rect 70180 5190 70203 6197
rect 69997 4190 70203 5190
rect 69997 3213 70020 4190
rect 66990 3190 70020 3213
rect 70180 3213 70203 4190
rect 73187 5190 73210 6197
rect 73370 6197 76400 6220
rect 73370 5190 73393 6197
rect 73187 4190 73393 5190
rect 73187 3213 73210 4190
rect 70180 3190 73210 3213
rect 73370 3213 73393 4190
rect 76377 5190 76400 6197
rect 76560 6197 79590 6220
rect 76560 5190 76583 6197
rect 76377 4190 76583 5190
rect 76377 3213 76400 4190
rect 73370 3190 76400 3213
rect 76560 3213 76583 4190
rect 79567 5190 79590 6197
rect 79750 6197 82780 6220
rect 79750 5190 79773 6197
rect 79567 4190 79773 5190
rect 79567 3213 79590 4190
rect 76560 3190 79590 3213
rect 79750 3213 79773 4190
rect 82757 5190 82780 6197
rect 82940 6197 85970 6220
rect 82940 5190 82963 6197
rect 82757 4190 82963 5190
rect 82757 3213 82780 4190
rect 79750 3190 82780 3213
rect 82940 3213 82963 4190
rect 85947 5190 85970 6197
rect 86130 6197 89160 6220
rect 86130 5190 86153 6197
rect 85947 4190 86153 5190
rect 85947 3213 85970 4190
rect 82940 3190 85970 3213
rect 86130 3213 86153 4190
rect 89137 5190 89160 6197
rect 89320 6197 92350 6220
rect 89320 5190 89343 6197
rect 89137 4190 89343 5190
rect 89137 3213 89160 4190
rect 86130 3190 89160 3213
rect 89320 3213 89343 4190
rect 92327 5190 92350 6197
rect 92510 6197 95540 6220
rect 92510 5190 92533 6197
rect 92327 4190 92533 5190
rect 92327 3213 92350 4190
rect 89320 3190 92350 3213
rect 92510 3213 92533 4190
rect 95517 5190 95540 6197
rect 95700 6197 98730 6220
rect 95700 5190 95723 6197
rect 95517 4190 95723 5190
rect 95517 3213 95540 4190
rect 92510 3190 95540 3213
rect 95700 3213 95723 4190
rect 98707 5190 98730 6197
rect 98890 6197 101920 6220
rect 98890 5190 98913 6197
rect 98707 4190 98913 5190
rect 98707 3213 98730 4190
rect 95700 3190 98730 3213
rect 98890 3213 98913 4190
rect 101897 5190 101920 6197
rect 102080 6197 105110 6220
rect 102080 5190 102103 6197
rect 101897 4190 102103 5190
rect 101897 3213 101920 4190
rect 98890 3190 101920 3213
rect 102080 3213 102103 4190
rect 105087 5190 105110 6197
rect 105270 6197 108300 6220
rect 105270 5190 105293 6197
rect 105087 4190 105293 5190
rect 105087 3213 105110 4190
rect 102080 3190 105110 3213
rect 105270 3213 105293 4190
rect 108277 5190 108300 6197
rect 108460 6197 111490 6220
rect 108460 5190 108483 6197
rect 108277 4190 108483 5190
rect 108277 3213 108300 4190
rect 105270 3190 108300 3213
rect 108460 3213 108483 4190
rect 111467 5190 111490 6197
rect 111650 6197 114680 6220
rect 111650 5190 111673 6197
rect 111467 4190 111673 5190
rect 111467 3213 111490 4190
rect 108460 3190 111490 3213
rect 111650 3213 111673 4190
rect 114657 5190 114680 6197
rect 114840 6197 117870 6220
rect 114840 5190 114863 6197
rect 114657 4190 114863 5190
rect 114657 3213 114680 4190
rect 111650 3190 114680 3213
rect 114840 3213 114863 4190
rect 117847 5190 117870 6197
rect 118030 6197 121060 6220
rect 118030 5190 118053 6197
rect 117847 4190 118053 5190
rect 117847 3213 117870 4190
rect 114840 3190 117870 3213
rect 118030 3213 118053 4190
rect 121037 5190 121060 6197
rect 121220 6197 124250 6220
rect 121220 5190 121243 6197
rect 121037 4190 121243 5190
rect 121037 3213 121060 4190
rect 118030 3190 121060 3213
rect 121220 3213 121243 4190
rect 124227 5190 124250 6197
rect 124410 6197 127440 6220
rect 124410 5190 124433 6197
rect 124227 4190 124433 5190
rect 124227 3213 124250 4190
rect 121220 3190 124250 3213
rect 124410 3213 124433 4190
rect 127417 5190 127440 6197
rect 127600 6197 130630 6220
rect 127600 5190 127623 6197
rect 127417 4190 127623 5190
rect 127417 3213 127440 4190
rect 124410 3190 127440 3213
rect 127600 3213 127623 4190
rect 130607 5190 130630 6197
rect 130790 6197 133820 6220
rect 130790 5190 130813 6197
rect 130607 4190 130813 5190
rect 130607 3213 130630 4190
rect 127600 3190 130630 3213
rect 130790 3213 130813 4190
rect 133797 5190 133820 6197
rect 133980 6197 137010 6220
rect 133980 5190 134003 6197
rect 133797 4190 134003 5190
rect 133797 3213 133820 4190
rect 130790 3190 133820 3213
rect 133980 3213 134003 4190
rect 136987 5190 137010 6197
rect 136987 4190 137170 5190
rect 136987 3213 137010 4190
rect 133980 3190 137010 3213
rect 1000 3030 2000 3190
rect 4190 3030 5190 3190
rect 7380 3030 8380 3190
rect 10570 3030 11570 3190
rect 13760 3030 14760 3190
rect 16950 3030 17950 3190
rect 20140 3030 21140 3190
rect 23330 3030 24330 3190
rect 26520 3030 27520 3190
rect 29710 3030 30710 3190
rect 32900 3030 33900 3190
rect 36090 3030 37090 3190
rect 39280 3030 40280 3190
rect 42470 3030 43470 3190
rect 45660 3030 46660 3190
rect 48850 3030 49850 3190
rect 52040 3030 53040 3190
rect 55230 3030 56230 3190
rect 58420 3030 59420 3190
rect 61610 3030 62610 3190
rect 64800 3030 65800 3190
rect 67990 3030 68990 3190
rect 71180 3030 72180 3190
rect 74370 3030 75370 3190
rect 77560 3030 78560 3190
rect 80750 3030 81750 3190
rect 83940 3030 84940 3190
rect 87130 3030 88130 3190
rect 90320 3030 91320 3190
rect 93510 3030 94510 3190
rect 96700 3030 97700 3190
rect 99890 3030 100890 3190
rect 103080 3030 104080 3190
rect 106270 3030 107270 3190
rect 109460 3030 110460 3190
rect 112650 3030 113650 3190
rect 115840 3030 116840 3190
rect 119030 3030 120030 3190
rect 122220 3030 123220 3190
rect 125410 3030 126410 3190
rect 128600 3030 129600 3190
rect 131790 3030 132790 3190
rect 134980 3030 135980 3190
rect 0 3007 3030 3030
rect 0 23 23 3007
rect 3007 2000 3030 3007
rect 3190 3007 6220 3030
rect 3190 2000 3213 3007
rect 3007 1000 3213 2000
rect 3007 23 3030 1000
rect 0 0 3030 23
rect 3190 23 3213 1000
rect 6197 2000 6220 3007
rect 6380 3007 9410 3030
rect 6380 2000 6403 3007
rect 6197 1000 6403 2000
rect 6197 23 6220 1000
rect 3190 0 6220 23
rect 6380 23 6403 1000
rect 9387 2000 9410 3007
rect 9570 3007 12600 3030
rect 9570 2000 9593 3007
rect 9387 1000 9593 2000
rect 9387 23 9410 1000
rect 6380 0 9410 23
rect 9570 23 9593 1000
rect 12577 2000 12600 3007
rect 12760 3007 15790 3030
rect 12760 2000 12783 3007
rect 12577 1000 12783 2000
rect 12577 23 12600 1000
rect 9570 0 12600 23
rect 12760 23 12783 1000
rect 15767 2000 15790 3007
rect 15950 3007 18980 3030
rect 15950 2000 15973 3007
rect 15767 1000 15973 2000
rect 15767 23 15790 1000
rect 12760 0 15790 23
rect 15950 23 15973 1000
rect 18957 2000 18980 3007
rect 19140 3007 22170 3030
rect 19140 2000 19163 3007
rect 18957 1000 19163 2000
rect 18957 23 18980 1000
rect 15950 0 18980 23
rect 19140 23 19163 1000
rect 22147 2000 22170 3007
rect 22330 3007 25360 3030
rect 22330 2000 22353 3007
rect 22147 1000 22353 2000
rect 22147 23 22170 1000
rect 19140 0 22170 23
rect 22330 23 22353 1000
rect 25337 2000 25360 3007
rect 25520 3007 28550 3030
rect 25520 2000 25543 3007
rect 25337 1000 25543 2000
rect 25337 23 25360 1000
rect 22330 0 25360 23
rect 25520 23 25543 1000
rect 28527 2000 28550 3007
rect 28710 3007 31740 3030
rect 28710 2000 28733 3007
rect 28527 1000 28733 2000
rect 28527 23 28550 1000
rect 25520 0 28550 23
rect 28710 23 28733 1000
rect 31717 2000 31740 3007
rect 31900 3007 34930 3030
rect 31900 2000 31923 3007
rect 31717 1000 31923 2000
rect 31717 23 31740 1000
rect 28710 0 31740 23
rect 31900 23 31923 1000
rect 34907 2000 34930 3007
rect 35090 3007 38120 3030
rect 35090 2000 35113 3007
rect 34907 1000 35113 2000
rect 34907 23 34930 1000
rect 31900 0 34930 23
rect 35090 23 35113 1000
rect 38097 2000 38120 3007
rect 38280 3007 41310 3030
rect 38280 2000 38303 3007
rect 38097 1000 38303 2000
rect 38097 23 38120 1000
rect 35090 0 38120 23
rect 38280 23 38303 1000
rect 41287 2000 41310 3007
rect 41470 3007 44500 3030
rect 41470 2000 41493 3007
rect 41287 1000 41493 2000
rect 41287 23 41310 1000
rect 38280 0 41310 23
rect 41470 23 41493 1000
rect 44477 2000 44500 3007
rect 44660 3007 47690 3030
rect 44660 2000 44683 3007
rect 44477 1000 44683 2000
rect 44477 23 44500 1000
rect 41470 0 44500 23
rect 44660 23 44683 1000
rect 47667 2000 47690 3007
rect 47850 3007 50880 3030
rect 47850 2000 47873 3007
rect 47667 1000 47873 2000
rect 47667 23 47690 1000
rect 44660 0 47690 23
rect 47850 23 47873 1000
rect 50857 2000 50880 3007
rect 51040 3007 54070 3030
rect 51040 2000 51063 3007
rect 50857 1000 51063 2000
rect 50857 23 50880 1000
rect 47850 0 50880 23
rect 51040 23 51063 1000
rect 54047 2000 54070 3007
rect 54230 3007 57260 3030
rect 54230 2000 54253 3007
rect 54047 1000 54253 2000
rect 54047 23 54070 1000
rect 51040 0 54070 23
rect 54230 23 54253 1000
rect 57237 2000 57260 3007
rect 57420 3007 60450 3030
rect 57420 2000 57443 3007
rect 57237 1000 57443 2000
rect 57237 23 57260 1000
rect 54230 0 57260 23
rect 57420 23 57443 1000
rect 60427 2000 60450 3007
rect 60610 3007 63640 3030
rect 60610 2000 60633 3007
rect 60427 1000 60633 2000
rect 60427 23 60450 1000
rect 57420 0 60450 23
rect 60610 23 60633 1000
rect 63617 2000 63640 3007
rect 63800 3007 66830 3030
rect 63800 2000 63823 3007
rect 63617 1000 63823 2000
rect 63617 23 63640 1000
rect 60610 0 63640 23
rect 63800 23 63823 1000
rect 66807 2000 66830 3007
rect 66990 3007 70020 3030
rect 66990 2000 67013 3007
rect 66807 1000 67013 2000
rect 66807 23 66830 1000
rect 63800 0 66830 23
rect 66990 23 67013 1000
rect 69997 2000 70020 3007
rect 70180 3007 73210 3030
rect 70180 2000 70203 3007
rect 69997 1000 70203 2000
rect 69997 23 70020 1000
rect 66990 0 70020 23
rect 70180 23 70203 1000
rect 73187 2000 73210 3007
rect 73370 3007 76400 3030
rect 73370 2000 73393 3007
rect 73187 1000 73393 2000
rect 73187 23 73210 1000
rect 70180 0 73210 23
rect 73370 23 73393 1000
rect 76377 2000 76400 3007
rect 76560 3007 79590 3030
rect 76560 2000 76583 3007
rect 76377 1000 76583 2000
rect 76377 23 76400 1000
rect 73370 0 76400 23
rect 76560 23 76583 1000
rect 79567 2000 79590 3007
rect 79750 3007 82780 3030
rect 79750 2000 79773 3007
rect 79567 1000 79773 2000
rect 79567 23 79590 1000
rect 76560 0 79590 23
rect 79750 23 79773 1000
rect 82757 2000 82780 3007
rect 82940 3007 85970 3030
rect 82940 2000 82963 3007
rect 82757 1000 82963 2000
rect 82757 23 82780 1000
rect 79750 0 82780 23
rect 82940 23 82963 1000
rect 85947 2000 85970 3007
rect 86130 3007 89160 3030
rect 86130 2000 86153 3007
rect 85947 1000 86153 2000
rect 85947 23 85970 1000
rect 82940 0 85970 23
rect 86130 23 86153 1000
rect 89137 2000 89160 3007
rect 89320 3007 92350 3030
rect 89320 2000 89343 3007
rect 89137 1000 89343 2000
rect 89137 23 89160 1000
rect 86130 0 89160 23
rect 89320 23 89343 1000
rect 92327 2000 92350 3007
rect 92510 3007 95540 3030
rect 92510 2000 92533 3007
rect 92327 1000 92533 2000
rect 92327 23 92350 1000
rect 89320 0 92350 23
rect 92510 23 92533 1000
rect 95517 2000 95540 3007
rect 95700 3007 98730 3030
rect 95700 2000 95723 3007
rect 95517 1000 95723 2000
rect 95517 23 95540 1000
rect 92510 0 95540 23
rect 95700 23 95723 1000
rect 98707 2000 98730 3007
rect 98890 3007 101920 3030
rect 98890 2000 98913 3007
rect 98707 1000 98913 2000
rect 98707 23 98730 1000
rect 95700 0 98730 23
rect 98890 23 98913 1000
rect 101897 2000 101920 3007
rect 102080 3007 105110 3030
rect 102080 2000 102103 3007
rect 101897 1000 102103 2000
rect 101897 23 101920 1000
rect 98890 0 101920 23
rect 102080 23 102103 1000
rect 105087 2000 105110 3007
rect 105270 3007 108300 3030
rect 105270 2000 105293 3007
rect 105087 1000 105293 2000
rect 105087 23 105110 1000
rect 102080 0 105110 23
rect 105270 23 105293 1000
rect 108277 2000 108300 3007
rect 108460 3007 111490 3030
rect 108460 2000 108483 3007
rect 108277 1000 108483 2000
rect 108277 23 108300 1000
rect 105270 0 108300 23
rect 108460 23 108483 1000
rect 111467 2000 111490 3007
rect 111650 3007 114680 3030
rect 111650 2000 111673 3007
rect 111467 1000 111673 2000
rect 111467 23 111490 1000
rect 108460 0 111490 23
rect 111650 23 111673 1000
rect 114657 2000 114680 3007
rect 114840 3007 117870 3030
rect 114840 2000 114863 3007
rect 114657 1000 114863 2000
rect 114657 23 114680 1000
rect 111650 0 114680 23
rect 114840 23 114863 1000
rect 117847 2000 117870 3007
rect 118030 3007 121060 3030
rect 118030 2000 118053 3007
rect 117847 1000 118053 2000
rect 117847 23 117870 1000
rect 114840 0 117870 23
rect 118030 23 118053 1000
rect 121037 2000 121060 3007
rect 121220 3007 124250 3030
rect 121220 2000 121243 3007
rect 121037 1000 121243 2000
rect 121037 23 121060 1000
rect 118030 0 121060 23
rect 121220 23 121243 1000
rect 124227 2000 124250 3007
rect 124410 3007 127440 3030
rect 124410 2000 124433 3007
rect 124227 1000 124433 2000
rect 124227 23 124250 1000
rect 121220 0 124250 23
rect 124410 23 124433 1000
rect 127417 2000 127440 3007
rect 127600 3007 130630 3030
rect 127600 2000 127623 3007
rect 127417 1000 127623 2000
rect 127417 23 127440 1000
rect 124410 0 127440 23
rect 127600 23 127623 1000
rect 130607 2000 130630 3007
rect 130790 3007 133820 3030
rect 130790 2000 130813 3007
rect 130607 1000 130813 2000
rect 130607 23 130630 1000
rect 127600 0 130630 23
rect 130790 23 130813 1000
rect 133797 2000 133820 3007
rect 133980 3007 137010 3030
rect 133980 2000 134003 3007
rect 133797 1000 134003 2000
rect 133797 23 133820 1000
rect 130790 0 133820 23
rect 133980 23 134003 1000
rect 136987 2000 137010 3007
rect 136987 1000 137170 2000
rect 136987 23 137010 1000
rect 133980 0 137010 23
<< via4 >>
rect 1020 166020 68970 166980
rect 71200 166020 135960 166980
rect 50 121310 9320 140110
rect 50 79839 9320 98639
<< mimcap2 >>
rect 15 165697 3015 165705
rect 15 162713 23 165697
rect 3007 162713 3015 165697
rect 15 162705 3015 162713
rect 3205 165697 6205 165705
rect 3205 162713 3213 165697
rect 6197 162713 6205 165697
rect 3205 162705 6205 162713
rect 6395 165697 9395 165705
rect 6395 162713 6403 165697
rect 9387 162713 9395 165697
rect 6395 162705 9395 162713
rect 9585 165697 12585 165705
rect 9585 162713 9593 165697
rect 12577 162713 12585 165697
rect 9585 162705 12585 162713
rect 12775 165697 15775 165705
rect 12775 162713 12783 165697
rect 15767 162713 15775 165697
rect 12775 162705 15775 162713
rect 15965 165697 18965 165705
rect 15965 162713 15973 165697
rect 18957 162713 18965 165697
rect 15965 162705 18965 162713
rect 19155 165697 22155 165705
rect 19155 162713 19163 165697
rect 22147 162713 22155 165697
rect 19155 162705 22155 162713
rect 22345 165697 25345 165705
rect 22345 162713 22353 165697
rect 25337 162713 25345 165697
rect 22345 162705 25345 162713
rect 25535 165697 28535 165705
rect 25535 162713 25543 165697
rect 28527 162713 28535 165697
rect 25535 162705 28535 162713
rect 28725 165697 31725 165705
rect 28725 162713 28733 165697
rect 31717 162713 31725 165697
rect 28725 162705 31725 162713
rect 31915 165697 34915 165705
rect 31915 162713 31923 165697
rect 34907 162713 34915 165697
rect 31915 162705 34915 162713
rect 35105 165697 38105 165705
rect 35105 162713 35113 165697
rect 38097 162713 38105 165697
rect 35105 162705 38105 162713
rect 38295 165697 41295 165705
rect 38295 162713 38303 165697
rect 41287 162713 41295 165697
rect 38295 162705 41295 162713
rect 41485 165697 44485 165705
rect 41485 162713 41493 165697
rect 44477 162713 44485 165697
rect 41485 162705 44485 162713
rect 44675 165697 47675 165705
rect 44675 162713 44683 165697
rect 47667 162713 47675 165697
rect 44675 162705 47675 162713
rect 47865 165697 50865 165705
rect 47865 162713 47873 165697
rect 50857 162713 50865 165697
rect 47865 162705 50865 162713
rect 51055 165697 54055 165705
rect 51055 162713 51063 165697
rect 54047 162713 54055 165697
rect 51055 162705 54055 162713
rect 54245 165697 57245 165705
rect 54245 162713 54253 165697
rect 57237 162713 57245 165697
rect 54245 162705 57245 162713
rect 57435 165697 60435 165705
rect 57435 162713 57443 165697
rect 60427 162713 60435 165697
rect 57435 162705 60435 162713
rect 60625 165697 63625 165705
rect 60625 162713 60633 165697
rect 63617 162713 63625 165697
rect 60625 162705 63625 162713
rect 63815 165697 66815 165705
rect 63815 162713 63823 165697
rect 66807 162713 66815 165697
rect 63815 162705 66815 162713
rect 67005 165697 70005 165705
rect 67005 162713 67013 165697
rect 69997 162713 70005 165697
rect 67005 162705 70005 162713
rect 70195 165697 73195 165705
rect 70195 162713 70203 165697
rect 73187 162713 73195 165697
rect 70195 162705 73195 162713
rect 73385 165697 76385 165705
rect 73385 162713 73393 165697
rect 76377 162713 76385 165697
rect 73385 162705 76385 162713
rect 76575 165697 79575 165705
rect 76575 162713 76583 165697
rect 79567 162713 79575 165697
rect 76575 162705 79575 162713
rect 79765 165697 82765 165705
rect 79765 162713 79773 165697
rect 82757 162713 82765 165697
rect 79765 162705 82765 162713
rect 82955 165697 85955 165705
rect 82955 162713 82963 165697
rect 85947 162713 85955 165697
rect 82955 162705 85955 162713
rect 86145 165697 89145 165705
rect 86145 162713 86153 165697
rect 89137 162713 89145 165697
rect 86145 162705 89145 162713
rect 89335 165697 92335 165705
rect 89335 162713 89343 165697
rect 92327 162713 92335 165697
rect 89335 162705 92335 162713
rect 92525 165697 95525 165705
rect 92525 162713 92533 165697
rect 95517 162713 95525 165697
rect 92525 162705 95525 162713
rect 95715 165697 98715 165705
rect 95715 162713 95723 165697
rect 98707 162713 98715 165697
rect 95715 162705 98715 162713
rect 98905 165697 101905 165705
rect 98905 162713 98913 165697
rect 101897 162713 101905 165697
rect 98905 162705 101905 162713
rect 102095 165697 105095 165705
rect 102095 162713 102103 165697
rect 105087 162713 105095 165697
rect 102095 162705 105095 162713
rect 105285 165697 108285 165705
rect 105285 162713 105293 165697
rect 108277 162713 108285 165697
rect 105285 162705 108285 162713
rect 108475 165697 111475 165705
rect 108475 162713 108483 165697
rect 111467 162713 111475 165697
rect 108475 162705 111475 162713
rect 111665 165697 114665 165705
rect 111665 162713 111673 165697
rect 114657 162713 114665 165697
rect 111665 162705 114665 162713
rect 114855 165697 117855 165705
rect 114855 162713 114863 165697
rect 117847 162713 117855 165697
rect 114855 162705 117855 162713
rect 118045 165697 121045 165705
rect 118045 162713 118053 165697
rect 121037 162713 121045 165697
rect 118045 162705 121045 162713
rect 121235 165697 124235 165705
rect 121235 162713 121243 165697
rect 124227 162713 124235 165697
rect 121235 162705 124235 162713
rect 124425 165697 127425 165705
rect 124425 162713 124433 165697
rect 127417 162713 127425 165697
rect 124425 162705 127425 162713
rect 127615 165697 130615 165705
rect 127615 162713 127623 165697
rect 130607 162713 130615 165697
rect 127615 162705 130615 162713
rect 130805 165697 133805 165705
rect 130805 162713 130813 165697
rect 133797 162713 133805 165697
rect 130805 162705 133805 162713
rect 133995 165697 136995 165705
rect 133995 162713 134003 165697
rect 136987 162713 136995 165697
rect 133995 162705 136995 162713
rect 15 162507 3015 162515
rect 15 159523 23 162507
rect 3007 159523 3015 162507
rect 15 159515 3015 159523
rect 3205 162507 6205 162515
rect 3205 159523 3213 162507
rect 6197 159523 6205 162507
rect 3205 159515 6205 159523
rect 6395 162507 9395 162515
rect 6395 159523 6403 162507
rect 9387 159523 9395 162507
rect 6395 159515 9395 159523
rect 9585 162507 12585 162515
rect 9585 159523 9593 162507
rect 12577 159523 12585 162507
rect 9585 159515 12585 159523
rect 12775 162507 15775 162515
rect 12775 159523 12783 162507
rect 15767 159523 15775 162507
rect 12775 159515 15775 159523
rect 15965 162507 18965 162515
rect 15965 159523 15973 162507
rect 18957 159523 18965 162507
rect 15965 159515 18965 159523
rect 19155 162507 22155 162515
rect 19155 159523 19163 162507
rect 22147 159523 22155 162507
rect 19155 159515 22155 159523
rect 22345 162507 25345 162515
rect 22345 159523 22353 162507
rect 25337 159523 25345 162507
rect 22345 159515 25345 159523
rect 25535 162507 28535 162515
rect 25535 159523 25543 162507
rect 28527 159523 28535 162507
rect 25535 159515 28535 159523
rect 28725 162507 31725 162515
rect 28725 159523 28733 162507
rect 31717 159523 31725 162507
rect 28725 159515 31725 159523
rect 31915 162507 34915 162515
rect 31915 159523 31923 162507
rect 34907 159523 34915 162507
rect 31915 159515 34915 159523
rect 35105 162507 38105 162515
rect 35105 159523 35113 162507
rect 38097 159523 38105 162507
rect 35105 159515 38105 159523
rect 38295 162507 41295 162515
rect 38295 159523 38303 162507
rect 41287 159523 41295 162507
rect 38295 159515 41295 159523
rect 41485 162507 44485 162515
rect 41485 159523 41493 162507
rect 44477 159523 44485 162507
rect 41485 159515 44485 159523
rect 44675 162507 47675 162515
rect 44675 159523 44683 162507
rect 47667 159523 47675 162507
rect 44675 159515 47675 159523
rect 47865 162507 50865 162515
rect 47865 159523 47873 162507
rect 50857 159523 50865 162507
rect 47865 159515 50865 159523
rect 51055 162507 54055 162515
rect 51055 159523 51063 162507
rect 54047 159523 54055 162507
rect 51055 159515 54055 159523
rect 54245 162507 57245 162515
rect 54245 159523 54253 162507
rect 57237 159523 57245 162507
rect 54245 159515 57245 159523
rect 57435 162507 60435 162515
rect 57435 159523 57443 162507
rect 60427 159523 60435 162507
rect 57435 159515 60435 159523
rect 60625 162507 63625 162515
rect 60625 159523 60633 162507
rect 63617 159523 63625 162507
rect 60625 159515 63625 159523
rect 63815 162507 66815 162515
rect 63815 159523 63823 162507
rect 66807 159523 66815 162507
rect 63815 159515 66815 159523
rect 67005 162507 70005 162515
rect 67005 159523 67013 162507
rect 69997 159523 70005 162507
rect 67005 159515 70005 159523
rect 70195 162507 73195 162515
rect 70195 159523 70203 162507
rect 73187 159523 73195 162507
rect 70195 159515 73195 159523
rect 73385 162507 76385 162515
rect 73385 159523 73393 162507
rect 76377 159523 76385 162507
rect 73385 159515 76385 159523
rect 76575 162507 79575 162515
rect 76575 159523 76583 162507
rect 79567 159523 79575 162507
rect 76575 159515 79575 159523
rect 79765 162507 82765 162515
rect 79765 159523 79773 162507
rect 82757 159523 82765 162507
rect 79765 159515 82765 159523
rect 82955 162507 85955 162515
rect 82955 159523 82963 162507
rect 85947 159523 85955 162507
rect 82955 159515 85955 159523
rect 86145 162507 89145 162515
rect 86145 159523 86153 162507
rect 89137 159523 89145 162507
rect 86145 159515 89145 159523
rect 89335 162507 92335 162515
rect 89335 159523 89343 162507
rect 92327 159523 92335 162507
rect 89335 159515 92335 159523
rect 92525 162507 95525 162515
rect 92525 159523 92533 162507
rect 95517 159523 95525 162507
rect 92525 159515 95525 159523
rect 95715 162507 98715 162515
rect 95715 159523 95723 162507
rect 98707 159523 98715 162507
rect 95715 159515 98715 159523
rect 98905 162507 101905 162515
rect 98905 159523 98913 162507
rect 101897 159523 101905 162507
rect 98905 159515 101905 159523
rect 102095 162507 105095 162515
rect 102095 159523 102103 162507
rect 105087 159523 105095 162507
rect 102095 159515 105095 159523
rect 105285 162507 108285 162515
rect 105285 159523 105293 162507
rect 108277 159523 108285 162507
rect 105285 159515 108285 159523
rect 108475 162507 111475 162515
rect 108475 159523 108483 162507
rect 111467 159523 111475 162507
rect 108475 159515 111475 159523
rect 111665 162507 114665 162515
rect 111665 159523 111673 162507
rect 114657 159523 114665 162507
rect 111665 159515 114665 159523
rect 114855 162507 117855 162515
rect 114855 159523 114863 162507
rect 117847 159523 117855 162507
rect 114855 159515 117855 159523
rect 118045 162507 121045 162515
rect 118045 159523 118053 162507
rect 121037 159523 121045 162507
rect 118045 159515 121045 159523
rect 121235 162507 124235 162515
rect 121235 159523 121243 162507
rect 124227 159523 124235 162507
rect 121235 159515 124235 159523
rect 124425 162507 127425 162515
rect 124425 159523 124433 162507
rect 127417 159523 127425 162507
rect 124425 159515 127425 159523
rect 127615 162507 130615 162515
rect 127615 159523 127623 162507
rect 130607 159523 130615 162507
rect 127615 159515 130615 159523
rect 130805 162507 133805 162515
rect 130805 159523 130813 162507
rect 133797 159523 133805 162507
rect 130805 159515 133805 159523
rect 133995 162507 136995 162515
rect 133995 159523 134003 162507
rect 136987 159523 136995 162507
rect 133995 159515 136995 159523
rect 15 159317 3015 159325
rect 15 156333 23 159317
rect 3007 156333 3015 159317
rect 15 156325 3015 156333
rect 3205 159317 6205 159325
rect 3205 156333 3213 159317
rect 6197 156333 6205 159317
rect 3205 156325 6205 156333
rect 6395 159317 9395 159325
rect 6395 156333 6403 159317
rect 9387 156333 9395 159317
rect 6395 156325 9395 156333
rect 9585 159317 12585 159325
rect 9585 156333 9593 159317
rect 12577 156333 12585 159317
rect 9585 156325 12585 156333
rect 12775 159317 15775 159325
rect 12775 156333 12783 159317
rect 15767 156333 15775 159317
rect 12775 156325 15775 156333
rect 15965 159317 18965 159325
rect 15965 156333 15973 159317
rect 18957 156333 18965 159317
rect 15965 156325 18965 156333
rect 19155 159317 22155 159325
rect 19155 156333 19163 159317
rect 22147 156333 22155 159317
rect 19155 156325 22155 156333
rect 22345 159317 25345 159325
rect 22345 156333 22353 159317
rect 25337 156333 25345 159317
rect 22345 156325 25345 156333
rect 25535 159317 28535 159325
rect 25535 156333 25543 159317
rect 28527 156333 28535 159317
rect 25535 156325 28535 156333
rect 28725 159317 31725 159325
rect 28725 156333 28733 159317
rect 31717 156333 31725 159317
rect 28725 156325 31725 156333
rect 31915 159317 34915 159325
rect 31915 156333 31923 159317
rect 34907 156333 34915 159317
rect 31915 156325 34915 156333
rect 35105 159317 38105 159325
rect 35105 156333 35113 159317
rect 38097 156333 38105 159317
rect 35105 156325 38105 156333
rect 38295 159317 41295 159325
rect 38295 156333 38303 159317
rect 41287 156333 41295 159317
rect 38295 156325 41295 156333
rect 41485 159317 44485 159325
rect 41485 156333 41493 159317
rect 44477 156333 44485 159317
rect 41485 156325 44485 156333
rect 44675 159317 47675 159325
rect 44675 156333 44683 159317
rect 47667 156333 47675 159317
rect 44675 156325 47675 156333
rect 47865 159317 50865 159325
rect 47865 156333 47873 159317
rect 50857 156333 50865 159317
rect 47865 156325 50865 156333
rect 51055 159317 54055 159325
rect 51055 156333 51063 159317
rect 54047 156333 54055 159317
rect 51055 156325 54055 156333
rect 54245 159317 57245 159325
rect 54245 156333 54253 159317
rect 57237 156333 57245 159317
rect 54245 156325 57245 156333
rect 57435 159317 60435 159325
rect 57435 156333 57443 159317
rect 60427 156333 60435 159317
rect 57435 156325 60435 156333
rect 60625 159317 63625 159325
rect 60625 156333 60633 159317
rect 63617 156333 63625 159317
rect 60625 156325 63625 156333
rect 63815 159317 66815 159325
rect 63815 156333 63823 159317
rect 66807 156333 66815 159317
rect 63815 156325 66815 156333
rect 67005 159317 70005 159325
rect 67005 156333 67013 159317
rect 69997 156333 70005 159317
rect 67005 156325 70005 156333
rect 70195 159317 73195 159325
rect 70195 156333 70203 159317
rect 73187 156333 73195 159317
rect 70195 156325 73195 156333
rect 73385 159317 76385 159325
rect 73385 156333 73393 159317
rect 76377 156333 76385 159317
rect 73385 156325 76385 156333
rect 76575 159317 79575 159325
rect 76575 156333 76583 159317
rect 79567 156333 79575 159317
rect 76575 156325 79575 156333
rect 79765 159317 82765 159325
rect 79765 156333 79773 159317
rect 82757 156333 82765 159317
rect 79765 156325 82765 156333
rect 82955 159317 85955 159325
rect 82955 156333 82963 159317
rect 85947 156333 85955 159317
rect 82955 156325 85955 156333
rect 86145 159317 89145 159325
rect 86145 156333 86153 159317
rect 89137 156333 89145 159317
rect 86145 156325 89145 156333
rect 89335 159317 92335 159325
rect 89335 156333 89343 159317
rect 92327 156333 92335 159317
rect 89335 156325 92335 156333
rect 92525 159317 95525 159325
rect 92525 156333 92533 159317
rect 95517 156333 95525 159317
rect 92525 156325 95525 156333
rect 95715 159317 98715 159325
rect 95715 156333 95723 159317
rect 98707 156333 98715 159317
rect 95715 156325 98715 156333
rect 98905 159317 101905 159325
rect 98905 156333 98913 159317
rect 101897 156333 101905 159317
rect 98905 156325 101905 156333
rect 102095 159317 105095 159325
rect 102095 156333 102103 159317
rect 105087 156333 105095 159317
rect 102095 156325 105095 156333
rect 105285 159317 108285 159325
rect 105285 156333 105293 159317
rect 108277 156333 108285 159317
rect 105285 156325 108285 156333
rect 108475 159317 111475 159325
rect 108475 156333 108483 159317
rect 111467 156333 111475 159317
rect 108475 156325 111475 156333
rect 111665 159317 114665 159325
rect 111665 156333 111673 159317
rect 114657 156333 114665 159317
rect 111665 156325 114665 156333
rect 114855 159317 117855 159325
rect 114855 156333 114863 159317
rect 117847 156333 117855 159317
rect 114855 156325 117855 156333
rect 118045 159317 121045 159325
rect 118045 156333 118053 159317
rect 121037 156333 121045 159317
rect 118045 156325 121045 156333
rect 121235 159317 124235 159325
rect 121235 156333 121243 159317
rect 124227 156333 124235 159317
rect 121235 156325 124235 156333
rect 124425 159317 127425 159325
rect 124425 156333 124433 159317
rect 127417 156333 127425 159317
rect 124425 156325 127425 156333
rect 127615 159317 130615 159325
rect 127615 156333 127623 159317
rect 130607 156333 130615 159317
rect 127615 156325 130615 156333
rect 130805 159317 133805 159325
rect 130805 156333 130813 159317
rect 133797 156333 133805 159317
rect 130805 156325 133805 156333
rect 133995 159317 136995 159325
rect 133995 156333 134003 159317
rect 136987 156333 136995 159317
rect 133995 156325 136995 156333
rect 15 156127 3015 156135
rect 15 153143 23 156127
rect 3007 153143 3015 156127
rect 15 153135 3015 153143
rect 3205 156127 6205 156135
rect 3205 153143 3213 156127
rect 6197 153143 6205 156127
rect 3205 153135 6205 153143
rect 6395 156127 9395 156135
rect 6395 153143 6403 156127
rect 9387 153143 9395 156127
rect 6395 153135 9395 153143
rect 9585 156127 12585 156135
rect 9585 153143 9593 156127
rect 12577 153143 12585 156127
rect 9585 153135 12585 153143
rect 12775 156127 15775 156135
rect 12775 153143 12783 156127
rect 15767 153143 15775 156127
rect 12775 153135 15775 153143
rect 15965 156127 18965 156135
rect 15965 153143 15973 156127
rect 18957 153143 18965 156127
rect 15965 153135 18965 153143
rect 19155 156127 22155 156135
rect 19155 153143 19163 156127
rect 22147 153143 22155 156127
rect 19155 153135 22155 153143
rect 22345 156127 25345 156135
rect 22345 153143 22353 156127
rect 25337 153143 25345 156127
rect 22345 153135 25345 153143
rect 25535 156127 28535 156135
rect 25535 153143 25543 156127
rect 28527 153143 28535 156127
rect 25535 153135 28535 153143
rect 28725 156127 31725 156135
rect 28725 153143 28733 156127
rect 31717 153143 31725 156127
rect 28725 153135 31725 153143
rect 31915 156127 34915 156135
rect 31915 153143 31923 156127
rect 34907 153143 34915 156127
rect 31915 153135 34915 153143
rect 35105 156127 38105 156135
rect 35105 153143 35113 156127
rect 38097 153143 38105 156127
rect 35105 153135 38105 153143
rect 38295 156127 41295 156135
rect 38295 153143 38303 156127
rect 41287 153143 41295 156127
rect 38295 153135 41295 153143
rect 41485 156127 44485 156135
rect 41485 153143 41493 156127
rect 44477 153143 44485 156127
rect 41485 153135 44485 153143
rect 44675 156127 47675 156135
rect 44675 153143 44683 156127
rect 47667 153143 47675 156127
rect 44675 153135 47675 153143
rect 47865 156127 50865 156135
rect 47865 153143 47873 156127
rect 50857 153143 50865 156127
rect 47865 153135 50865 153143
rect 51055 156127 54055 156135
rect 51055 153143 51063 156127
rect 54047 153143 54055 156127
rect 51055 153135 54055 153143
rect 54245 156127 57245 156135
rect 54245 153143 54253 156127
rect 57237 153143 57245 156127
rect 54245 153135 57245 153143
rect 57435 156127 60435 156135
rect 57435 153143 57443 156127
rect 60427 153143 60435 156127
rect 57435 153135 60435 153143
rect 60625 156127 63625 156135
rect 60625 153143 60633 156127
rect 63617 153143 63625 156127
rect 60625 153135 63625 153143
rect 63815 156127 66815 156135
rect 63815 153143 63823 156127
rect 66807 153143 66815 156127
rect 63815 153135 66815 153143
rect 67005 156127 70005 156135
rect 67005 153143 67013 156127
rect 69997 153143 70005 156127
rect 67005 153135 70005 153143
rect 70195 156127 73195 156135
rect 70195 153143 70203 156127
rect 73187 153143 73195 156127
rect 70195 153135 73195 153143
rect 73385 156127 76385 156135
rect 73385 153143 73393 156127
rect 76377 153143 76385 156127
rect 73385 153135 76385 153143
rect 76575 156127 79575 156135
rect 76575 153143 76583 156127
rect 79567 153143 79575 156127
rect 76575 153135 79575 153143
rect 79765 156127 82765 156135
rect 79765 153143 79773 156127
rect 82757 153143 82765 156127
rect 79765 153135 82765 153143
rect 82955 156127 85955 156135
rect 82955 153143 82963 156127
rect 85947 153143 85955 156127
rect 82955 153135 85955 153143
rect 86145 156127 89145 156135
rect 86145 153143 86153 156127
rect 89137 153143 89145 156127
rect 86145 153135 89145 153143
rect 89335 156127 92335 156135
rect 89335 153143 89343 156127
rect 92327 153143 92335 156127
rect 89335 153135 92335 153143
rect 92525 156127 95525 156135
rect 92525 153143 92533 156127
rect 95517 153143 95525 156127
rect 92525 153135 95525 153143
rect 95715 156127 98715 156135
rect 95715 153143 95723 156127
rect 98707 153143 98715 156127
rect 95715 153135 98715 153143
rect 98905 156127 101905 156135
rect 98905 153143 98913 156127
rect 101897 153143 101905 156127
rect 98905 153135 101905 153143
rect 102095 156127 105095 156135
rect 102095 153143 102103 156127
rect 105087 153143 105095 156127
rect 102095 153135 105095 153143
rect 105285 156127 108285 156135
rect 105285 153143 105293 156127
rect 108277 153143 108285 156127
rect 105285 153135 108285 153143
rect 108475 156127 111475 156135
rect 108475 153143 108483 156127
rect 111467 153143 111475 156127
rect 108475 153135 111475 153143
rect 111665 156127 114665 156135
rect 111665 153143 111673 156127
rect 114657 153143 114665 156127
rect 111665 153135 114665 153143
rect 114855 156127 117855 156135
rect 114855 153143 114863 156127
rect 117847 153143 117855 156127
rect 114855 153135 117855 153143
rect 118045 156127 121045 156135
rect 118045 153143 118053 156127
rect 121037 153143 121045 156127
rect 118045 153135 121045 153143
rect 121235 156127 124235 156135
rect 121235 153143 121243 156127
rect 124227 153143 124235 156127
rect 121235 153135 124235 153143
rect 124425 156127 127425 156135
rect 124425 153143 124433 156127
rect 127417 153143 127425 156127
rect 124425 153135 127425 153143
rect 127615 156127 130615 156135
rect 127615 153143 127623 156127
rect 130607 153143 130615 156127
rect 127615 153135 130615 153143
rect 130805 156127 133805 156135
rect 130805 153143 130813 156127
rect 133797 153143 133805 156127
rect 130805 153135 133805 153143
rect 133995 156127 136995 156135
rect 133995 153143 134003 156127
rect 136987 153143 136995 156127
rect 133995 153135 136995 153143
rect 15 152937 3015 152945
rect 15 149953 23 152937
rect 3007 149953 3015 152937
rect 15 149945 3015 149953
rect 3205 152937 6205 152945
rect 3205 149953 3213 152937
rect 6197 149953 6205 152937
rect 3205 149945 6205 149953
rect 6395 152937 9395 152945
rect 6395 149953 6403 152937
rect 9387 149953 9395 152937
rect 6395 149945 9395 149953
rect 9585 152937 12585 152945
rect 9585 149953 9593 152937
rect 12577 149953 12585 152937
rect 9585 149945 12585 149953
rect 12775 152937 15775 152945
rect 12775 149953 12783 152937
rect 15767 149953 15775 152937
rect 12775 149945 15775 149953
rect 15965 152937 18965 152945
rect 15965 149953 15973 152937
rect 18957 149953 18965 152937
rect 15965 149945 18965 149953
rect 19155 152937 22155 152945
rect 19155 149953 19163 152937
rect 22147 149953 22155 152937
rect 19155 149945 22155 149953
rect 22345 152937 25345 152945
rect 22345 149953 22353 152937
rect 25337 149953 25345 152937
rect 22345 149945 25345 149953
rect 25535 152937 28535 152945
rect 25535 149953 25543 152937
rect 28527 149953 28535 152937
rect 25535 149945 28535 149953
rect 28725 152937 31725 152945
rect 28725 149953 28733 152937
rect 31717 149953 31725 152937
rect 28725 149945 31725 149953
rect 31915 152937 34915 152945
rect 31915 149953 31923 152937
rect 34907 149953 34915 152937
rect 31915 149945 34915 149953
rect 35105 152937 38105 152945
rect 35105 149953 35113 152937
rect 38097 149953 38105 152937
rect 35105 149945 38105 149953
rect 38295 152937 41295 152945
rect 38295 149953 38303 152937
rect 41287 149953 41295 152937
rect 38295 149945 41295 149953
rect 41485 152937 44485 152945
rect 41485 149953 41493 152937
rect 44477 149953 44485 152937
rect 41485 149945 44485 149953
rect 44675 152937 47675 152945
rect 44675 149953 44683 152937
rect 47667 149953 47675 152937
rect 44675 149945 47675 149953
rect 47865 152937 50865 152945
rect 47865 149953 47873 152937
rect 50857 149953 50865 152937
rect 47865 149945 50865 149953
rect 51055 152937 54055 152945
rect 51055 149953 51063 152937
rect 54047 149953 54055 152937
rect 51055 149945 54055 149953
rect 54245 152937 57245 152945
rect 54245 149953 54253 152937
rect 57237 149953 57245 152937
rect 54245 149945 57245 149953
rect 57435 152937 60435 152945
rect 57435 149953 57443 152937
rect 60427 149953 60435 152937
rect 57435 149945 60435 149953
rect 60625 152937 63625 152945
rect 60625 149953 60633 152937
rect 63617 149953 63625 152937
rect 60625 149945 63625 149953
rect 63815 152937 66815 152945
rect 63815 149953 63823 152937
rect 66807 149953 66815 152937
rect 63815 149945 66815 149953
rect 67005 152937 70005 152945
rect 67005 149953 67013 152937
rect 69997 149953 70005 152937
rect 67005 149945 70005 149953
rect 70195 152937 73195 152945
rect 70195 149953 70203 152937
rect 73187 149953 73195 152937
rect 70195 149945 73195 149953
rect 73385 152937 76385 152945
rect 73385 149953 73393 152937
rect 76377 149953 76385 152937
rect 73385 149945 76385 149953
rect 76575 152937 79575 152945
rect 76575 149953 76583 152937
rect 79567 149953 79575 152937
rect 76575 149945 79575 149953
rect 79765 152937 82765 152945
rect 79765 149953 79773 152937
rect 82757 149953 82765 152937
rect 79765 149945 82765 149953
rect 82955 152937 85955 152945
rect 82955 149953 82963 152937
rect 85947 149953 85955 152937
rect 82955 149945 85955 149953
rect 86145 152937 89145 152945
rect 86145 149953 86153 152937
rect 89137 149953 89145 152937
rect 86145 149945 89145 149953
rect 89335 152937 92335 152945
rect 89335 149953 89343 152937
rect 92327 149953 92335 152937
rect 89335 149945 92335 149953
rect 92525 152937 95525 152945
rect 92525 149953 92533 152937
rect 95517 149953 95525 152937
rect 92525 149945 95525 149953
rect 95715 152937 98715 152945
rect 95715 149953 95723 152937
rect 98707 149953 98715 152937
rect 95715 149945 98715 149953
rect 98905 152937 101905 152945
rect 98905 149953 98913 152937
rect 101897 149953 101905 152937
rect 98905 149945 101905 149953
rect 102095 152937 105095 152945
rect 102095 149953 102103 152937
rect 105087 149953 105095 152937
rect 102095 149945 105095 149953
rect 105285 152937 108285 152945
rect 105285 149953 105293 152937
rect 108277 149953 108285 152937
rect 105285 149945 108285 149953
rect 108475 152937 111475 152945
rect 108475 149953 108483 152937
rect 111467 149953 111475 152937
rect 108475 149945 111475 149953
rect 111665 152937 114665 152945
rect 111665 149953 111673 152937
rect 114657 149953 114665 152937
rect 111665 149945 114665 149953
rect 114855 152937 117855 152945
rect 114855 149953 114863 152937
rect 117847 149953 117855 152937
rect 114855 149945 117855 149953
rect 118045 152937 121045 152945
rect 118045 149953 118053 152937
rect 121037 149953 121045 152937
rect 118045 149945 121045 149953
rect 121235 152937 124235 152945
rect 121235 149953 121243 152937
rect 124227 149953 124235 152937
rect 121235 149945 124235 149953
rect 124425 152937 127425 152945
rect 124425 149953 124433 152937
rect 127417 149953 127425 152937
rect 124425 149945 127425 149953
rect 127615 152937 130615 152945
rect 127615 149953 127623 152937
rect 130607 149953 130615 152937
rect 127615 149945 130615 149953
rect 130805 152937 133805 152945
rect 130805 149953 130813 152937
rect 133797 149953 133805 152937
rect 130805 149945 133805 149953
rect 133995 152937 136995 152945
rect 133995 149953 134003 152937
rect 136987 149953 136995 152937
rect 133995 149945 136995 149953
rect 15 149747 3015 149755
rect 15 146763 23 149747
rect 3007 146763 3015 149747
rect 15 146755 3015 146763
rect 3205 149747 6205 149755
rect 3205 146763 3213 149747
rect 6197 146763 6205 149747
rect 3205 146755 6205 146763
rect 6395 149747 9395 149755
rect 6395 146763 6403 149747
rect 9387 146763 9395 149747
rect 6395 146755 9395 146763
rect 9585 149747 12585 149755
rect 9585 146763 9593 149747
rect 12577 146763 12585 149747
rect 9585 146755 12585 146763
rect 12775 149747 15775 149755
rect 12775 146763 12783 149747
rect 15767 146763 15775 149747
rect 12775 146755 15775 146763
rect 15965 149747 18965 149755
rect 15965 146763 15973 149747
rect 18957 146763 18965 149747
rect 15965 146755 18965 146763
rect 19155 149747 22155 149755
rect 19155 146763 19163 149747
rect 22147 146763 22155 149747
rect 19155 146755 22155 146763
rect 22345 149747 25345 149755
rect 22345 146763 22353 149747
rect 25337 146763 25345 149747
rect 22345 146755 25345 146763
rect 25535 149747 28535 149755
rect 25535 146763 25543 149747
rect 28527 146763 28535 149747
rect 25535 146755 28535 146763
rect 28725 149747 31725 149755
rect 28725 146763 28733 149747
rect 31717 146763 31725 149747
rect 28725 146755 31725 146763
rect 31915 149747 34915 149755
rect 31915 146763 31923 149747
rect 34907 146763 34915 149747
rect 31915 146755 34915 146763
rect 35105 149747 38105 149755
rect 35105 146763 35113 149747
rect 38097 146763 38105 149747
rect 35105 146755 38105 146763
rect 38295 149747 41295 149755
rect 38295 146763 38303 149747
rect 41287 146763 41295 149747
rect 38295 146755 41295 146763
rect 41485 149747 44485 149755
rect 41485 146763 41493 149747
rect 44477 146763 44485 149747
rect 41485 146755 44485 146763
rect 44675 149747 47675 149755
rect 44675 146763 44683 149747
rect 47667 146763 47675 149747
rect 44675 146755 47675 146763
rect 47865 149747 50865 149755
rect 47865 146763 47873 149747
rect 50857 146763 50865 149747
rect 47865 146755 50865 146763
rect 51055 149747 54055 149755
rect 51055 146763 51063 149747
rect 54047 146763 54055 149747
rect 51055 146755 54055 146763
rect 54245 149747 57245 149755
rect 54245 146763 54253 149747
rect 57237 146763 57245 149747
rect 54245 146755 57245 146763
rect 57435 149747 60435 149755
rect 57435 146763 57443 149747
rect 60427 146763 60435 149747
rect 57435 146755 60435 146763
rect 60625 149747 63625 149755
rect 60625 146763 60633 149747
rect 63617 146763 63625 149747
rect 60625 146755 63625 146763
rect 63815 149747 66815 149755
rect 63815 146763 63823 149747
rect 66807 146763 66815 149747
rect 63815 146755 66815 146763
rect 67005 149747 70005 149755
rect 67005 146763 67013 149747
rect 69997 146763 70005 149747
rect 67005 146755 70005 146763
rect 70195 149747 73195 149755
rect 70195 146763 70203 149747
rect 73187 146763 73195 149747
rect 70195 146755 73195 146763
rect 73385 149747 76385 149755
rect 73385 146763 73393 149747
rect 76377 146763 76385 149747
rect 73385 146755 76385 146763
rect 76575 149747 79575 149755
rect 76575 146763 76583 149747
rect 79567 146763 79575 149747
rect 76575 146755 79575 146763
rect 79765 149747 82765 149755
rect 79765 146763 79773 149747
rect 82757 146763 82765 149747
rect 79765 146755 82765 146763
rect 82955 149747 85955 149755
rect 82955 146763 82963 149747
rect 85947 146763 85955 149747
rect 82955 146755 85955 146763
rect 86145 149747 89145 149755
rect 86145 146763 86153 149747
rect 89137 146763 89145 149747
rect 86145 146755 89145 146763
rect 89335 149747 92335 149755
rect 89335 146763 89343 149747
rect 92327 146763 92335 149747
rect 89335 146755 92335 146763
rect 92525 149747 95525 149755
rect 92525 146763 92533 149747
rect 95517 146763 95525 149747
rect 92525 146755 95525 146763
rect 95715 149747 98715 149755
rect 95715 146763 95723 149747
rect 98707 146763 98715 149747
rect 95715 146755 98715 146763
rect 98905 149747 101905 149755
rect 98905 146763 98913 149747
rect 101897 146763 101905 149747
rect 98905 146755 101905 146763
rect 102095 149747 105095 149755
rect 102095 146763 102103 149747
rect 105087 146763 105095 149747
rect 102095 146755 105095 146763
rect 105285 149747 108285 149755
rect 105285 146763 105293 149747
rect 108277 146763 108285 149747
rect 105285 146755 108285 146763
rect 108475 149747 111475 149755
rect 108475 146763 108483 149747
rect 111467 146763 111475 149747
rect 108475 146755 111475 146763
rect 111665 149747 114665 149755
rect 111665 146763 111673 149747
rect 114657 146763 114665 149747
rect 111665 146755 114665 146763
rect 114855 149747 117855 149755
rect 114855 146763 114863 149747
rect 117847 146763 117855 149747
rect 114855 146755 117855 146763
rect 118045 149747 121045 149755
rect 118045 146763 118053 149747
rect 121037 146763 121045 149747
rect 118045 146755 121045 146763
rect 121235 149747 124235 149755
rect 121235 146763 121243 149747
rect 124227 146763 124235 149747
rect 121235 146755 124235 146763
rect 124425 149747 127425 149755
rect 124425 146763 124433 149747
rect 127417 146763 127425 149747
rect 124425 146755 127425 146763
rect 127615 149747 130615 149755
rect 127615 146763 127623 149747
rect 130607 146763 130615 149747
rect 127615 146755 130615 146763
rect 130805 149747 133805 149755
rect 130805 146763 130813 149747
rect 133797 146763 133805 149747
rect 130805 146755 133805 146763
rect 133995 149747 136995 149755
rect 133995 146763 134003 149747
rect 136987 146763 136995 149747
rect 133995 146755 136995 146763
rect 15 146557 3015 146565
rect 15 143573 23 146557
rect 3007 143573 3015 146557
rect 15 143565 3015 143573
rect 3205 146557 6205 146565
rect 3205 143573 3213 146557
rect 6197 143573 6205 146557
rect 3205 143565 6205 143573
rect 6395 146557 9395 146565
rect 6395 143573 6403 146557
rect 9387 143573 9395 146557
rect 6395 143565 9395 143573
rect 9585 146557 12585 146565
rect 9585 143573 9593 146557
rect 12577 143573 12585 146557
rect 9585 143565 12585 143573
rect 12775 146557 15775 146565
rect 12775 143573 12783 146557
rect 15767 143573 15775 146557
rect 12775 143565 15775 143573
rect 15965 146557 18965 146565
rect 15965 143573 15973 146557
rect 18957 143573 18965 146557
rect 15965 143565 18965 143573
rect 19155 146557 22155 146565
rect 19155 143573 19163 146557
rect 22147 143573 22155 146557
rect 19155 143565 22155 143573
rect 22345 146557 25345 146565
rect 22345 143573 22353 146557
rect 25337 143573 25345 146557
rect 22345 143565 25345 143573
rect 25535 146557 28535 146565
rect 25535 143573 25543 146557
rect 28527 143573 28535 146557
rect 25535 143565 28535 143573
rect 28725 146557 31725 146565
rect 28725 143573 28733 146557
rect 31717 143573 31725 146557
rect 28725 143565 31725 143573
rect 31915 146557 34915 146565
rect 31915 143573 31923 146557
rect 34907 143573 34915 146557
rect 31915 143565 34915 143573
rect 35105 146557 38105 146565
rect 35105 143573 35113 146557
rect 38097 143573 38105 146557
rect 35105 143565 38105 143573
rect 38295 146557 41295 146565
rect 38295 143573 38303 146557
rect 41287 143573 41295 146557
rect 38295 143565 41295 143573
rect 41485 146557 44485 146565
rect 41485 143573 41493 146557
rect 44477 143573 44485 146557
rect 41485 143565 44485 143573
rect 44675 146557 47675 146565
rect 44675 143573 44683 146557
rect 47667 143573 47675 146557
rect 44675 143565 47675 143573
rect 47865 146557 50865 146565
rect 47865 143573 47873 146557
rect 50857 143573 50865 146557
rect 47865 143565 50865 143573
rect 51055 146557 54055 146565
rect 51055 143573 51063 146557
rect 54047 143573 54055 146557
rect 51055 143565 54055 143573
rect 54245 146557 57245 146565
rect 54245 143573 54253 146557
rect 57237 143573 57245 146557
rect 54245 143565 57245 143573
rect 57435 146557 60435 146565
rect 57435 143573 57443 146557
rect 60427 143573 60435 146557
rect 57435 143565 60435 143573
rect 60625 146557 63625 146565
rect 60625 143573 60633 146557
rect 63617 143573 63625 146557
rect 60625 143565 63625 143573
rect 63815 146557 66815 146565
rect 63815 143573 63823 146557
rect 66807 143573 66815 146557
rect 63815 143565 66815 143573
rect 67005 146557 70005 146565
rect 67005 143573 67013 146557
rect 69997 143573 70005 146557
rect 67005 143565 70005 143573
rect 70195 146557 73195 146565
rect 70195 143573 70203 146557
rect 73187 143573 73195 146557
rect 70195 143565 73195 143573
rect 73385 146557 76385 146565
rect 73385 143573 73393 146557
rect 76377 143573 76385 146557
rect 73385 143565 76385 143573
rect 76575 146557 79575 146565
rect 76575 143573 76583 146557
rect 79567 143573 79575 146557
rect 76575 143565 79575 143573
rect 79765 146557 82765 146565
rect 79765 143573 79773 146557
rect 82757 143573 82765 146557
rect 79765 143565 82765 143573
rect 82955 146557 85955 146565
rect 82955 143573 82963 146557
rect 85947 143573 85955 146557
rect 82955 143565 85955 143573
rect 86145 146557 89145 146565
rect 86145 143573 86153 146557
rect 89137 143573 89145 146557
rect 86145 143565 89145 143573
rect 89335 146557 92335 146565
rect 89335 143573 89343 146557
rect 92327 143573 92335 146557
rect 89335 143565 92335 143573
rect 92525 146557 95525 146565
rect 92525 143573 92533 146557
rect 95517 143573 95525 146557
rect 92525 143565 95525 143573
rect 95715 146557 98715 146565
rect 95715 143573 95723 146557
rect 98707 143573 98715 146557
rect 95715 143565 98715 143573
rect 98905 146557 101905 146565
rect 98905 143573 98913 146557
rect 101897 143573 101905 146557
rect 98905 143565 101905 143573
rect 102095 146557 105095 146565
rect 102095 143573 102103 146557
rect 105087 143573 105095 146557
rect 102095 143565 105095 143573
rect 105285 146557 108285 146565
rect 105285 143573 105293 146557
rect 108277 143573 108285 146557
rect 105285 143565 108285 143573
rect 108475 146557 111475 146565
rect 108475 143573 108483 146557
rect 111467 143573 111475 146557
rect 108475 143565 111475 143573
rect 111665 146557 114665 146565
rect 111665 143573 111673 146557
rect 114657 143573 114665 146557
rect 111665 143565 114665 143573
rect 114855 146557 117855 146565
rect 114855 143573 114863 146557
rect 117847 143573 117855 146557
rect 114855 143565 117855 143573
rect 118045 146557 121045 146565
rect 118045 143573 118053 146557
rect 121037 143573 121045 146557
rect 118045 143565 121045 143573
rect 121235 146557 124235 146565
rect 121235 143573 121243 146557
rect 124227 143573 124235 146557
rect 121235 143565 124235 143573
rect 124425 146557 127425 146565
rect 124425 143573 124433 146557
rect 127417 143573 127425 146557
rect 124425 143565 127425 143573
rect 127615 146557 130615 146565
rect 127615 143573 127623 146557
rect 130607 143573 130615 146557
rect 127615 143565 130615 143573
rect 130805 146557 133805 146565
rect 130805 143573 130813 146557
rect 133797 143573 133805 146557
rect 130805 143565 133805 143573
rect 133995 146557 136995 146565
rect 133995 143573 134003 146557
rect 136987 143573 136995 146557
rect 133995 143565 136995 143573
rect 15 143367 3015 143375
rect 15 140383 23 143367
rect 3007 140383 3015 143367
rect 15 140375 3015 140383
rect 3205 143367 6205 143375
rect 3205 140383 3213 143367
rect 6197 140383 6205 143367
rect 3205 140375 6205 140383
rect 6395 143367 9395 143375
rect 6395 140383 6403 143367
rect 9387 140383 9395 143367
rect 6395 140375 9395 140383
rect 9585 143367 12585 143375
rect 9585 140383 9593 143367
rect 12577 140383 12585 143367
rect 9585 140375 12585 140383
rect 12775 143367 15775 143375
rect 12775 140383 12783 143367
rect 15767 140383 15775 143367
rect 12775 140375 15775 140383
rect 15965 143367 18965 143375
rect 15965 140383 15973 143367
rect 18957 140383 18965 143367
rect 15965 140375 18965 140383
rect 19155 143367 22155 143375
rect 19155 140383 19163 143367
rect 22147 140383 22155 143367
rect 19155 140375 22155 140383
rect 22345 143367 25345 143375
rect 22345 140383 22353 143367
rect 25337 140383 25345 143367
rect 22345 140375 25345 140383
rect 25535 143367 28535 143375
rect 25535 140383 25543 143367
rect 28527 140383 28535 143367
rect 25535 140375 28535 140383
rect 28725 143367 31725 143375
rect 28725 140383 28733 143367
rect 31717 140383 31725 143367
rect 28725 140375 31725 140383
rect 31915 143367 34915 143375
rect 31915 140383 31923 143367
rect 34907 140383 34915 143367
rect 31915 140375 34915 140383
rect 35105 143367 38105 143375
rect 35105 140383 35113 143367
rect 38097 140383 38105 143367
rect 35105 140375 38105 140383
rect 38295 143367 41295 143375
rect 38295 140383 38303 143367
rect 41287 140383 41295 143367
rect 38295 140375 41295 140383
rect 41485 143367 44485 143375
rect 41485 140383 41493 143367
rect 44477 140383 44485 143367
rect 41485 140375 44485 140383
rect 44675 143367 47675 143375
rect 44675 140383 44683 143367
rect 47667 140383 47675 143367
rect 44675 140375 47675 140383
rect 47865 143367 50865 143375
rect 47865 140383 47873 143367
rect 50857 140383 50865 143367
rect 47865 140375 50865 140383
rect 51055 143367 54055 143375
rect 51055 140383 51063 143367
rect 54047 140383 54055 143367
rect 51055 140375 54055 140383
rect 54245 143367 57245 143375
rect 54245 140383 54253 143367
rect 57237 140383 57245 143367
rect 54245 140375 57245 140383
rect 57435 143367 60435 143375
rect 57435 140383 57443 143367
rect 60427 140383 60435 143367
rect 57435 140375 60435 140383
rect 60625 143367 63625 143375
rect 60625 140383 60633 143367
rect 63617 140383 63625 143367
rect 60625 140375 63625 140383
rect 63815 143367 66815 143375
rect 63815 140383 63823 143367
rect 66807 140383 66815 143367
rect 63815 140375 66815 140383
rect 67005 143367 70005 143375
rect 67005 140383 67013 143367
rect 69997 140383 70005 143367
rect 67005 140375 70005 140383
rect 70195 143367 73195 143375
rect 70195 140383 70203 143367
rect 73187 140383 73195 143367
rect 70195 140375 73195 140383
rect 73385 143367 76385 143375
rect 73385 140383 73393 143367
rect 76377 140383 76385 143367
rect 73385 140375 76385 140383
rect 76575 143367 79575 143375
rect 76575 140383 76583 143367
rect 79567 140383 79575 143367
rect 76575 140375 79575 140383
rect 79765 143367 82765 143375
rect 79765 140383 79773 143367
rect 82757 140383 82765 143367
rect 79765 140375 82765 140383
rect 82955 143367 85955 143375
rect 82955 140383 82963 143367
rect 85947 140383 85955 143367
rect 82955 140375 85955 140383
rect 86145 143367 89145 143375
rect 86145 140383 86153 143367
rect 89137 140383 89145 143367
rect 86145 140375 89145 140383
rect 89335 143367 92335 143375
rect 89335 140383 89343 143367
rect 92327 140383 92335 143367
rect 89335 140375 92335 140383
rect 92525 143367 95525 143375
rect 92525 140383 92533 143367
rect 95517 140383 95525 143367
rect 92525 140375 95525 140383
rect 95715 143367 98715 143375
rect 95715 140383 95723 143367
rect 98707 140383 98715 143367
rect 95715 140375 98715 140383
rect 98905 143367 101905 143375
rect 98905 140383 98913 143367
rect 101897 140383 101905 143367
rect 98905 140375 101905 140383
rect 102095 143367 105095 143375
rect 102095 140383 102103 143367
rect 105087 140383 105095 143367
rect 102095 140375 105095 140383
rect 105285 143367 108285 143375
rect 105285 140383 105293 143367
rect 108277 140383 108285 143367
rect 105285 140375 108285 140383
rect 108475 143367 111475 143375
rect 108475 140383 108483 143367
rect 111467 140383 111475 143367
rect 108475 140375 111475 140383
rect 111665 143367 114665 143375
rect 111665 140383 111673 143367
rect 114657 140383 114665 143367
rect 111665 140375 114665 140383
rect 114855 143367 117855 143375
rect 114855 140383 114863 143367
rect 117847 140383 117855 143367
rect 114855 140375 117855 140383
rect 118045 143367 121045 143375
rect 118045 140383 118053 143367
rect 121037 140383 121045 143367
rect 118045 140375 121045 140383
rect 121235 143367 124235 143375
rect 121235 140383 121243 143367
rect 124227 140383 124235 143367
rect 121235 140375 124235 140383
rect 124425 143367 127425 143375
rect 124425 140383 124433 143367
rect 127417 140383 127425 143367
rect 124425 140375 127425 140383
rect 127615 143367 130615 143375
rect 127615 140383 127623 143367
rect 130607 140383 130615 143367
rect 127615 140375 130615 140383
rect 130805 143367 133805 143375
rect 130805 140383 130813 143367
rect 133797 140383 133805 143367
rect 130805 140375 133805 140383
rect 133995 143367 136995 143375
rect 133995 140383 134003 143367
rect 136987 140383 136995 143367
rect 133995 140375 136995 140383
rect 9585 140177 12585 140185
rect 9585 137193 9593 140177
rect 12577 137193 12585 140177
rect 9585 137185 12585 137193
rect 12775 140177 15775 140185
rect 12775 137193 12783 140177
rect 15767 137193 15775 140177
rect 12775 137185 15775 137193
rect 15965 140177 18965 140185
rect 15965 137193 15973 140177
rect 18957 137193 18965 140177
rect 15965 137185 18965 137193
rect 19155 140177 22155 140185
rect 19155 137193 19163 140177
rect 22147 137193 22155 140177
rect 19155 137185 22155 137193
rect 22345 140177 25345 140185
rect 22345 137193 22353 140177
rect 25337 137193 25345 140177
rect 22345 137185 25345 137193
rect 25535 140177 28535 140185
rect 25535 137193 25543 140177
rect 28527 137193 28535 140177
rect 25535 137185 28535 137193
rect 28725 140177 31725 140185
rect 28725 137193 28733 140177
rect 31717 137193 31725 140177
rect 28725 137185 31725 137193
rect 31915 140177 34915 140185
rect 31915 137193 31923 140177
rect 34907 137193 34915 140177
rect 31915 137185 34915 137193
rect 35105 140177 38105 140185
rect 35105 137193 35113 140177
rect 38097 137193 38105 140177
rect 35105 137185 38105 137193
rect 38295 140177 41295 140185
rect 38295 137193 38303 140177
rect 41287 137193 41295 140177
rect 38295 137185 41295 137193
rect 41485 140177 44485 140185
rect 41485 137193 41493 140177
rect 44477 137193 44485 140177
rect 41485 137185 44485 137193
rect 44675 140177 47675 140185
rect 44675 137193 44683 140177
rect 47667 137193 47675 140177
rect 44675 137185 47675 137193
rect 47865 140177 50865 140185
rect 47865 137193 47873 140177
rect 50857 137193 50865 140177
rect 47865 137185 50865 137193
rect 51055 140177 54055 140185
rect 51055 137193 51063 140177
rect 54047 137193 54055 140177
rect 51055 137185 54055 137193
rect 54245 140177 57245 140185
rect 54245 137193 54253 140177
rect 57237 137193 57245 140177
rect 54245 137185 57245 137193
rect 57435 140177 60435 140185
rect 57435 137193 57443 140177
rect 60427 137193 60435 140177
rect 57435 137185 60435 137193
rect 60625 140177 63625 140185
rect 60625 137193 60633 140177
rect 63617 137193 63625 140177
rect 60625 137185 63625 137193
rect 63815 140177 66815 140185
rect 63815 137193 63823 140177
rect 66807 137193 66815 140177
rect 63815 137185 66815 137193
rect 67005 140177 70005 140185
rect 67005 137193 67013 140177
rect 69997 137193 70005 140177
rect 67005 137185 70005 137193
rect 70195 140177 73195 140185
rect 70195 137193 70203 140177
rect 73187 137193 73195 140177
rect 70195 137185 73195 137193
rect 73385 140177 76385 140185
rect 73385 137193 73393 140177
rect 76377 137193 76385 140177
rect 73385 137185 76385 137193
rect 76575 140177 79575 140185
rect 76575 137193 76583 140177
rect 79567 137193 79575 140177
rect 76575 137185 79575 137193
rect 79765 140177 82765 140185
rect 79765 137193 79773 140177
rect 82757 137193 82765 140177
rect 79765 137185 82765 137193
rect 82955 140177 85955 140185
rect 82955 137193 82963 140177
rect 85947 137193 85955 140177
rect 82955 137185 85955 137193
rect 86145 140177 89145 140185
rect 86145 137193 86153 140177
rect 89137 137193 89145 140177
rect 86145 137185 89145 137193
rect 89335 140177 92335 140185
rect 89335 137193 89343 140177
rect 92327 137193 92335 140177
rect 89335 137185 92335 137193
rect 92525 140177 95525 140185
rect 92525 137193 92533 140177
rect 95517 137193 95525 140177
rect 92525 137185 95525 137193
rect 95715 140177 98715 140185
rect 95715 137193 95723 140177
rect 98707 137193 98715 140177
rect 95715 137185 98715 137193
rect 98905 140177 101905 140185
rect 98905 137193 98913 140177
rect 101897 137193 101905 140177
rect 98905 137185 101905 137193
rect 102095 140177 105095 140185
rect 102095 137193 102103 140177
rect 105087 137193 105095 140177
rect 102095 137185 105095 137193
rect 105285 140177 108285 140185
rect 105285 137193 105293 140177
rect 108277 137193 108285 140177
rect 105285 137185 108285 137193
rect 108475 140177 111475 140185
rect 108475 137193 108483 140177
rect 111467 137193 111475 140177
rect 108475 137185 111475 137193
rect 111665 140177 114665 140185
rect 111665 137193 111673 140177
rect 114657 137193 114665 140177
rect 111665 137185 114665 137193
rect 114855 140177 117855 140185
rect 114855 137193 114863 140177
rect 117847 137193 117855 140177
rect 114855 137185 117855 137193
rect 118045 140177 121045 140185
rect 118045 137193 118053 140177
rect 121037 137193 121045 140177
rect 118045 137185 121045 137193
rect 121235 140177 124235 140185
rect 121235 137193 121243 140177
rect 124227 137193 124235 140177
rect 121235 137185 124235 137193
rect 124425 140177 127425 140185
rect 124425 137193 124433 140177
rect 127417 137193 127425 140177
rect 124425 137185 127425 137193
rect 127615 140177 130615 140185
rect 127615 137193 127623 140177
rect 130607 137193 130615 140177
rect 127615 137185 130615 137193
rect 130805 140177 133805 140185
rect 130805 137193 130813 140177
rect 133797 137193 133805 140177
rect 130805 137185 133805 137193
rect 133995 140177 136995 140185
rect 133995 137193 134003 140177
rect 136987 137193 136995 140177
rect 133995 137185 136995 137193
rect 9585 136987 12585 136995
rect 9585 134003 9593 136987
rect 12577 134003 12585 136987
rect 9585 133995 12585 134003
rect 12775 136987 15775 136995
rect 12775 134003 12783 136987
rect 15767 134003 15775 136987
rect 12775 133995 15775 134003
rect 15965 136987 18965 136995
rect 15965 134003 15973 136987
rect 18957 134003 18965 136987
rect 15965 133995 18965 134003
rect 19155 136987 22155 136995
rect 19155 134003 19163 136987
rect 22147 134003 22155 136987
rect 19155 133995 22155 134003
rect 22345 136987 25345 136995
rect 22345 134003 22353 136987
rect 25337 134003 25345 136987
rect 22345 133995 25345 134003
rect 25535 136987 28535 136995
rect 25535 134003 25543 136987
rect 28527 134003 28535 136987
rect 25535 133995 28535 134003
rect 28725 136987 31725 136995
rect 28725 134003 28733 136987
rect 31717 134003 31725 136987
rect 28725 133995 31725 134003
rect 31915 136987 34915 136995
rect 31915 134003 31923 136987
rect 34907 134003 34915 136987
rect 31915 133995 34915 134003
rect 35105 136987 38105 136995
rect 35105 134003 35113 136987
rect 38097 134003 38105 136987
rect 35105 133995 38105 134003
rect 38295 136987 41295 136995
rect 38295 134003 38303 136987
rect 41287 134003 41295 136987
rect 38295 133995 41295 134003
rect 41485 136987 44485 136995
rect 41485 134003 41493 136987
rect 44477 134003 44485 136987
rect 41485 133995 44485 134003
rect 44675 136987 47675 136995
rect 44675 134003 44683 136987
rect 47667 134003 47675 136987
rect 44675 133995 47675 134003
rect 47865 136987 50865 136995
rect 47865 134003 47873 136987
rect 50857 134003 50865 136987
rect 47865 133995 50865 134003
rect 51055 136987 54055 136995
rect 51055 134003 51063 136987
rect 54047 134003 54055 136987
rect 51055 133995 54055 134003
rect 54245 136987 57245 136995
rect 54245 134003 54253 136987
rect 57237 134003 57245 136987
rect 54245 133995 57245 134003
rect 57435 136987 60435 136995
rect 57435 134003 57443 136987
rect 60427 134003 60435 136987
rect 57435 133995 60435 134003
rect 60625 136987 63625 136995
rect 60625 134003 60633 136987
rect 63617 134003 63625 136987
rect 60625 133995 63625 134003
rect 63815 136987 66815 136995
rect 63815 134003 63823 136987
rect 66807 134003 66815 136987
rect 63815 133995 66815 134003
rect 67005 136987 70005 136995
rect 67005 134003 67013 136987
rect 69997 134003 70005 136987
rect 67005 133995 70005 134003
rect 70195 136987 73195 136995
rect 70195 134003 70203 136987
rect 73187 134003 73195 136987
rect 70195 133995 73195 134003
rect 73385 136987 76385 136995
rect 73385 134003 73393 136987
rect 76377 134003 76385 136987
rect 73385 133995 76385 134003
rect 76575 136987 79575 136995
rect 76575 134003 76583 136987
rect 79567 134003 79575 136987
rect 76575 133995 79575 134003
rect 79765 136987 82765 136995
rect 79765 134003 79773 136987
rect 82757 134003 82765 136987
rect 79765 133995 82765 134003
rect 82955 136987 85955 136995
rect 82955 134003 82963 136987
rect 85947 134003 85955 136987
rect 82955 133995 85955 134003
rect 86145 136987 89145 136995
rect 86145 134003 86153 136987
rect 89137 134003 89145 136987
rect 86145 133995 89145 134003
rect 89335 136987 92335 136995
rect 89335 134003 89343 136987
rect 92327 134003 92335 136987
rect 89335 133995 92335 134003
rect 92525 136987 95525 136995
rect 92525 134003 92533 136987
rect 95517 134003 95525 136987
rect 92525 133995 95525 134003
rect 95715 136987 98715 136995
rect 95715 134003 95723 136987
rect 98707 134003 98715 136987
rect 95715 133995 98715 134003
rect 98905 136987 101905 136995
rect 98905 134003 98913 136987
rect 101897 134003 101905 136987
rect 98905 133995 101905 134003
rect 102095 136987 105095 136995
rect 102095 134003 102103 136987
rect 105087 134003 105095 136987
rect 102095 133995 105095 134003
rect 105285 136987 108285 136995
rect 105285 134003 105293 136987
rect 108277 134003 108285 136987
rect 105285 133995 108285 134003
rect 108475 136987 111475 136995
rect 108475 134003 108483 136987
rect 111467 134003 111475 136987
rect 108475 133995 111475 134003
rect 111665 136987 114665 136995
rect 111665 134003 111673 136987
rect 114657 134003 114665 136987
rect 111665 133995 114665 134003
rect 114855 136987 117855 136995
rect 114855 134003 114863 136987
rect 117847 134003 117855 136987
rect 114855 133995 117855 134003
rect 118045 136987 121045 136995
rect 118045 134003 118053 136987
rect 121037 134003 121045 136987
rect 118045 133995 121045 134003
rect 121235 136987 124235 136995
rect 121235 134003 121243 136987
rect 124227 134003 124235 136987
rect 121235 133995 124235 134003
rect 124425 136987 127425 136995
rect 124425 134003 124433 136987
rect 127417 134003 127425 136987
rect 124425 133995 127425 134003
rect 127615 136987 130615 136995
rect 127615 134003 127623 136987
rect 130607 134003 130615 136987
rect 127615 133995 130615 134003
rect 130805 136987 133805 136995
rect 130805 134003 130813 136987
rect 133797 134003 133805 136987
rect 130805 133995 133805 134003
rect 133995 136987 136995 136995
rect 133995 134003 134003 136987
rect 136987 134003 136995 136987
rect 133995 133995 136995 134003
rect 9585 133797 12585 133805
rect 9585 130813 9593 133797
rect 12577 130813 12585 133797
rect 9585 130805 12585 130813
rect 12775 133797 15775 133805
rect 12775 130813 12783 133797
rect 15767 130813 15775 133797
rect 12775 130805 15775 130813
rect 15965 133797 18965 133805
rect 15965 130813 15973 133797
rect 18957 130813 18965 133797
rect 15965 130805 18965 130813
rect 19155 133797 22155 133805
rect 19155 130813 19163 133797
rect 22147 130813 22155 133797
rect 19155 130805 22155 130813
rect 22345 133797 25345 133805
rect 22345 130813 22353 133797
rect 25337 130813 25345 133797
rect 22345 130805 25345 130813
rect 25535 133797 28535 133805
rect 25535 130813 25543 133797
rect 28527 130813 28535 133797
rect 25535 130805 28535 130813
rect 28725 133797 31725 133805
rect 28725 130813 28733 133797
rect 31717 130813 31725 133797
rect 28725 130805 31725 130813
rect 31915 133797 34915 133805
rect 31915 130813 31923 133797
rect 34907 130813 34915 133797
rect 31915 130805 34915 130813
rect 35105 133797 38105 133805
rect 35105 130813 35113 133797
rect 38097 130813 38105 133797
rect 35105 130805 38105 130813
rect 38295 133797 41295 133805
rect 38295 130813 38303 133797
rect 41287 130813 41295 133797
rect 38295 130805 41295 130813
rect 41485 133797 44485 133805
rect 41485 130813 41493 133797
rect 44477 130813 44485 133797
rect 41485 130805 44485 130813
rect 44675 133797 47675 133805
rect 44675 130813 44683 133797
rect 47667 130813 47675 133797
rect 44675 130805 47675 130813
rect 47865 133797 50865 133805
rect 47865 130813 47873 133797
rect 50857 130813 50865 133797
rect 47865 130805 50865 130813
rect 51055 133797 54055 133805
rect 51055 130813 51063 133797
rect 54047 130813 54055 133797
rect 51055 130805 54055 130813
rect 54245 133797 57245 133805
rect 54245 130813 54253 133797
rect 57237 130813 57245 133797
rect 54245 130805 57245 130813
rect 57435 133797 60435 133805
rect 57435 130813 57443 133797
rect 60427 130813 60435 133797
rect 57435 130805 60435 130813
rect 60625 133797 63625 133805
rect 60625 130813 60633 133797
rect 63617 130813 63625 133797
rect 60625 130805 63625 130813
rect 63815 133797 66815 133805
rect 63815 130813 63823 133797
rect 66807 130813 66815 133797
rect 63815 130805 66815 130813
rect 67005 133797 70005 133805
rect 67005 130813 67013 133797
rect 69997 130813 70005 133797
rect 67005 130805 70005 130813
rect 70195 133797 73195 133805
rect 70195 130813 70203 133797
rect 73187 130813 73195 133797
rect 70195 130805 73195 130813
rect 73385 133797 76385 133805
rect 73385 130813 73393 133797
rect 76377 130813 76385 133797
rect 73385 130805 76385 130813
rect 76575 133797 79575 133805
rect 76575 130813 76583 133797
rect 79567 130813 79575 133797
rect 76575 130805 79575 130813
rect 79765 133797 82765 133805
rect 79765 130813 79773 133797
rect 82757 130813 82765 133797
rect 79765 130805 82765 130813
rect 82955 133797 85955 133805
rect 82955 130813 82963 133797
rect 85947 130813 85955 133797
rect 82955 130805 85955 130813
rect 86145 133797 89145 133805
rect 86145 130813 86153 133797
rect 89137 130813 89145 133797
rect 86145 130805 89145 130813
rect 89335 133797 92335 133805
rect 89335 130813 89343 133797
rect 92327 130813 92335 133797
rect 89335 130805 92335 130813
rect 92525 133797 95525 133805
rect 92525 130813 92533 133797
rect 95517 130813 95525 133797
rect 92525 130805 95525 130813
rect 95715 133797 98715 133805
rect 95715 130813 95723 133797
rect 98707 130813 98715 133797
rect 95715 130805 98715 130813
rect 98905 133797 101905 133805
rect 98905 130813 98913 133797
rect 101897 130813 101905 133797
rect 98905 130805 101905 130813
rect 102095 133797 105095 133805
rect 102095 130813 102103 133797
rect 105087 130813 105095 133797
rect 102095 130805 105095 130813
rect 105285 133797 108285 133805
rect 105285 130813 105293 133797
rect 108277 130813 108285 133797
rect 105285 130805 108285 130813
rect 108475 133797 111475 133805
rect 108475 130813 108483 133797
rect 111467 130813 111475 133797
rect 108475 130805 111475 130813
rect 111665 133797 114665 133805
rect 111665 130813 111673 133797
rect 114657 130813 114665 133797
rect 111665 130805 114665 130813
rect 114855 133797 117855 133805
rect 114855 130813 114863 133797
rect 117847 130813 117855 133797
rect 114855 130805 117855 130813
rect 118045 133797 121045 133805
rect 118045 130813 118053 133797
rect 121037 130813 121045 133797
rect 118045 130805 121045 130813
rect 121235 133797 124235 133805
rect 121235 130813 121243 133797
rect 124227 130813 124235 133797
rect 121235 130805 124235 130813
rect 124425 133797 127425 133805
rect 124425 130813 124433 133797
rect 127417 130813 127425 133797
rect 124425 130805 127425 130813
rect 127615 133797 130615 133805
rect 127615 130813 127623 133797
rect 130607 130813 130615 133797
rect 127615 130805 130615 130813
rect 130805 133797 133805 133805
rect 130805 130813 130813 133797
rect 133797 130813 133805 133797
rect 130805 130805 133805 130813
rect 133995 133797 136995 133805
rect 133995 130813 134003 133797
rect 136987 130813 136995 133797
rect 133995 130805 136995 130813
rect 9585 130607 12585 130615
rect 9585 127623 9593 130607
rect 12577 127623 12585 130607
rect 9585 127615 12585 127623
rect 12775 130607 15775 130615
rect 12775 127623 12783 130607
rect 15767 127623 15775 130607
rect 12775 127615 15775 127623
rect 15965 130607 18965 130615
rect 15965 127623 15973 130607
rect 18957 127623 18965 130607
rect 15965 127615 18965 127623
rect 19155 130607 22155 130615
rect 19155 127623 19163 130607
rect 22147 127623 22155 130607
rect 19155 127615 22155 127623
rect 22345 130607 25345 130615
rect 22345 127623 22353 130607
rect 25337 127623 25345 130607
rect 22345 127615 25345 127623
rect 25535 130607 28535 130615
rect 25535 127623 25543 130607
rect 28527 127623 28535 130607
rect 25535 127615 28535 127623
rect 28725 130607 31725 130615
rect 28725 127623 28733 130607
rect 31717 127623 31725 130607
rect 28725 127615 31725 127623
rect 31915 130607 34915 130615
rect 31915 127623 31923 130607
rect 34907 127623 34915 130607
rect 31915 127615 34915 127623
rect 35105 130607 38105 130615
rect 35105 127623 35113 130607
rect 38097 127623 38105 130607
rect 35105 127615 38105 127623
rect 38295 130607 41295 130615
rect 38295 127623 38303 130607
rect 41287 127623 41295 130607
rect 38295 127615 41295 127623
rect 41485 130607 44485 130615
rect 41485 127623 41493 130607
rect 44477 127623 44485 130607
rect 41485 127615 44485 127623
rect 44675 130607 47675 130615
rect 44675 127623 44683 130607
rect 47667 127623 47675 130607
rect 44675 127615 47675 127623
rect 47865 130607 50865 130615
rect 47865 127623 47873 130607
rect 50857 127623 50865 130607
rect 47865 127615 50865 127623
rect 51055 130607 54055 130615
rect 51055 127623 51063 130607
rect 54047 127623 54055 130607
rect 51055 127615 54055 127623
rect 54245 130607 57245 130615
rect 54245 127623 54253 130607
rect 57237 127623 57245 130607
rect 54245 127615 57245 127623
rect 57435 130607 60435 130615
rect 57435 127623 57443 130607
rect 60427 127623 60435 130607
rect 57435 127615 60435 127623
rect 60625 130607 63625 130615
rect 60625 127623 60633 130607
rect 63617 127623 63625 130607
rect 60625 127615 63625 127623
rect 63815 130607 66815 130615
rect 63815 127623 63823 130607
rect 66807 127623 66815 130607
rect 63815 127615 66815 127623
rect 67005 130607 70005 130615
rect 67005 127623 67013 130607
rect 69997 127623 70005 130607
rect 67005 127615 70005 127623
rect 70195 130607 73195 130615
rect 70195 127623 70203 130607
rect 73187 127623 73195 130607
rect 70195 127615 73195 127623
rect 73385 130607 76385 130615
rect 73385 127623 73393 130607
rect 76377 127623 76385 130607
rect 73385 127615 76385 127623
rect 76575 130607 79575 130615
rect 76575 127623 76583 130607
rect 79567 127623 79575 130607
rect 76575 127615 79575 127623
rect 79765 130607 82765 130615
rect 79765 127623 79773 130607
rect 82757 127623 82765 130607
rect 79765 127615 82765 127623
rect 82955 130607 85955 130615
rect 82955 127623 82963 130607
rect 85947 127623 85955 130607
rect 82955 127615 85955 127623
rect 86145 130607 89145 130615
rect 86145 127623 86153 130607
rect 89137 127623 89145 130607
rect 86145 127615 89145 127623
rect 89335 130607 92335 130615
rect 89335 127623 89343 130607
rect 92327 127623 92335 130607
rect 89335 127615 92335 127623
rect 92525 130607 95525 130615
rect 92525 127623 92533 130607
rect 95517 127623 95525 130607
rect 92525 127615 95525 127623
rect 95715 130607 98715 130615
rect 95715 127623 95723 130607
rect 98707 127623 98715 130607
rect 95715 127615 98715 127623
rect 98905 130607 101905 130615
rect 98905 127623 98913 130607
rect 101897 127623 101905 130607
rect 98905 127615 101905 127623
rect 102095 130607 105095 130615
rect 102095 127623 102103 130607
rect 105087 127623 105095 130607
rect 102095 127615 105095 127623
rect 105285 130607 108285 130615
rect 105285 127623 105293 130607
rect 108277 127623 108285 130607
rect 105285 127615 108285 127623
rect 108475 130607 111475 130615
rect 108475 127623 108483 130607
rect 111467 127623 111475 130607
rect 108475 127615 111475 127623
rect 111665 130607 114665 130615
rect 111665 127623 111673 130607
rect 114657 127623 114665 130607
rect 111665 127615 114665 127623
rect 114855 130607 117855 130615
rect 114855 127623 114863 130607
rect 117847 127623 117855 130607
rect 114855 127615 117855 127623
rect 118045 130607 121045 130615
rect 118045 127623 118053 130607
rect 121037 127623 121045 130607
rect 118045 127615 121045 127623
rect 121235 130607 124235 130615
rect 121235 127623 121243 130607
rect 124227 127623 124235 130607
rect 121235 127615 124235 127623
rect 124425 130607 127425 130615
rect 124425 127623 124433 130607
rect 127417 127623 127425 130607
rect 124425 127615 127425 127623
rect 127615 130607 130615 130615
rect 127615 127623 127623 130607
rect 130607 127623 130615 130607
rect 127615 127615 130615 127623
rect 130805 130607 133805 130615
rect 130805 127623 130813 130607
rect 133797 127623 133805 130607
rect 130805 127615 133805 127623
rect 133995 130607 136995 130615
rect 133995 127623 134003 130607
rect 136987 127623 136995 130607
rect 133995 127615 136995 127623
rect 9585 127417 12585 127425
rect 9585 124433 9593 127417
rect 12577 124433 12585 127417
rect 9585 124425 12585 124433
rect 12775 127417 15775 127425
rect 12775 124433 12783 127417
rect 15767 124433 15775 127417
rect 12775 124425 15775 124433
rect 15965 127417 18965 127425
rect 15965 124433 15973 127417
rect 18957 124433 18965 127417
rect 15965 124425 18965 124433
rect 19155 127417 22155 127425
rect 19155 124433 19163 127417
rect 22147 124433 22155 127417
rect 19155 124425 22155 124433
rect 22345 127417 25345 127425
rect 22345 124433 22353 127417
rect 25337 124433 25345 127417
rect 22345 124425 25345 124433
rect 25535 127417 28535 127425
rect 25535 124433 25543 127417
rect 28527 124433 28535 127417
rect 25535 124425 28535 124433
rect 28725 127417 31725 127425
rect 28725 124433 28733 127417
rect 31717 124433 31725 127417
rect 28725 124425 31725 124433
rect 31915 127417 34915 127425
rect 31915 124433 31923 127417
rect 34907 124433 34915 127417
rect 31915 124425 34915 124433
rect 35105 127417 38105 127425
rect 35105 124433 35113 127417
rect 38097 124433 38105 127417
rect 35105 124425 38105 124433
rect 38295 127417 41295 127425
rect 38295 124433 38303 127417
rect 41287 124433 41295 127417
rect 38295 124425 41295 124433
rect 41485 127417 44485 127425
rect 41485 124433 41493 127417
rect 44477 124433 44485 127417
rect 41485 124425 44485 124433
rect 44675 127417 47675 127425
rect 44675 124433 44683 127417
rect 47667 124433 47675 127417
rect 44675 124425 47675 124433
rect 47865 127417 50865 127425
rect 47865 124433 47873 127417
rect 50857 124433 50865 127417
rect 47865 124425 50865 124433
rect 51055 127417 54055 127425
rect 51055 124433 51063 127417
rect 54047 124433 54055 127417
rect 51055 124425 54055 124433
rect 54245 127417 57245 127425
rect 54245 124433 54253 127417
rect 57237 124433 57245 127417
rect 54245 124425 57245 124433
rect 57435 127417 60435 127425
rect 57435 124433 57443 127417
rect 60427 124433 60435 127417
rect 57435 124425 60435 124433
rect 60625 127417 63625 127425
rect 60625 124433 60633 127417
rect 63617 124433 63625 127417
rect 60625 124425 63625 124433
rect 63815 127417 66815 127425
rect 63815 124433 63823 127417
rect 66807 124433 66815 127417
rect 63815 124425 66815 124433
rect 67005 127417 70005 127425
rect 67005 124433 67013 127417
rect 69997 124433 70005 127417
rect 67005 124425 70005 124433
rect 70195 127417 73195 127425
rect 70195 124433 70203 127417
rect 73187 124433 73195 127417
rect 70195 124425 73195 124433
rect 73385 127417 76385 127425
rect 73385 124433 73393 127417
rect 76377 124433 76385 127417
rect 73385 124425 76385 124433
rect 76575 127417 79575 127425
rect 76575 124433 76583 127417
rect 79567 124433 79575 127417
rect 76575 124425 79575 124433
rect 79765 127417 82765 127425
rect 79765 124433 79773 127417
rect 82757 124433 82765 127417
rect 79765 124425 82765 124433
rect 82955 127417 85955 127425
rect 82955 124433 82963 127417
rect 85947 124433 85955 127417
rect 82955 124425 85955 124433
rect 86145 127417 89145 127425
rect 86145 124433 86153 127417
rect 89137 124433 89145 127417
rect 86145 124425 89145 124433
rect 89335 127417 92335 127425
rect 89335 124433 89343 127417
rect 92327 124433 92335 127417
rect 89335 124425 92335 124433
rect 92525 127417 95525 127425
rect 92525 124433 92533 127417
rect 95517 124433 95525 127417
rect 92525 124425 95525 124433
rect 95715 127417 98715 127425
rect 95715 124433 95723 127417
rect 98707 124433 98715 127417
rect 95715 124425 98715 124433
rect 98905 127417 101905 127425
rect 98905 124433 98913 127417
rect 101897 124433 101905 127417
rect 98905 124425 101905 124433
rect 102095 127417 105095 127425
rect 102095 124433 102103 127417
rect 105087 124433 105095 127417
rect 102095 124425 105095 124433
rect 105285 127417 108285 127425
rect 105285 124433 105293 127417
rect 108277 124433 108285 127417
rect 105285 124425 108285 124433
rect 108475 127417 111475 127425
rect 108475 124433 108483 127417
rect 111467 124433 111475 127417
rect 108475 124425 111475 124433
rect 111665 127417 114665 127425
rect 111665 124433 111673 127417
rect 114657 124433 114665 127417
rect 111665 124425 114665 124433
rect 114855 127417 117855 127425
rect 114855 124433 114863 127417
rect 117847 124433 117855 127417
rect 114855 124425 117855 124433
rect 118045 127417 121045 127425
rect 118045 124433 118053 127417
rect 121037 124433 121045 127417
rect 118045 124425 121045 124433
rect 121235 127417 124235 127425
rect 121235 124433 121243 127417
rect 124227 124433 124235 127417
rect 121235 124425 124235 124433
rect 124425 127417 127425 127425
rect 124425 124433 124433 127417
rect 127417 124433 127425 127417
rect 124425 124425 127425 124433
rect 127615 127417 130615 127425
rect 127615 124433 127623 127417
rect 130607 124433 130615 127417
rect 127615 124425 130615 124433
rect 130805 127417 133805 127425
rect 130805 124433 130813 127417
rect 133797 124433 133805 127417
rect 130805 124425 133805 124433
rect 133995 127417 136995 127425
rect 133995 124433 134003 127417
rect 136987 124433 136995 127417
rect 133995 124425 136995 124433
rect 9585 124227 12585 124235
rect 9585 121243 9593 124227
rect 12577 121243 12585 124227
rect 9585 121235 12585 121243
rect 12775 124227 15775 124235
rect 12775 121243 12783 124227
rect 15767 121243 15775 124227
rect 12775 121235 15775 121243
rect 15965 124227 18965 124235
rect 15965 121243 15973 124227
rect 18957 121243 18965 124227
rect 15965 121235 18965 121243
rect 19155 124227 22155 124235
rect 19155 121243 19163 124227
rect 22147 121243 22155 124227
rect 19155 121235 22155 121243
rect 22345 124227 25345 124235
rect 22345 121243 22353 124227
rect 25337 121243 25345 124227
rect 22345 121235 25345 121243
rect 25535 124227 28535 124235
rect 25535 121243 25543 124227
rect 28527 121243 28535 124227
rect 25535 121235 28535 121243
rect 28725 124227 31725 124235
rect 28725 121243 28733 124227
rect 31717 121243 31725 124227
rect 28725 121235 31725 121243
rect 31915 124227 34915 124235
rect 31915 121243 31923 124227
rect 34907 121243 34915 124227
rect 31915 121235 34915 121243
rect 35105 124227 38105 124235
rect 35105 121243 35113 124227
rect 38097 121243 38105 124227
rect 35105 121235 38105 121243
rect 38295 124227 41295 124235
rect 38295 121243 38303 124227
rect 41287 121243 41295 124227
rect 38295 121235 41295 121243
rect 41485 124227 44485 124235
rect 41485 121243 41493 124227
rect 44477 121243 44485 124227
rect 41485 121235 44485 121243
rect 44675 124227 47675 124235
rect 44675 121243 44683 124227
rect 47667 121243 47675 124227
rect 44675 121235 47675 121243
rect 47865 124227 50865 124235
rect 47865 121243 47873 124227
rect 50857 121243 50865 124227
rect 47865 121235 50865 121243
rect 51055 124227 54055 124235
rect 51055 121243 51063 124227
rect 54047 121243 54055 124227
rect 51055 121235 54055 121243
rect 54245 124227 57245 124235
rect 54245 121243 54253 124227
rect 57237 121243 57245 124227
rect 54245 121235 57245 121243
rect 57435 124227 60435 124235
rect 57435 121243 57443 124227
rect 60427 121243 60435 124227
rect 57435 121235 60435 121243
rect 60625 124227 63625 124235
rect 60625 121243 60633 124227
rect 63617 121243 63625 124227
rect 60625 121235 63625 121243
rect 63815 124227 66815 124235
rect 63815 121243 63823 124227
rect 66807 121243 66815 124227
rect 63815 121235 66815 121243
rect 67005 124227 70005 124235
rect 67005 121243 67013 124227
rect 69997 121243 70005 124227
rect 67005 121235 70005 121243
rect 70195 124227 73195 124235
rect 70195 121243 70203 124227
rect 73187 121243 73195 124227
rect 70195 121235 73195 121243
rect 73385 124227 76385 124235
rect 73385 121243 73393 124227
rect 76377 121243 76385 124227
rect 73385 121235 76385 121243
rect 76575 124227 79575 124235
rect 76575 121243 76583 124227
rect 79567 121243 79575 124227
rect 76575 121235 79575 121243
rect 79765 124227 82765 124235
rect 79765 121243 79773 124227
rect 82757 121243 82765 124227
rect 79765 121235 82765 121243
rect 82955 124227 85955 124235
rect 82955 121243 82963 124227
rect 85947 121243 85955 124227
rect 82955 121235 85955 121243
rect 86145 124227 89145 124235
rect 86145 121243 86153 124227
rect 89137 121243 89145 124227
rect 86145 121235 89145 121243
rect 89335 124227 92335 124235
rect 89335 121243 89343 124227
rect 92327 121243 92335 124227
rect 89335 121235 92335 121243
rect 92525 124227 95525 124235
rect 92525 121243 92533 124227
rect 95517 121243 95525 124227
rect 92525 121235 95525 121243
rect 95715 124227 98715 124235
rect 95715 121243 95723 124227
rect 98707 121243 98715 124227
rect 95715 121235 98715 121243
rect 98905 124227 101905 124235
rect 98905 121243 98913 124227
rect 101897 121243 101905 124227
rect 98905 121235 101905 121243
rect 102095 124227 105095 124235
rect 102095 121243 102103 124227
rect 105087 121243 105095 124227
rect 102095 121235 105095 121243
rect 105285 124227 108285 124235
rect 105285 121243 105293 124227
rect 108277 121243 108285 124227
rect 105285 121235 108285 121243
rect 108475 124227 111475 124235
rect 108475 121243 108483 124227
rect 111467 121243 111475 124227
rect 108475 121235 111475 121243
rect 111665 124227 114665 124235
rect 111665 121243 111673 124227
rect 114657 121243 114665 124227
rect 111665 121235 114665 121243
rect 114855 124227 117855 124235
rect 114855 121243 114863 124227
rect 117847 121243 117855 124227
rect 114855 121235 117855 121243
rect 118045 124227 121045 124235
rect 118045 121243 118053 124227
rect 121037 121243 121045 124227
rect 118045 121235 121045 121243
rect 121235 124227 124235 124235
rect 121235 121243 121243 124227
rect 124227 121243 124235 124227
rect 121235 121235 124235 121243
rect 124425 124227 127425 124235
rect 124425 121243 124433 124227
rect 127417 121243 127425 124227
rect 124425 121235 127425 121243
rect 127615 124227 130615 124235
rect 127615 121243 127623 124227
rect 130607 121243 130615 124227
rect 127615 121235 130615 121243
rect 130805 124227 133805 124235
rect 130805 121243 130813 124227
rect 133797 121243 133805 124227
rect 130805 121235 133805 121243
rect 133995 124227 136995 124235
rect 133995 121243 134003 124227
rect 136987 121243 136995 124227
rect 133995 121235 136995 121243
rect 15 121037 3015 121045
rect 15 118053 23 121037
rect 3007 118053 3015 121037
rect 15 118045 3015 118053
rect 3205 121037 6205 121045
rect 3205 118053 3213 121037
rect 6197 118053 6205 121037
rect 3205 118045 6205 118053
rect 6395 121037 9395 121045
rect 6395 118053 6403 121037
rect 9387 118053 9395 121037
rect 6395 118045 9395 118053
rect 9585 121037 12585 121045
rect 9585 118053 9593 121037
rect 12577 118053 12585 121037
rect 9585 118045 12585 118053
rect 12775 121037 15775 121045
rect 12775 118053 12783 121037
rect 15767 118053 15775 121037
rect 12775 118045 15775 118053
rect 15965 121037 18965 121045
rect 15965 118053 15973 121037
rect 18957 118053 18965 121037
rect 15965 118045 18965 118053
rect 19155 121037 22155 121045
rect 19155 118053 19163 121037
rect 22147 118053 22155 121037
rect 19155 118045 22155 118053
rect 22345 121037 25345 121045
rect 22345 118053 22353 121037
rect 25337 118053 25345 121037
rect 22345 118045 25345 118053
rect 25535 121037 28535 121045
rect 25535 118053 25543 121037
rect 28527 118053 28535 121037
rect 25535 118045 28535 118053
rect 28725 121037 31725 121045
rect 28725 118053 28733 121037
rect 31717 118053 31725 121037
rect 28725 118045 31725 118053
rect 31915 121037 34915 121045
rect 31915 118053 31923 121037
rect 34907 118053 34915 121037
rect 31915 118045 34915 118053
rect 35105 121037 38105 121045
rect 35105 118053 35113 121037
rect 38097 118053 38105 121037
rect 35105 118045 38105 118053
rect 38295 121037 41295 121045
rect 38295 118053 38303 121037
rect 41287 118053 41295 121037
rect 38295 118045 41295 118053
rect 41485 121037 44485 121045
rect 41485 118053 41493 121037
rect 44477 118053 44485 121037
rect 41485 118045 44485 118053
rect 44675 121037 47675 121045
rect 44675 118053 44683 121037
rect 47667 118053 47675 121037
rect 44675 118045 47675 118053
rect 47865 121037 50865 121045
rect 47865 118053 47873 121037
rect 50857 118053 50865 121037
rect 47865 118045 50865 118053
rect 51055 121037 54055 121045
rect 51055 118053 51063 121037
rect 54047 118053 54055 121037
rect 51055 118045 54055 118053
rect 54245 121037 57245 121045
rect 54245 118053 54253 121037
rect 57237 118053 57245 121037
rect 54245 118045 57245 118053
rect 57435 121037 60435 121045
rect 57435 118053 57443 121037
rect 60427 118053 60435 121037
rect 57435 118045 60435 118053
rect 60625 121037 63625 121045
rect 60625 118053 60633 121037
rect 63617 118053 63625 121037
rect 60625 118045 63625 118053
rect 63815 121037 66815 121045
rect 63815 118053 63823 121037
rect 66807 118053 66815 121037
rect 63815 118045 66815 118053
rect 67005 121037 70005 121045
rect 67005 118053 67013 121037
rect 69997 118053 70005 121037
rect 67005 118045 70005 118053
rect 70195 121037 73195 121045
rect 70195 118053 70203 121037
rect 73187 118053 73195 121037
rect 70195 118045 73195 118053
rect 73385 121037 76385 121045
rect 73385 118053 73393 121037
rect 76377 118053 76385 121037
rect 73385 118045 76385 118053
rect 76575 121037 79575 121045
rect 76575 118053 76583 121037
rect 79567 118053 79575 121037
rect 76575 118045 79575 118053
rect 79765 121037 82765 121045
rect 79765 118053 79773 121037
rect 82757 118053 82765 121037
rect 79765 118045 82765 118053
rect 82955 121037 85955 121045
rect 82955 118053 82963 121037
rect 85947 118053 85955 121037
rect 82955 118045 85955 118053
rect 86145 121037 89145 121045
rect 86145 118053 86153 121037
rect 89137 118053 89145 121037
rect 86145 118045 89145 118053
rect 89335 121037 92335 121045
rect 89335 118053 89343 121037
rect 92327 118053 92335 121037
rect 89335 118045 92335 118053
rect 92525 121037 95525 121045
rect 92525 118053 92533 121037
rect 95517 118053 95525 121037
rect 92525 118045 95525 118053
rect 95715 121037 98715 121045
rect 95715 118053 95723 121037
rect 98707 118053 98715 121037
rect 95715 118045 98715 118053
rect 98905 121037 101905 121045
rect 98905 118053 98913 121037
rect 101897 118053 101905 121037
rect 98905 118045 101905 118053
rect 102095 121037 105095 121045
rect 102095 118053 102103 121037
rect 105087 118053 105095 121037
rect 102095 118045 105095 118053
rect 105285 121037 108285 121045
rect 105285 118053 105293 121037
rect 108277 118053 108285 121037
rect 105285 118045 108285 118053
rect 108475 121037 111475 121045
rect 108475 118053 108483 121037
rect 111467 118053 111475 121037
rect 108475 118045 111475 118053
rect 111665 121037 114665 121045
rect 111665 118053 111673 121037
rect 114657 118053 114665 121037
rect 111665 118045 114665 118053
rect 114855 121037 117855 121045
rect 114855 118053 114863 121037
rect 117847 118053 117855 121037
rect 114855 118045 117855 118053
rect 118045 121037 121045 121045
rect 118045 118053 118053 121037
rect 121037 118053 121045 121037
rect 118045 118045 121045 118053
rect 121235 121037 124235 121045
rect 121235 118053 121243 121037
rect 124227 118053 124235 121037
rect 121235 118045 124235 118053
rect 124425 121037 127425 121045
rect 124425 118053 124433 121037
rect 127417 118053 127425 121037
rect 124425 118045 127425 118053
rect 127615 121037 130615 121045
rect 127615 118053 127623 121037
rect 130607 118053 130615 121037
rect 127615 118045 130615 118053
rect 130805 121037 133805 121045
rect 130805 118053 130813 121037
rect 133797 118053 133805 121037
rect 130805 118045 133805 118053
rect 133995 121037 136995 121045
rect 133995 118053 134003 121037
rect 136987 118053 136995 121037
rect 133995 118045 136995 118053
rect 15 117847 3015 117855
rect 15 114863 23 117847
rect 3007 114863 3015 117847
rect 15 114855 3015 114863
rect 3205 117847 6205 117855
rect 3205 114863 3213 117847
rect 6197 114863 6205 117847
rect 3205 114855 6205 114863
rect 6395 117847 9395 117855
rect 6395 114863 6403 117847
rect 9387 114863 9395 117847
rect 6395 114855 9395 114863
rect 9585 117847 12585 117855
rect 9585 114863 9593 117847
rect 12577 114863 12585 117847
rect 9585 114855 12585 114863
rect 12775 117847 15775 117855
rect 12775 114863 12783 117847
rect 15767 114863 15775 117847
rect 12775 114855 15775 114863
rect 15965 117847 18965 117855
rect 15965 114863 15973 117847
rect 18957 114863 18965 117847
rect 15965 114855 18965 114863
rect 19155 117847 22155 117855
rect 19155 114863 19163 117847
rect 22147 114863 22155 117847
rect 19155 114855 22155 114863
rect 22345 117847 25345 117855
rect 22345 114863 22353 117847
rect 25337 114863 25345 117847
rect 22345 114855 25345 114863
rect 25535 117847 28535 117855
rect 25535 114863 25543 117847
rect 28527 114863 28535 117847
rect 25535 114855 28535 114863
rect 28725 117847 31725 117855
rect 28725 114863 28733 117847
rect 31717 114863 31725 117847
rect 28725 114855 31725 114863
rect 31915 117847 34915 117855
rect 31915 114863 31923 117847
rect 34907 114863 34915 117847
rect 31915 114855 34915 114863
rect 35105 117847 38105 117855
rect 35105 114863 35113 117847
rect 38097 114863 38105 117847
rect 35105 114855 38105 114863
rect 38295 117847 41295 117855
rect 38295 114863 38303 117847
rect 41287 114863 41295 117847
rect 38295 114855 41295 114863
rect 41485 117847 44485 117855
rect 41485 114863 41493 117847
rect 44477 114863 44485 117847
rect 41485 114855 44485 114863
rect 44675 117847 47675 117855
rect 44675 114863 44683 117847
rect 47667 114863 47675 117847
rect 44675 114855 47675 114863
rect 47865 117847 50865 117855
rect 47865 114863 47873 117847
rect 50857 114863 50865 117847
rect 47865 114855 50865 114863
rect 51055 117847 54055 117855
rect 51055 114863 51063 117847
rect 54047 114863 54055 117847
rect 51055 114855 54055 114863
rect 54245 117847 57245 117855
rect 54245 114863 54253 117847
rect 57237 114863 57245 117847
rect 54245 114855 57245 114863
rect 57435 117847 60435 117855
rect 57435 114863 57443 117847
rect 60427 114863 60435 117847
rect 57435 114855 60435 114863
rect 60625 117847 63625 117855
rect 60625 114863 60633 117847
rect 63617 114863 63625 117847
rect 60625 114855 63625 114863
rect 63815 117847 66815 117855
rect 63815 114863 63823 117847
rect 66807 114863 66815 117847
rect 63815 114855 66815 114863
rect 67005 117847 70005 117855
rect 67005 114863 67013 117847
rect 69997 114863 70005 117847
rect 67005 114855 70005 114863
rect 70195 117847 73195 117855
rect 70195 114863 70203 117847
rect 73187 114863 73195 117847
rect 70195 114855 73195 114863
rect 73385 117847 76385 117855
rect 73385 114863 73393 117847
rect 76377 114863 76385 117847
rect 73385 114855 76385 114863
rect 76575 117847 79575 117855
rect 76575 114863 76583 117847
rect 79567 114863 79575 117847
rect 76575 114855 79575 114863
rect 79765 117847 82765 117855
rect 79765 114863 79773 117847
rect 82757 114863 82765 117847
rect 79765 114855 82765 114863
rect 82955 117847 85955 117855
rect 82955 114863 82963 117847
rect 85947 114863 85955 117847
rect 82955 114855 85955 114863
rect 86145 117847 89145 117855
rect 86145 114863 86153 117847
rect 89137 114863 89145 117847
rect 86145 114855 89145 114863
rect 89335 117847 92335 117855
rect 89335 114863 89343 117847
rect 92327 114863 92335 117847
rect 89335 114855 92335 114863
rect 92525 117847 95525 117855
rect 92525 114863 92533 117847
rect 95517 114863 95525 117847
rect 92525 114855 95525 114863
rect 95715 117847 98715 117855
rect 95715 114863 95723 117847
rect 98707 114863 98715 117847
rect 95715 114855 98715 114863
rect 98905 117847 101905 117855
rect 98905 114863 98913 117847
rect 101897 114863 101905 117847
rect 98905 114855 101905 114863
rect 102095 117847 105095 117855
rect 102095 114863 102103 117847
rect 105087 114863 105095 117847
rect 102095 114855 105095 114863
rect 105285 117847 108285 117855
rect 105285 114863 105293 117847
rect 108277 114863 108285 117847
rect 105285 114855 108285 114863
rect 108475 117847 111475 117855
rect 108475 114863 108483 117847
rect 111467 114863 111475 117847
rect 108475 114855 111475 114863
rect 111665 117847 114665 117855
rect 111665 114863 111673 117847
rect 114657 114863 114665 117847
rect 111665 114855 114665 114863
rect 114855 117847 117855 117855
rect 114855 114863 114863 117847
rect 117847 114863 117855 117847
rect 114855 114855 117855 114863
rect 118045 117847 121045 117855
rect 118045 114863 118053 117847
rect 121037 114863 121045 117847
rect 118045 114855 121045 114863
rect 121235 117847 124235 117855
rect 121235 114863 121243 117847
rect 124227 114863 124235 117847
rect 121235 114855 124235 114863
rect 124425 117847 127425 117855
rect 124425 114863 124433 117847
rect 127417 114863 127425 117847
rect 124425 114855 127425 114863
rect 127615 117847 130615 117855
rect 127615 114863 127623 117847
rect 130607 114863 130615 117847
rect 127615 114855 130615 114863
rect 130805 117847 133805 117855
rect 130805 114863 130813 117847
rect 133797 114863 133805 117847
rect 130805 114855 133805 114863
rect 133995 117847 136995 117855
rect 133995 114863 134003 117847
rect 136987 114863 136995 117847
rect 133995 114855 136995 114863
rect 15 114657 3015 114665
rect 15 111673 23 114657
rect 3007 111673 3015 114657
rect 15 111665 3015 111673
rect 3205 114657 6205 114665
rect 3205 111673 3213 114657
rect 6197 111673 6205 114657
rect 3205 111665 6205 111673
rect 6395 114657 9395 114665
rect 6395 111673 6403 114657
rect 9387 111673 9395 114657
rect 6395 111665 9395 111673
rect 9585 114657 12585 114665
rect 9585 111673 9593 114657
rect 12577 111673 12585 114657
rect 9585 111665 12585 111673
rect 12775 114657 15775 114665
rect 12775 111673 12783 114657
rect 15767 111673 15775 114657
rect 12775 111665 15775 111673
rect 15965 114657 18965 114665
rect 15965 111673 15973 114657
rect 18957 111673 18965 114657
rect 15965 111665 18965 111673
rect 19155 114657 22155 114665
rect 19155 111673 19163 114657
rect 22147 111673 22155 114657
rect 19155 111665 22155 111673
rect 22345 114657 25345 114665
rect 22345 111673 22353 114657
rect 25337 111673 25345 114657
rect 22345 111665 25345 111673
rect 25535 114657 28535 114665
rect 25535 111673 25543 114657
rect 28527 111673 28535 114657
rect 25535 111665 28535 111673
rect 28725 114657 31725 114665
rect 28725 111673 28733 114657
rect 31717 111673 31725 114657
rect 28725 111665 31725 111673
rect 31915 114657 34915 114665
rect 31915 111673 31923 114657
rect 34907 111673 34915 114657
rect 31915 111665 34915 111673
rect 35105 114657 38105 114665
rect 35105 111673 35113 114657
rect 38097 111673 38105 114657
rect 35105 111665 38105 111673
rect 38295 114657 41295 114665
rect 38295 111673 38303 114657
rect 41287 111673 41295 114657
rect 38295 111665 41295 111673
rect 41485 114657 44485 114665
rect 41485 111673 41493 114657
rect 44477 111673 44485 114657
rect 41485 111665 44485 111673
rect 44675 114657 47675 114665
rect 44675 111673 44683 114657
rect 47667 111673 47675 114657
rect 44675 111665 47675 111673
rect 47865 114657 50865 114665
rect 47865 111673 47873 114657
rect 50857 111673 50865 114657
rect 47865 111665 50865 111673
rect 51055 114657 54055 114665
rect 51055 111673 51063 114657
rect 54047 111673 54055 114657
rect 51055 111665 54055 111673
rect 54245 114657 57245 114665
rect 54245 111673 54253 114657
rect 57237 111673 57245 114657
rect 54245 111665 57245 111673
rect 57435 114657 60435 114665
rect 57435 111673 57443 114657
rect 60427 111673 60435 114657
rect 57435 111665 60435 111673
rect 60625 114657 63625 114665
rect 60625 111673 60633 114657
rect 63617 111673 63625 114657
rect 60625 111665 63625 111673
rect 63815 114657 66815 114665
rect 63815 111673 63823 114657
rect 66807 111673 66815 114657
rect 63815 111665 66815 111673
rect 67005 114657 70005 114665
rect 67005 111673 67013 114657
rect 69997 111673 70005 114657
rect 67005 111665 70005 111673
rect 70195 114657 73195 114665
rect 70195 111673 70203 114657
rect 73187 111673 73195 114657
rect 70195 111665 73195 111673
rect 73385 114657 76385 114665
rect 73385 111673 73393 114657
rect 76377 111673 76385 114657
rect 73385 111665 76385 111673
rect 76575 114657 79575 114665
rect 76575 111673 76583 114657
rect 79567 111673 79575 114657
rect 76575 111665 79575 111673
rect 79765 114657 82765 114665
rect 79765 111673 79773 114657
rect 82757 111673 82765 114657
rect 79765 111665 82765 111673
rect 82955 114657 85955 114665
rect 82955 111673 82963 114657
rect 85947 111673 85955 114657
rect 82955 111665 85955 111673
rect 86145 114657 89145 114665
rect 86145 111673 86153 114657
rect 89137 111673 89145 114657
rect 86145 111665 89145 111673
rect 89335 114657 92335 114665
rect 89335 111673 89343 114657
rect 92327 111673 92335 114657
rect 89335 111665 92335 111673
rect 92525 114657 95525 114665
rect 92525 111673 92533 114657
rect 95517 111673 95525 114657
rect 92525 111665 95525 111673
rect 95715 114657 98715 114665
rect 95715 111673 95723 114657
rect 98707 111673 98715 114657
rect 95715 111665 98715 111673
rect 98905 114657 101905 114665
rect 98905 111673 98913 114657
rect 101897 111673 101905 114657
rect 98905 111665 101905 111673
rect 102095 114657 105095 114665
rect 102095 111673 102103 114657
rect 105087 111673 105095 114657
rect 102095 111665 105095 111673
rect 105285 114657 108285 114665
rect 105285 111673 105293 114657
rect 108277 111673 108285 114657
rect 105285 111665 108285 111673
rect 108475 114657 111475 114665
rect 108475 111673 108483 114657
rect 111467 111673 111475 114657
rect 108475 111665 111475 111673
rect 111665 114657 114665 114665
rect 111665 111673 111673 114657
rect 114657 111673 114665 114657
rect 111665 111665 114665 111673
rect 114855 114657 117855 114665
rect 114855 111673 114863 114657
rect 117847 111673 117855 114657
rect 114855 111665 117855 111673
rect 118045 114657 121045 114665
rect 118045 111673 118053 114657
rect 121037 111673 121045 114657
rect 118045 111665 121045 111673
rect 121235 114657 124235 114665
rect 121235 111673 121243 114657
rect 124227 111673 124235 114657
rect 121235 111665 124235 111673
rect 124425 114657 127425 114665
rect 124425 111673 124433 114657
rect 127417 111673 127425 114657
rect 124425 111665 127425 111673
rect 127615 114657 130615 114665
rect 127615 111673 127623 114657
rect 130607 111673 130615 114657
rect 127615 111665 130615 111673
rect 130805 114657 133805 114665
rect 130805 111673 130813 114657
rect 133797 111673 133805 114657
rect 130805 111665 133805 111673
rect 133995 114657 136995 114665
rect 133995 111673 134003 114657
rect 136987 111673 136995 114657
rect 133995 111665 136995 111673
rect 15 111467 3015 111475
rect 15 108483 23 111467
rect 3007 108483 3015 111467
rect 15 108475 3015 108483
rect 3205 111467 6205 111475
rect 3205 108483 3213 111467
rect 6197 108483 6205 111467
rect 3205 108475 6205 108483
rect 6395 111467 9395 111475
rect 6395 108483 6403 111467
rect 9387 108483 9395 111467
rect 6395 108475 9395 108483
rect 9585 111467 12585 111475
rect 9585 108483 9593 111467
rect 12577 108483 12585 111467
rect 9585 108475 12585 108483
rect 12775 111467 15775 111475
rect 12775 108483 12783 111467
rect 15767 108483 15775 111467
rect 12775 108475 15775 108483
rect 15965 111467 18965 111475
rect 15965 108483 15973 111467
rect 18957 108483 18965 111467
rect 15965 108475 18965 108483
rect 19155 111467 22155 111475
rect 19155 108483 19163 111467
rect 22147 108483 22155 111467
rect 19155 108475 22155 108483
rect 22345 111467 25345 111475
rect 22345 108483 22353 111467
rect 25337 108483 25345 111467
rect 22345 108475 25345 108483
rect 25535 111467 28535 111475
rect 25535 108483 25543 111467
rect 28527 108483 28535 111467
rect 25535 108475 28535 108483
rect 28725 111467 31725 111475
rect 28725 108483 28733 111467
rect 31717 108483 31725 111467
rect 28725 108475 31725 108483
rect 31915 111467 34915 111475
rect 31915 108483 31923 111467
rect 34907 108483 34915 111467
rect 31915 108475 34915 108483
rect 35105 111467 38105 111475
rect 35105 108483 35113 111467
rect 38097 108483 38105 111467
rect 35105 108475 38105 108483
rect 38295 111467 41295 111475
rect 38295 108483 38303 111467
rect 41287 108483 41295 111467
rect 38295 108475 41295 108483
rect 41485 111467 44485 111475
rect 41485 108483 41493 111467
rect 44477 108483 44485 111467
rect 41485 108475 44485 108483
rect 44675 111467 47675 111475
rect 44675 108483 44683 111467
rect 47667 108483 47675 111467
rect 44675 108475 47675 108483
rect 47865 111467 50865 111475
rect 47865 108483 47873 111467
rect 50857 108483 50865 111467
rect 47865 108475 50865 108483
rect 51055 111467 54055 111475
rect 51055 108483 51063 111467
rect 54047 108483 54055 111467
rect 51055 108475 54055 108483
rect 54245 111467 57245 111475
rect 54245 108483 54253 111467
rect 57237 108483 57245 111467
rect 54245 108475 57245 108483
rect 57435 111467 60435 111475
rect 57435 108483 57443 111467
rect 60427 108483 60435 111467
rect 57435 108475 60435 108483
rect 60625 111467 63625 111475
rect 60625 108483 60633 111467
rect 63617 108483 63625 111467
rect 60625 108475 63625 108483
rect 63815 111467 66815 111475
rect 63815 108483 63823 111467
rect 66807 108483 66815 111467
rect 63815 108475 66815 108483
rect 67005 111467 70005 111475
rect 67005 108483 67013 111467
rect 69997 108483 70005 111467
rect 67005 108475 70005 108483
rect 70195 111467 73195 111475
rect 70195 108483 70203 111467
rect 73187 108483 73195 111467
rect 70195 108475 73195 108483
rect 73385 111467 76385 111475
rect 73385 108483 73393 111467
rect 76377 108483 76385 111467
rect 73385 108475 76385 108483
rect 76575 111467 79575 111475
rect 76575 108483 76583 111467
rect 79567 108483 79575 111467
rect 76575 108475 79575 108483
rect 79765 111467 82765 111475
rect 79765 108483 79773 111467
rect 82757 108483 82765 111467
rect 79765 108475 82765 108483
rect 82955 111467 85955 111475
rect 82955 108483 82963 111467
rect 85947 108483 85955 111467
rect 82955 108475 85955 108483
rect 86145 111467 89145 111475
rect 86145 108483 86153 111467
rect 89137 108483 89145 111467
rect 86145 108475 89145 108483
rect 89335 111467 92335 111475
rect 89335 108483 89343 111467
rect 92327 108483 92335 111467
rect 89335 108475 92335 108483
rect 92525 111467 95525 111475
rect 92525 108483 92533 111467
rect 95517 108483 95525 111467
rect 92525 108475 95525 108483
rect 95715 111467 98715 111475
rect 95715 108483 95723 111467
rect 98707 108483 98715 111467
rect 95715 108475 98715 108483
rect 98905 111467 101905 111475
rect 98905 108483 98913 111467
rect 101897 108483 101905 111467
rect 98905 108475 101905 108483
rect 102095 111467 105095 111475
rect 102095 108483 102103 111467
rect 105087 108483 105095 111467
rect 102095 108475 105095 108483
rect 105285 111467 108285 111475
rect 105285 108483 105293 111467
rect 108277 108483 108285 111467
rect 105285 108475 108285 108483
rect 108475 111467 111475 111475
rect 108475 108483 108483 111467
rect 111467 108483 111475 111467
rect 108475 108475 111475 108483
rect 111665 111467 114665 111475
rect 111665 108483 111673 111467
rect 114657 108483 114665 111467
rect 111665 108475 114665 108483
rect 114855 111467 117855 111475
rect 114855 108483 114863 111467
rect 117847 108483 117855 111467
rect 114855 108475 117855 108483
rect 118045 111467 121045 111475
rect 118045 108483 118053 111467
rect 121037 108483 121045 111467
rect 118045 108475 121045 108483
rect 121235 111467 124235 111475
rect 121235 108483 121243 111467
rect 124227 108483 124235 111467
rect 121235 108475 124235 108483
rect 124425 111467 127425 111475
rect 124425 108483 124433 111467
rect 127417 108483 127425 111467
rect 124425 108475 127425 108483
rect 127615 111467 130615 111475
rect 127615 108483 127623 111467
rect 130607 108483 130615 111467
rect 127615 108475 130615 108483
rect 130805 111467 133805 111475
rect 130805 108483 130813 111467
rect 133797 108483 133805 111467
rect 130805 108475 133805 108483
rect 133995 111467 136995 111475
rect 133995 108483 134003 111467
rect 136987 108483 136995 111467
rect 133995 108475 136995 108483
rect 15 108277 3015 108285
rect 15 105293 23 108277
rect 3007 105293 3015 108277
rect 15 105285 3015 105293
rect 3205 108277 6205 108285
rect 3205 105293 3213 108277
rect 6197 105293 6205 108277
rect 3205 105285 6205 105293
rect 6395 108277 9395 108285
rect 6395 105293 6403 108277
rect 9387 105293 9395 108277
rect 6395 105285 9395 105293
rect 9585 108277 12585 108285
rect 9585 105293 9593 108277
rect 12577 105293 12585 108277
rect 9585 105285 12585 105293
rect 12775 108277 15775 108285
rect 12775 105293 12783 108277
rect 15767 105293 15775 108277
rect 12775 105285 15775 105293
rect 15965 108277 18965 108285
rect 15965 105293 15973 108277
rect 18957 105293 18965 108277
rect 15965 105285 18965 105293
rect 19155 108277 22155 108285
rect 19155 105293 19163 108277
rect 22147 105293 22155 108277
rect 19155 105285 22155 105293
rect 22345 108277 25345 108285
rect 22345 105293 22353 108277
rect 25337 105293 25345 108277
rect 22345 105285 25345 105293
rect 25535 108277 28535 108285
rect 25535 105293 25543 108277
rect 28527 105293 28535 108277
rect 25535 105285 28535 105293
rect 28725 108277 31725 108285
rect 28725 105293 28733 108277
rect 31717 105293 31725 108277
rect 28725 105285 31725 105293
rect 31915 108277 34915 108285
rect 31915 105293 31923 108277
rect 34907 105293 34915 108277
rect 31915 105285 34915 105293
rect 35105 108277 38105 108285
rect 35105 105293 35113 108277
rect 38097 105293 38105 108277
rect 35105 105285 38105 105293
rect 38295 108277 41295 108285
rect 38295 105293 38303 108277
rect 41287 105293 41295 108277
rect 38295 105285 41295 105293
rect 41485 108277 44485 108285
rect 41485 105293 41493 108277
rect 44477 105293 44485 108277
rect 41485 105285 44485 105293
rect 44675 108277 47675 108285
rect 44675 105293 44683 108277
rect 47667 105293 47675 108277
rect 44675 105285 47675 105293
rect 47865 108277 50865 108285
rect 47865 105293 47873 108277
rect 50857 105293 50865 108277
rect 47865 105285 50865 105293
rect 51055 108277 54055 108285
rect 51055 105293 51063 108277
rect 54047 105293 54055 108277
rect 51055 105285 54055 105293
rect 54245 108277 57245 108285
rect 54245 105293 54253 108277
rect 57237 105293 57245 108277
rect 54245 105285 57245 105293
rect 57435 108277 60435 108285
rect 57435 105293 57443 108277
rect 60427 105293 60435 108277
rect 57435 105285 60435 105293
rect 60625 108277 63625 108285
rect 60625 105293 60633 108277
rect 63617 105293 63625 108277
rect 60625 105285 63625 105293
rect 63815 108277 66815 108285
rect 63815 105293 63823 108277
rect 66807 105293 66815 108277
rect 63815 105285 66815 105293
rect 67005 108277 70005 108285
rect 67005 105293 67013 108277
rect 69997 105293 70005 108277
rect 67005 105285 70005 105293
rect 70195 108277 73195 108285
rect 70195 105293 70203 108277
rect 73187 105293 73195 108277
rect 70195 105285 73195 105293
rect 73385 108277 76385 108285
rect 73385 105293 73393 108277
rect 76377 105293 76385 108277
rect 73385 105285 76385 105293
rect 76575 108277 79575 108285
rect 76575 105293 76583 108277
rect 79567 105293 79575 108277
rect 76575 105285 79575 105293
rect 79765 108277 82765 108285
rect 79765 105293 79773 108277
rect 82757 105293 82765 108277
rect 79765 105285 82765 105293
rect 82955 108277 85955 108285
rect 82955 105293 82963 108277
rect 85947 105293 85955 108277
rect 82955 105285 85955 105293
rect 86145 108277 89145 108285
rect 86145 105293 86153 108277
rect 89137 105293 89145 108277
rect 86145 105285 89145 105293
rect 89335 108277 92335 108285
rect 89335 105293 89343 108277
rect 92327 105293 92335 108277
rect 89335 105285 92335 105293
rect 92525 108277 95525 108285
rect 92525 105293 92533 108277
rect 95517 105293 95525 108277
rect 92525 105285 95525 105293
rect 95715 108277 98715 108285
rect 95715 105293 95723 108277
rect 98707 105293 98715 108277
rect 95715 105285 98715 105293
rect 98905 108277 101905 108285
rect 98905 105293 98913 108277
rect 101897 105293 101905 108277
rect 98905 105285 101905 105293
rect 102095 108277 105095 108285
rect 102095 105293 102103 108277
rect 105087 105293 105095 108277
rect 102095 105285 105095 105293
rect 105285 108277 108285 108285
rect 105285 105293 105293 108277
rect 108277 105293 108285 108277
rect 105285 105285 108285 105293
rect 108475 108277 111475 108285
rect 108475 105293 108483 108277
rect 111467 105293 111475 108277
rect 108475 105285 111475 105293
rect 111665 108277 114665 108285
rect 111665 105293 111673 108277
rect 114657 105293 114665 108277
rect 111665 105285 114665 105293
rect 114855 108277 117855 108285
rect 114855 105293 114863 108277
rect 117847 105293 117855 108277
rect 114855 105285 117855 105293
rect 118045 108277 121045 108285
rect 118045 105293 118053 108277
rect 121037 105293 121045 108277
rect 118045 105285 121045 105293
rect 121235 108277 124235 108285
rect 121235 105293 121243 108277
rect 124227 105293 124235 108277
rect 121235 105285 124235 105293
rect 124425 108277 127425 108285
rect 124425 105293 124433 108277
rect 127417 105293 127425 108277
rect 124425 105285 127425 105293
rect 127615 108277 130615 108285
rect 127615 105293 127623 108277
rect 130607 105293 130615 108277
rect 127615 105285 130615 105293
rect 130805 108277 133805 108285
rect 130805 105293 130813 108277
rect 133797 105293 133805 108277
rect 130805 105285 133805 105293
rect 133995 108277 136995 108285
rect 133995 105293 134003 108277
rect 136987 105293 136995 108277
rect 133995 105285 136995 105293
rect 15 105087 3015 105095
rect 15 102103 23 105087
rect 3007 102103 3015 105087
rect 15 102095 3015 102103
rect 3205 105087 6205 105095
rect 3205 102103 3213 105087
rect 6197 102103 6205 105087
rect 3205 102095 6205 102103
rect 6395 105087 9395 105095
rect 6395 102103 6403 105087
rect 9387 102103 9395 105087
rect 6395 102095 9395 102103
rect 9585 105087 12585 105095
rect 9585 102103 9593 105087
rect 12577 102103 12585 105087
rect 9585 102095 12585 102103
rect 12775 105087 15775 105095
rect 12775 102103 12783 105087
rect 15767 102103 15775 105087
rect 12775 102095 15775 102103
rect 15965 105087 18965 105095
rect 15965 102103 15973 105087
rect 18957 102103 18965 105087
rect 15965 102095 18965 102103
rect 19155 105087 22155 105095
rect 19155 102103 19163 105087
rect 22147 102103 22155 105087
rect 19155 102095 22155 102103
rect 22345 105087 25345 105095
rect 22345 102103 22353 105087
rect 25337 102103 25345 105087
rect 22345 102095 25345 102103
rect 25535 105087 28535 105095
rect 25535 102103 25543 105087
rect 28527 102103 28535 105087
rect 25535 102095 28535 102103
rect 28725 105087 31725 105095
rect 28725 102103 28733 105087
rect 31717 102103 31725 105087
rect 28725 102095 31725 102103
rect 31915 105087 34915 105095
rect 31915 102103 31923 105087
rect 34907 102103 34915 105087
rect 31915 102095 34915 102103
rect 35105 105087 38105 105095
rect 35105 102103 35113 105087
rect 38097 102103 38105 105087
rect 35105 102095 38105 102103
rect 38295 105087 41295 105095
rect 38295 102103 38303 105087
rect 41287 102103 41295 105087
rect 38295 102095 41295 102103
rect 41485 105087 44485 105095
rect 41485 102103 41493 105087
rect 44477 102103 44485 105087
rect 41485 102095 44485 102103
rect 44675 105087 47675 105095
rect 44675 102103 44683 105087
rect 47667 102103 47675 105087
rect 44675 102095 47675 102103
rect 47865 105087 50865 105095
rect 47865 102103 47873 105087
rect 50857 102103 50865 105087
rect 47865 102095 50865 102103
rect 51055 105087 54055 105095
rect 51055 102103 51063 105087
rect 54047 102103 54055 105087
rect 51055 102095 54055 102103
rect 54245 105087 57245 105095
rect 54245 102103 54253 105087
rect 57237 102103 57245 105087
rect 54245 102095 57245 102103
rect 57435 105087 60435 105095
rect 57435 102103 57443 105087
rect 60427 102103 60435 105087
rect 57435 102095 60435 102103
rect 60625 105087 63625 105095
rect 60625 102103 60633 105087
rect 63617 102103 63625 105087
rect 60625 102095 63625 102103
rect 63815 105087 66815 105095
rect 63815 102103 63823 105087
rect 66807 102103 66815 105087
rect 63815 102095 66815 102103
rect 67005 105087 70005 105095
rect 67005 102103 67013 105087
rect 69997 102103 70005 105087
rect 67005 102095 70005 102103
rect 70195 105087 73195 105095
rect 70195 102103 70203 105087
rect 73187 102103 73195 105087
rect 70195 102095 73195 102103
rect 73385 105087 76385 105095
rect 73385 102103 73393 105087
rect 76377 102103 76385 105087
rect 73385 102095 76385 102103
rect 76575 105087 79575 105095
rect 76575 102103 76583 105087
rect 79567 102103 79575 105087
rect 76575 102095 79575 102103
rect 79765 105087 82765 105095
rect 79765 102103 79773 105087
rect 82757 102103 82765 105087
rect 79765 102095 82765 102103
rect 82955 105087 85955 105095
rect 82955 102103 82963 105087
rect 85947 102103 85955 105087
rect 82955 102095 85955 102103
rect 86145 105087 89145 105095
rect 86145 102103 86153 105087
rect 89137 102103 89145 105087
rect 86145 102095 89145 102103
rect 89335 105087 92335 105095
rect 89335 102103 89343 105087
rect 92327 102103 92335 105087
rect 89335 102095 92335 102103
rect 92525 105087 95525 105095
rect 92525 102103 92533 105087
rect 95517 102103 95525 105087
rect 92525 102095 95525 102103
rect 95715 105087 98715 105095
rect 95715 102103 95723 105087
rect 98707 102103 98715 105087
rect 95715 102095 98715 102103
rect 98905 105087 101905 105095
rect 98905 102103 98913 105087
rect 101897 102103 101905 105087
rect 98905 102095 101905 102103
rect 102095 105087 105095 105095
rect 102095 102103 102103 105087
rect 105087 102103 105095 105087
rect 102095 102095 105095 102103
rect 105285 105087 108285 105095
rect 105285 102103 105293 105087
rect 108277 102103 108285 105087
rect 105285 102095 108285 102103
rect 108475 105087 111475 105095
rect 108475 102103 108483 105087
rect 111467 102103 111475 105087
rect 108475 102095 111475 102103
rect 111665 105087 114665 105095
rect 111665 102103 111673 105087
rect 114657 102103 114665 105087
rect 111665 102095 114665 102103
rect 114855 105087 117855 105095
rect 114855 102103 114863 105087
rect 117847 102103 117855 105087
rect 114855 102095 117855 102103
rect 118045 105087 121045 105095
rect 118045 102103 118053 105087
rect 121037 102103 121045 105087
rect 118045 102095 121045 102103
rect 121235 105087 124235 105095
rect 121235 102103 121243 105087
rect 124227 102103 124235 105087
rect 121235 102095 124235 102103
rect 124425 105087 127425 105095
rect 124425 102103 124433 105087
rect 127417 102103 127425 105087
rect 124425 102095 127425 102103
rect 127615 105087 130615 105095
rect 127615 102103 127623 105087
rect 130607 102103 130615 105087
rect 127615 102095 130615 102103
rect 130805 105087 133805 105095
rect 130805 102103 130813 105087
rect 133797 102103 133805 105087
rect 130805 102095 133805 102103
rect 133995 105087 136995 105095
rect 133995 102103 134003 105087
rect 136987 102103 136995 105087
rect 133995 102095 136995 102103
rect 15 101897 3015 101905
rect 15 98913 23 101897
rect 3007 98913 3015 101897
rect 15 98905 3015 98913
rect 3205 101897 6205 101905
rect 3205 98913 3213 101897
rect 6197 98913 6205 101897
rect 3205 98905 6205 98913
rect 6395 101897 9395 101905
rect 6395 98913 6403 101897
rect 9387 98913 9395 101897
rect 6395 98905 9395 98913
rect 9585 101897 12585 101905
rect 9585 98913 9593 101897
rect 12577 98913 12585 101897
rect 9585 98905 12585 98913
rect 12775 101897 15775 101905
rect 12775 98913 12783 101897
rect 15767 98913 15775 101897
rect 12775 98905 15775 98913
rect 15965 101897 18965 101905
rect 15965 98913 15973 101897
rect 18957 98913 18965 101897
rect 15965 98905 18965 98913
rect 19155 101897 22155 101905
rect 19155 98913 19163 101897
rect 22147 98913 22155 101897
rect 19155 98905 22155 98913
rect 22345 101897 25345 101905
rect 22345 98913 22353 101897
rect 25337 98913 25345 101897
rect 22345 98905 25345 98913
rect 25535 101897 28535 101905
rect 25535 98913 25543 101897
rect 28527 98913 28535 101897
rect 25535 98905 28535 98913
rect 28725 101897 31725 101905
rect 28725 98913 28733 101897
rect 31717 98913 31725 101897
rect 28725 98905 31725 98913
rect 31915 101897 34915 101905
rect 31915 98913 31923 101897
rect 34907 98913 34915 101897
rect 31915 98905 34915 98913
rect 35105 101897 38105 101905
rect 35105 98913 35113 101897
rect 38097 98913 38105 101897
rect 35105 98905 38105 98913
rect 38295 101897 41295 101905
rect 38295 98913 38303 101897
rect 41287 98913 41295 101897
rect 38295 98905 41295 98913
rect 41485 101897 44485 101905
rect 41485 98913 41493 101897
rect 44477 98913 44485 101897
rect 41485 98905 44485 98913
rect 44675 101897 47675 101905
rect 44675 98913 44683 101897
rect 47667 98913 47675 101897
rect 44675 98905 47675 98913
rect 47865 101897 50865 101905
rect 47865 98913 47873 101897
rect 50857 98913 50865 101897
rect 47865 98905 50865 98913
rect 51055 101897 54055 101905
rect 51055 98913 51063 101897
rect 54047 98913 54055 101897
rect 51055 98905 54055 98913
rect 54245 101897 57245 101905
rect 54245 98913 54253 101897
rect 57237 98913 57245 101897
rect 54245 98905 57245 98913
rect 57435 101897 60435 101905
rect 57435 98913 57443 101897
rect 60427 98913 60435 101897
rect 57435 98905 60435 98913
rect 60625 101897 63625 101905
rect 60625 98913 60633 101897
rect 63617 98913 63625 101897
rect 60625 98905 63625 98913
rect 63815 101897 66815 101905
rect 63815 98913 63823 101897
rect 66807 98913 66815 101897
rect 63815 98905 66815 98913
rect 67005 101897 70005 101905
rect 67005 98913 67013 101897
rect 69997 98913 70005 101897
rect 67005 98905 70005 98913
rect 70195 101897 73195 101905
rect 70195 98913 70203 101897
rect 73187 98913 73195 101897
rect 70195 98905 73195 98913
rect 73385 101897 76385 101905
rect 73385 98913 73393 101897
rect 76377 98913 76385 101897
rect 73385 98905 76385 98913
rect 76575 101897 79575 101905
rect 76575 98913 76583 101897
rect 79567 98913 79575 101897
rect 76575 98905 79575 98913
rect 79765 101897 82765 101905
rect 79765 98913 79773 101897
rect 82757 98913 82765 101897
rect 79765 98905 82765 98913
rect 82955 101897 85955 101905
rect 82955 98913 82963 101897
rect 85947 98913 85955 101897
rect 82955 98905 85955 98913
rect 86145 101897 89145 101905
rect 86145 98913 86153 101897
rect 89137 98913 89145 101897
rect 86145 98905 89145 98913
rect 89335 101897 92335 101905
rect 89335 98913 89343 101897
rect 92327 98913 92335 101897
rect 89335 98905 92335 98913
rect 92525 101897 95525 101905
rect 92525 98913 92533 101897
rect 95517 98913 95525 101897
rect 92525 98905 95525 98913
rect 95715 101897 98715 101905
rect 95715 98913 95723 101897
rect 98707 98913 98715 101897
rect 95715 98905 98715 98913
rect 98905 101897 101905 101905
rect 98905 98913 98913 101897
rect 101897 98913 101905 101897
rect 98905 98905 101905 98913
rect 102095 101897 105095 101905
rect 102095 98913 102103 101897
rect 105087 98913 105095 101897
rect 102095 98905 105095 98913
rect 105285 101897 108285 101905
rect 105285 98913 105293 101897
rect 108277 98913 108285 101897
rect 105285 98905 108285 98913
rect 108475 101897 111475 101905
rect 108475 98913 108483 101897
rect 111467 98913 111475 101897
rect 108475 98905 111475 98913
rect 111665 101897 114665 101905
rect 111665 98913 111673 101897
rect 114657 98913 114665 101897
rect 111665 98905 114665 98913
rect 114855 101897 117855 101905
rect 114855 98913 114863 101897
rect 117847 98913 117855 101897
rect 114855 98905 117855 98913
rect 118045 101897 121045 101905
rect 118045 98913 118053 101897
rect 121037 98913 121045 101897
rect 118045 98905 121045 98913
rect 121235 101897 124235 101905
rect 121235 98913 121243 101897
rect 124227 98913 124235 101897
rect 121235 98905 124235 98913
rect 124425 101897 127425 101905
rect 124425 98913 124433 101897
rect 127417 98913 127425 101897
rect 124425 98905 127425 98913
rect 127615 101897 130615 101905
rect 127615 98913 127623 101897
rect 130607 98913 130615 101897
rect 127615 98905 130615 98913
rect 130805 101897 133805 101905
rect 130805 98913 130813 101897
rect 133797 98913 133805 101897
rect 130805 98905 133805 98913
rect 133995 101897 136995 101905
rect 133995 98913 134003 101897
rect 136987 98913 136995 101897
rect 133995 98905 136995 98913
rect 9585 98707 12585 98715
rect 9585 95723 9593 98707
rect 12577 95723 12585 98707
rect 9585 95715 12585 95723
rect 12775 98707 15775 98715
rect 12775 95723 12783 98707
rect 15767 95723 15775 98707
rect 12775 95715 15775 95723
rect 15965 98707 18965 98715
rect 15965 95723 15973 98707
rect 18957 95723 18965 98707
rect 15965 95715 18965 95723
rect 19155 98707 22155 98715
rect 19155 95723 19163 98707
rect 22147 95723 22155 98707
rect 19155 95715 22155 95723
rect 22345 98707 25345 98715
rect 22345 95723 22353 98707
rect 25337 95723 25345 98707
rect 22345 95715 25345 95723
rect 25535 98707 28535 98715
rect 25535 95723 25543 98707
rect 28527 95723 28535 98707
rect 25535 95715 28535 95723
rect 28725 98707 31725 98715
rect 28725 95723 28733 98707
rect 31717 95723 31725 98707
rect 28725 95715 31725 95723
rect 31915 98707 34915 98715
rect 31915 95723 31923 98707
rect 34907 95723 34915 98707
rect 31915 95715 34915 95723
rect 35105 98707 38105 98715
rect 35105 95723 35113 98707
rect 38097 95723 38105 98707
rect 35105 95715 38105 95723
rect 38295 98707 41295 98715
rect 38295 95723 38303 98707
rect 41287 95723 41295 98707
rect 38295 95715 41295 95723
rect 41485 98707 44485 98715
rect 41485 95723 41493 98707
rect 44477 95723 44485 98707
rect 41485 95715 44485 95723
rect 44675 98707 47675 98715
rect 44675 95723 44683 98707
rect 47667 95723 47675 98707
rect 44675 95715 47675 95723
rect 47865 98707 50865 98715
rect 47865 95723 47873 98707
rect 50857 95723 50865 98707
rect 47865 95715 50865 95723
rect 51055 98707 54055 98715
rect 51055 95723 51063 98707
rect 54047 95723 54055 98707
rect 51055 95715 54055 95723
rect 54245 98707 57245 98715
rect 54245 95723 54253 98707
rect 57237 95723 57245 98707
rect 54245 95715 57245 95723
rect 57435 98707 60435 98715
rect 57435 95723 57443 98707
rect 60427 95723 60435 98707
rect 57435 95715 60435 95723
rect 60625 98707 63625 98715
rect 60625 95723 60633 98707
rect 63617 95723 63625 98707
rect 60625 95715 63625 95723
rect 63815 98707 66815 98715
rect 63815 95723 63823 98707
rect 66807 95723 66815 98707
rect 63815 95715 66815 95723
rect 67005 98707 70005 98715
rect 67005 95723 67013 98707
rect 69997 95723 70005 98707
rect 67005 95715 70005 95723
rect 70195 98707 73195 98715
rect 70195 95723 70203 98707
rect 73187 95723 73195 98707
rect 70195 95715 73195 95723
rect 73385 98707 76385 98715
rect 73385 95723 73393 98707
rect 76377 95723 76385 98707
rect 73385 95715 76385 95723
rect 76575 98707 79575 98715
rect 76575 95723 76583 98707
rect 79567 95723 79575 98707
rect 76575 95715 79575 95723
rect 79765 98707 82765 98715
rect 79765 95723 79773 98707
rect 82757 95723 82765 98707
rect 79765 95715 82765 95723
rect 82955 98707 85955 98715
rect 82955 95723 82963 98707
rect 85947 95723 85955 98707
rect 82955 95715 85955 95723
rect 86145 98707 89145 98715
rect 86145 95723 86153 98707
rect 89137 95723 89145 98707
rect 86145 95715 89145 95723
rect 89335 98707 92335 98715
rect 89335 95723 89343 98707
rect 92327 95723 92335 98707
rect 89335 95715 92335 95723
rect 92525 98707 95525 98715
rect 92525 95723 92533 98707
rect 95517 95723 95525 98707
rect 92525 95715 95525 95723
rect 95715 98707 98715 98715
rect 95715 95723 95723 98707
rect 98707 95723 98715 98707
rect 95715 95715 98715 95723
rect 98905 98707 101905 98715
rect 98905 95723 98913 98707
rect 101897 95723 101905 98707
rect 98905 95715 101905 95723
rect 102095 98707 105095 98715
rect 102095 95723 102103 98707
rect 105087 95723 105095 98707
rect 102095 95715 105095 95723
rect 105285 98707 108285 98715
rect 105285 95723 105293 98707
rect 108277 95723 108285 98707
rect 105285 95715 108285 95723
rect 108475 98707 111475 98715
rect 108475 95723 108483 98707
rect 111467 95723 111475 98707
rect 108475 95715 111475 95723
rect 111665 98707 114665 98715
rect 111665 95723 111673 98707
rect 114657 95723 114665 98707
rect 111665 95715 114665 95723
rect 114855 98707 117855 98715
rect 114855 95723 114863 98707
rect 117847 95723 117855 98707
rect 114855 95715 117855 95723
rect 118045 98707 121045 98715
rect 118045 95723 118053 98707
rect 121037 95723 121045 98707
rect 118045 95715 121045 95723
rect 121235 98707 124235 98715
rect 121235 95723 121243 98707
rect 124227 95723 124235 98707
rect 121235 95715 124235 95723
rect 124425 98707 127425 98715
rect 124425 95723 124433 98707
rect 127417 95723 127425 98707
rect 124425 95715 127425 95723
rect 127615 98707 130615 98715
rect 127615 95723 127623 98707
rect 130607 95723 130615 98707
rect 127615 95715 130615 95723
rect 130805 98707 133805 98715
rect 130805 95723 130813 98707
rect 133797 95723 133805 98707
rect 130805 95715 133805 95723
rect 133995 98707 136995 98715
rect 133995 95723 134003 98707
rect 136987 95723 136995 98707
rect 133995 95715 136995 95723
rect 9585 95517 12585 95525
rect 9585 92533 9593 95517
rect 12577 92533 12585 95517
rect 9585 92525 12585 92533
rect 12775 95517 15775 95525
rect 12775 92533 12783 95517
rect 15767 92533 15775 95517
rect 12775 92525 15775 92533
rect 15965 95517 18965 95525
rect 15965 92533 15973 95517
rect 18957 92533 18965 95517
rect 15965 92525 18965 92533
rect 19155 95517 22155 95525
rect 19155 92533 19163 95517
rect 22147 92533 22155 95517
rect 19155 92525 22155 92533
rect 22345 95517 25345 95525
rect 22345 92533 22353 95517
rect 25337 92533 25345 95517
rect 22345 92525 25345 92533
rect 25535 95517 28535 95525
rect 25535 92533 25543 95517
rect 28527 92533 28535 95517
rect 25535 92525 28535 92533
rect 28725 95517 31725 95525
rect 28725 92533 28733 95517
rect 31717 92533 31725 95517
rect 28725 92525 31725 92533
rect 31915 95517 34915 95525
rect 31915 92533 31923 95517
rect 34907 92533 34915 95517
rect 31915 92525 34915 92533
rect 35105 95517 38105 95525
rect 35105 92533 35113 95517
rect 38097 92533 38105 95517
rect 35105 92525 38105 92533
rect 38295 95517 41295 95525
rect 38295 92533 38303 95517
rect 41287 92533 41295 95517
rect 38295 92525 41295 92533
rect 41485 95517 44485 95525
rect 41485 92533 41493 95517
rect 44477 92533 44485 95517
rect 41485 92525 44485 92533
rect 44675 95517 47675 95525
rect 44675 92533 44683 95517
rect 47667 92533 47675 95517
rect 44675 92525 47675 92533
rect 47865 95517 50865 95525
rect 47865 92533 47873 95517
rect 50857 92533 50865 95517
rect 47865 92525 50865 92533
rect 51055 95517 54055 95525
rect 51055 92533 51063 95517
rect 54047 92533 54055 95517
rect 51055 92525 54055 92533
rect 54245 95517 57245 95525
rect 54245 92533 54253 95517
rect 57237 92533 57245 95517
rect 54245 92525 57245 92533
rect 57435 95517 60435 95525
rect 57435 92533 57443 95517
rect 60427 92533 60435 95517
rect 57435 92525 60435 92533
rect 60625 95517 63625 95525
rect 60625 92533 60633 95517
rect 63617 92533 63625 95517
rect 60625 92525 63625 92533
rect 63815 95517 66815 95525
rect 63815 92533 63823 95517
rect 66807 92533 66815 95517
rect 63815 92525 66815 92533
rect 67005 95517 70005 95525
rect 67005 92533 67013 95517
rect 69997 92533 70005 95517
rect 67005 92525 70005 92533
rect 70195 95517 73195 95525
rect 70195 92533 70203 95517
rect 73187 92533 73195 95517
rect 70195 92525 73195 92533
rect 73385 95517 76385 95525
rect 73385 92533 73393 95517
rect 76377 92533 76385 95517
rect 73385 92525 76385 92533
rect 76575 95517 79575 95525
rect 76575 92533 76583 95517
rect 79567 92533 79575 95517
rect 76575 92525 79575 92533
rect 79765 95517 82765 95525
rect 79765 92533 79773 95517
rect 82757 92533 82765 95517
rect 79765 92525 82765 92533
rect 82955 95517 85955 95525
rect 82955 92533 82963 95517
rect 85947 92533 85955 95517
rect 82955 92525 85955 92533
rect 86145 95517 89145 95525
rect 86145 92533 86153 95517
rect 89137 92533 89145 95517
rect 86145 92525 89145 92533
rect 89335 95517 92335 95525
rect 89335 92533 89343 95517
rect 92327 92533 92335 95517
rect 89335 92525 92335 92533
rect 92525 95517 95525 95525
rect 92525 92533 92533 95517
rect 95517 92533 95525 95517
rect 92525 92525 95525 92533
rect 95715 95517 98715 95525
rect 95715 92533 95723 95517
rect 98707 92533 98715 95517
rect 95715 92525 98715 92533
rect 98905 95517 101905 95525
rect 98905 92533 98913 95517
rect 101897 92533 101905 95517
rect 98905 92525 101905 92533
rect 102095 95517 105095 95525
rect 102095 92533 102103 95517
rect 105087 92533 105095 95517
rect 102095 92525 105095 92533
rect 105285 95517 108285 95525
rect 105285 92533 105293 95517
rect 108277 92533 108285 95517
rect 105285 92525 108285 92533
rect 108475 95517 111475 95525
rect 108475 92533 108483 95517
rect 111467 92533 111475 95517
rect 108475 92525 111475 92533
rect 111665 95517 114665 95525
rect 111665 92533 111673 95517
rect 114657 92533 114665 95517
rect 111665 92525 114665 92533
rect 114855 95517 117855 95525
rect 114855 92533 114863 95517
rect 117847 92533 117855 95517
rect 114855 92525 117855 92533
rect 118045 95517 121045 95525
rect 118045 92533 118053 95517
rect 121037 92533 121045 95517
rect 118045 92525 121045 92533
rect 121235 95517 124235 95525
rect 121235 92533 121243 95517
rect 124227 92533 124235 95517
rect 121235 92525 124235 92533
rect 124425 95517 127425 95525
rect 124425 92533 124433 95517
rect 127417 92533 127425 95517
rect 124425 92525 127425 92533
rect 127615 95517 130615 95525
rect 127615 92533 127623 95517
rect 130607 92533 130615 95517
rect 127615 92525 130615 92533
rect 130805 95517 133805 95525
rect 130805 92533 130813 95517
rect 133797 92533 133805 95517
rect 130805 92525 133805 92533
rect 133995 95517 136995 95525
rect 133995 92533 134003 95517
rect 136987 92533 136995 95517
rect 133995 92525 136995 92533
rect 9585 92327 12585 92335
rect 9585 89343 9593 92327
rect 12577 89343 12585 92327
rect 9585 89335 12585 89343
rect 12775 92327 15775 92335
rect 12775 89343 12783 92327
rect 15767 89343 15775 92327
rect 12775 89335 15775 89343
rect 15965 92327 18965 92335
rect 15965 89343 15973 92327
rect 18957 89343 18965 92327
rect 15965 89335 18965 89343
rect 19155 92327 22155 92335
rect 19155 89343 19163 92327
rect 22147 89343 22155 92327
rect 19155 89335 22155 89343
rect 22345 92327 25345 92335
rect 22345 89343 22353 92327
rect 25337 89343 25345 92327
rect 22345 89335 25345 89343
rect 25535 92327 28535 92335
rect 25535 89343 25543 92327
rect 28527 89343 28535 92327
rect 25535 89335 28535 89343
rect 28725 92327 31725 92335
rect 28725 89343 28733 92327
rect 31717 89343 31725 92327
rect 28725 89335 31725 89343
rect 31915 92327 34915 92335
rect 31915 89343 31923 92327
rect 34907 89343 34915 92327
rect 31915 89335 34915 89343
rect 35105 92327 38105 92335
rect 35105 89343 35113 92327
rect 38097 89343 38105 92327
rect 35105 89335 38105 89343
rect 38295 92327 41295 92335
rect 38295 89343 38303 92327
rect 41287 89343 41295 92327
rect 38295 89335 41295 89343
rect 41485 92327 44485 92335
rect 41485 89343 41493 92327
rect 44477 89343 44485 92327
rect 41485 89335 44485 89343
rect 44675 92327 47675 92335
rect 44675 89343 44683 92327
rect 47667 89343 47675 92327
rect 44675 89335 47675 89343
rect 47865 92327 50865 92335
rect 47865 89343 47873 92327
rect 50857 89343 50865 92327
rect 47865 89335 50865 89343
rect 51055 92327 54055 92335
rect 51055 89343 51063 92327
rect 54047 89343 54055 92327
rect 51055 89335 54055 89343
rect 54245 92327 57245 92335
rect 54245 89343 54253 92327
rect 57237 89343 57245 92327
rect 54245 89335 57245 89343
rect 57435 92327 60435 92335
rect 57435 89343 57443 92327
rect 60427 89343 60435 92327
rect 57435 89335 60435 89343
rect 60625 92327 63625 92335
rect 60625 89343 60633 92327
rect 63617 89343 63625 92327
rect 60625 89335 63625 89343
rect 63815 92327 66815 92335
rect 63815 89343 63823 92327
rect 66807 89343 66815 92327
rect 63815 89335 66815 89343
rect 67005 92327 70005 92335
rect 67005 89343 67013 92327
rect 69997 89343 70005 92327
rect 67005 89335 70005 89343
rect 70195 92327 73195 92335
rect 70195 89343 70203 92327
rect 73187 89343 73195 92327
rect 70195 89335 73195 89343
rect 73385 92327 76385 92335
rect 73385 89343 73393 92327
rect 76377 89343 76385 92327
rect 73385 89335 76385 89343
rect 76575 92327 79575 92335
rect 76575 89343 76583 92327
rect 79567 89343 79575 92327
rect 76575 89335 79575 89343
rect 79765 92327 82765 92335
rect 79765 89343 79773 92327
rect 82757 89343 82765 92327
rect 79765 89335 82765 89343
rect 82955 92327 85955 92335
rect 82955 89343 82963 92327
rect 85947 89343 85955 92327
rect 82955 89335 85955 89343
rect 86145 92327 89145 92335
rect 86145 89343 86153 92327
rect 89137 89343 89145 92327
rect 86145 89335 89145 89343
rect 89335 92327 92335 92335
rect 89335 89343 89343 92327
rect 92327 89343 92335 92327
rect 89335 89335 92335 89343
rect 92525 92327 95525 92335
rect 92525 89343 92533 92327
rect 95517 89343 95525 92327
rect 92525 89335 95525 89343
rect 95715 92327 98715 92335
rect 95715 89343 95723 92327
rect 98707 89343 98715 92327
rect 95715 89335 98715 89343
rect 98905 92327 101905 92335
rect 98905 89343 98913 92327
rect 101897 89343 101905 92327
rect 98905 89335 101905 89343
rect 102095 92327 105095 92335
rect 102095 89343 102103 92327
rect 105087 89343 105095 92327
rect 102095 89335 105095 89343
rect 105285 92327 108285 92335
rect 105285 89343 105293 92327
rect 108277 89343 108285 92327
rect 105285 89335 108285 89343
rect 108475 92327 111475 92335
rect 108475 89343 108483 92327
rect 111467 89343 111475 92327
rect 108475 89335 111475 89343
rect 111665 92327 114665 92335
rect 111665 89343 111673 92327
rect 114657 89343 114665 92327
rect 111665 89335 114665 89343
rect 114855 92327 117855 92335
rect 114855 89343 114863 92327
rect 117847 89343 117855 92327
rect 114855 89335 117855 89343
rect 118045 92327 121045 92335
rect 118045 89343 118053 92327
rect 121037 89343 121045 92327
rect 118045 89335 121045 89343
rect 121235 92327 124235 92335
rect 121235 89343 121243 92327
rect 124227 89343 124235 92327
rect 121235 89335 124235 89343
rect 124425 92327 127425 92335
rect 124425 89343 124433 92327
rect 127417 89343 127425 92327
rect 124425 89335 127425 89343
rect 127615 92327 130615 92335
rect 127615 89343 127623 92327
rect 130607 89343 130615 92327
rect 127615 89335 130615 89343
rect 130805 92327 133805 92335
rect 130805 89343 130813 92327
rect 133797 89343 133805 92327
rect 130805 89335 133805 89343
rect 133995 92327 136995 92335
rect 133995 89343 134003 92327
rect 136987 89343 136995 92327
rect 133995 89335 136995 89343
rect 9585 89137 12585 89145
rect 9585 86153 9593 89137
rect 12577 86153 12585 89137
rect 9585 86145 12585 86153
rect 12775 89137 15775 89145
rect 12775 86153 12783 89137
rect 15767 86153 15775 89137
rect 12775 86145 15775 86153
rect 15965 89137 18965 89145
rect 15965 86153 15973 89137
rect 18957 86153 18965 89137
rect 15965 86145 18965 86153
rect 19155 89137 22155 89145
rect 19155 86153 19163 89137
rect 22147 86153 22155 89137
rect 19155 86145 22155 86153
rect 22345 89137 25345 89145
rect 22345 86153 22353 89137
rect 25337 86153 25345 89137
rect 22345 86145 25345 86153
rect 25535 89137 28535 89145
rect 25535 86153 25543 89137
rect 28527 86153 28535 89137
rect 25535 86145 28535 86153
rect 28725 89137 31725 89145
rect 28725 86153 28733 89137
rect 31717 86153 31725 89137
rect 28725 86145 31725 86153
rect 31915 89137 34915 89145
rect 31915 86153 31923 89137
rect 34907 86153 34915 89137
rect 31915 86145 34915 86153
rect 35105 89137 38105 89145
rect 35105 86153 35113 89137
rect 38097 86153 38105 89137
rect 35105 86145 38105 86153
rect 38295 89137 41295 89145
rect 38295 86153 38303 89137
rect 41287 86153 41295 89137
rect 38295 86145 41295 86153
rect 41485 89137 44485 89145
rect 41485 86153 41493 89137
rect 44477 86153 44485 89137
rect 41485 86145 44485 86153
rect 44675 89137 47675 89145
rect 44675 86153 44683 89137
rect 47667 86153 47675 89137
rect 44675 86145 47675 86153
rect 47865 89137 50865 89145
rect 47865 86153 47873 89137
rect 50857 86153 50865 89137
rect 47865 86145 50865 86153
rect 51055 89137 54055 89145
rect 51055 86153 51063 89137
rect 54047 86153 54055 89137
rect 51055 86145 54055 86153
rect 54245 89137 57245 89145
rect 54245 86153 54253 89137
rect 57237 86153 57245 89137
rect 54245 86145 57245 86153
rect 57435 89137 60435 89145
rect 57435 86153 57443 89137
rect 60427 86153 60435 89137
rect 57435 86145 60435 86153
rect 60625 89137 63625 89145
rect 60625 86153 60633 89137
rect 63617 86153 63625 89137
rect 60625 86145 63625 86153
rect 63815 89137 66815 89145
rect 63815 86153 63823 89137
rect 66807 86153 66815 89137
rect 63815 86145 66815 86153
rect 67005 89137 70005 89145
rect 67005 86153 67013 89137
rect 69997 86153 70005 89137
rect 67005 86145 70005 86153
rect 70195 89137 73195 89145
rect 70195 86153 70203 89137
rect 73187 86153 73195 89137
rect 70195 86145 73195 86153
rect 73385 89137 76385 89145
rect 73385 86153 73393 89137
rect 76377 86153 76385 89137
rect 73385 86145 76385 86153
rect 76575 89137 79575 89145
rect 76575 86153 76583 89137
rect 79567 86153 79575 89137
rect 76575 86145 79575 86153
rect 79765 89137 82765 89145
rect 79765 86153 79773 89137
rect 82757 86153 82765 89137
rect 79765 86145 82765 86153
rect 82955 89137 85955 89145
rect 82955 86153 82963 89137
rect 85947 86153 85955 89137
rect 82955 86145 85955 86153
rect 86145 89137 89145 89145
rect 86145 86153 86153 89137
rect 89137 86153 89145 89137
rect 86145 86145 89145 86153
rect 89335 89137 92335 89145
rect 89335 86153 89343 89137
rect 92327 86153 92335 89137
rect 89335 86145 92335 86153
rect 92525 89137 95525 89145
rect 92525 86153 92533 89137
rect 95517 86153 95525 89137
rect 92525 86145 95525 86153
rect 95715 89137 98715 89145
rect 95715 86153 95723 89137
rect 98707 86153 98715 89137
rect 95715 86145 98715 86153
rect 98905 89137 101905 89145
rect 98905 86153 98913 89137
rect 101897 86153 101905 89137
rect 98905 86145 101905 86153
rect 102095 89137 105095 89145
rect 102095 86153 102103 89137
rect 105087 86153 105095 89137
rect 102095 86145 105095 86153
rect 105285 89137 108285 89145
rect 105285 86153 105293 89137
rect 108277 86153 108285 89137
rect 105285 86145 108285 86153
rect 108475 89137 111475 89145
rect 108475 86153 108483 89137
rect 111467 86153 111475 89137
rect 108475 86145 111475 86153
rect 111665 89137 114665 89145
rect 111665 86153 111673 89137
rect 114657 86153 114665 89137
rect 111665 86145 114665 86153
rect 114855 89137 117855 89145
rect 114855 86153 114863 89137
rect 117847 86153 117855 89137
rect 114855 86145 117855 86153
rect 118045 89137 121045 89145
rect 118045 86153 118053 89137
rect 121037 86153 121045 89137
rect 118045 86145 121045 86153
rect 121235 89137 124235 89145
rect 121235 86153 121243 89137
rect 124227 86153 124235 89137
rect 121235 86145 124235 86153
rect 124425 89137 127425 89145
rect 124425 86153 124433 89137
rect 127417 86153 127425 89137
rect 124425 86145 127425 86153
rect 127615 89137 130615 89145
rect 127615 86153 127623 89137
rect 130607 86153 130615 89137
rect 127615 86145 130615 86153
rect 130805 89137 133805 89145
rect 130805 86153 130813 89137
rect 133797 86153 133805 89137
rect 130805 86145 133805 86153
rect 133995 89137 136995 89145
rect 133995 86153 134003 89137
rect 136987 86153 136995 89137
rect 133995 86145 136995 86153
rect 9585 85947 12585 85955
rect 9585 82963 9593 85947
rect 12577 82963 12585 85947
rect 9585 82955 12585 82963
rect 12775 85947 15775 85955
rect 12775 82963 12783 85947
rect 15767 82963 15775 85947
rect 12775 82955 15775 82963
rect 15965 85947 18965 85955
rect 15965 82963 15973 85947
rect 18957 82963 18965 85947
rect 15965 82955 18965 82963
rect 19155 85947 22155 85955
rect 19155 82963 19163 85947
rect 22147 82963 22155 85947
rect 19155 82955 22155 82963
rect 22345 85947 25345 85955
rect 22345 82963 22353 85947
rect 25337 82963 25345 85947
rect 22345 82955 25345 82963
rect 25535 85947 28535 85955
rect 25535 82963 25543 85947
rect 28527 82963 28535 85947
rect 25535 82955 28535 82963
rect 28725 85947 31725 85955
rect 28725 82963 28733 85947
rect 31717 82963 31725 85947
rect 28725 82955 31725 82963
rect 31915 85947 34915 85955
rect 31915 82963 31923 85947
rect 34907 82963 34915 85947
rect 31915 82955 34915 82963
rect 35105 85947 38105 85955
rect 35105 82963 35113 85947
rect 38097 82963 38105 85947
rect 35105 82955 38105 82963
rect 38295 85947 41295 85955
rect 38295 82963 38303 85947
rect 41287 82963 41295 85947
rect 38295 82955 41295 82963
rect 41485 85947 44485 85955
rect 41485 82963 41493 85947
rect 44477 82963 44485 85947
rect 41485 82955 44485 82963
rect 44675 85947 47675 85955
rect 44675 82963 44683 85947
rect 47667 82963 47675 85947
rect 44675 82955 47675 82963
rect 47865 85947 50865 85955
rect 47865 82963 47873 85947
rect 50857 82963 50865 85947
rect 47865 82955 50865 82963
rect 51055 85947 54055 85955
rect 51055 82963 51063 85947
rect 54047 82963 54055 85947
rect 51055 82955 54055 82963
rect 54245 85947 57245 85955
rect 54245 82963 54253 85947
rect 57237 82963 57245 85947
rect 54245 82955 57245 82963
rect 57435 85947 60435 85955
rect 57435 82963 57443 85947
rect 60427 82963 60435 85947
rect 57435 82955 60435 82963
rect 60625 85947 63625 85955
rect 60625 82963 60633 85947
rect 63617 82963 63625 85947
rect 60625 82955 63625 82963
rect 63815 85947 66815 85955
rect 63815 82963 63823 85947
rect 66807 82963 66815 85947
rect 63815 82955 66815 82963
rect 67005 85947 70005 85955
rect 67005 82963 67013 85947
rect 69997 82963 70005 85947
rect 67005 82955 70005 82963
rect 70195 85947 73195 85955
rect 70195 82963 70203 85947
rect 73187 82963 73195 85947
rect 70195 82955 73195 82963
rect 73385 85947 76385 85955
rect 73385 82963 73393 85947
rect 76377 82963 76385 85947
rect 73385 82955 76385 82963
rect 76575 85947 79575 85955
rect 76575 82963 76583 85947
rect 79567 82963 79575 85947
rect 76575 82955 79575 82963
rect 79765 85947 82765 85955
rect 79765 82963 79773 85947
rect 82757 82963 82765 85947
rect 79765 82955 82765 82963
rect 82955 85947 85955 85955
rect 82955 82963 82963 85947
rect 85947 82963 85955 85947
rect 82955 82955 85955 82963
rect 86145 85947 89145 85955
rect 86145 82963 86153 85947
rect 89137 82963 89145 85947
rect 86145 82955 89145 82963
rect 89335 85947 92335 85955
rect 89335 82963 89343 85947
rect 92327 82963 92335 85947
rect 89335 82955 92335 82963
rect 92525 85947 95525 85955
rect 92525 82963 92533 85947
rect 95517 82963 95525 85947
rect 92525 82955 95525 82963
rect 95715 85947 98715 85955
rect 95715 82963 95723 85947
rect 98707 82963 98715 85947
rect 95715 82955 98715 82963
rect 98905 85947 101905 85955
rect 98905 82963 98913 85947
rect 101897 82963 101905 85947
rect 98905 82955 101905 82963
rect 102095 85947 105095 85955
rect 102095 82963 102103 85947
rect 105087 82963 105095 85947
rect 102095 82955 105095 82963
rect 105285 85947 108285 85955
rect 105285 82963 105293 85947
rect 108277 82963 108285 85947
rect 105285 82955 108285 82963
rect 108475 85947 111475 85955
rect 108475 82963 108483 85947
rect 111467 82963 111475 85947
rect 108475 82955 111475 82963
rect 111665 85947 114665 85955
rect 111665 82963 111673 85947
rect 114657 82963 114665 85947
rect 111665 82955 114665 82963
rect 114855 85947 117855 85955
rect 114855 82963 114863 85947
rect 117847 82963 117855 85947
rect 114855 82955 117855 82963
rect 118045 85947 121045 85955
rect 118045 82963 118053 85947
rect 121037 82963 121045 85947
rect 118045 82955 121045 82963
rect 121235 85947 124235 85955
rect 121235 82963 121243 85947
rect 124227 82963 124235 85947
rect 121235 82955 124235 82963
rect 124425 85947 127425 85955
rect 124425 82963 124433 85947
rect 127417 82963 127425 85947
rect 124425 82955 127425 82963
rect 127615 85947 130615 85955
rect 127615 82963 127623 85947
rect 130607 82963 130615 85947
rect 127615 82955 130615 82963
rect 130805 85947 133805 85955
rect 130805 82963 130813 85947
rect 133797 82963 133805 85947
rect 130805 82955 133805 82963
rect 133995 85947 136995 85955
rect 133995 82963 134003 85947
rect 136987 82963 136995 85947
rect 133995 82955 136995 82963
rect 9585 82757 12585 82765
rect 9585 79773 9593 82757
rect 12577 79773 12585 82757
rect 9585 79765 12585 79773
rect 12775 82757 15775 82765
rect 12775 79773 12783 82757
rect 15767 79773 15775 82757
rect 12775 79765 15775 79773
rect 15965 82757 18965 82765
rect 15965 79773 15973 82757
rect 18957 79773 18965 82757
rect 15965 79765 18965 79773
rect 19155 82757 22155 82765
rect 19155 79773 19163 82757
rect 22147 79773 22155 82757
rect 19155 79765 22155 79773
rect 22345 82757 25345 82765
rect 22345 79773 22353 82757
rect 25337 79773 25345 82757
rect 22345 79765 25345 79773
rect 25535 82757 28535 82765
rect 25535 79773 25543 82757
rect 28527 79773 28535 82757
rect 25535 79765 28535 79773
rect 28725 82757 31725 82765
rect 28725 79773 28733 82757
rect 31717 79773 31725 82757
rect 28725 79765 31725 79773
rect 31915 82757 34915 82765
rect 31915 79773 31923 82757
rect 34907 79773 34915 82757
rect 31915 79765 34915 79773
rect 35105 82757 38105 82765
rect 35105 79773 35113 82757
rect 38097 79773 38105 82757
rect 35105 79765 38105 79773
rect 38295 82757 41295 82765
rect 38295 79773 38303 82757
rect 41287 79773 41295 82757
rect 38295 79765 41295 79773
rect 41485 82757 44485 82765
rect 41485 79773 41493 82757
rect 44477 79773 44485 82757
rect 41485 79765 44485 79773
rect 44675 82757 47675 82765
rect 44675 79773 44683 82757
rect 47667 79773 47675 82757
rect 44675 79765 47675 79773
rect 47865 82757 50865 82765
rect 47865 79773 47873 82757
rect 50857 79773 50865 82757
rect 47865 79765 50865 79773
rect 51055 82757 54055 82765
rect 51055 79773 51063 82757
rect 54047 79773 54055 82757
rect 51055 79765 54055 79773
rect 54245 82757 57245 82765
rect 54245 79773 54253 82757
rect 57237 79773 57245 82757
rect 54245 79765 57245 79773
rect 57435 82757 60435 82765
rect 57435 79773 57443 82757
rect 60427 79773 60435 82757
rect 57435 79765 60435 79773
rect 60625 82757 63625 82765
rect 60625 79773 60633 82757
rect 63617 79773 63625 82757
rect 60625 79765 63625 79773
rect 63815 82757 66815 82765
rect 63815 79773 63823 82757
rect 66807 79773 66815 82757
rect 63815 79765 66815 79773
rect 67005 82757 70005 82765
rect 67005 79773 67013 82757
rect 69997 79773 70005 82757
rect 67005 79765 70005 79773
rect 70195 82757 73195 82765
rect 70195 79773 70203 82757
rect 73187 79773 73195 82757
rect 70195 79765 73195 79773
rect 73385 82757 76385 82765
rect 73385 79773 73393 82757
rect 76377 79773 76385 82757
rect 73385 79765 76385 79773
rect 76575 82757 79575 82765
rect 76575 79773 76583 82757
rect 79567 79773 79575 82757
rect 76575 79765 79575 79773
rect 79765 82757 82765 82765
rect 79765 79773 79773 82757
rect 82757 79773 82765 82757
rect 79765 79765 82765 79773
rect 82955 82757 85955 82765
rect 82955 79773 82963 82757
rect 85947 79773 85955 82757
rect 82955 79765 85955 79773
rect 86145 82757 89145 82765
rect 86145 79773 86153 82757
rect 89137 79773 89145 82757
rect 86145 79765 89145 79773
rect 89335 82757 92335 82765
rect 89335 79773 89343 82757
rect 92327 79773 92335 82757
rect 89335 79765 92335 79773
rect 92525 82757 95525 82765
rect 92525 79773 92533 82757
rect 95517 79773 95525 82757
rect 92525 79765 95525 79773
rect 95715 82757 98715 82765
rect 95715 79773 95723 82757
rect 98707 79773 98715 82757
rect 95715 79765 98715 79773
rect 98905 82757 101905 82765
rect 98905 79773 98913 82757
rect 101897 79773 101905 82757
rect 98905 79765 101905 79773
rect 102095 82757 105095 82765
rect 102095 79773 102103 82757
rect 105087 79773 105095 82757
rect 102095 79765 105095 79773
rect 105285 82757 108285 82765
rect 105285 79773 105293 82757
rect 108277 79773 108285 82757
rect 105285 79765 108285 79773
rect 108475 82757 111475 82765
rect 108475 79773 108483 82757
rect 111467 79773 111475 82757
rect 108475 79765 111475 79773
rect 111665 82757 114665 82765
rect 111665 79773 111673 82757
rect 114657 79773 114665 82757
rect 111665 79765 114665 79773
rect 114855 82757 117855 82765
rect 114855 79773 114863 82757
rect 117847 79773 117855 82757
rect 114855 79765 117855 79773
rect 118045 82757 121045 82765
rect 118045 79773 118053 82757
rect 121037 79773 121045 82757
rect 118045 79765 121045 79773
rect 121235 82757 124235 82765
rect 121235 79773 121243 82757
rect 124227 79773 124235 82757
rect 121235 79765 124235 79773
rect 124425 82757 127425 82765
rect 124425 79773 124433 82757
rect 127417 79773 127425 82757
rect 124425 79765 127425 79773
rect 127615 82757 130615 82765
rect 127615 79773 127623 82757
rect 130607 79773 130615 82757
rect 127615 79765 130615 79773
rect 130805 82757 133805 82765
rect 130805 79773 130813 82757
rect 133797 79773 133805 82757
rect 130805 79765 133805 79773
rect 133995 82757 136995 82765
rect 133995 79773 134003 82757
rect 136987 79773 136995 82757
rect 133995 79765 136995 79773
rect 15 79567 3015 79575
rect 15 76583 23 79567
rect 3007 76583 3015 79567
rect 15 76575 3015 76583
rect 3205 79567 6205 79575
rect 3205 76583 3213 79567
rect 6197 76583 6205 79567
rect 3205 76575 6205 76583
rect 6395 79567 9395 79575
rect 6395 76583 6403 79567
rect 9387 76583 9395 79567
rect 6395 76575 9395 76583
rect 9585 79567 12585 79575
rect 9585 76583 9593 79567
rect 12577 76583 12585 79567
rect 9585 76575 12585 76583
rect 12775 79567 15775 79575
rect 12775 76583 12783 79567
rect 15767 76583 15775 79567
rect 12775 76575 15775 76583
rect 15965 79567 18965 79575
rect 15965 76583 15973 79567
rect 18957 76583 18965 79567
rect 15965 76575 18965 76583
rect 19155 79567 22155 79575
rect 19155 76583 19163 79567
rect 22147 76583 22155 79567
rect 19155 76575 22155 76583
rect 22345 79567 25345 79575
rect 22345 76583 22353 79567
rect 25337 76583 25345 79567
rect 22345 76575 25345 76583
rect 25535 79567 28535 79575
rect 25535 76583 25543 79567
rect 28527 76583 28535 79567
rect 25535 76575 28535 76583
rect 28725 79567 31725 79575
rect 28725 76583 28733 79567
rect 31717 76583 31725 79567
rect 28725 76575 31725 76583
rect 31915 79567 34915 79575
rect 31915 76583 31923 79567
rect 34907 76583 34915 79567
rect 31915 76575 34915 76583
rect 35105 79567 38105 79575
rect 35105 76583 35113 79567
rect 38097 76583 38105 79567
rect 35105 76575 38105 76583
rect 38295 79567 41295 79575
rect 38295 76583 38303 79567
rect 41287 76583 41295 79567
rect 38295 76575 41295 76583
rect 41485 79567 44485 79575
rect 41485 76583 41493 79567
rect 44477 76583 44485 79567
rect 41485 76575 44485 76583
rect 44675 79567 47675 79575
rect 44675 76583 44683 79567
rect 47667 76583 47675 79567
rect 44675 76575 47675 76583
rect 47865 79567 50865 79575
rect 47865 76583 47873 79567
rect 50857 76583 50865 79567
rect 47865 76575 50865 76583
rect 51055 79567 54055 79575
rect 51055 76583 51063 79567
rect 54047 76583 54055 79567
rect 51055 76575 54055 76583
rect 54245 79567 57245 79575
rect 54245 76583 54253 79567
rect 57237 76583 57245 79567
rect 54245 76575 57245 76583
rect 57435 79567 60435 79575
rect 57435 76583 57443 79567
rect 60427 76583 60435 79567
rect 57435 76575 60435 76583
rect 60625 79567 63625 79575
rect 60625 76583 60633 79567
rect 63617 76583 63625 79567
rect 60625 76575 63625 76583
rect 63815 79567 66815 79575
rect 63815 76583 63823 79567
rect 66807 76583 66815 79567
rect 63815 76575 66815 76583
rect 67005 79567 70005 79575
rect 67005 76583 67013 79567
rect 69997 76583 70005 79567
rect 67005 76575 70005 76583
rect 70195 79567 73195 79575
rect 70195 76583 70203 79567
rect 73187 76583 73195 79567
rect 70195 76575 73195 76583
rect 73385 79567 76385 79575
rect 73385 76583 73393 79567
rect 76377 76583 76385 79567
rect 73385 76575 76385 76583
rect 76575 79567 79575 79575
rect 76575 76583 76583 79567
rect 79567 76583 79575 79567
rect 76575 76575 79575 76583
rect 79765 79567 82765 79575
rect 79765 76583 79773 79567
rect 82757 76583 82765 79567
rect 79765 76575 82765 76583
rect 82955 79567 85955 79575
rect 82955 76583 82963 79567
rect 85947 76583 85955 79567
rect 82955 76575 85955 76583
rect 86145 79567 89145 79575
rect 86145 76583 86153 79567
rect 89137 76583 89145 79567
rect 86145 76575 89145 76583
rect 89335 79567 92335 79575
rect 89335 76583 89343 79567
rect 92327 76583 92335 79567
rect 89335 76575 92335 76583
rect 92525 79567 95525 79575
rect 92525 76583 92533 79567
rect 95517 76583 95525 79567
rect 92525 76575 95525 76583
rect 95715 79567 98715 79575
rect 95715 76583 95723 79567
rect 98707 76583 98715 79567
rect 95715 76575 98715 76583
rect 98905 79567 101905 79575
rect 98905 76583 98913 79567
rect 101897 76583 101905 79567
rect 98905 76575 101905 76583
rect 102095 79567 105095 79575
rect 102095 76583 102103 79567
rect 105087 76583 105095 79567
rect 102095 76575 105095 76583
rect 105285 79567 108285 79575
rect 105285 76583 105293 79567
rect 108277 76583 108285 79567
rect 105285 76575 108285 76583
rect 108475 79567 111475 79575
rect 108475 76583 108483 79567
rect 111467 76583 111475 79567
rect 108475 76575 111475 76583
rect 111665 79567 114665 79575
rect 111665 76583 111673 79567
rect 114657 76583 114665 79567
rect 111665 76575 114665 76583
rect 114855 79567 117855 79575
rect 114855 76583 114863 79567
rect 117847 76583 117855 79567
rect 114855 76575 117855 76583
rect 118045 79567 121045 79575
rect 118045 76583 118053 79567
rect 121037 76583 121045 79567
rect 118045 76575 121045 76583
rect 121235 79567 124235 79575
rect 121235 76583 121243 79567
rect 124227 76583 124235 79567
rect 121235 76575 124235 76583
rect 124425 79567 127425 79575
rect 124425 76583 124433 79567
rect 127417 76583 127425 79567
rect 124425 76575 127425 76583
rect 127615 79567 130615 79575
rect 127615 76583 127623 79567
rect 130607 76583 130615 79567
rect 127615 76575 130615 76583
rect 130805 79567 133805 79575
rect 130805 76583 130813 79567
rect 133797 76583 133805 79567
rect 130805 76575 133805 76583
rect 133995 79567 136995 79575
rect 133995 76583 134003 79567
rect 136987 76583 136995 79567
rect 133995 76575 136995 76583
rect 15 76377 3015 76385
rect 15 73393 23 76377
rect 3007 73393 3015 76377
rect 15 73385 3015 73393
rect 3205 76377 6205 76385
rect 3205 73393 3213 76377
rect 6197 73393 6205 76377
rect 3205 73385 6205 73393
rect 6395 76377 9395 76385
rect 6395 73393 6403 76377
rect 9387 73393 9395 76377
rect 6395 73385 9395 73393
rect 9585 76377 12585 76385
rect 9585 73393 9593 76377
rect 12577 73393 12585 76377
rect 9585 73385 12585 73393
rect 12775 76377 15775 76385
rect 12775 73393 12783 76377
rect 15767 73393 15775 76377
rect 12775 73385 15775 73393
rect 15965 76377 18965 76385
rect 15965 73393 15973 76377
rect 18957 73393 18965 76377
rect 15965 73385 18965 73393
rect 19155 76377 22155 76385
rect 19155 73393 19163 76377
rect 22147 73393 22155 76377
rect 19155 73385 22155 73393
rect 22345 76377 25345 76385
rect 22345 73393 22353 76377
rect 25337 73393 25345 76377
rect 22345 73385 25345 73393
rect 25535 76377 28535 76385
rect 25535 73393 25543 76377
rect 28527 73393 28535 76377
rect 25535 73385 28535 73393
rect 28725 76377 31725 76385
rect 28725 73393 28733 76377
rect 31717 73393 31725 76377
rect 28725 73385 31725 73393
rect 31915 76377 34915 76385
rect 31915 73393 31923 76377
rect 34907 73393 34915 76377
rect 31915 73385 34915 73393
rect 35105 76377 38105 76385
rect 35105 73393 35113 76377
rect 38097 73393 38105 76377
rect 35105 73385 38105 73393
rect 38295 76377 41295 76385
rect 38295 73393 38303 76377
rect 41287 73393 41295 76377
rect 38295 73385 41295 73393
rect 41485 76377 44485 76385
rect 41485 73393 41493 76377
rect 44477 73393 44485 76377
rect 41485 73385 44485 73393
rect 44675 76377 47675 76385
rect 44675 73393 44683 76377
rect 47667 73393 47675 76377
rect 44675 73385 47675 73393
rect 47865 76377 50865 76385
rect 47865 73393 47873 76377
rect 50857 73393 50865 76377
rect 47865 73385 50865 73393
rect 51055 76377 54055 76385
rect 51055 73393 51063 76377
rect 54047 73393 54055 76377
rect 51055 73385 54055 73393
rect 54245 76377 57245 76385
rect 54245 73393 54253 76377
rect 57237 73393 57245 76377
rect 54245 73385 57245 73393
rect 57435 76377 60435 76385
rect 57435 73393 57443 76377
rect 60427 73393 60435 76377
rect 57435 73385 60435 73393
rect 60625 76377 63625 76385
rect 60625 73393 60633 76377
rect 63617 73393 63625 76377
rect 60625 73385 63625 73393
rect 63815 76377 66815 76385
rect 63815 73393 63823 76377
rect 66807 73393 66815 76377
rect 63815 73385 66815 73393
rect 67005 76377 70005 76385
rect 67005 73393 67013 76377
rect 69997 73393 70005 76377
rect 67005 73385 70005 73393
rect 70195 76377 73195 76385
rect 70195 73393 70203 76377
rect 73187 73393 73195 76377
rect 70195 73385 73195 73393
rect 73385 76377 76385 76385
rect 73385 73393 73393 76377
rect 76377 73393 76385 76377
rect 73385 73385 76385 73393
rect 76575 76377 79575 76385
rect 76575 73393 76583 76377
rect 79567 73393 79575 76377
rect 76575 73385 79575 73393
rect 79765 76377 82765 76385
rect 79765 73393 79773 76377
rect 82757 73393 82765 76377
rect 79765 73385 82765 73393
rect 82955 76377 85955 76385
rect 82955 73393 82963 76377
rect 85947 73393 85955 76377
rect 82955 73385 85955 73393
rect 86145 76377 89145 76385
rect 86145 73393 86153 76377
rect 89137 73393 89145 76377
rect 86145 73385 89145 73393
rect 89335 76377 92335 76385
rect 89335 73393 89343 76377
rect 92327 73393 92335 76377
rect 89335 73385 92335 73393
rect 92525 76377 95525 76385
rect 92525 73393 92533 76377
rect 95517 73393 95525 76377
rect 92525 73385 95525 73393
rect 95715 76377 98715 76385
rect 95715 73393 95723 76377
rect 98707 73393 98715 76377
rect 95715 73385 98715 73393
rect 98905 76377 101905 76385
rect 98905 73393 98913 76377
rect 101897 73393 101905 76377
rect 98905 73385 101905 73393
rect 102095 76377 105095 76385
rect 102095 73393 102103 76377
rect 105087 73393 105095 76377
rect 102095 73385 105095 73393
rect 105285 76377 108285 76385
rect 105285 73393 105293 76377
rect 108277 73393 108285 76377
rect 105285 73385 108285 73393
rect 108475 76377 111475 76385
rect 108475 73393 108483 76377
rect 111467 73393 111475 76377
rect 108475 73385 111475 73393
rect 111665 76377 114665 76385
rect 111665 73393 111673 76377
rect 114657 73393 114665 76377
rect 111665 73385 114665 73393
rect 114855 76377 117855 76385
rect 114855 73393 114863 76377
rect 117847 73393 117855 76377
rect 114855 73385 117855 73393
rect 118045 76377 121045 76385
rect 118045 73393 118053 76377
rect 121037 73393 121045 76377
rect 118045 73385 121045 73393
rect 121235 76377 124235 76385
rect 121235 73393 121243 76377
rect 124227 73393 124235 76377
rect 121235 73385 124235 73393
rect 124425 76377 127425 76385
rect 124425 73393 124433 76377
rect 127417 73393 127425 76377
rect 124425 73385 127425 73393
rect 127615 76377 130615 76385
rect 127615 73393 127623 76377
rect 130607 73393 130615 76377
rect 127615 73385 130615 73393
rect 130805 76377 133805 76385
rect 130805 73393 130813 76377
rect 133797 73393 133805 76377
rect 130805 73385 133805 73393
rect 133995 76377 136995 76385
rect 133995 73393 134003 76377
rect 136987 73393 136995 76377
rect 133995 73385 136995 73393
rect 15 73187 3015 73195
rect 15 70203 23 73187
rect 3007 70203 3015 73187
rect 15 70195 3015 70203
rect 3205 73187 6205 73195
rect 3205 70203 3213 73187
rect 6197 70203 6205 73187
rect 3205 70195 6205 70203
rect 6395 73187 9395 73195
rect 6395 70203 6403 73187
rect 9387 70203 9395 73187
rect 6395 70195 9395 70203
rect 9585 73187 12585 73195
rect 9585 70203 9593 73187
rect 12577 70203 12585 73187
rect 9585 70195 12585 70203
rect 12775 73187 15775 73195
rect 12775 70203 12783 73187
rect 15767 70203 15775 73187
rect 12775 70195 15775 70203
rect 15965 73187 18965 73195
rect 15965 70203 15973 73187
rect 18957 70203 18965 73187
rect 15965 70195 18965 70203
rect 19155 73187 22155 73195
rect 19155 70203 19163 73187
rect 22147 70203 22155 73187
rect 19155 70195 22155 70203
rect 22345 73187 25345 73195
rect 22345 70203 22353 73187
rect 25337 70203 25345 73187
rect 22345 70195 25345 70203
rect 25535 73187 28535 73195
rect 25535 70203 25543 73187
rect 28527 70203 28535 73187
rect 25535 70195 28535 70203
rect 28725 73187 31725 73195
rect 28725 70203 28733 73187
rect 31717 70203 31725 73187
rect 28725 70195 31725 70203
rect 31915 73187 34915 73195
rect 31915 70203 31923 73187
rect 34907 70203 34915 73187
rect 31915 70195 34915 70203
rect 35105 73187 38105 73195
rect 35105 70203 35113 73187
rect 38097 70203 38105 73187
rect 35105 70195 38105 70203
rect 38295 73187 41295 73195
rect 38295 70203 38303 73187
rect 41287 70203 41295 73187
rect 38295 70195 41295 70203
rect 41485 73187 44485 73195
rect 41485 70203 41493 73187
rect 44477 70203 44485 73187
rect 41485 70195 44485 70203
rect 44675 73187 47675 73195
rect 44675 70203 44683 73187
rect 47667 70203 47675 73187
rect 44675 70195 47675 70203
rect 47865 73187 50865 73195
rect 47865 70203 47873 73187
rect 50857 70203 50865 73187
rect 47865 70195 50865 70203
rect 51055 73187 54055 73195
rect 51055 70203 51063 73187
rect 54047 70203 54055 73187
rect 51055 70195 54055 70203
rect 54245 73187 57245 73195
rect 54245 70203 54253 73187
rect 57237 70203 57245 73187
rect 54245 70195 57245 70203
rect 57435 73187 60435 73195
rect 57435 70203 57443 73187
rect 60427 70203 60435 73187
rect 57435 70195 60435 70203
rect 60625 73187 63625 73195
rect 60625 70203 60633 73187
rect 63617 70203 63625 73187
rect 60625 70195 63625 70203
rect 63815 73187 66815 73195
rect 63815 70203 63823 73187
rect 66807 70203 66815 73187
rect 63815 70195 66815 70203
rect 67005 73187 70005 73195
rect 67005 70203 67013 73187
rect 69997 70203 70005 73187
rect 67005 70195 70005 70203
rect 70195 73187 73195 73195
rect 70195 70203 70203 73187
rect 73187 70203 73195 73187
rect 70195 70195 73195 70203
rect 73385 73187 76385 73195
rect 73385 70203 73393 73187
rect 76377 70203 76385 73187
rect 73385 70195 76385 70203
rect 76575 73187 79575 73195
rect 76575 70203 76583 73187
rect 79567 70203 79575 73187
rect 76575 70195 79575 70203
rect 79765 73187 82765 73195
rect 79765 70203 79773 73187
rect 82757 70203 82765 73187
rect 79765 70195 82765 70203
rect 82955 73187 85955 73195
rect 82955 70203 82963 73187
rect 85947 70203 85955 73187
rect 82955 70195 85955 70203
rect 86145 73187 89145 73195
rect 86145 70203 86153 73187
rect 89137 70203 89145 73187
rect 86145 70195 89145 70203
rect 89335 73187 92335 73195
rect 89335 70203 89343 73187
rect 92327 70203 92335 73187
rect 89335 70195 92335 70203
rect 92525 73187 95525 73195
rect 92525 70203 92533 73187
rect 95517 70203 95525 73187
rect 92525 70195 95525 70203
rect 95715 73187 98715 73195
rect 95715 70203 95723 73187
rect 98707 70203 98715 73187
rect 95715 70195 98715 70203
rect 98905 73187 101905 73195
rect 98905 70203 98913 73187
rect 101897 70203 101905 73187
rect 98905 70195 101905 70203
rect 102095 73187 105095 73195
rect 102095 70203 102103 73187
rect 105087 70203 105095 73187
rect 102095 70195 105095 70203
rect 105285 73187 108285 73195
rect 105285 70203 105293 73187
rect 108277 70203 108285 73187
rect 105285 70195 108285 70203
rect 108475 73187 111475 73195
rect 108475 70203 108483 73187
rect 111467 70203 111475 73187
rect 108475 70195 111475 70203
rect 111665 73187 114665 73195
rect 111665 70203 111673 73187
rect 114657 70203 114665 73187
rect 111665 70195 114665 70203
rect 114855 73187 117855 73195
rect 114855 70203 114863 73187
rect 117847 70203 117855 73187
rect 114855 70195 117855 70203
rect 118045 73187 121045 73195
rect 118045 70203 118053 73187
rect 121037 70203 121045 73187
rect 118045 70195 121045 70203
rect 121235 73187 124235 73195
rect 121235 70203 121243 73187
rect 124227 70203 124235 73187
rect 121235 70195 124235 70203
rect 124425 73187 127425 73195
rect 124425 70203 124433 73187
rect 127417 70203 127425 73187
rect 124425 70195 127425 70203
rect 127615 73187 130615 73195
rect 127615 70203 127623 73187
rect 130607 70203 130615 73187
rect 127615 70195 130615 70203
rect 130805 73187 133805 73195
rect 130805 70203 130813 73187
rect 133797 70203 133805 73187
rect 130805 70195 133805 70203
rect 133995 73187 136995 73195
rect 133995 70203 134003 73187
rect 136987 70203 136995 73187
rect 133995 70195 136995 70203
rect 15 69997 3015 70005
rect 15 67013 23 69997
rect 3007 67013 3015 69997
rect 15 67005 3015 67013
rect 3205 69997 6205 70005
rect 3205 67013 3213 69997
rect 6197 67013 6205 69997
rect 3205 67005 6205 67013
rect 6395 69997 9395 70005
rect 6395 67013 6403 69997
rect 9387 67013 9395 69997
rect 6395 67005 9395 67013
rect 9585 69997 12585 70005
rect 9585 67013 9593 69997
rect 12577 67013 12585 69997
rect 9585 67005 12585 67013
rect 12775 69997 15775 70005
rect 12775 67013 12783 69997
rect 15767 67013 15775 69997
rect 12775 67005 15775 67013
rect 15965 69997 18965 70005
rect 15965 67013 15973 69997
rect 18957 67013 18965 69997
rect 15965 67005 18965 67013
rect 19155 69997 22155 70005
rect 19155 67013 19163 69997
rect 22147 67013 22155 69997
rect 19155 67005 22155 67013
rect 22345 69997 25345 70005
rect 22345 67013 22353 69997
rect 25337 67013 25345 69997
rect 22345 67005 25345 67013
rect 25535 69997 28535 70005
rect 25535 67013 25543 69997
rect 28527 67013 28535 69997
rect 25535 67005 28535 67013
rect 28725 69997 31725 70005
rect 28725 67013 28733 69997
rect 31717 67013 31725 69997
rect 28725 67005 31725 67013
rect 31915 69997 34915 70005
rect 31915 67013 31923 69997
rect 34907 67013 34915 69997
rect 31915 67005 34915 67013
rect 35105 69997 38105 70005
rect 35105 67013 35113 69997
rect 38097 67013 38105 69997
rect 35105 67005 38105 67013
rect 38295 69997 41295 70005
rect 38295 67013 38303 69997
rect 41287 67013 41295 69997
rect 38295 67005 41295 67013
rect 41485 69997 44485 70005
rect 41485 67013 41493 69997
rect 44477 67013 44485 69997
rect 41485 67005 44485 67013
rect 44675 69997 47675 70005
rect 44675 67013 44683 69997
rect 47667 67013 47675 69997
rect 44675 67005 47675 67013
rect 47865 69997 50865 70005
rect 47865 67013 47873 69997
rect 50857 67013 50865 69997
rect 47865 67005 50865 67013
rect 51055 69997 54055 70005
rect 51055 67013 51063 69997
rect 54047 67013 54055 69997
rect 51055 67005 54055 67013
rect 54245 69997 57245 70005
rect 54245 67013 54253 69997
rect 57237 67013 57245 69997
rect 54245 67005 57245 67013
rect 57435 69997 60435 70005
rect 57435 67013 57443 69997
rect 60427 67013 60435 69997
rect 57435 67005 60435 67013
rect 60625 69997 63625 70005
rect 60625 67013 60633 69997
rect 63617 67013 63625 69997
rect 60625 67005 63625 67013
rect 63815 69997 66815 70005
rect 63815 67013 63823 69997
rect 66807 67013 66815 69997
rect 63815 67005 66815 67013
rect 67005 69997 70005 70005
rect 67005 67013 67013 69997
rect 69997 67013 70005 69997
rect 67005 67005 70005 67013
rect 70195 69997 73195 70005
rect 70195 67013 70203 69997
rect 73187 67013 73195 69997
rect 70195 67005 73195 67013
rect 73385 69997 76385 70005
rect 73385 67013 73393 69997
rect 76377 67013 76385 69997
rect 73385 67005 76385 67013
rect 76575 69997 79575 70005
rect 76575 67013 76583 69997
rect 79567 67013 79575 69997
rect 76575 67005 79575 67013
rect 79765 69997 82765 70005
rect 79765 67013 79773 69997
rect 82757 67013 82765 69997
rect 79765 67005 82765 67013
rect 82955 69997 85955 70005
rect 82955 67013 82963 69997
rect 85947 67013 85955 69997
rect 82955 67005 85955 67013
rect 86145 69997 89145 70005
rect 86145 67013 86153 69997
rect 89137 67013 89145 69997
rect 86145 67005 89145 67013
rect 89335 69997 92335 70005
rect 89335 67013 89343 69997
rect 92327 67013 92335 69997
rect 89335 67005 92335 67013
rect 92525 69997 95525 70005
rect 92525 67013 92533 69997
rect 95517 67013 95525 69997
rect 92525 67005 95525 67013
rect 95715 69997 98715 70005
rect 95715 67013 95723 69997
rect 98707 67013 98715 69997
rect 95715 67005 98715 67013
rect 98905 69997 101905 70005
rect 98905 67013 98913 69997
rect 101897 67013 101905 69997
rect 98905 67005 101905 67013
rect 102095 69997 105095 70005
rect 102095 67013 102103 69997
rect 105087 67013 105095 69997
rect 102095 67005 105095 67013
rect 105285 69997 108285 70005
rect 105285 67013 105293 69997
rect 108277 67013 108285 69997
rect 105285 67005 108285 67013
rect 108475 69997 111475 70005
rect 108475 67013 108483 69997
rect 111467 67013 111475 69997
rect 108475 67005 111475 67013
rect 111665 69997 114665 70005
rect 111665 67013 111673 69997
rect 114657 67013 114665 69997
rect 111665 67005 114665 67013
rect 114855 69997 117855 70005
rect 114855 67013 114863 69997
rect 117847 67013 117855 69997
rect 114855 67005 117855 67013
rect 118045 69997 121045 70005
rect 118045 67013 118053 69997
rect 121037 67013 121045 69997
rect 118045 67005 121045 67013
rect 121235 69997 124235 70005
rect 121235 67013 121243 69997
rect 124227 67013 124235 69997
rect 121235 67005 124235 67013
rect 124425 69997 127425 70005
rect 124425 67013 124433 69997
rect 127417 67013 127425 69997
rect 124425 67005 127425 67013
rect 127615 69997 130615 70005
rect 127615 67013 127623 69997
rect 130607 67013 130615 69997
rect 127615 67005 130615 67013
rect 130805 69997 133805 70005
rect 130805 67013 130813 69997
rect 133797 67013 133805 69997
rect 130805 67005 133805 67013
rect 133995 69997 136995 70005
rect 133995 67013 134003 69997
rect 136987 67013 136995 69997
rect 133995 67005 136995 67013
rect 15 66807 3015 66815
rect 15 63823 23 66807
rect 3007 63823 3015 66807
rect 15 63815 3015 63823
rect 3205 66807 6205 66815
rect 3205 63823 3213 66807
rect 6197 63823 6205 66807
rect 3205 63815 6205 63823
rect 6395 66807 9395 66815
rect 6395 63823 6403 66807
rect 9387 63823 9395 66807
rect 6395 63815 9395 63823
rect 9585 66807 12585 66815
rect 9585 63823 9593 66807
rect 12577 63823 12585 66807
rect 9585 63815 12585 63823
rect 12775 66807 15775 66815
rect 12775 63823 12783 66807
rect 15767 63823 15775 66807
rect 12775 63815 15775 63823
rect 15965 66807 18965 66815
rect 15965 63823 15973 66807
rect 18957 63823 18965 66807
rect 15965 63815 18965 63823
rect 19155 66807 22155 66815
rect 19155 63823 19163 66807
rect 22147 63823 22155 66807
rect 19155 63815 22155 63823
rect 22345 66807 25345 66815
rect 22345 63823 22353 66807
rect 25337 63823 25345 66807
rect 22345 63815 25345 63823
rect 25535 66807 28535 66815
rect 25535 63823 25543 66807
rect 28527 63823 28535 66807
rect 25535 63815 28535 63823
rect 28725 66807 31725 66815
rect 28725 63823 28733 66807
rect 31717 63823 31725 66807
rect 28725 63815 31725 63823
rect 31915 66807 34915 66815
rect 31915 63823 31923 66807
rect 34907 63823 34915 66807
rect 31915 63815 34915 63823
rect 35105 66807 38105 66815
rect 35105 63823 35113 66807
rect 38097 63823 38105 66807
rect 35105 63815 38105 63823
rect 38295 66807 41295 66815
rect 38295 63823 38303 66807
rect 41287 63823 41295 66807
rect 38295 63815 41295 63823
rect 41485 66807 44485 66815
rect 41485 63823 41493 66807
rect 44477 63823 44485 66807
rect 41485 63815 44485 63823
rect 44675 66807 47675 66815
rect 44675 63823 44683 66807
rect 47667 63823 47675 66807
rect 44675 63815 47675 63823
rect 47865 66807 50865 66815
rect 47865 63823 47873 66807
rect 50857 63823 50865 66807
rect 47865 63815 50865 63823
rect 51055 66807 54055 66815
rect 51055 63823 51063 66807
rect 54047 63823 54055 66807
rect 51055 63815 54055 63823
rect 54245 66807 57245 66815
rect 54245 63823 54253 66807
rect 57237 63823 57245 66807
rect 54245 63815 57245 63823
rect 57435 66807 60435 66815
rect 57435 63823 57443 66807
rect 60427 63823 60435 66807
rect 57435 63815 60435 63823
rect 60625 66807 63625 66815
rect 60625 63823 60633 66807
rect 63617 63823 63625 66807
rect 60625 63815 63625 63823
rect 63815 66807 66815 66815
rect 63815 63823 63823 66807
rect 66807 63823 66815 66807
rect 63815 63815 66815 63823
rect 67005 66807 70005 66815
rect 67005 63823 67013 66807
rect 69997 63823 70005 66807
rect 67005 63815 70005 63823
rect 70195 66807 73195 66815
rect 70195 63823 70203 66807
rect 73187 63823 73195 66807
rect 70195 63815 73195 63823
rect 73385 66807 76385 66815
rect 73385 63823 73393 66807
rect 76377 63823 76385 66807
rect 73385 63815 76385 63823
rect 76575 66807 79575 66815
rect 76575 63823 76583 66807
rect 79567 63823 79575 66807
rect 76575 63815 79575 63823
rect 79765 66807 82765 66815
rect 79765 63823 79773 66807
rect 82757 63823 82765 66807
rect 79765 63815 82765 63823
rect 82955 66807 85955 66815
rect 82955 63823 82963 66807
rect 85947 63823 85955 66807
rect 82955 63815 85955 63823
rect 86145 66807 89145 66815
rect 86145 63823 86153 66807
rect 89137 63823 89145 66807
rect 86145 63815 89145 63823
rect 89335 66807 92335 66815
rect 89335 63823 89343 66807
rect 92327 63823 92335 66807
rect 89335 63815 92335 63823
rect 92525 66807 95525 66815
rect 92525 63823 92533 66807
rect 95517 63823 95525 66807
rect 92525 63815 95525 63823
rect 95715 66807 98715 66815
rect 95715 63823 95723 66807
rect 98707 63823 98715 66807
rect 95715 63815 98715 63823
rect 98905 66807 101905 66815
rect 98905 63823 98913 66807
rect 101897 63823 101905 66807
rect 98905 63815 101905 63823
rect 102095 66807 105095 66815
rect 102095 63823 102103 66807
rect 105087 63823 105095 66807
rect 102095 63815 105095 63823
rect 105285 66807 108285 66815
rect 105285 63823 105293 66807
rect 108277 63823 108285 66807
rect 105285 63815 108285 63823
rect 108475 66807 111475 66815
rect 108475 63823 108483 66807
rect 111467 63823 111475 66807
rect 108475 63815 111475 63823
rect 111665 66807 114665 66815
rect 111665 63823 111673 66807
rect 114657 63823 114665 66807
rect 111665 63815 114665 63823
rect 114855 66807 117855 66815
rect 114855 63823 114863 66807
rect 117847 63823 117855 66807
rect 114855 63815 117855 63823
rect 118045 66807 121045 66815
rect 118045 63823 118053 66807
rect 121037 63823 121045 66807
rect 118045 63815 121045 63823
rect 121235 66807 124235 66815
rect 121235 63823 121243 66807
rect 124227 63823 124235 66807
rect 121235 63815 124235 63823
rect 124425 66807 127425 66815
rect 124425 63823 124433 66807
rect 127417 63823 127425 66807
rect 124425 63815 127425 63823
rect 127615 66807 130615 66815
rect 127615 63823 127623 66807
rect 130607 63823 130615 66807
rect 127615 63815 130615 63823
rect 130805 66807 133805 66815
rect 130805 63823 130813 66807
rect 133797 63823 133805 66807
rect 130805 63815 133805 63823
rect 133995 66807 136995 66815
rect 133995 63823 134003 66807
rect 136987 63823 136995 66807
rect 133995 63815 136995 63823
rect 15 63617 3015 63625
rect 15 60633 23 63617
rect 3007 60633 3015 63617
rect 15 60625 3015 60633
rect 3205 63617 6205 63625
rect 3205 60633 3213 63617
rect 6197 60633 6205 63617
rect 3205 60625 6205 60633
rect 6395 63617 9395 63625
rect 6395 60633 6403 63617
rect 9387 60633 9395 63617
rect 6395 60625 9395 60633
rect 9585 63617 12585 63625
rect 9585 60633 9593 63617
rect 12577 60633 12585 63617
rect 9585 60625 12585 60633
rect 12775 63617 15775 63625
rect 12775 60633 12783 63617
rect 15767 60633 15775 63617
rect 12775 60625 15775 60633
rect 15965 63617 18965 63625
rect 15965 60633 15973 63617
rect 18957 60633 18965 63617
rect 15965 60625 18965 60633
rect 19155 63617 22155 63625
rect 19155 60633 19163 63617
rect 22147 60633 22155 63617
rect 19155 60625 22155 60633
rect 22345 63617 25345 63625
rect 22345 60633 22353 63617
rect 25337 60633 25345 63617
rect 22345 60625 25345 60633
rect 25535 63617 28535 63625
rect 25535 60633 25543 63617
rect 28527 60633 28535 63617
rect 25535 60625 28535 60633
rect 28725 63617 31725 63625
rect 28725 60633 28733 63617
rect 31717 60633 31725 63617
rect 28725 60625 31725 60633
rect 31915 63617 34915 63625
rect 31915 60633 31923 63617
rect 34907 60633 34915 63617
rect 31915 60625 34915 60633
rect 35105 63617 38105 63625
rect 35105 60633 35113 63617
rect 38097 60633 38105 63617
rect 35105 60625 38105 60633
rect 38295 63617 41295 63625
rect 38295 60633 38303 63617
rect 41287 60633 41295 63617
rect 38295 60625 41295 60633
rect 41485 63617 44485 63625
rect 41485 60633 41493 63617
rect 44477 60633 44485 63617
rect 41485 60625 44485 60633
rect 44675 63617 47675 63625
rect 44675 60633 44683 63617
rect 47667 60633 47675 63617
rect 44675 60625 47675 60633
rect 47865 63617 50865 63625
rect 47865 60633 47873 63617
rect 50857 60633 50865 63617
rect 47865 60625 50865 60633
rect 51055 63617 54055 63625
rect 51055 60633 51063 63617
rect 54047 60633 54055 63617
rect 51055 60625 54055 60633
rect 54245 63617 57245 63625
rect 54245 60633 54253 63617
rect 57237 60633 57245 63617
rect 54245 60625 57245 60633
rect 57435 63617 60435 63625
rect 57435 60633 57443 63617
rect 60427 60633 60435 63617
rect 57435 60625 60435 60633
rect 60625 63617 63625 63625
rect 60625 60633 60633 63617
rect 63617 60633 63625 63617
rect 60625 60625 63625 60633
rect 63815 63617 66815 63625
rect 63815 60633 63823 63617
rect 66807 60633 66815 63617
rect 63815 60625 66815 60633
rect 67005 63617 70005 63625
rect 67005 60633 67013 63617
rect 69997 60633 70005 63617
rect 67005 60625 70005 60633
rect 70195 63617 73195 63625
rect 70195 60633 70203 63617
rect 73187 60633 73195 63617
rect 70195 60625 73195 60633
rect 73385 63617 76385 63625
rect 73385 60633 73393 63617
rect 76377 60633 76385 63617
rect 73385 60625 76385 60633
rect 76575 63617 79575 63625
rect 76575 60633 76583 63617
rect 79567 60633 79575 63617
rect 76575 60625 79575 60633
rect 79765 63617 82765 63625
rect 79765 60633 79773 63617
rect 82757 60633 82765 63617
rect 79765 60625 82765 60633
rect 82955 63617 85955 63625
rect 82955 60633 82963 63617
rect 85947 60633 85955 63617
rect 82955 60625 85955 60633
rect 86145 63617 89145 63625
rect 86145 60633 86153 63617
rect 89137 60633 89145 63617
rect 86145 60625 89145 60633
rect 89335 63617 92335 63625
rect 89335 60633 89343 63617
rect 92327 60633 92335 63617
rect 89335 60625 92335 60633
rect 92525 63617 95525 63625
rect 92525 60633 92533 63617
rect 95517 60633 95525 63617
rect 92525 60625 95525 60633
rect 95715 63617 98715 63625
rect 95715 60633 95723 63617
rect 98707 60633 98715 63617
rect 95715 60625 98715 60633
rect 98905 63617 101905 63625
rect 98905 60633 98913 63617
rect 101897 60633 101905 63617
rect 98905 60625 101905 60633
rect 102095 63617 105095 63625
rect 102095 60633 102103 63617
rect 105087 60633 105095 63617
rect 102095 60625 105095 60633
rect 105285 63617 108285 63625
rect 105285 60633 105293 63617
rect 108277 60633 108285 63617
rect 105285 60625 108285 60633
rect 108475 63617 111475 63625
rect 108475 60633 108483 63617
rect 111467 60633 111475 63617
rect 108475 60625 111475 60633
rect 111665 63617 114665 63625
rect 111665 60633 111673 63617
rect 114657 60633 114665 63617
rect 111665 60625 114665 60633
rect 114855 63617 117855 63625
rect 114855 60633 114863 63617
rect 117847 60633 117855 63617
rect 114855 60625 117855 60633
rect 118045 63617 121045 63625
rect 118045 60633 118053 63617
rect 121037 60633 121045 63617
rect 118045 60625 121045 60633
rect 121235 63617 124235 63625
rect 121235 60633 121243 63617
rect 124227 60633 124235 63617
rect 121235 60625 124235 60633
rect 124425 63617 127425 63625
rect 124425 60633 124433 63617
rect 127417 60633 127425 63617
rect 124425 60625 127425 60633
rect 127615 63617 130615 63625
rect 127615 60633 127623 63617
rect 130607 60633 130615 63617
rect 127615 60625 130615 60633
rect 130805 63617 133805 63625
rect 130805 60633 130813 63617
rect 133797 60633 133805 63617
rect 130805 60625 133805 60633
rect 133995 63617 136995 63625
rect 133995 60633 134003 63617
rect 136987 60633 136995 63617
rect 133995 60625 136995 60633
rect 15 60427 3015 60435
rect 15 57443 23 60427
rect 3007 57443 3015 60427
rect 15 57435 3015 57443
rect 3205 60427 6205 60435
rect 3205 57443 3213 60427
rect 6197 57443 6205 60427
rect 3205 57435 6205 57443
rect 6395 60427 9395 60435
rect 6395 57443 6403 60427
rect 9387 57443 9395 60427
rect 6395 57435 9395 57443
rect 9585 60427 12585 60435
rect 9585 57443 9593 60427
rect 12577 57443 12585 60427
rect 9585 57435 12585 57443
rect 12775 60427 15775 60435
rect 12775 57443 12783 60427
rect 15767 57443 15775 60427
rect 12775 57435 15775 57443
rect 15965 60427 18965 60435
rect 15965 57443 15973 60427
rect 18957 57443 18965 60427
rect 15965 57435 18965 57443
rect 19155 60427 22155 60435
rect 19155 57443 19163 60427
rect 22147 57443 22155 60427
rect 19155 57435 22155 57443
rect 22345 60427 25345 60435
rect 22345 57443 22353 60427
rect 25337 57443 25345 60427
rect 22345 57435 25345 57443
rect 25535 60427 28535 60435
rect 25535 57443 25543 60427
rect 28527 57443 28535 60427
rect 25535 57435 28535 57443
rect 28725 60427 31725 60435
rect 28725 57443 28733 60427
rect 31717 57443 31725 60427
rect 28725 57435 31725 57443
rect 31915 60427 34915 60435
rect 31915 57443 31923 60427
rect 34907 57443 34915 60427
rect 31915 57435 34915 57443
rect 35105 60427 38105 60435
rect 35105 57443 35113 60427
rect 38097 57443 38105 60427
rect 35105 57435 38105 57443
rect 38295 60427 41295 60435
rect 38295 57443 38303 60427
rect 41287 57443 41295 60427
rect 38295 57435 41295 57443
rect 41485 60427 44485 60435
rect 41485 57443 41493 60427
rect 44477 57443 44485 60427
rect 41485 57435 44485 57443
rect 44675 60427 47675 60435
rect 44675 57443 44683 60427
rect 47667 57443 47675 60427
rect 44675 57435 47675 57443
rect 47865 60427 50865 60435
rect 47865 57443 47873 60427
rect 50857 57443 50865 60427
rect 47865 57435 50865 57443
rect 51055 60427 54055 60435
rect 51055 57443 51063 60427
rect 54047 57443 54055 60427
rect 51055 57435 54055 57443
rect 54245 60427 57245 60435
rect 54245 57443 54253 60427
rect 57237 57443 57245 60427
rect 54245 57435 57245 57443
rect 57435 60427 60435 60435
rect 57435 57443 57443 60427
rect 60427 57443 60435 60427
rect 57435 57435 60435 57443
rect 60625 60427 63625 60435
rect 60625 57443 60633 60427
rect 63617 57443 63625 60427
rect 60625 57435 63625 57443
rect 63815 60427 66815 60435
rect 63815 57443 63823 60427
rect 66807 57443 66815 60427
rect 63815 57435 66815 57443
rect 67005 60427 70005 60435
rect 67005 57443 67013 60427
rect 69997 57443 70005 60427
rect 67005 57435 70005 57443
rect 70195 60427 73195 60435
rect 70195 57443 70203 60427
rect 73187 57443 73195 60427
rect 70195 57435 73195 57443
rect 73385 60427 76385 60435
rect 73385 57443 73393 60427
rect 76377 57443 76385 60427
rect 73385 57435 76385 57443
rect 76575 60427 79575 60435
rect 76575 57443 76583 60427
rect 79567 57443 79575 60427
rect 76575 57435 79575 57443
rect 79765 60427 82765 60435
rect 79765 57443 79773 60427
rect 82757 57443 82765 60427
rect 79765 57435 82765 57443
rect 82955 60427 85955 60435
rect 82955 57443 82963 60427
rect 85947 57443 85955 60427
rect 82955 57435 85955 57443
rect 86145 60427 89145 60435
rect 86145 57443 86153 60427
rect 89137 57443 89145 60427
rect 86145 57435 89145 57443
rect 89335 60427 92335 60435
rect 89335 57443 89343 60427
rect 92327 57443 92335 60427
rect 89335 57435 92335 57443
rect 92525 60427 95525 60435
rect 92525 57443 92533 60427
rect 95517 57443 95525 60427
rect 92525 57435 95525 57443
rect 95715 60427 98715 60435
rect 95715 57443 95723 60427
rect 98707 57443 98715 60427
rect 95715 57435 98715 57443
rect 98905 60427 101905 60435
rect 98905 57443 98913 60427
rect 101897 57443 101905 60427
rect 98905 57435 101905 57443
rect 102095 60427 105095 60435
rect 102095 57443 102103 60427
rect 105087 57443 105095 60427
rect 102095 57435 105095 57443
rect 105285 60427 108285 60435
rect 105285 57443 105293 60427
rect 108277 57443 108285 60427
rect 105285 57435 108285 57443
rect 108475 60427 111475 60435
rect 108475 57443 108483 60427
rect 111467 57443 111475 60427
rect 108475 57435 111475 57443
rect 111665 60427 114665 60435
rect 111665 57443 111673 60427
rect 114657 57443 114665 60427
rect 111665 57435 114665 57443
rect 114855 60427 117855 60435
rect 114855 57443 114863 60427
rect 117847 57443 117855 60427
rect 114855 57435 117855 57443
rect 118045 60427 121045 60435
rect 118045 57443 118053 60427
rect 121037 57443 121045 60427
rect 118045 57435 121045 57443
rect 121235 60427 124235 60435
rect 121235 57443 121243 60427
rect 124227 57443 124235 60427
rect 121235 57435 124235 57443
rect 124425 60427 127425 60435
rect 124425 57443 124433 60427
rect 127417 57443 127425 60427
rect 124425 57435 127425 57443
rect 127615 60427 130615 60435
rect 127615 57443 127623 60427
rect 130607 57443 130615 60427
rect 127615 57435 130615 57443
rect 130805 60427 133805 60435
rect 130805 57443 130813 60427
rect 133797 57443 133805 60427
rect 130805 57435 133805 57443
rect 133995 60427 136995 60435
rect 133995 57443 134003 60427
rect 136987 57443 136995 60427
rect 133995 57435 136995 57443
rect 15 57237 3015 57245
rect 15 54253 23 57237
rect 3007 54253 3015 57237
rect 15 54245 3015 54253
rect 3205 57237 6205 57245
rect 3205 54253 3213 57237
rect 6197 54253 6205 57237
rect 3205 54245 6205 54253
rect 6395 57237 9395 57245
rect 6395 54253 6403 57237
rect 9387 54253 9395 57237
rect 6395 54245 9395 54253
rect 9585 57237 12585 57245
rect 9585 54253 9593 57237
rect 12577 54253 12585 57237
rect 9585 54245 12585 54253
rect 12775 57237 15775 57245
rect 12775 54253 12783 57237
rect 15767 54253 15775 57237
rect 12775 54245 15775 54253
rect 15965 57237 18965 57245
rect 15965 54253 15973 57237
rect 18957 54253 18965 57237
rect 15965 54245 18965 54253
rect 19155 57237 22155 57245
rect 19155 54253 19163 57237
rect 22147 54253 22155 57237
rect 19155 54245 22155 54253
rect 22345 57237 25345 57245
rect 22345 54253 22353 57237
rect 25337 54253 25345 57237
rect 22345 54245 25345 54253
rect 25535 57237 28535 57245
rect 25535 54253 25543 57237
rect 28527 54253 28535 57237
rect 25535 54245 28535 54253
rect 28725 57237 31725 57245
rect 28725 54253 28733 57237
rect 31717 54253 31725 57237
rect 28725 54245 31725 54253
rect 31915 57237 34915 57245
rect 31915 54253 31923 57237
rect 34907 54253 34915 57237
rect 31915 54245 34915 54253
rect 35105 57237 38105 57245
rect 35105 54253 35113 57237
rect 38097 54253 38105 57237
rect 35105 54245 38105 54253
rect 38295 57237 41295 57245
rect 38295 54253 38303 57237
rect 41287 54253 41295 57237
rect 38295 54245 41295 54253
rect 41485 57237 44485 57245
rect 41485 54253 41493 57237
rect 44477 54253 44485 57237
rect 41485 54245 44485 54253
rect 44675 57237 47675 57245
rect 44675 54253 44683 57237
rect 47667 54253 47675 57237
rect 44675 54245 47675 54253
rect 47865 57237 50865 57245
rect 47865 54253 47873 57237
rect 50857 54253 50865 57237
rect 47865 54245 50865 54253
rect 51055 57237 54055 57245
rect 51055 54253 51063 57237
rect 54047 54253 54055 57237
rect 51055 54245 54055 54253
rect 54245 57237 57245 57245
rect 54245 54253 54253 57237
rect 57237 54253 57245 57237
rect 54245 54245 57245 54253
rect 57435 57237 60435 57245
rect 57435 54253 57443 57237
rect 60427 54253 60435 57237
rect 57435 54245 60435 54253
rect 60625 57237 63625 57245
rect 60625 54253 60633 57237
rect 63617 54253 63625 57237
rect 60625 54245 63625 54253
rect 63815 57237 66815 57245
rect 63815 54253 63823 57237
rect 66807 54253 66815 57237
rect 63815 54245 66815 54253
rect 67005 57237 70005 57245
rect 67005 54253 67013 57237
rect 69997 54253 70005 57237
rect 67005 54245 70005 54253
rect 70195 57237 73195 57245
rect 70195 54253 70203 57237
rect 73187 54253 73195 57237
rect 70195 54245 73195 54253
rect 73385 57237 76385 57245
rect 73385 54253 73393 57237
rect 76377 54253 76385 57237
rect 73385 54245 76385 54253
rect 76575 57237 79575 57245
rect 76575 54253 76583 57237
rect 79567 54253 79575 57237
rect 76575 54245 79575 54253
rect 79765 57237 82765 57245
rect 79765 54253 79773 57237
rect 82757 54253 82765 57237
rect 79765 54245 82765 54253
rect 82955 57237 85955 57245
rect 82955 54253 82963 57237
rect 85947 54253 85955 57237
rect 82955 54245 85955 54253
rect 86145 57237 89145 57245
rect 86145 54253 86153 57237
rect 89137 54253 89145 57237
rect 86145 54245 89145 54253
rect 89335 57237 92335 57245
rect 89335 54253 89343 57237
rect 92327 54253 92335 57237
rect 89335 54245 92335 54253
rect 92525 57237 95525 57245
rect 92525 54253 92533 57237
rect 95517 54253 95525 57237
rect 92525 54245 95525 54253
rect 95715 57237 98715 57245
rect 95715 54253 95723 57237
rect 98707 54253 98715 57237
rect 95715 54245 98715 54253
rect 98905 57237 101905 57245
rect 98905 54253 98913 57237
rect 101897 54253 101905 57237
rect 98905 54245 101905 54253
rect 102095 57237 105095 57245
rect 102095 54253 102103 57237
rect 105087 54253 105095 57237
rect 102095 54245 105095 54253
rect 105285 57237 108285 57245
rect 105285 54253 105293 57237
rect 108277 54253 108285 57237
rect 105285 54245 108285 54253
rect 108475 57237 111475 57245
rect 108475 54253 108483 57237
rect 111467 54253 111475 57237
rect 108475 54245 111475 54253
rect 111665 57237 114665 57245
rect 111665 54253 111673 57237
rect 114657 54253 114665 57237
rect 111665 54245 114665 54253
rect 114855 57237 117855 57245
rect 114855 54253 114863 57237
rect 117847 54253 117855 57237
rect 114855 54245 117855 54253
rect 118045 57237 121045 57245
rect 118045 54253 118053 57237
rect 121037 54253 121045 57237
rect 118045 54245 121045 54253
rect 121235 57237 124235 57245
rect 121235 54253 121243 57237
rect 124227 54253 124235 57237
rect 121235 54245 124235 54253
rect 124425 57237 127425 57245
rect 124425 54253 124433 57237
rect 127417 54253 127425 57237
rect 124425 54245 127425 54253
rect 127615 57237 130615 57245
rect 127615 54253 127623 57237
rect 130607 54253 130615 57237
rect 127615 54245 130615 54253
rect 130805 57237 133805 57245
rect 130805 54253 130813 57237
rect 133797 54253 133805 57237
rect 130805 54245 133805 54253
rect 133995 57237 136995 57245
rect 133995 54253 134003 57237
rect 136987 54253 136995 57237
rect 133995 54245 136995 54253
rect 15 54047 3015 54055
rect 15 51063 23 54047
rect 3007 51063 3015 54047
rect 15 51055 3015 51063
rect 3205 54047 6205 54055
rect 3205 51063 3213 54047
rect 6197 51063 6205 54047
rect 3205 51055 6205 51063
rect 6395 54047 9395 54055
rect 6395 51063 6403 54047
rect 9387 51063 9395 54047
rect 6395 51055 9395 51063
rect 9585 54047 12585 54055
rect 9585 51063 9593 54047
rect 12577 51063 12585 54047
rect 9585 51055 12585 51063
rect 12775 54047 15775 54055
rect 12775 51063 12783 54047
rect 15767 51063 15775 54047
rect 12775 51055 15775 51063
rect 15965 54047 18965 54055
rect 15965 51063 15973 54047
rect 18957 51063 18965 54047
rect 15965 51055 18965 51063
rect 19155 54047 22155 54055
rect 19155 51063 19163 54047
rect 22147 51063 22155 54047
rect 19155 51055 22155 51063
rect 22345 54047 25345 54055
rect 22345 51063 22353 54047
rect 25337 51063 25345 54047
rect 22345 51055 25345 51063
rect 25535 54047 28535 54055
rect 25535 51063 25543 54047
rect 28527 51063 28535 54047
rect 25535 51055 28535 51063
rect 28725 54047 31725 54055
rect 28725 51063 28733 54047
rect 31717 51063 31725 54047
rect 28725 51055 31725 51063
rect 31915 54047 34915 54055
rect 31915 51063 31923 54047
rect 34907 51063 34915 54047
rect 31915 51055 34915 51063
rect 35105 54047 38105 54055
rect 35105 51063 35113 54047
rect 38097 51063 38105 54047
rect 35105 51055 38105 51063
rect 38295 54047 41295 54055
rect 38295 51063 38303 54047
rect 41287 51063 41295 54047
rect 38295 51055 41295 51063
rect 41485 54047 44485 54055
rect 41485 51063 41493 54047
rect 44477 51063 44485 54047
rect 41485 51055 44485 51063
rect 44675 54047 47675 54055
rect 44675 51063 44683 54047
rect 47667 51063 47675 54047
rect 44675 51055 47675 51063
rect 47865 54047 50865 54055
rect 47865 51063 47873 54047
rect 50857 51063 50865 54047
rect 47865 51055 50865 51063
rect 51055 54047 54055 54055
rect 51055 51063 51063 54047
rect 54047 51063 54055 54047
rect 51055 51055 54055 51063
rect 54245 54047 57245 54055
rect 54245 51063 54253 54047
rect 57237 51063 57245 54047
rect 54245 51055 57245 51063
rect 57435 54047 60435 54055
rect 57435 51063 57443 54047
rect 60427 51063 60435 54047
rect 57435 51055 60435 51063
rect 60625 54047 63625 54055
rect 60625 51063 60633 54047
rect 63617 51063 63625 54047
rect 60625 51055 63625 51063
rect 63815 54047 66815 54055
rect 63815 51063 63823 54047
rect 66807 51063 66815 54047
rect 63815 51055 66815 51063
rect 67005 54047 70005 54055
rect 67005 51063 67013 54047
rect 69997 51063 70005 54047
rect 67005 51055 70005 51063
rect 70195 54047 73195 54055
rect 70195 51063 70203 54047
rect 73187 51063 73195 54047
rect 70195 51055 73195 51063
rect 73385 54047 76385 54055
rect 73385 51063 73393 54047
rect 76377 51063 76385 54047
rect 73385 51055 76385 51063
rect 76575 54047 79575 54055
rect 76575 51063 76583 54047
rect 79567 51063 79575 54047
rect 76575 51055 79575 51063
rect 79765 54047 82765 54055
rect 79765 51063 79773 54047
rect 82757 51063 82765 54047
rect 79765 51055 82765 51063
rect 82955 54047 85955 54055
rect 82955 51063 82963 54047
rect 85947 51063 85955 54047
rect 82955 51055 85955 51063
rect 86145 54047 89145 54055
rect 86145 51063 86153 54047
rect 89137 51063 89145 54047
rect 86145 51055 89145 51063
rect 89335 54047 92335 54055
rect 89335 51063 89343 54047
rect 92327 51063 92335 54047
rect 89335 51055 92335 51063
rect 92525 54047 95525 54055
rect 92525 51063 92533 54047
rect 95517 51063 95525 54047
rect 92525 51055 95525 51063
rect 95715 54047 98715 54055
rect 95715 51063 95723 54047
rect 98707 51063 98715 54047
rect 95715 51055 98715 51063
rect 98905 54047 101905 54055
rect 98905 51063 98913 54047
rect 101897 51063 101905 54047
rect 98905 51055 101905 51063
rect 102095 54047 105095 54055
rect 102095 51063 102103 54047
rect 105087 51063 105095 54047
rect 102095 51055 105095 51063
rect 105285 54047 108285 54055
rect 105285 51063 105293 54047
rect 108277 51063 108285 54047
rect 105285 51055 108285 51063
rect 108475 54047 111475 54055
rect 108475 51063 108483 54047
rect 111467 51063 111475 54047
rect 108475 51055 111475 51063
rect 111665 54047 114665 54055
rect 111665 51063 111673 54047
rect 114657 51063 114665 54047
rect 111665 51055 114665 51063
rect 114855 54047 117855 54055
rect 114855 51063 114863 54047
rect 117847 51063 117855 54047
rect 114855 51055 117855 51063
rect 118045 54047 121045 54055
rect 118045 51063 118053 54047
rect 121037 51063 121045 54047
rect 118045 51055 121045 51063
rect 121235 54047 124235 54055
rect 121235 51063 121243 54047
rect 124227 51063 124235 54047
rect 121235 51055 124235 51063
rect 124425 54047 127425 54055
rect 124425 51063 124433 54047
rect 127417 51063 127425 54047
rect 124425 51055 127425 51063
rect 127615 54047 130615 54055
rect 127615 51063 127623 54047
rect 130607 51063 130615 54047
rect 127615 51055 130615 51063
rect 130805 54047 133805 54055
rect 130805 51063 130813 54047
rect 133797 51063 133805 54047
rect 130805 51055 133805 51063
rect 133995 54047 136995 54055
rect 133995 51063 134003 54047
rect 136987 51063 136995 54047
rect 133995 51055 136995 51063
rect 15 50857 3015 50865
rect 15 47873 23 50857
rect 3007 47873 3015 50857
rect 15 47865 3015 47873
rect 3205 50857 6205 50865
rect 3205 47873 3213 50857
rect 6197 47873 6205 50857
rect 3205 47865 6205 47873
rect 6395 50857 9395 50865
rect 6395 47873 6403 50857
rect 9387 47873 9395 50857
rect 6395 47865 9395 47873
rect 9585 50857 12585 50865
rect 9585 47873 9593 50857
rect 12577 47873 12585 50857
rect 9585 47865 12585 47873
rect 12775 50857 15775 50865
rect 12775 47873 12783 50857
rect 15767 47873 15775 50857
rect 12775 47865 15775 47873
rect 15965 50857 18965 50865
rect 15965 47873 15973 50857
rect 18957 47873 18965 50857
rect 15965 47865 18965 47873
rect 19155 50857 22155 50865
rect 19155 47873 19163 50857
rect 22147 47873 22155 50857
rect 19155 47865 22155 47873
rect 22345 50857 25345 50865
rect 22345 47873 22353 50857
rect 25337 47873 25345 50857
rect 22345 47865 25345 47873
rect 25535 50857 28535 50865
rect 25535 47873 25543 50857
rect 28527 47873 28535 50857
rect 25535 47865 28535 47873
rect 28725 50857 31725 50865
rect 28725 47873 28733 50857
rect 31717 47873 31725 50857
rect 28725 47865 31725 47873
rect 31915 50857 34915 50865
rect 31915 47873 31923 50857
rect 34907 47873 34915 50857
rect 31915 47865 34915 47873
rect 35105 50857 38105 50865
rect 35105 47873 35113 50857
rect 38097 47873 38105 50857
rect 35105 47865 38105 47873
rect 38295 50857 41295 50865
rect 38295 47873 38303 50857
rect 41287 47873 41295 50857
rect 38295 47865 41295 47873
rect 41485 50857 44485 50865
rect 41485 47873 41493 50857
rect 44477 47873 44485 50857
rect 41485 47865 44485 47873
rect 44675 50857 47675 50865
rect 44675 47873 44683 50857
rect 47667 47873 47675 50857
rect 44675 47865 47675 47873
rect 47865 50857 50865 50865
rect 47865 47873 47873 50857
rect 50857 47873 50865 50857
rect 47865 47865 50865 47873
rect 51055 50857 54055 50865
rect 51055 47873 51063 50857
rect 54047 47873 54055 50857
rect 51055 47865 54055 47873
rect 54245 50857 57245 50865
rect 54245 47873 54253 50857
rect 57237 47873 57245 50857
rect 54245 47865 57245 47873
rect 57435 50857 60435 50865
rect 57435 47873 57443 50857
rect 60427 47873 60435 50857
rect 57435 47865 60435 47873
rect 60625 50857 63625 50865
rect 60625 47873 60633 50857
rect 63617 47873 63625 50857
rect 60625 47865 63625 47873
rect 63815 50857 66815 50865
rect 63815 47873 63823 50857
rect 66807 47873 66815 50857
rect 63815 47865 66815 47873
rect 67005 50857 70005 50865
rect 67005 47873 67013 50857
rect 69997 47873 70005 50857
rect 67005 47865 70005 47873
rect 70195 50857 73195 50865
rect 70195 47873 70203 50857
rect 73187 47873 73195 50857
rect 70195 47865 73195 47873
rect 73385 50857 76385 50865
rect 73385 47873 73393 50857
rect 76377 47873 76385 50857
rect 73385 47865 76385 47873
rect 76575 50857 79575 50865
rect 76575 47873 76583 50857
rect 79567 47873 79575 50857
rect 76575 47865 79575 47873
rect 79765 50857 82765 50865
rect 79765 47873 79773 50857
rect 82757 47873 82765 50857
rect 79765 47865 82765 47873
rect 82955 50857 85955 50865
rect 82955 47873 82963 50857
rect 85947 47873 85955 50857
rect 82955 47865 85955 47873
rect 86145 50857 89145 50865
rect 86145 47873 86153 50857
rect 89137 47873 89145 50857
rect 86145 47865 89145 47873
rect 89335 50857 92335 50865
rect 89335 47873 89343 50857
rect 92327 47873 92335 50857
rect 89335 47865 92335 47873
rect 92525 50857 95525 50865
rect 92525 47873 92533 50857
rect 95517 47873 95525 50857
rect 92525 47865 95525 47873
rect 95715 50857 98715 50865
rect 95715 47873 95723 50857
rect 98707 47873 98715 50857
rect 95715 47865 98715 47873
rect 98905 50857 101905 50865
rect 98905 47873 98913 50857
rect 101897 47873 101905 50857
rect 98905 47865 101905 47873
rect 102095 50857 105095 50865
rect 102095 47873 102103 50857
rect 105087 47873 105095 50857
rect 102095 47865 105095 47873
rect 105285 50857 108285 50865
rect 105285 47873 105293 50857
rect 108277 47873 108285 50857
rect 105285 47865 108285 47873
rect 108475 50857 111475 50865
rect 108475 47873 108483 50857
rect 111467 47873 111475 50857
rect 108475 47865 111475 47873
rect 111665 50857 114665 50865
rect 111665 47873 111673 50857
rect 114657 47873 114665 50857
rect 111665 47865 114665 47873
rect 114855 50857 117855 50865
rect 114855 47873 114863 50857
rect 117847 47873 117855 50857
rect 114855 47865 117855 47873
rect 118045 50857 121045 50865
rect 118045 47873 118053 50857
rect 121037 47873 121045 50857
rect 118045 47865 121045 47873
rect 121235 50857 124235 50865
rect 121235 47873 121243 50857
rect 124227 47873 124235 50857
rect 121235 47865 124235 47873
rect 124425 50857 127425 50865
rect 124425 47873 124433 50857
rect 127417 47873 127425 50857
rect 124425 47865 127425 47873
rect 127615 50857 130615 50865
rect 127615 47873 127623 50857
rect 130607 47873 130615 50857
rect 127615 47865 130615 47873
rect 130805 50857 133805 50865
rect 130805 47873 130813 50857
rect 133797 47873 133805 50857
rect 130805 47865 133805 47873
rect 133995 50857 136995 50865
rect 133995 47873 134003 50857
rect 136987 47873 136995 50857
rect 133995 47865 136995 47873
rect 15 47667 3015 47675
rect 15 44683 23 47667
rect 3007 44683 3015 47667
rect 15 44675 3015 44683
rect 3205 47667 6205 47675
rect 3205 44683 3213 47667
rect 6197 44683 6205 47667
rect 3205 44675 6205 44683
rect 6395 47667 9395 47675
rect 6395 44683 6403 47667
rect 9387 44683 9395 47667
rect 6395 44675 9395 44683
rect 9585 47667 12585 47675
rect 9585 44683 9593 47667
rect 12577 44683 12585 47667
rect 9585 44675 12585 44683
rect 12775 47667 15775 47675
rect 12775 44683 12783 47667
rect 15767 44683 15775 47667
rect 12775 44675 15775 44683
rect 15965 47667 18965 47675
rect 15965 44683 15973 47667
rect 18957 44683 18965 47667
rect 15965 44675 18965 44683
rect 19155 47667 22155 47675
rect 19155 44683 19163 47667
rect 22147 44683 22155 47667
rect 19155 44675 22155 44683
rect 22345 47667 25345 47675
rect 22345 44683 22353 47667
rect 25337 44683 25345 47667
rect 22345 44675 25345 44683
rect 25535 47667 28535 47675
rect 25535 44683 25543 47667
rect 28527 44683 28535 47667
rect 25535 44675 28535 44683
rect 28725 47667 31725 47675
rect 28725 44683 28733 47667
rect 31717 44683 31725 47667
rect 28725 44675 31725 44683
rect 31915 47667 34915 47675
rect 31915 44683 31923 47667
rect 34907 44683 34915 47667
rect 31915 44675 34915 44683
rect 35105 47667 38105 47675
rect 35105 44683 35113 47667
rect 38097 44683 38105 47667
rect 35105 44675 38105 44683
rect 38295 47667 41295 47675
rect 38295 44683 38303 47667
rect 41287 44683 41295 47667
rect 38295 44675 41295 44683
rect 41485 47667 44485 47675
rect 41485 44683 41493 47667
rect 44477 44683 44485 47667
rect 41485 44675 44485 44683
rect 44675 47667 47675 47675
rect 44675 44683 44683 47667
rect 47667 44683 47675 47667
rect 44675 44675 47675 44683
rect 47865 47667 50865 47675
rect 47865 44683 47873 47667
rect 50857 44683 50865 47667
rect 47865 44675 50865 44683
rect 51055 47667 54055 47675
rect 51055 44683 51063 47667
rect 54047 44683 54055 47667
rect 51055 44675 54055 44683
rect 54245 47667 57245 47675
rect 54245 44683 54253 47667
rect 57237 44683 57245 47667
rect 54245 44675 57245 44683
rect 57435 47667 60435 47675
rect 57435 44683 57443 47667
rect 60427 44683 60435 47667
rect 57435 44675 60435 44683
rect 60625 47667 63625 47675
rect 60625 44683 60633 47667
rect 63617 44683 63625 47667
rect 60625 44675 63625 44683
rect 63815 47667 66815 47675
rect 63815 44683 63823 47667
rect 66807 44683 66815 47667
rect 63815 44675 66815 44683
rect 67005 47667 70005 47675
rect 67005 44683 67013 47667
rect 69997 44683 70005 47667
rect 67005 44675 70005 44683
rect 70195 47667 73195 47675
rect 70195 44683 70203 47667
rect 73187 44683 73195 47667
rect 70195 44675 73195 44683
rect 73385 47667 76385 47675
rect 73385 44683 73393 47667
rect 76377 44683 76385 47667
rect 73385 44675 76385 44683
rect 76575 47667 79575 47675
rect 76575 44683 76583 47667
rect 79567 44683 79575 47667
rect 76575 44675 79575 44683
rect 79765 47667 82765 47675
rect 79765 44683 79773 47667
rect 82757 44683 82765 47667
rect 79765 44675 82765 44683
rect 82955 47667 85955 47675
rect 82955 44683 82963 47667
rect 85947 44683 85955 47667
rect 82955 44675 85955 44683
rect 86145 47667 89145 47675
rect 86145 44683 86153 47667
rect 89137 44683 89145 47667
rect 86145 44675 89145 44683
rect 89335 47667 92335 47675
rect 89335 44683 89343 47667
rect 92327 44683 92335 47667
rect 89335 44675 92335 44683
rect 92525 47667 95525 47675
rect 92525 44683 92533 47667
rect 95517 44683 95525 47667
rect 92525 44675 95525 44683
rect 95715 47667 98715 47675
rect 95715 44683 95723 47667
rect 98707 44683 98715 47667
rect 95715 44675 98715 44683
rect 98905 47667 101905 47675
rect 98905 44683 98913 47667
rect 101897 44683 101905 47667
rect 98905 44675 101905 44683
rect 102095 47667 105095 47675
rect 102095 44683 102103 47667
rect 105087 44683 105095 47667
rect 102095 44675 105095 44683
rect 105285 47667 108285 47675
rect 105285 44683 105293 47667
rect 108277 44683 108285 47667
rect 105285 44675 108285 44683
rect 108475 47667 111475 47675
rect 108475 44683 108483 47667
rect 111467 44683 111475 47667
rect 108475 44675 111475 44683
rect 111665 47667 114665 47675
rect 111665 44683 111673 47667
rect 114657 44683 114665 47667
rect 111665 44675 114665 44683
rect 114855 47667 117855 47675
rect 114855 44683 114863 47667
rect 117847 44683 117855 47667
rect 114855 44675 117855 44683
rect 118045 47667 121045 47675
rect 118045 44683 118053 47667
rect 121037 44683 121045 47667
rect 118045 44675 121045 44683
rect 121235 47667 124235 47675
rect 121235 44683 121243 47667
rect 124227 44683 124235 47667
rect 121235 44675 124235 44683
rect 124425 47667 127425 47675
rect 124425 44683 124433 47667
rect 127417 44683 127425 47667
rect 124425 44675 127425 44683
rect 127615 47667 130615 47675
rect 127615 44683 127623 47667
rect 130607 44683 130615 47667
rect 127615 44675 130615 44683
rect 130805 47667 133805 47675
rect 130805 44683 130813 47667
rect 133797 44683 133805 47667
rect 130805 44675 133805 44683
rect 133995 47667 136995 47675
rect 133995 44683 134003 47667
rect 136987 44683 136995 47667
rect 133995 44675 136995 44683
rect 15 44477 3015 44485
rect 15 41493 23 44477
rect 3007 41493 3015 44477
rect 15 41485 3015 41493
rect 3205 44477 6205 44485
rect 3205 41493 3213 44477
rect 6197 41493 6205 44477
rect 3205 41485 6205 41493
rect 6395 44477 9395 44485
rect 6395 41493 6403 44477
rect 9387 41493 9395 44477
rect 6395 41485 9395 41493
rect 9585 44477 12585 44485
rect 9585 41493 9593 44477
rect 12577 41493 12585 44477
rect 9585 41485 12585 41493
rect 12775 44477 15775 44485
rect 12775 41493 12783 44477
rect 15767 41493 15775 44477
rect 12775 41485 15775 41493
rect 15965 44477 18965 44485
rect 15965 41493 15973 44477
rect 18957 41493 18965 44477
rect 15965 41485 18965 41493
rect 19155 44477 22155 44485
rect 19155 41493 19163 44477
rect 22147 41493 22155 44477
rect 19155 41485 22155 41493
rect 22345 44477 25345 44485
rect 22345 41493 22353 44477
rect 25337 41493 25345 44477
rect 22345 41485 25345 41493
rect 25535 44477 28535 44485
rect 25535 41493 25543 44477
rect 28527 41493 28535 44477
rect 25535 41485 28535 41493
rect 28725 44477 31725 44485
rect 28725 41493 28733 44477
rect 31717 41493 31725 44477
rect 28725 41485 31725 41493
rect 31915 44477 34915 44485
rect 31915 41493 31923 44477
rect 34907 41493 34915 44477
rect 31915 41485 34915 41493
rect 35105 44477 38105 44485
rect 35105 41493 35113 44477
rect 38097 41493 38105 44477
rect 35105 41485 38105 41493
rect 38295 44477 41295 44485
rect 38295 41493 38303 44477
rect 41287 41493 41295 44477
rect 38295 41485 41295 41493
rect 41485 44477 44485 44485
rect 41485 41493 41493 44477
rect 44477 41493 44485 44477
rect 41485 41485 44485 41493
rect 44675 44477 47675 44485
rect 44675 41493 44683 44477
rect 47667 41493 47675 44477
rect 44675 41485 47675 41493
rect 47865 44477 50865 44485
rect 47865 41493 47873 44477
rect 50857 41493 50865 44477
rect 47865 41485 50865 41493
rect 51055 44477 54055 44485
rect 51055 41493 51063 44477
rect 54047 41493 54055 44477
rect 51055 41485 54055 41493
rect 54245 44477 57245 44485
rect 54245 41493 54253 44477
rect 57237 41493 57245 44477
rect 54245 41485 57245 41493
rect 57435 44477 60435 44485
rect 57435 41493 57443 44477
rect 60427 41493 60435 44477
rect 57435 41485 60435 41493
rect 60625 44477 63625 44485
rect 60625 41493 60633 44477
rect 63617 41493 63625 44477
rect 60625 41485 63625 41493
rect 63815 44477 66815 44485
rect 63815 41493 63823 44477
rect 66807 41493 66815 44477
rect 63815 41485 66815 41493
rect 67005 44477 70005 44485
rect 67005 41493 67013 44477
rect 69997 41493 70005 44477
rect 67005 41485 70005 41493
rect 70195 44477 73195 44485
rect 70195 41493 70203 44477
rect 73187 41493 73195 44477
rect 70195 41485 73195 41493
rect 73385 44477 76385 44485
rect 73385 41493 73393 44477
rect 76377 41493 76385 44477
rect 73385 41485 76385 41493
rect 76575 44477 79575 44485
rect 76575 41493 76583 44477
rect 79567 41493 79575 44477
rect 76575 41485 79575 41493
rect 79765 44477 82765 44485
rect 79765 41493 79773 44477
rect 82757 41493 82765 44477
rect 79765 41485 82765 41493
rect 82955 44477 85955 44485
rect 82955 41493 82963 44477
rect 85947 41493 85955 44477
rect 82955 41485 85955 41493
rect 86145 44477 89145 44485
rect 86145 41493 86153 44477
rect 89137 41493 89145 44477
rect 86145 41485 89145 41493
rect 89335 44477 92335 44485
rect 89335 41493 89343 44477
rect 92327 41493 92335 44477
rect 89335 41485 92335 41493
rect 92525 44477 95525 44485
rect 92525 41493 92533 44477
rect 95517 41493 95525 44477
rect 92525 41485 95525 41493
rect 95715 44477 98715 44485
rect 95715 41493 95723 44477
rect 98707 41493 98715 44477
rect 95715 41485 98715 41493
rect 98905 44477 101905 44485
rect 98905 41493 98913 44477
rect 101897 41493 101905 44477
rect 98905 41485 101905 41493
rect 102095 44477 105095 44485
rect 102095 41493 102103 44477
rect 105087 41493 105095 44477
rect 102095 41485 105095 41493
rect 105285 44477 108285 44485
rect 105285 41493 105293 44477
rect 108277 41493 108285 44477
rect 105285 41485 108285 41493
rect 108475 44477 111475 44485
rect 108475 41493 108483 44477
rect 111467 41493 111475 44477
rect 108475 41485 111475 41493
rect 111665 44477 114665 44485
rect 111665 41493 111673 44477
rect 114657 41493 114665 44477
rect 111665 41485 114665 41493
rect 114855 44477 117855 44485
rect 114855 41493 114863 44477
rect 117847 41493 117855 44477
rect 114855 41485 117855 41493
rect 118045 44477 121045 44485
rect 118045 41493 118053 44477
rect 121037 41493 121045 44477
rect 118045 41485 121045 41493
rect 121235 44477 124235 44485
rect 121235 41493 121243 44477
rect 124227 41493 124235 44477
rect 121235 41485 124235 41493
rect 124425 44477 127425 44485
rect 124425 41493 124433 44477
rect 127417 41493 127425 44477
rect 124425 41485 127425 41493
rect 127615 44477 130615 44485
rect 127615 41493 127623 44477
rect 130607 41493 130615 44477
rect 127615 41485 130615 41493
rect 130805 44477 133805 44485
rect 130805 41493 130813 44477
rect 133797 41493 133805 44477
rect 130805 41485 133805 41493
rect 133995 44477 136995 44485
rect 133995 41493 134003 44477
rect 136987 41493 136995 44477
rect 133995 41485 136995 41493
rect 15 41287 3015 41295
rect 15 38303 23 41287
rect 3007 38303 3015 41287
rect 15 38295 3015 38303
rect 3205 41287 6205 41295
rect 3205 38303 3213 41287
rect 6197 38303 6205 41287
rect 3205 38295 6205 38303
rect 6395 41287 9395 41295
rect 6395 38303 6403 41287
rect 9387 38303 9395 41287
rect 6395 38295 9395 38303
rect 9585 41287 12585 41295
rect 9585 38303 9593 41287
rect 12577 38303 12585 41287
rect 9585 38295 12585 38303
rect 12775 41287 15775 41295
rect 12775 38303 12783 41287
rect 15767 38303 15775 41287
rect 12775 38295 15775 38303
rect 15965 41287 18965 41295
rect 15965 38303 15973 41287
rect 18957 38303 18965 41287
rect 15965 38295 18965 38303
rect 19155 41287 22155 41295
rect 19155 38303 19163 41287
rect 22147 38303 22155 41287
rect 19155 38295 22155 38303
rect 22345 41287 25345 41295
rect 22345 38303 22353 41287
rect 25337 38303 25345 41287
rect 22345 38295 25345 38303
rect 25535 41287 28535 41295
rect 25535 38303 25543 41287
rect 28527 38303 28535 41287
rect 25535 38295 28535 38303
rect 28725 41287 31725 41295
rect 28725 38303 28733 41287
rect 31717 38303 31725 41287
rect 28725 38295 31725 38303
rect 31915 41287 34915 41295
rect 31915 38303 31923 41287
rect 34907 38303 34915 41287
rect 31915 38295 34915 38303
rect 35105 41287 38105 41295
rect 35105 38303 35113 41287
rect 38097 38303 38105 41287
rect 35105 38295 38105 38303
rect 38295 41287 41295 41295
rect 38295 38303 38303 41287
rect 41287 38303 41295 41287
rect 38295 38295 41295 38303
rect 41485 41287 44485 41295
rect 41485 38303 41493 41287
rect 44477 38303 44485 41287
rect 41485 38295 44485 38303
rect 44675 41287 47675 41295
rect 44675 38303 44683 41287
rect 47667 38303 47675 41287
rect 44675 38295 47675 38303
rect 47865 41287 50865 41295
rect 47865 38303 47873 41287
rect 50857 38303 50865 41287
rect 47865 38295 50865 38303
rect 51055 41287 54055 41295
rect 51055 38303 51063 41287
rect 54047 38303 54055 41287
rect 51055 38295 54055 38303
rect 54245 41287 57245 41295
rect 54245 38303 54253 41287
rect 57237 38303 57245 41287
rect 54245 38295 57245 38303
rect 57435 41287 60435 41295
rect 57435 38303 57443 41287
rect 60427 38303 60435 41287
rect 57435 38295 60435 38303
rect 60625 41287 63625 41295
rect 60625 38303 60633 41287
rect 63617 38303 63625 41287
rect 60625 38295 63625 38303
rect 63815 41287 66815 41295
rect 63815 38303 63823 41287
rect 66807 38303 66815 41287
rect 63815 38295 66815 38303
rect 67005 41287 70005 41295
rect 67005 38303 67013 41287
rect 69997 38303 70005 41287
rect 67005 38295 70005 38303
rect 70195 41287 73195 41295
rect 70195 38303 70203 41287
rect 73187 38303 73195 41287
rect 70195 38295 73195 38303
rect 73385 41287 76385 41295
rect 73385 38303 73393 41287
rect 76377 38303 76385 41287
rect 73385 38295 76385 38303
rect 76575 41287 79575 41295
rect 76575 38303 76583 41287
rect 79567 38303 79575 41287
rect 76575 38295 79575 38303
rect 79765 41287 82765 41295
rect 79765 38303 79773 41287
rect 82757 38303 82765 41287
rect 79765 38295 82765 38303
rect 82955 41287 85955 41295
rect 82955 38303 82963 41287
rect 85947 38303 85955 41287
rect 82955 38295 85955 38303
rect 86145 41287 89145 41295
rect 86145 38303 86153 41287
rect 89137 38303 89145 41287
rect 86145 38295 89145 38303
rect 89335 41287 92335 41295
rect 89335 38303 89343 41287
rect 92327 38303 92335 41287
rect 89335 38295 92335 38303
rect 92525 41287 95525 41295
rect 92525 38303 92533 41287
rect 95517 38303 95525 41287
rect 92525 38295 95525 38303
rect 95715 41287 98715 41295
rect 95715 38303 95723 41287
rect 98707 38303 98715 41287
rect 95715 38295 98715 38303
rect 98905 41287 101905 41295
rect 98905 38303 98913 41287
rect 101897 38303 101905 41287
rect 98905 38295 101905 38303
rect 102095 41287 105095 41295
rect 102095 38303 102103 41287
rect 105087 38303 105095 41287
rect 102095 38295 105095 38303
rect 105285 41287 108285 41295
rect 105285 38303 105293 41287
rect 108277 38303 108285 41287
rect 105285 38295 108285 38303
rect 108475 41287 111475 41295
rect 108475 38303 108483 41287
rect 111467 38303 111475 41287
rect 108475 38295 111475 38303
rect 111665 41287 114665 41295
rect 111665 38303 111673 41287
rect 114657 38303 114665 41287
rect 111665 38295 114665 38303
rect 114855 41287 117855 41295
rect 114855 38303 114863 41287
rect 117847 38303 117855 41287
rect 114855 38295 117855 38303
rect 118045 41287 121045 41295
rect 118045 38303 118053 41287
rect 121037 38303 121045 41287
rect 118045 38295 121045 38303
rect 121235 41287 124235 41295
rect 121235 38303 121243 41287
rect 124227 38303 124235 41287
rect 121235 38295 124235 38303
rect 124425 41287 127425 41295
rect 124425 38303 124433 41287
rect 127417 38303 127425 41287
rect 124425 38295 127425 38303
rect 127615 41287 130615 41295
rect 127615 38303 127623 41287
rect 130607 38303 130615 41287
rect 127615 38295 130615 38303
rect 130805 41287 133805 41295
rect 130805 38303 130813 41287
rect 133797 38303 133805 41287
rect 130805 38295 133805 38303
rect 133995 41287 136995 41295
rect 133995 38303 134003 41287
rect 136987 38303 136995 41287
rect 133995 38295 136995 38303
rect 15 38097 3015 38105
rect 15 35113 23 38097
rect 3007 35113 3015 38097
rect 15 35105 3015 35113
rect 3205 38097 6205 38105
rect 3205 35113 3213 38097
rect 6197 35113 6205 38097
rect 3205 35105 6205 35113
rect 6395 38097 9395 38105
rect 6395 35113 6403 38097
rect 9387 35113 9395 38097
rect 6395 35105 9395 35113
rect 9585 38097 12585 38105
rect 9585 35113 9593 38097
rect 12577 35113 12585 38097
rect 9585 35105 12585 35113
rect 12775 38097 15775 38105
rect 12775 35113 12783 38097
rect 15767 35113 15775 38097
rect 12775 35105 15775 35113
rect 15965 38097 18965 38105
rect 15965 35113 15973 38097
rect 18957 35113 18965 38097
rect 15965 35105 18965 35113
rect 19155 38097 22155 38105
rect 19155 35113 19163 38097
rect 22147 35113 22155 38097
rect 19155 35105 22155 35113
rect 22345 38097 25345 38105
rect 22345 35113 22353 38097
rect 25337 35113 25345 38097
rect 22345 35105 25345 35113
rect 25535 38097 28535 38105
rect 25535 35113 25543 38097
rect 28527 35113 28535 38097
rect 25535 35105 28535 35113
rect 28725 38097 31725 38105
rect 28725 35113 28733 38097
rect 31717 35113 31725 38097
rect 28725 35105 31725 35113
rect 31915 38097 34915 38105
rect 31915 35113 31923 38097
rect 34907 35113 34915 38097
rect 31915 35105 34915 35113
rect 35105 38097 38105 38105
rect 35105 35113 35113 38097
rect 38097 35113 38105 38097
rect 35105 35105 38105 35113
rect 38295 38097 41295 38105
rect 38295 35113 38303 38097
rect 41287 35113 41295 38097
rect 38295 35105 41295 35113
rect 41485 38097 44485 38105
rect 41485 35113 41493 38097
rect 44477 35113 44485 38097
rect 41485 35105 44485 35113
rect 44675 38097 47675 38105
rect 44675 35113 44683 38097
rect 47667 35113 47675 38097
rect 44675 35105 47675 35113
rect 47865 38097 50865 38105
rect 47865 35113 47873 38097
rect 50857 35113 50865 38097
rect 47865 35105 50865 35113
rect 51055 38097 54055 38105
rect 51055 35113 51063 38097
rect 54047 35113 54055 38097
rect 51055 35105 54055 35113
rect 54245 38097 57245 38105
rect 54245 35113 54253 38097
rect 57237 35113 57245 38097
rect 54245 35105 57245 35113
rect 57435 38097 60435 38105
rect 57435 35113 57443 38097
rect 60427 35113 60435 38097
rect 57435 35105 60435 35113
rect 60625 38097 63625 38105
rect 60625 35113 60633 38097
rect 63617 35113 63625 38097
rect 60625 35105 63625 35113
rect 63815 38097 66815 38105
rect 63815 35113 63823 38097
rect 66807 35113 66815 38097
rect 63815 35105 66815 35113
rect 67005 38097 70005 38105
rect 67005 35113 67013 38097
rect 69997 35113 70005 38097
rect 67005 35105 70005 35113
rect 70195 38097 73195 38105
rect 70195 35113 70203 38097
rect 73187 35113 73195 38097
rect 70195 35105 73195 35113
rect 73385 38097 76385 38105
rect 73385 35113 73393 38097
rect 76377 35113 76385 38097
rect 73385 35105 76385 35113
rect 76575 38097 79575 38105
rect 76575 35113 76583 38097
rect 79567 35113 79575 38097
rect 76575 35105 79575 35113
rect 79765 38097 82765 38105
rect 79765 35113 79773 38097
rect 82757 35113 82765 38097
rect 79765 35105 82765 35113
rect 82955 38097 85955 38105
rect 82955 35113 82963 38097
rect 85947 35113 85955 38097
rect 82955 35105 85955 35113
rect 86145 38097 89145 38105
rect 86145 35113 86153 38097
rect 89137 35113 89145 38097
rect 86145 35105 89145 35113
rect 89335 38097 92335 38105
rect 89335 35113 89343 38097
rect 92327 35113 92335 38097
rect 89335 35105 92335 35113
rect 92525 38097 95525 38105
rect 92525 35113 92533 38097
rect 95517 35113 95525 38097
rect 92525 35105 95525 35113
rect 95715 38097 98715 38105
rect 95715 35113 95723 38097
rect 98707 35113 98715 38097
rect 95715 35105 98715 35113
rect 98905 38097 101905 38105
rect 98905 35113 98913 38097
rect 101897 35113 101905 38097
rect 98905 35105 101905 35113
rect 102095 38097 105095 38105
rect 102095 35113 102103 38097
rect 105087 35113 105095 38097
rect 102095 35105 105095 35113
rect 105285 38097 108285 38105
rect 105285 35113 105293 38097
rect 108277 35113 108285 38097
rect 105285 35105 108285 35113
rect 108475 38097 111475 38105
rect 108475 35113 108483 38097
rect 111467 35113 111475 38097
rect 108475 35105 111475 35113
rect 111665 38097 114665 38105
rect 111665 35113 111673 38097
rect 114657 35113 114665 38097
rect 111665 35105 114665 35113
rect 114855 38097 117855 38105
rect 114855 35113 114863 38097
rect 117847 35113 117855 38097
rect 114855 35105 117855 35113
rect 118045 38097 121045 38105
rect 118045 35113 118053 38097
rect 121037 35113 121045 38097
rect 118045 35105 121045 35113
rect 121235 38097 124235 38105
rect 121235 35113 121243 38097
rect 124227 35113 124235 38097
rect 121235 35105 124235 35113
rect 124425 38097 127425 38105
rect 124425 35113 124433 38097
rect 127417 35113 127425 38097
rect 124425 35105 127425 35113
rect 127615 38097 130615 38105
rect 127615 35113 127623 38097
rect 130607 35113 130615 38097
rect 127615 35105 130615 35113
rect 130805 38097 133805 38105
rect 130805 35113 130813 38097
rect 133797 35113 133805 38097
rect 130805 35105 133805 35113
rect 133995 38097 136995 38105
rect 133995 35113 134003 38097
rect 136987 35113 136995 38097
rect 133995 35105 136995 35113
rect 15 34907 3015 34915
rect 15 31923 23 34907
rect 3007 31923 3015 34907
rect 15 31915 3015 31923
rect 3205 34907 6205 34915
rect 3205 31923 3213 34907
rect 6197 31923 6205 34907
rect 3205 31915 6205 31923
rect 6395 34907 9395 34915
rect 6395 31923 6403 34907
rect 9387 31923 9395 34907
rect 6395 31915 9395 31923
rect 9585 34907 12585 34915
rect 9585 31923 9593 34907
rect 12577 31923 12585 34907
rect 9585 31915 12585 31923
rect 12775 34907 15775 34915
rect 12775 31923 12783 34907
rect 15767 31923 15775 34907
rect 12775 31915 15775 31923
rect 15965 34907 18965 34915
rect 15965 31923 15973 34907
rect 18957 31923 18965 34907
rect 15965 31915 18965 31923
rect 19155 34907 22155 34915
rect 19155 31923 19163 34907
rect 22147 31923 22155 34907
rect 19155 31915 22155 31923
rect 22345 34907 25345 34915
rect 22345 31923 22353 34907
rect 25337 31923 25345 34907
rect 22345 31915 25345 31923
rect 25535 34907 28535 34915
rect 25535 31923 25543 34907
rect 28527 31923 28535 34907
rect 25535 31915 28535 31923
rect 28725 34907 31725 34915
rect 28725 31923 28733 34907
rect 31717 31923 31725 34907
rect 28725 31915 31725 31923
rect 31915 34907 34915 34915
rect 31915 31923 31923 34907
rect 34907 31923 34915 34907
rect 31915 31915 34915 31923
rect 35105 34907 38105 34915
rect 35105 31923 35113 34907
rect 38097 31923 38105 34907
rect 35105 31915 38105 31923
rect 38295 34907 41295 34915
rect 38295 31923 38303 34907
rect 41287 31923 41295 34907
rect 38295 31915 41295 31923
rect 41485 34907 44485 34915
rect 41485 31923 41493 34907
rect 44477 31923 44485 34907
rect 41485 31915 44485 31923
rect 44675 34907 47675 34915
rect 44675 31923 44683 34907
rect 47667 31923 47675 34907
rect 44675 31915 47675 31923
rect 47865 34907 50865 34915
rect 47865 31923 47873 34907
rect 50857 31923 50865 34907
rect 47865 31915 50865 31923
rect 51055 34907 54055 34915
rect 51055 31923 51063 34907
rect 54047 31923 54055 34907
rect 51055 31915 54055 31923
rect 54245 34907 57245 34915
rect 54245 31923 54253 34907
rect 57237 31923 57245 34907
rect 54245 31915 57245 31923
rect 57435 34907 60435 34915
rect 57435 31923 57443 34907
rect 60427 31923 60435 34907
rect 57435 31915 60435 31923
rect 60625 34907 63625 34915
rect 60625 31923 60633 34907
rect 63617 31923 63625 34907
rect 60625 31915 63625 31923
rect 63815 34907 66815 34915
rect 63815 31923 63823 34907
rect 66807 31923 66815 34907
rect 63815 31915 66815 31923
rect 67005 34907 70005 34915
rect 67005 31923 67013 34907
rect 69997 31923 70005 34907
rect 67005 31915 70005 31923
rect 70195 34907 73195 34915
rect 70195 31923 70203 34907
rect 73187 31923 73195 34907
rect 70195 31915 73195 31923
rect 73385 34907 76385 34915
rect 73385 31923 73393 34907
rect 76377 31923 76385 34907
rect 73385 31915 76385 31923
rect 76575 34907 79575 34915
rect 76575 31923 76583 34907
rect 79567 31923 79575 34907
rect 76575 31915 79575 31923
rect 79765 34907 82765 34915
rect 79765 31923 79773 34907
rect 82757 31923 82765 34907
rect 79765 31915 82765 31923
rect 82955 34907 85955 34915
rect 82955 31923 82963 34907
rect 85947 31923 85955 34907
rect 82955 31915 85955 31923
rect 86145 34907 89145 34915
rect 86145 31923 86153 34907
rect 89137 31923 89145 34907
rect 86145 31915 89145 31923
rect 89335 34907 92335 34915
rect 89335 31923 89343 34907
rect 92327 31923 92335 34907
rect 89335 31915 92335 31923
rect 92525 34907 95525 34915
rect 92525 31923 92533 34907
rect 95517 31923 95525 34907
rect 92525 31915 95525 31923
rect 95715 34907 98715 34915
rect 95715 31923 95723 34907
rect 98707 31923 98715 34907
rect 95715 31915 98715 31923
rect 98905 34907 101905 34915
rect 98905 31923 98913 34907
rect 101897 31923 101905 34907
rect 98905 31915 101905 31923
rect 102095 34907 105095 34915
rect 102095 31923 102103 34907
rect 105087 31923 105095 34907
rect 102095 31915 105095 31923
rect 105285 34907 108285 34915
rect 105285 31923 105293 34907
rect 108277 31923 108285 34907
rect 105285 31915 108285 31923
rect 108475 34907 111475 34915
rect 108475 31923 108483 34907
rect 111467 31923 111475 34907
rect 108475 31915 111475 31923
rect 111665 34907 114665 34915
rect 111665 31923 111673 34907
rect 114657 31923 114665 34907
rect 111665 31915 114665 31923
rect 114855 34907 117855 34915
rect 114855 31923 114863 34907
rect 117847 31923 117855 34907
rect 114855 31915 117855 31923
rect 118045 34907 121045 34915
rect 118045 31923 118053 34907
rect 121037 31923 121045 34907
rect 118045 31915 121045 31923
rect 121235 34907 124235 34915
rect 121235 31923 121243 34907
rect 124227 31923 124235 34907
rect 121235 31915 124235 31923
rect 124425 34907 127425 34915
rect 124425 31923 124433 34907
rect 127417 31923 127425 34907
rect 124425 31915 127425 31923
rect 127615 34907 130615 34915
rect 127615 31923 127623 34907
rect 130607 31923 130615 34907
rect 127615 31915 130615 31923
rect 130805 34907 133805 34915
rect 130805 31923 130813 34907
rect 133797 31923 133805 34907
rect 130805 31915 133805 31923
rect 133995 34907 136995 34915
rect 133995 31923 134003 34907
rect 136987 31923 136995 34907
rect 133995 31915 136995 31923
rect 15 31717 3015 31725
rect 15 28733 23 31717
rect 3007 28733 3015 31717
rect 15 28725 3015 28733
rect 3205 31717 6205 31725
rect 3205 28733 3213 31717
rect 6197 28733 6205 31717
rect 3205 28725 6205 28733
rect 6395 31717 9395 31725
rect 6395 28733 6403 31717
rect 9387 28733 9395 31717
rect 6395 28725 9395 28733
rect 9585 31717 12585 31725
rect 9585 28733 9593 31717
rect 12577 28733 12585 31717
rect 9585 28725 12585 28733
rect 12775 31717 15775 31725
rect 12775 28733 12783 31717
rect 15767 28733 15775 31717
rect 12775 28725 15775 28733
rect 15965 31717 18965 31725
rect 15965 28733 15973 31717
rect 18957 28733 18965 31717
rect 15965 28725 18965 28733
rect 19155 31717 22155 31725
rect 19155 28733 19163 31717
rect 22147 28733 22155 31717
rect 19155 28725 22155 28733
rect 22345 31717 25345 31725
rect 22345 28733 22353 31717
rect 25337 28733 25345 31717
rect 22345 28725 25345 28733
rect 25535 31717 28535 31725
rect 25535 28733 25543 31717
rect 28527 28733 28535 31717
rect 25535 28725 28535 28733
rect 28725 31717 31725 31725
rect 28725 28733 28733 31717
rect 31717 28733 31725 31717
rect 28725 28725 31725 28733
rect 31915 31717 34915 31725
rect 31915 28733 31923 31717
rect 34907 28733 34915 31717
rect 31915 28725 34915 28733
rect 35105 31717 38105 31725
rect 35105 28733 35113 31717
rect 38097 28733 38105 31717
rect 35105 28725 38105 28733
rect 38295 31717 41295 31725
rect 38295 28733 38303 31717
rect 41287 28733 41295 31717
rect 38295 28725 41295 28733
rect 41485 31717 44485 31725
rect 41485 28733 41493 31717
rect 44477 28733 44485 31717
rect 41485 28725 44485 28733
rect 44675 31717 47675 31725
rect 44675 28733 44683 31717
rect 47667 28733 47675 31717
rect 44675 28725 47675 28733
rect 47865 31717 50865 31725
rect 47865 28733 47873 31717
rect 50857 28733 50865 31717
rect 47865 28725 50865 28733
rect 51055 31717 54055 31725
rect 51055 28733 51063 31717
rect 54047 28733 54055 31717
rect 51055 28725 54055 28733
rect 54245 31717 57245 31725
rect 54245 28733 54253 31717
rect 57237 28733 57245 31717
rect 54245 28725 57245 28733
rect 57435 31717 60435 31725
rect 57435 28733 57443 31717
rect 60427 28733 60435 31717
rect 57435 28725 60435 28733
rect 60625 31717 63625 31725
rect 60625 28733 60633 31717
rect 63617 28733 63625 31717
rect 60625 28725 63625 28733
rect 63815 31717 66815 31725
rect 63815 28733 63823 31717
rect 66807 28733 66815 31717
rect 63815 28725 66815 28733
rect 67005 31717 70005 31725
rect 67005 28733 67013 31717
rect 69997 28733 70005 31717
rect 67005 28725 70005 28733
rect 70195 31717 73195 31725
rect 70195 28733 70203 31717
rect 73187 28733 73195 31717
rect 70195 28725 73195 28733
rect 73385 31717 76385 31725
rect 73385 28733 73393 31717
rect 76377 28733 76385 31717
rect 73385 28725 76385 28733
rect 76575 31717 79575 31725
rect 76575 28733 76583 31717
rect 79567 28733 79575 31717
rect 76575 28725 79575 28733
rect 79765 31717 82765 31725
rect 79765 28733 79773 31717
rect 82757 28733 82765 31717
rect 79765 28725 82765 28733
rect 82955 31717 85955 31725
rect 82955 28733 82963 31717
rect 85947 28733 85955 31717
rect 82955 28725 85955 28733
rect 86145 31717 89145 31725
rect 86145 28733 86153 31717
rect 89137 28733 89145 31717
rect 86145 28725 89145 28733
rect 89335 31717 92335 31725
rect 89335 28733 89343 31717
rect 92327 28733 92335 31717
rect 89335 28725 92335 28733
rect 92525 31717 95525 31725
rect 92525 28733 92533 31717
rect 95517 28733 95525 31717
rect 92525 28725 95525 28733
rect 95715 31717 98715 31725
rect 95715 28733 95723 31717
rect 98707 28733 98715 31717
rect 95715 28725 98715 28733
rect 98905 31717 101905 31725
rect 98905 28733 98913 31717
rect 101897 28733 101905 31717
rect 98905 28725 101905 28733
rect 102095 31717 105095 31725
rect 102095 28733 102103 31717
rect 105087 28733 105095 31717
rect 102095 28725 105095 28733
rect 105285 31717 108285 31725
rect 105285 28733 105293 31717
rect 108277 28733 108285 31717
rect 105285 28725 108285 28733
rect 108475 31717 111475 31725
rect 108475 28733 108483 31717
rect 111467 28733 111475 31717
rect 108475 28725 111475 28733
rect 111665 31717 114665 31725
rect 111665 28733 111673 31717
rect 114657 28733 114665 31717
rect 111665 28725 114665 28733
rect 114855 31717 117855 31725
rect 114855 28733 114863 31717
rect 117847 28733 117855 31717
rect 114855 28725 117855 28733
rect 118045 31717 121045 31725
rect 118045 28733 118053 31717
rect 121037 28733 121045 31717
rect 118045 28725 121045 28733
rect 121235 31717 124235 31725
rect 121235 28733 121243 31717
rect 124227 28733 124235 31717
rect 121235 28725 124235 28733
rect 124425 31717 127425 31725
rect 124425 28733 124433 31717
rect 127417 28733 127425 31717
rect 124425 28725 127425 28733
rect 127615 31717 130615 31725
rect 127615 28733 127623 31717
rect 130607 28733 130615 31717
rect 127615 28725 130615 28733
rect 130805 31717 133805 31725
rect 130805 28733 130813 31717
rect 133797 28733 133805 31717
rect 130805 28725 133805 28733
rect 133995 31717 136995 31725
rect 133995 28733 134003 31717
rect 136987 28733 136995 31717
rect 133995 28725 136995 28733
rect 15 28527 3015 28535
rect 15 25543 23 28527
rect 3007 25543 3015 28527
rect 15 25535 3015 25543
rect 3205 28527 6205 28535
rect 3205 25543 3213 28527
rect 6197 25543 6205 28527
rect 3205 25535 6205 25543
rect 6395 28527 9395 28535
rect 6395 25543 6403 28527
rect 9387 25543 9395 28527
rect 6395 25535 9395 25543
rect 9585 28527 12585 28535
rect 9585 25543 9593 28527
rect 12577 25543 12585 28527
rect 9585 25535 12585 25543
rect 12775 28527 15775 28535
rect 12775 25543 12783 28527
rect 15767 25543 15775 28527
rect 12775 25535 15775 25543
rect 15965 28527 18965 28535
rect 15965 25543 15973 28527
rect 18957 25543 18965 28527
rect 15965 25535 18965 25543
rect 19155 28527 22155 28535
rect 19155 25543 19163 28527
rect 22147 25543 22155 28527
rect 19155 25535 22155 25543
rect 22345 28527 25345 28535
rect 22345 25543 22353 28527
rect 25337 25543 25345 28527
rect 22345 25535 25345 25543
rect 25535 28527 28535 28535
rect 25535 25543 25543 28527
rect 28527 25543 28535 28527
rect 25535 25535 28535 25543
rect 28725 28527 31725 28535
rect 28725 25543 28733 28527
rect 31717 25543 31725 28527
rect 28725 25535 31725 25543
rect 31915 28527 34915 28535
rect 31915 25543 31923 28527
rect 34907 25543 34915 28527
rect 31915 25535 34915 25543
rect 35105 28527 38105 28535
rect 35105 25543 35113 28527
rect 38097 25543 38105 28527
rect 35105 25535 38105 25543
rect 38295 28527 41295 28535
rect 38295 25543 38303 28527
rect 41287 25543 41295 28527
rect 38295 25535 41295 25543
rect 41485 28527 44485 28535
rect 41485 25543 41493 28527
rect 44477 25543 44485 28527
rect 41485 25535 44485 25543
rect 44675 28527 47675 28535
rect 44675 25543 44683 28527
rect 47667 25543 47675 28527
rect 44675 25535 47675 25543
rect 47865 28527 50865 28535
rect 47865 25543 47873 28527
rect 50857 25543 50865 28527
rect 47865 25535 50865 25543
rect 51055 28527 54055 28535
rect 51055 25543 51063 28527
rect 54047 25543 54055 28527
rect 51055 25535 54055 25543
rect 54245 28527 57245 28535
rect 54245 25543 54253 28527
rect 57237 25543 57245 28527
rect 54245 25535 57245 25543
rect 57435 28527 60435 28535
rect 57435 25543 57443 28527
rect 60427 25543 60435 28527
rect 57435 25535 60435 25543
rect 60625 28527 63625 28535
rect 60625 25543 60633 28527
rect 63617 25543 63625 28527
rect 60625 25535 63625 25543
rect 63815 28527 66815 28535
rect 63815 25543 63823 28527
rect 66807 25543 66815 28527
rect 63815 25535 66815 25543
rect 67005 28527 70005 28535
rect 67005 25543 67013 28527
rect 69997 25543 70005 28527
rect 67005 25535 70005 25543
rect 70195 28527 73195 28535
rect 70195 25543 70203 28527
rect 73187 25543 73195 28527
rect 70195 25535 73195 25543
rect 73385 28527 76385 28535
rect 73385 25543 73393 28527
rect 76377 25543 76385 28527
rect 73385 25535 76385 25543
rect 76575 28527 79575 28535
rect 76575 25543 76583 28527
rect 79567 25543 79575 28527
rect 76575 25535 79575 25543
rect 79765 28527 82765 28535
rect 79765 25543 79773 28527
rect 82757 25543 82765 28527
rect 79765 25535 82765 25543
rect 82955 28527 85955 28535
rect 82955 25543 82963 28527
rect 85947 25543 85955 28527
rect 82955 25535 85955 25543
rect 86145 28527 89145 28535
rect 86145 25543 86153 28527
rect 89137 25543 89145 28527
rect 86145 25535 89145 25543
rect 89335 28527 92335 28535
rect 89335 25543 89343 28527
rect 92327 25543 92335 28527
rect 89335 25535 92335 25543
rect 92525 28527 95525 28535
rect 92525 25543 92533 28527
rect 95517 25543 95525 28527
rect 92525 25535 95525 25543
rect 95715 28527 98715 28535
rect 95715 25543 95723 28527
rect 98707 25543 98715 28527
rect 95715 25535 98715 25543
rect 98905 28527 101905 28535
rect 98905 25543 98913 28527
rect 101897 25543 101905 28527
rect 98905 25535 101905 25543
rect 102095 28527 105095 28535
rect 102095 25543 102103 28527
rect 105087 25543 105095 28527
rect 102095 25535 105095 25543
rect 105285 28527 108285 28535
rect 105285 25543 105293 28527
rect 108277 25543 108285 28527
rect 105285 25535 108285 25543
rect 108475 28527 111475 28535
rect 108475 25543 108483 28527
rect 111467 25543 111475 28527
rect 108475 25535 111475 25543
rect 111665 28527 114665 28535
rect 111665 25543 111673 28527
rect 114657 25543 114665 28527
rect 111665 25535 114665 25543
rect 114855 28527 117855 28535
rect 114855 25543 114863 28527
rect 117847 25543 117855 28527
rect 114855 25535 117855 25543
rect 118045 28527 121045 28535
rect 118045 25543 118053 28527
rect 121037 25543 121045 28527
rect 118045 25535 121045 25543
rect 121235 28527 124235 28535
rect 121235 25543 121243 28527
rect 124227 25543 124235 28527
rect 121235 25535 124235 25543
rect 124425 28527 127425 28535
rect 124425 25543 124433 28527
rect 127417 25543 127425 28527
rect 124425 25535 127425 25543
rect 127615 28527 130615 28535
rect 127615 25543 127623 28527
rect 130607 25543 130615 28527
rect 127615 25535 130615 25543
rect 130805 28527 133805 28535
rect 130805 25543 130813 28527
rect 133797 25543 133805 28527
rect 130805 25535 133805 25543
rect 133995 28527 136995 28535
rect 133995 25543 134003 28527
rect 136987 25543 136995 28527
rect 133995 25535 136995 25543
rect 15 25337 3015 25345
rect 15 22353 23 25337
rect 3007 22353 3015 25337
rect 15 22345 3015 22353
rect 3205 25337 6205 25345
rect 3205 22353 3213 25337
rect 6197 22353 6205 25337
rect 3205 22345 6205 22353
rect 6395 25337 9395 25345
rect 6395 22353 6403 25337
rect 9387 22353 9395 25337
rect 6395 22345 9395 22353
rect 9585 25337 12585 25345
rect 9585 22353 9593 25337
rect 12577 22353 12585 25337
rect 9585 22345 12585 22353
rect 12775 25337 15775 25345
rect 12775 22353 12783 25337
rect 15767 22353 15775 25337
rect 12775 22345 15775 22353
rect 15965 25337 18965 25345
rect 15965 22353 15973 25337
rect 18957 22353 18965 25337
rect 15965 22345 18965 22353
rect 19155 25337 22155 25345
rect 19155 22353 19163 25337
rect 22147 22353 22155 25337
rect 19155 22345 22155 22353
rect 22345 25337 25345 25345
rect 22345 22353 22353 25337
rect 25337 22353 25345 25337
rect 22345 22345 25345 22353
rect 25535 25337 28535 25345
rect 25535 22353 25543 25337
rect 28527 22353 28535 25337
rect 25535 22345 28535 22353
rect 28725 25337 31725 25345
rect 28725 22353 28733 25337
rect 31717 22353 31725 25337
rect 28725 22345 31725 22353
rect 31915 25337 34915 25345
rect 31915 22353 31923 25337
rect 34907 22353 34915 25337
rect 31915 22345 34915 22353
rect 35105 25337 38105 25345
rect 35105 22353 35113 25337
rect 38097 22353 38105 25337
rect 35105 22345 38105 22353
rect 38295 25337 41295 25345
rect 38295 22353 38303 25337
rect 41287 22353 41295 25337
rect 38295 22345 41295 22353
rect 41485 25337 44485 25345
rect 41485 22353 41493 25337
rect 44477 22353 44485 25337
rect 41485 22345 44485 22353
rect 44675 25337 47675 25345
rect 44675 22353 44683 25337
rect 47667 22353 47675 25337
rect 44675 22345 47675 22353
rect 47865 25337 50865 25345
rect 47865 22353 47873 25337
rect 50857 22353 50865 25337
rect 47865 22345 50865 22353
rect 51055 25337 54055 25345
rect 51055 22353 51063 25337
rect 54047 22353 54055 25337
rect 51055 22345 54055 22353
rect 54245 25337 57245 25345
rect 54245 22353 54253 25337
rect 57237 22353 57245 25337
rect 54245 22345 57245 22353
rect 57435 25337 60435 25345
rect 57435 22353 57443 25337
rect 60427 22353 60435 25337
rect 57435 22345 60435 22353
rect 60625 25337 63625 25345
rect 60625 22353 60633 25337
rect 63617 22353 63625 25337
rect 60625 22345 63625 22353
rect 63815 25337 66815 25345
rect 63815 22353 63823 25337
rect 66807 22353 66815 25337
rect 63815 22345 66815 22353
rect 67005 25337 70005 25345
rect 67005 22353 67013 25337
rect 69997 22353 70005 25337
rect 67005 22345 70005 22353
rect 70195 25337 73195 25345
rect 70195 22353 70203 25337
rect 73187 22353 73195 25337
rect 70195 22345 73195 22353
rect 73385 25337 76385 25345
rect 73385 22353 73393 25337
rect 76377 22353 76385 25337
rect 73385 22345 76385 22353
rect 76575 25337 79575 25345
rect 76575 22353 76583 25337
rect 79567 22353 79575 25337
rect 76575 22345 79575 22353
rect 79765 25337 82765 25345
rect 79765 22353 79773 25337
rect 82757 22353 82765 25337
rect 79765 22345 82765 22353
rect 82955 25337 85955 25345
rect 82955 22353 82963 25337
rect 85947 22353 85955 25337
rect 82955 22345 85955 22353
rect 86145 25337 89145 25345
rect 86145 22353 86153 25337
rect 89137 22353 89145 25337
rect 86145 22345 89145 22353
rect 89335 25337 92335 25345
rect 89335 22353 89343 25337
rect 92327 22353 92335 25337
rect 89335 22345 92335 22353
rect 92525 25337 95525 25345
rect 92525 22353 92533 25337
rect 95517 22353 95525 25337
rect 92525 22345 95525 22353
rect 95715 25337 98715 25345
rect 95715 22353 95723 25337
rect 98707 22353 98715 25337
rect 95715 22345 98715 22353
rect 98905 25337 101905 25345
rect 98905 22353 98913 25337
rect 101897 22353 101905 25337
rect 98905 22345 101905 22353
rect 102095 25337 105095 25345
rect 102095 22353 102103 25337
rect 105087 22353 105095 25337
rect 102095 22345 105095 22353
rect 105285 25337 108285 25345
rect 105285 22353 105293 25337
rect 108277 22353 108285 25337
rect 105285 22345 108285 22353
rect 108475 25337 111475 25345
rect 108475 22353 108483 25337
rect 111467 22353 111475 25337
rect 108475 22345 111475 22353
rect 111665 25337 114665 25345
rect 111665 22353 111673 25337
rect 114657 22353 114665 25337
rect 111665 22345 114665 22353
rect 114855 25337 117855 25345
rect 114855 22353 114863 25337
rect 117847 22353 117855 25337
rect 114855 22345 117855 22353
rect 118045 25337 121045 25345
rect 118045 22353 118053 25337
rect 121037 22353 121045 25337
rect 118045 22345 121045 22353
rect 121235 25337 124235 25345
rect 121235 22353 121243 25337
rect 124227 22353 124235 25337
rect 121235 22345 124235 22353
rect 124425 25337 127425 25345
rect 124425 22353 124433 25337
rect 127417 22353 127425 25337
rect 124425 22345 127425 22353
rect 127615 25337 130615 25345
rect 127615 22353 127623 25337
rect 130607 22353 130615 25337
rect 127615 22345 130615 22353
rect 130805 25337 133805 25345
rect 130805 22353 130813 25337
rect 133797 22353 133805 25337
rect 130805 22345 133805 22353
rect 133995 25337 136995 25345
rect 133995 22353 134003 25337
rect 136987 22353 136995 25337
rect 133995 22345 136995 22353
rect 15 22147 3015 22155
rect 15 19163 23 22147
rect 3007 19163 3015 22147
rect 15 19155 3015 19163
rect 3205 22147 6205 22155
rect 3205 19163 3213 22147
rect 6197 19163 6205 22147
rect 3205 19155 6205 19163
rect 6395 22147 9395 22155
rect 6395 19163 6403 22147
rect 9387 19163 9395 22147
rect 6395 19155 9395 19163
rect 9585 22147 12585 22155
rect 9585 19163 9593 22147
rect 12577 19163 12585 22147
rect 9585 19155 12585 19163
rect 12775 22147 15775 22155
rect 12775 19163 12783 22147
rect 15767 19163 15775 22147
rect 12775 19155 15775 19163
rect 15965 22147 18965 22155
rect 15965 19163 15973 22147
rect 18957 19163 18965 22147
rect 15965 19155 18965 19163
rect 19155 22147 22155 22155
rect 19155 19163 19163 22147
rect 22147 19163 22155 22147
rect 19155 19155 22155 19163
rect 22345 22147 25345 22155
rect 22345 19163 22353 22147
rect 25337 19163 25345 22147
rect 22345 19155 25345 19163
rect 25535 22147 28535 22155
rect 25535 19163 25543 22147
rect 28527 19163 28535 22147
rect 25535 19155 28535 19163
rect 28725 22147 31725 22155
rect 28725 19163 28733 22147
rect 31717 19163 31725 22147
rect 28725 19155 31725 19163
rect 31915 22147 34915 22155
rect 31915 19163 31923 22147
rect 34907 19163 34915 22147
rect 31915 19155 34915 19163
rect 35105 22147 38105 22155
rect 35105 19163 35113 22147
rect 38097 19163 38105 22147
rect 35105 19155 38105 19163
rect 38295 22147 41295 22155
rect 38295 19163 38303 22147
rect 41287 19163 41295 22147
rect 38295 19155 41295 19163
rect 41485 22147 44485 22155
rect 41485 19163 41493 22147
rect 44477 19163 44485 22147
rect 41485 19155 44485 19163
rect 44675 22147 47675 22155
rect 44675 19163 44683 22147
rect 47667 19163 47675 22147
rect 44675 19155 47675 19163
rect 47865 22147 50865 22155
rect 47865 19163 47873 22147
rect 50857 19163 50865 22147
rect 47865 19155 50865 19163
rect 51055 22147 54055 22155
rect 51055 19163 51063 22147
rect 54047 19163 54055 22147
rect 51055 19155 54055 19163
rect 54245 22147 57245 22155
rect 54245 19163 54253 22147
rect 57237 19163 57245 22147
rect 54245 19155 57245 19163
rect 57435 22147 60435 22155
rect 57435 19163 57443 22147
rect 60427 19163 60435 22147
rect 57435 19155 60435 19163
rect 60625 22147 63625 22155
rect 60625 19163 60633 22147
rect 63617 19163 63625 22147
rect 60625 19155 63625 19163
rect 63815 22147 66815 22155
rect 63815 19163 63823 22147
rect 66807 19163 66815 22147
rect 63815 19155 66815 19163
rect 67005 22147 70005 22155
rect 67005 19163 67013 22147
rect 69997 19163 70005 22147
rect 67005 19155 70005 19163
rect 70195 22147 73195 22155
rect 70195 19163 70203 22147
rect 73187 19163 73195 22147
rect 70195 19155 73195 19163
rect 73385 22147 76385 22155
rect 73385 19163 73393 22147
rect 76377 19163 76385 22147
rect 73385 19155 76385 19163
rect 76575 22147 79575 22155
rect 76575 19163 76583 22147
rect 79567 19163 79575 22147
rect 76575 19155 79575 19163
rect 79765 22147 82765 22155
rect 79765 19163 79773 22147
rect 82757 19163 82765 22147
rect 79765 19155 82765 19163
rect 82955 22147 85955 22155
rect 82955 19163 82963 22147
rect 85947 19163 85955 22147
rect 82955 19155 85955 19163
rect 86145 22147 89145 22155
rect 86145 19163 86153 22147
rect 89137 19163 89145 22147
rect 86145 19155 89145 19163
rect 89335 22147 92335 22155
rect 89335 19163 89343 22147
rect 92327 19163 92335 22147
rect 89335 19155 92335 19163
rect 92525 22147 95525 22155
rect 92525 19163 92533 22147
rect 95517 19163 95525 22147
rect 92525 19155 95525 19163
rect 95715 22147 98715 22155
rect 95715 19163 95723 22147
rect 98707 19163 98715 22147
rect 95715 19155 98715 19163
rect 98905 22147 101905 22155
rect 98905 19163 98913 22147
rect 101897 19163 101905 22147
rect 98905 19155 101905 19163
rect 102095 22147 105095 22155
rect 102095 19163 102103 22147
rect 105087 19163 105095 22147
rect 102095 19155 105095 19163
rect 105285 22147 108285 22155
rect 105285 19163 105293 22147
rect 108277 19163 108285 22147
rect 105285 19155 108285 19163
rect 108475 22147 111475 22155
rect 108475 19163 108483 22147
rect 111467 19163 111475 22147
rect 108475 19155 111475 19163
rect 111665 22147 114665 22155
rect 111665 19163 111673 22147
rect 114657 19163 114665 22147
rect 111665 19155 114665 19163
rect 114855 22147 117855 22155
rect 114855 19163 114863 22147
rect 117847 19163 117855 22147
rect 114855 19155 117855 19163
rect 118045 22147 121045 22155
rect 118045 19163 118053 22147
rect 121037 19163 121045 22147
rect 118045 19155 121045 19163
rect 121235 22147 124235 22155
rect 121235 19163 121243 22147
rect 124227 19163 124235 22147
rect 121235 19155 124235 19163
rect 124425 22147 127425 22155
rect 124425 19163 124433 22147
rect 127417 19163 127425 22147
rect 124425 19155 127425 19163
rect 127615 22147 130615 22155
rect 127615 19163 127623 22147
rect 130607 19163 130615 22147
rect 127615 19155 130615 19163
rect 130805 22147 133805 22155
rect 130805 19163 130813 22147
rect 133797 19163 133805 22147
rect 130805 19155 133805 19163
rect 133995 22147 136995 22155
rect 133995 19163 134003 22147
rect 136987 19163 136995 22147
rect 133995 19155 136995 19163
rect 15 18957 3015 18965
rect 15 15973 23 18957
rect 3007 15973 3015 18957
rect 15 15965 3015 15973
rect 3205 18957 6205 18965
rect 3205 15973 3213 18957
rect 6197 15973 6205 18957
rect 3205 15965 6205 15973
rect 6395 18957 9395 18965
rect 6395 15973 6403 18957
rect 9387 15973 9395 18957
rect 6395 15965 9395 15973
rect 9585 18957 12585 18965
rect 9585 15973 9593 18957
rect 12577 15973 12585 18957
rect 9585 15965 12585 15973
rect 12775 18957 15775 18965
rect 12775 15973 12783 18957
rect 15767 15973 15775 18957
rect 12775 15965 15775 15973
rect 15965 18957 18965 18965
rect 15965 15973 15973 18957
rect 18957 15973 18965 18957
rect 15965 15965 18965 15973
rect 19155 18957 22155 18965
rect 19155 15973 19163 18957
rect 22147 15973 22155 18957
rect 19155 15965 22155 15973
rect 22345 18957 25345 18965
rect 22345 15973 22353 18957
rect 25337 15973 25345 18957
rect 22345 15965 25345 15973
rect 25535 18957 28535 18965
rect 25535 15973 25543 18957
rect 28527 15973 28535 18957
rect 25535 15965 28535 15973
rect 28725 18957 31725 18965
rect 28725 15973 28733 18957
rect 31717 15973 31725 18957
rect 28725 15965 31725 15973
rect 31915 18957 34915 18965
rect 31915 15973 31923 18957
rect 34907 15973 34915 18957
rect 31915 15965 34915 15973
rect 35105 18957 38105 18965
rect 35105 15973 35113 18957
rect 38097 15973 38105 18957
rect 35105 15965 38105 15973
rect 38295 18957 41295 18965
rect 38295 15973 38303 18957
rect 41287 15973 41295 18957
rect 38295 15965 41295 15973
rect 41485 18957 44485 18965
rect 41485 15973 41493 18957
rect 44477 15973 44485 18957
rect 41485 15965 44485 15973
rect 44675 18957 47675 18965
rect 44675 15973 44683 18957
rect 47667 15973 47675 18957
rect 44675 15965 47675 15973
rect 47865 18957 50865 18965
rect 47865 15973 47873 18957
rect 50857 15973 50865 18957
rect 47865 15965 50865 15973
rect 51055 18957 54055 18965
rect 51055 15973 51063 18957
rect 54047 15973 54055 18957
rect 51055 15965 54055 15973
rect 54245 18957 57245 18965
rect 54245 15973 54253 18957
rect 57237 15973 57245 18957
rect 54245 15965 57245 15973
rect 57435 18957 60435 18965
rect 57435 15973 57443 18957
rect 60427 15973 60435 18957
rect 57435 15965 60435 15973
rect 60625 18957 63625 18965
rect 60625 15973 60633 18957
rect 63617 15973 63625 18957
rect 60625 15965 63625 15973
rect 63815 18957 66815 18965
rect 63815 15973 63823 18957
rect 66807 15973 66815 18957
rect 63815 15965 66815 15973
rect 67005 18957 70005 18965
rect 67005 15973 67013 18957
rect 69997 15973 70005 18957
rect 67005 15965 70005 15973
rect 70195 18957 73195 18965
rect 70195 15973 70203 18957
rect 73187 15973 73195 18957
rect 70195 15965 73195 15973
rect 73385 18957 76385 18965
rect 73385 15973 73393 18957
rect 76377 15973 76385 18957
rect 73385 15965 76385 15973
rect 76575 18957 79575 18965
rect 76575 15973 76583 18957
rect 79567 15973 79575 18957
rect 76575 15965 79575 15973
rect 79765 18957 82765 18965
rect 79765 15973 79773 18957
rect 82757 15973 82765 18957
rect 79765 15965 82765 15973
rect 82955 18957 85955 18965
rect 82955 15973 82963 18957
rect 85947 15973 85955 18957
rect 82955 15965 85955 15973
rect 86145 18957 89145 18965
rect 86145 15973 86153 18957
rect 89137 15973 89145 18957
rect 86145 15965 89145 15973
rect 89335 18957 92335 18965
rect 89335 15973 89343 18957
rect 92327 15973 92335 18957
rect 89335 15965 92335 15973
rect 92525 18957 95525 18965
rect 92525 15973 92533 18957
rect 95517 15973 95525 18957
rect 92525 15965 95525 15973
rect 95715 18957 98715 18965
rect 95715 15973 95723 18957
rect 98707 15973 98715 18957
rect 95715 15965 98715 15973
rect 98905 18957 101905 18965
rect 98905 15973 98913 18957
rect 101897 15973 101905 18957
rect 98905 15965 101905 15973
rect 102095 18957 105095 18965
rect 102095 15973 102103 18957
rect 105087 15973 105095 18957
rect 102095 15965 105095 15973
rect 105285 18957 108285 18965
rect 105285 15973 105293 18957
rect 108277 15973 108285 18957
rect 105285 15965 108285 15973
rect 108475 18957 111475 18965
rect 108475 15973 108483 18957
rect 111467 15973 111475 18957
rect 108475 15965 111475 15973
rect 111665 18957 114665 18965
rect 111665 15973 111673 18957
rect 114657 15973 114665 18957
rect 111665 15965 114665 15973
rect 114855 18957 117855 18965
rect 114855 15973 114863 18957
rect 117847 15973 117855 18957
rect 114855 15965 117855 15973
rect 118045 18957 121045 18965
rect 118045 15973 118053 18957
rect 121037 15973 121045 18957
rect 118045 15965 121045 15973
rect 121235 18957 124235 18965
rect 121235 15973 121243 18957
rect 124227 15973 124235 18957
rect 121235 15965 124235 15973
rect 124425 18957 127425 18965
rect 124425 15973 124433 18957
rect 127417 15973 127425 18957
rect 124425 15965 127425 15973
rect 127615 18957 130615 18965
rect 127615 15973 127623 18957
rect 130607 15973 130615 18957
rect 127615 15965 130615 15973
rect 130805 18957 133805 18965
rect 130805 15973 130813 18957
rect 133797 15973 133805 18957
rect 130805 15965 133805 15973
rect 133995 18957 136995 18965
rect 133995 15973 134003 18957
rect 136987 15973 136995 18957
rect 133995 15965 136995 15973
rect 15 15767 3015 15775
rect 15 12783 23 15767
rect 3007 12783 3015 15767
rect 15 12775 3015 12783
rect 3205 15767 6205 15775
rect 3205 12783 3213 15767
rect 6197 12783 6205 15767
rect 3205 12775 6205 12783
rect 6395 15767 9395 15775
rect 6395 12783 6403 15767
rect 9387 12783 9395 15767
rect 6395 12775 9395 12783
rect 9585 15767 12585 15775
rect 9585 12783 9593 15767
rect 12577 12783 12585 15767
rect 9585 12775 12585 12783
rect 12775 15767 15775 15775
rect 12775 12783 12783 15767
rect 15767 12783 15775 15767
rect 12775 12775 15775 12783
rect 15965 15767 18965 15775
rect 15965 12783 15973 15767
rect 18957 12783 18965 15767
rect 15965 12775 18965 12783
rect 19155 15767 22155 15775
rect 19155 12783 19163 15767
rect 22147 12783 22155 15767
rect 19155 12775 22155 12783
rect 22345 15767 25345 15775
rect 22345 12783 22353 15767
rect 25337 12783 25345 15767
rect 22345 12775 25345 12783
rect 25535 15767 28535 15775
rect 25535 12783 25543 15767
rect 28527 12783 28535 15767
rect 25535 12775 28535 12783
rect 28725 15767 31725 15775
rect 28725 12783 28733 15767
rect 31717 12783 31725 15767
rect 28725 12775 31725 12783
rect 31915 15767 34915 15775
rect 31915 12783 31923 15767
rect 34907 12783 34915 15767
rect 31915 12775 34915 12783
rect 35105 15767 38105 15775
rect 35105 12783 35113 15767
rect 38097 12783 38105 15767
rect 35105 12775 38105 12783
rect 38295 15767 41295 15775
rect 38295 12783 38303 15767
rect 41287 12783 41295 15767
rect 38295 12775 41295 12783
rect 41485 15767 44485 15775
rect 41485 12783 41493 15767
rect 44477 12783 44485 15767
rect 41485 12775 44485 12783
rect 44675 15767 47675 15775
rect 44675 12783 44683 15767
rect 47667 12783 47675 15767
rect 44675 12775 47675 12783
rect 47865 15767 50865 15775
rect 47865 12783 47873 15767
rect 50857 12783 50865 15767
rect 47865 12775 50865 12783
rect 51055 15767 54055 15775
rect 51055 12783 51063 15767
rect 54047 12783 54055 15767
rect 51055 12775 54055 12783
rect 54245 15767 57245 15775
rect 54245 12783 54253 15767
rect 57237 12783 57245 15767
rect 54245 12775 57245 12783
rect 57435 15767 60435 15775
rect 57435 12783 57443 15767
rect 60427 12783 60435 15767
rect 57435 12775 60435 12783
rect 60625 15767 63625 15775
rect 60625 12783 60633 15767
rect 63617 12783 63625 15767
rect 60625 12775 63625 12783
rect 63815 15767 66815 15775
rect 63815 12783 63823 15767
rect 66807 12783 66815 15767
rect 63815 12775 66815 12783
rect 67005 15767 70005 15775
rect 67005 12783 67013 15767
rect 69997 12783 70005 15767
rect 67005 12775 70005 12783
rect 70195 15767 73195 15775
rect 70195 12783 70203 15767
rect 73187 12783 73195 15767
rect 70195 12775 73195 12783
rect 73385 15767 76385 15775
rect 73385 12783 73393 15767
rect 76377 12783 76385 15767
rect 73385 12775 76385 12783
rect 76575 15767 79575 15775
rect 76575 12783 76583 15767
rect 79567 12783 79575 15767
rect 76575 12775 79575 12783
rect 79765 15767 82765 15775
rect 79765 12783 79773 15767
rect 82757 12783 82765 15767
rect 79765 12775 82765 12783
rect 82955 15767 85955 15775
rect 82955 12783 82963 15767
rect 85947 12783 85955 15767
rect 82955 12775 85955 12783
rect 86145 15767 89145 15775
rect 86145 12783 86153 15767
rect 89137 12783 89145 15767
rect 86145 12775 89145 12783
rect 89335 15767 92335 15775
rect 89335 12783 89343 15767
rect 92327 12783 92335 15767
rect 89335 12775 92335 12783
rect 92525 15767 95525 15775
rect 92525 12783 92533 15767
rect 95517 12783 95525 15767
rect 92525 12775 95525 12783
rect 95715 15767 98715 15775
rect 95715 12783 95723 15767
rect 98707 12783 98715 15767
rect 95715 12775 98715 12783
rect 98905 15767 101905 15775
rect 98905 12783 98913 15767
rect 101897 12783 101905 15767
rect 98905 12775 101905 12783
rect 102095 15767 105095 15775
rect 102095 12783 102103 15767
rect 105087 12783 105095 15767
rect 102095 12775 105095 12783
rect 105285 15767 108285 15775
rect 105285 12783 105293 15767
rect 108277 12783 108285 15767
rect 105285 12775 108285 12783
rect 108475 15767 111475 15775
rect 108475 12783 108483 15767
rect 111467 12783 111475 15767
rect 108475 12775 111475 12783
rect 111665 15767 114665 15775
rect 111665 12783 111673 15767
rect 114657 12783 114665 15767
rect 111665 12775 114665 12783
rect 114855 15767 117855 15775
rect 114855 12783 114863 15767
rect 117847 12783 117855 15767
rect 114855 12775 117855 12783
rect 118045 15767 121045 15775
rect 118045 12783 118053 15767
rect 121037 12783 121045 15767
rect 118045 12775 121045 12783
rect 121235 15767 124235 15775
rect 121235 12783 121243 15767
rect 124227 12783 124235 15767
rect 121235 12775 124235 12783
rect 124425 15767 127425 15775
rect 124425 12783 124433 15767
rect 127417 12783 127425 15767
rect 124425 12775 127425 12783
rect 127615 15767 130615 15775
rect 127615 12783 127623 15767
rect 130607 12783 130615 15767
rect 127615 12775 130615 12783
rect 130805 15767 133805 15775
rect 130805 12783 130813 15767
rect 133797 12783 133805 15767
rect 130805 12775 133805 12783
rect 133995 15767 136995 15775
rect 133995 12783 134003 15767
rect 136987 12783 136995 15767
rect 133995 12775 136995 12783
rect 15 12577 3015 12585
rect 15 9593 23 12577
rect 3007 9593 3015 12577
rect 15 9585 3015 9593
rect 3205 12577 6205 12585
rect 3205 9593 3213 12577
rect 6197 9593 6205 12577
rect 3205 9585 6205 9593
rect 6395 12577 9395 12585
rect 6395 9593 6403 12577
rect 9387 9593 9395 12577
rect 6395 9585 9395 9593
rect 9585 12577 12585 12585
rect 9585 9593 9593 12577
rect 12577 9593 12585 12577
rect 9585 9585 12585 9593
rect 12775 12577 15775 12585
rect 12775 9593 12783 12577
rect 15767 9593 15775 12577
rect 12775 9585 15775 9593
rect 15965 12577 18965 12585
rect 15965 9593 15973 12577
rect 18957 9593 18965 12577
rect 15965 9585 18965 9593
rect 19155 12577 22155 12585
rect 19155 9593 19163 12577
rect 22147 9593 22155 12577
rect 19155 9585 22155 9593
rect 22345 12577 25345 12585
rect 22345 9593 22353 12577
rect 25337 9593 25345 12577
rect 22345 9585 25345 9593
rect 25535 12577 28535 12585
rect 25535 9593 25543 12577
rect 28527 9593 28535 12577
rect 25535 9585 28535 9593
rect 28725 12577 31725 12585
rect 28725 9593 28733 12577
rect 31717 9593 31725 12577
rect 28725 9585 31725 9593
rect 31915 12577 34915 12585
rect 31915 9593 31923 12577
rect 34907 9593 34915 12577
rect 31915 9585 34915 9593
rect 35105 12577 38105 12585
rect 35105 9593 35113 12577
rect 38097 9593 38105 12577
rect 35105 9585 38105 9593
rect 38295 12577 41295 12585
rect 38295 9593 38303 12577
rect 41287 9593 41295 12577
rect 38295 9585 41295 9593
rect 41485 12577 44485 12585
rect 41485 9593 41493 12577
rect 44477 9593 44485 12577
rect 41485 9585 44485 9593
rect 44675 12577 47675 12585
rect 44675 9593 44683 12577
rect 47667 9593 47675 12577
rect 44675 9585 47675 9593
rect 47865 12577 50865 12585
rect 47865 9593 47873 12577
rect 50857 9593 50865 12577
rect 47865 9585 50865 9593
rect 51055 12577 54055 12585
rect 51055 9593 51063 12577
rect 54047 9593 54055 12577
rect 51055 9585 54055 9593
rect 54245 12577 57245 12585
rect 54245 9593 54253 12577
rect 57237 9593 57245 12577
rect 54245 9585 57245 9593
rect 57435 12577 60435 12585
rect 57435 9593 57443 12577
rect 60427 9593 60435 12577
rect 57435 9585 60435 9593
rect 60625 12577 63625 12585
rect 60625 9593 60633 12577
rect 63617 9593 63625 12577
rect 60625 9585 63625 9593
rect 63815 12577 66815 12585
rect 63815 9593 63823 12577
rect 66807 9593 66815 12577
rect 63815 9585 66815 9593
rect 67005 12577 70005 12585
rect 67005 9593 67013 12577
rect 69997 9593 70005 12577
rect 67005 9585 70005 9593
rect 70195 12577 73195 12585
rect 70195 9593 70203 12577
rect 73187 9593 73195 12577
rect 70195 9585 73195 9593
rect 73385 12577 76385 12585
rect 73385 9593 73393 12577
rect 76377 9593 76385 12577
rect 73385 9585 76385 9593
rect 76575 12577 79575 12585
rect 76575 9593 76583 12577
rect 79567 9593 79575 12577
rect 76575 9585 79575 9593
rect 79765 12577 82765 12585
rect 79765 9593 79773 12577
rect 82757 9593 82765 12577
rect 79765 9585 82765 9593
rect 82955 12577 85955 12585
rect 82955 9593 82963 12577
rect 85947 9593 85955 12577
rect 82955 9585 85955 9593
rect 86145 12577 89145 12585
rect 86145 9593 86153 12577
rect 89137 9593 89145 12577
rect 86145 9585 89145 9593
rect 89335 12577 92335 12585
rect 89335 9593 89343 12577
rect 92327 9593 92335 12577
rect 89335 9585 92335 9593
rect 92525 12577 95525 12585
rect 92525 9593 92533 12577
rect 95517 9593 95525 12577
rect 92525 9585 95525 9593
rect 95715 12577 98715 12585
rect 95715 9593 95723 12577
rect 98707 9593 98715 12577
rect 95715 9585 98715 9593
rect 98905 12577 101905 12585
rect 98905 9593 98913 12577
rect 101897 9593 101905 12577
rect 98905 9585 101905 9593
rect 102095 12577 105095 12585
rect 102095 9593 102103 12577
rect 105087 9593 105095 12577
rect 102095 9585 105095 9593
rect 105285 12577 108285 12585
rect 105285 9593 105293 12577
rect 108277 9593 108285 12577
rect 105285 9585 108285 9593
rect 108475 12577 111475 12585
rect 108475 9593 108483 12577
rect 111467 9593 111475 12577
rect 108475 9585 111475 9593
rect 111665 12577 114665 12585
rect 111665 9593 111673 12577
rect 114657 9593 114665 12577
rect 111665 9585 114665 9593
rect 114855 12577 117855 12585
rect 114855 9593 114863 12577
rect 117847 9593 117855 12577
rect 114855 9585 117855 9593
rect 118045 12577 121045 12585
rect 118045 9593 118053 12577
rect 121037 9593 121045 12577
rect 118045 9585 121045 9593
rect 121235 12577 124235 12585
rect 121235 9593 121243 12577
rect 124227 9593 124235 12577
rect 121235 9585 124235 9593
rect 124425 12577 127425 12585
rect 124425 9593 124433 12577
rect 127417 9593 127425 12577
rect 124425 9585 127425 9593
rect 127615 12577 130615 12585
rect 127615 9593 127623 12577
rect 130607 9593 130615 12577
rect 127615 9585 130615 9593
rect 130805 12577 133805 12585
rect 130805 9593 130813 12577
rect 133797 9593 133805 12577
rect 130805 9585 133805 9593
rect 133995 12577 136995 12585
rect 133995 9593 134003 12577
rect 136987 9593 136995 12577
rect 133995 9585 136995 9593
rect 15 9387 3015 9395
rect 15 6403 23 9387
rect 3007 6403 3015 9387
rect 15 6395 3015 6403
rect 3205 9387 6205 9395
rect 3205 6403 3213 9387
rect 6197 6403 6205 9387
rect 3205 6395 6205 6403
rect 6395 9387 9395 9395
rect 6395 6403 6403 9387
rect 9387 6403 9395 9387
rect 6395 6395 9395 6403
rect 9585 9387 12585 9395
rect 9585 6403 9593 9387
rect 12577 6403 12585 9387
rect 9585 6395 12585 6403
rect 12775 9387 15775 9395
rect 12775 6403 12783 9387
rect 15767 6403 15775 9387
rect 12775 6395 15775 6403
rect 15965 9387 18965 9395
rect 15965 6403 15973 9387
rect 18957 6403 18965 9387
rect 15965 6395 18965 6403
rect 19155 9387 22155 9395
rect 19155 6403 19163 9387
rect 22147 6403 22155 9387
rect 19155 6395 22155 6403
rect 22345 9387 25345 9395
rect 22345 6403 22353 9387
rect 25337 6403 25345 9387
rect 22345 6395 25345 6403
rect 25535 9387 28535 9395
rect 25535 6403 25543 9387
rect 28527 6403 28535 9387
rect 25535 6395 28535 6403
rect 28725 9387 31725 9395
rect 28725 6403 28733 9387
rect 31717 6403 31725 9387
rect 28725 6395 31725 6403
rect 31915 9387 34915 9395
rect 31915 6403 31923 9387
rect 34907 6403 34915 9387
rect 31915 6395 34915 6403
rect 35105 9387 38105 9395
rect 35105 6403 35113 9387
rect 38097 6403 38105 9387
rect 35105 6395 38105 6403
rect 38295 9387 41295 9395
rect 38295 6403 38303 9387
rect 41287 6403 41295 9387
rect 38295 6395 41295 6403
rect 41485 9387 44485 9395
rect 41485 6403 41493 9387
rect 44477 6403 44485 9387
rect 41485 6395 44485 6403
rect 44675 9387 47675 9395
rect 44675 6403 44683 9387
rect 47667 6403 47675 9387
rect 44675 6395 47675 6403
rect 47865 9387 50865 9395
rect 47865 6403 47873 9387
rect 50857 6403 50865 9387
rect 47865 6395 50865 6403
rect 51055 9387 54055 9395
rect 51055 6403 51063 9387
rect 54047 6403 54055 9387
rect 51055 6395 54055 6403
rect 54245 9387 57245 9395
rect 54245 6403 54253 9387
rect 57237 6403 57245 9387
rect 54245 6395 57245 6403
rect 57435 9387 60435 9395
rect 57435 6403 57443 9387
rect 60427 6403 60435 9387
rect 57435 6395 60435 6403
rect 60625 9387 63625 9395
rect 60625 6403 60633 9387
rect 63617 6403 63625 9387
rect 60625 6395 63625 6403
rect 63815 9387 66815 9395
rect 63815 6403 63823 9387
rect 66807 6403 66815 9387
rect 63815 6395 66815 6403
rect 67005 9387 70005 9395
rect 67005 6403 67013 9387
rect 69997 6403 70005 9387
rect 67005 6395 70005 6403
rect 70195 9387 73195 9395
rect 70195 6403 70203 9387
rect 73187 6403 73195 9387
rect 70195 6395 73195 6403
rect 73385 9387 76385 9395
rect 73385 6403 73393 9387
rect 76377 6403 76385 9387
rect 73385 6395 76385 6403
rect 76575 9387 79575 9395
rect 76575 6403 76583 9387
rect 79567 6403 79575 9387
rect 76575 6395 79575 6403
rect 79765 9387 82765 9395
rect 79765 6403 79773 9387
rect 82757 6403 82765 9387
rect 79765 6395 82765 6403
rect 82955 9387 85955 9395
rect 82955 6403 82963 9387
rect 85947 6403 85955 9387
rect 82955 6395 85955 6403
rect 86145 9387 89145 9395
rect 86145 6403 86153 9387
rect 89137 6403 89145 9387
rect 86145 6395 89145 6403
rect 89335 9387 92335 9395
rect 89335 6403 89343 9387
rect 92327 6403 92335 9387
rect 89335 6395 92335 6403
rect 92525 9387 95525 9395
rect 92525 6403 92533 9387
rect 95517 6403 95525 9387
rect 92525 6395 95525 6403
rect 95715 9387 98715 9395
rect 95715 6403 95723 9387
rect 98707 6403 98715 9387
rect 95715 6395 98715 6403
rect 98905 9387 101905 9395
rect 98905 6403 98913 9387
rect 101897 6403 101905 9387
rect 98905 6395 101905 6403
rect 102095 9387 105095 9395
rect 102095 6403 102103 9387
rect 105087 6403 105095 9387
rect 102095 6395 105095 6403
rect 105285 9387 108285 9395
rect 105285 6403 105293 9387
rect 108277 6403 108285 9387
rect 105285 6395 108285 6403
rect 108475 9387 111475 9395
rect 108475 6403 108483 9387
rect 111467 6403 111475 9387
rect 108475 6395 111475 6403
rect 111665 9387 114665 9395
rect 111665 6403 111673 9387
rect 114657 6403 114665 9387
rect 111665 6395 114665 6403
rect 114855 9387 117855 9395
rect 114855 6403 114863 9387
rect 117847 6403 117855 9387
rect 114855 6395 117855 6403
rect 118045 9387 121045 9395
rect 118045 6403 118053 9387
rect 121037 6403 121045 9387
rect 118045 6395 121045 6403
rect 121235 9387 124235 9395
rect 121235 6403 121243 9387
rect 124227 6403 124235 9387
rect 121235 6395 124235 6403
rect 124425 9387 127425 9395
rect 124425 6403 124433 9387
rect 127417 6403 127425 9387
rect 124425 6395 127425 6403
rect 127615 9387 130615 9395
rect 127615 6403 127623 9387
rect 130607 6403 130615 9387
rect 127615 6395 130615 6403
rect 130805 9387 133805 9395
rect 130805 6403 130813 9387
rect 133797 6403 133805 9387
rect 130805 6395 133805 6403
rect 133995 9387 136995 9395
rect 133995 6403 134003 9387
rect 136987 6403 136995 9387
rect 133995 6395 136995 6403
rect 15 6197 3015 6205
rect 15 3213 23 6197
rect 3007 3213 3015 6197
rect 15 3205 3015 3213
rect 3205 6197 6205 6205
rect 3205 3213 3213 6197
rect 6197 3213 6205 6197
rect 3205 3205 6205 3213
rect 6395 6197 9395 6205
rect 6395 3213 6403 6197
rect 9387 3213 9395 6197
rect 6395 3205 9395 3213
rect 9585 6197 12585 6205
rect 9585 3213 9593 6197
rect 12577 3213 12585 6197
rect 9585 3205 12585 3213
rect 12775 6197 15775 6205
rect 12775 3213 12783 6197
rect 15767 3213 15775 6197
rect 12775 3205 15775 3213
rect 15965 6197 18965 6205
rect 15965 3213 15973 6197
rect 18957 3213 18965 6197
rect 15965 3205 18965 3213
rect 19155 6197 22155 6205
rect 19155 3213 19163 6197
rect 22147 3213 22155 6197
rect 19155 3205 22155 3213
rect 22345 6197 25345 6205
rect 22345 3213 22353 6197
rect 25337 3213 25345 6197
rect 22345 3205 25345 3213
rect 25535 6197 28535 6205
rect 25535 3213 25543 6197
rect 28527 3213 28535 6197
rect 25535 3205 28535 3213
rect 28725 6197 31725 6205
rect 28725 3213 28733 6197
rect 31717 3213 31725 6197
rect 28725 3205 31725 3213
rect 31915 6197 34915 6205
rect 31915 3213 31923 6197
rect 34907 3213 34915 6197
rect 31915 3205 34915 3213
rect 35105 6197 38105 6205
rect 35105 3213 35113 6197
rect 38097 3213 38105 6197
rect 35105 3205 38105 3213
rect 38295 6197 41295 6205
rect 38295 3213 38303 6197
rect 41287 3213 41295 6197
rect 38295 3205 41295 3213
rect 41485 6197 44485 6205
rect 41485 3213 41493 6197
rect 44477 3213 44485 6197
rect 41485 3205 44485 3213
rect 44675 6197 47675 6205
rect 44675 3213 44683 6197
rect 47667 3213 47675 6197
rect 44675 3205 47675 3213
rect 47865 6197 50865 6205
rect 47865 3213 47873 6197
rect 50857 3213 50865 6197
rect 47865 3205 50865 3213
rect 51055 6197 54055 6205
rect 51055 3213 51063 6197
rect 54047 3213 54055 6197
rect 51055 3205 54055 3213
rect 54245 6197 57245 6205
rect 54245 3213 54253 6197
rect 57237 3213 57245 6197
rect 54245 3205 57245 3213
rect 57435 6197 60435 6205
rect 57435 3213 57443 6197
rect 60427 3213 60435 6197
rect 57435 3205 60435 3213
rect 60625 6197 63625 6205
rect 60625 3213 60633 6197
rect 63617 3213 63625 6197
rect 60625 3205 63625 3213
rect 63815 6197 66815 6205
rect 63815 3213 63823 6197
rect 66807 3213 66815 6197
rect 63815 3205 66815 3213
rect 67005 6197 70005 6205
rect 67005 3213 67013 6197
rect 69997 3213 70005 6197
rect 67005 3205 70005 3213
rect 70195 6197 73195 6205
rect 70195 3213 70203 6197
rect 73187 3213 73195 6197
rect 70195 3205 73195 3213
rect 73385 6197 76385 6205
rect 73385 3213 73393 6197
rect 76377 3213 76385 6197
rect 73385 3205 76385 3213
rect 76575 6197 79575 6205
rect 76575 3213 76583 6197
rect 79567 3213 79575 6197
rect 76575 3205 79575 3213
rect 79765 6197 82765 6205
rect 79765 3213 79773 6197
rect 82757 3213 82765 6197
rect 79765 3205 82765 3213
rect 82955 6197 85955 6205
rect 82955 3213 82963 6197
rect 85947 3213 85955 6197
rect 82955 3205 85955 3213
rect 86145 6197 89145 6205
rect 86145 3213 86153 6197
rect 89137 3213 89145 6197
rect 86145 3205 89145 3213
rect 89335 6197 92335 6205
rect 89335 3213 89343 6197
rect 92327 3213 92335 6197
rect 89335 3205 92335 3213
rect 92525 6197 95525 6205
rect 92525 3213 92533 6197
rect 95517 3213 95525 6197
rect 92525 3205 95525 3213
rect 95715 6197 98715 6205
rect 95715 3213 95723 6197
rect 98707 3213 98715 6197
rect 95715 3205 98715 3213
rect 98905 6197 101905 6205
rect 98905 3213 98913 6197
rect 101897 3213 101905 6197
rect 98905 3205 101905 3213
rect 102095 6197 105095 6205
rect 102095 3213 102103 6197
rect 105087 3213 105095 6197
rect 102095 3205 105095 3213
rect 105285 6197 108285 6205
rect 105285 3213 105293 6197
rect 108277 3213 108285 6197
rect 105285 3205 108285 3213
rect 108475 6197 111475 6205
rect 108475 3213 108483 6197
rect 111467 3213 111475 6197
rect 108475 3205 111475 3213
rect 111665 6197 114665 6205
rect 111665 3213 111673 6197
rect 114657 3213 114665 6197
rect 111665 3205 114665 3213
rect 114855 6197 117855 6205
rect 114855 3213 114863 6197
rect 117847 3213 117855 6197
rect 114855 3205 117855 3213
rect 118045 6197 121045 6205
rect 118045 3213 118053 6197
rect 121037 3213 121045 6197
rect 118045 3205 121045 3213
rect 121235 6197 124235 6205
rect 121235 3213 121243 6197
rect 124227 3213 124235 6197
rect 121235 3205 124235 3213
rect 124425 6197 127425 6205
rect 124425 3213 124433 6197
rect 127417 3213 127425 6197
rect 124425 3205 127425 3213
rect 127615 6197 130615 6205
rect 127615 3213 127623 6197
rect 130607 3213 130615 6197
rect 127615 3205 130615 3213
rect 130805 6197 133805 6205
rect 130805 3213 130813 6197
rect 133797 3213 133805 6197
rect 130805 3205 133805 3213
rect 133995 6197 136995 6205
rect 133995 3213 134003 6197
rect 136987 3213 136995 6197
rect 133995 3205 136995 3213
rect 15 3007 3015 3015
rect 15 23 23 3007
rect 3007 23 3015 3007
rect 15 15 3015 23
rect 3205 3007 6205 3015
rect 3205 23 3213 3007
rect 6197 23 6205 3007
rect 3205 15 6205 23
rect 6395 3007 9395 3015
rect 6395 23 6403 3007
rect 9387 23 9395 3007
rect 6395 15 9395 23
rect 9585 3007 12585 3015
rect 9585 23 9593 3007
rect 12577 23 12585 3007
rect 9585 15 12585 23
rect 12775 3007 15775 3015
rect 12775 23 12783 3007
rect 15767 23 15775 3007
rect 12775 15 15775 23
rect 15965 3007 18965 3015
rect 15965 23 15973 3007
rect 18957 23 18965 3007
rect 15965 15 18965 23
rect 19155 3007 22155 3015
rect 19155 23 19163 3007
rect 22147 23 22155 3007
rect 19155 15 22155 23
rect 22345 3007 25345 3015
rect 22345 23 22353 3007
rect 25337 23 25345 3007
rect 22345 15 25345 23
rect 25535 3007 28535 3015
rect 25535 23 25543 3007
rect 28527 23 28535 3007
rect 25535 15 28535 23
rect 28725 3007 31725 3015
rect 28725 23 28733 3007
rect 31717 23 31725 3007
rect 28725 15 31725 23
rect 31915 3007 34915 3015
rect 31915 23 31923 3007
rect 34907 23 34915 3007
rect 31915 15 34915 23
rect 35105 3007 38105 3015
rect 35105 23 35113 3007
rect 38097 23 38105 3007
rect 35105 15 38105 23
rect 38295 3007 41295 3015
rect 38295 23 38303 3007
rect 41287 23 41295 3007
rect 38295 15 41295 23
rect 41485 3007 44485 3015
rect 41485 23 41493 3007
rect 44477 23 44485 3007
rect 41485 15 44485 23
rect 44675 3007 47675 3015
rect 44675 23 44683 3007
rect 47667 23 47675 3007
rect 44675 15 47675 23
rect 47865 3007 50865 3015
rect 47865 23 47873 3007
rect 50857 23 50865 3007
rect 47865 15 50865 23
rect 51055 3007 54055 3015
rect 51055 23 51063 3007
rect 54047 23 54055 3007
rect 51055 15 54055 23
rect 54245 3007 57245 3015
rect 54245 23 54253 3007
rect 57237 23 57245 3007
rect 54245 15 57245 23
rect 57435 3007 60435 3015
rect 57435 23 57443 3007
rect 60427 23 60435 3007
rect 57435 15 60435 23
rect 60625 3007 63625 3015
rect 60625 23 60633 3007
rect 63617 23 63625 3007
rect 60625 15 63625 23
rect 63815 3007 66815 3015
rect 63815 23 63823 3007
rect 66807 23 66815 3007
rect 63815 15 66815 23
rect 67005 3007 70005 3015
rect 67005 23 67013 3007
rect 69997 23 70005 3007
rect 67005 15 70005 23
rect 70195 3007 73195 3015
rect 70195 23 70203 3007
rect 73187 23 73195 3007
rect 70195 15 73195 23
rect 73385 3007 76385 3015
rect 73385 23 73393 3007
rect 76377 23 76385 3007
rect 73385 15 76385 23
rect 76575 3007 79575 3015
rect 76575 23 76583 3007
rect 79567 23 79575 3007
rect 76575 15 79575 23
rect 79765 3007 82765 3015
rect 79765 23 79773 3007
rect 82757 23 82765 3007
rect 79765 15 82765 23
rect 82955 3007 85955 3015
rect 82955 23 82963 3007
rect 85947 23 85955 3007
rect 82955 15 85955 23
rect 86145 3007 89145 3015
rect 86145 23 86153 3007
rect 89137 23 89145 3007
rect 86145 15 89145 23
rect 89335 3007 92335 3015
rect 89335 23 89343 3007
rect 92327 23 92335 3007
rect 89335 15 92335 23
rect 92525 3007 95525 3015
rect 92525 23 92533 3007
rect 95517 23 95525 3007
rect 92525 15 95525 23
rect 95715 3007 98715 3015
rect 95715 23 95723 3007
rect 98707 23 98715 3007
rect 95715 15 98715 23
rect 98905 3007 101905 3015
rect 98905 23 98913 3007
rect 101897 23 101905 3007
rect 98905 15 101905 23
rect 102095 3007 105095 3015
rect 102095 23 102103 3007
rect 105087 23 105095 3007
rect 102095 15 105095 23
rect 105285 3007 108285 3015
rect 105285 23 105293 3007
rect 108277 23 108285 3007
rect 105285 15 108285 23
rect 108475 3007 111475 3015
rect 108475 23 108483 3007
rect 111467 23 111475 3007
rect 108475 15 111475 23
rect 111665 3007 114665 3015
rect 111665 23 111673 3007
rect 114657 23 114665 3007
rect 111665 15 114665 23
rect 114855 3007 117855 3015
rect 114855 23 114863 3007
rect 117847 23 117855 3007
rect 114855 15 117855 23
rect 118045 3007 121045 3015
rect 118045 23 118053 3007
rect 121037 23 121045 3007
rect 118045 15 121045 23
rect 121235 3007 124235 3015
rect 121235 23 121243 3007
rect 124227 23 124235 3007
rect 121235 15 124235 23
rect 124425 3007 127425 3015
rect 124425 23 124433 3007
rect 127417 23 127425 3007
rect 124425 15 127425 23
rect 127615 3007 130615 3015
rect 127615 23 127623 3007
rect 130607 23 130615 3007
rect 127615 15 130615 23
rect 130805 3007 133805 3015
rect 130805 23 130813 3007
rect 133797 23 133805 3007
rect 130805 15 133805 23
rect 133995 3007 136995 3015
rect 133995 23 134003 3007
rect 136987 23 136995 3007
rect 133995 15 136995 23
<< mimcap2contact >>
rect 23 162713 3007 165697
rect 3213 162713 6197 165697
rect 6403 162713 9387 165697
rect 9593 162713 12577 165697
rect 12783 162713 15767 165697
rect 15973 162713 18957 165697
rect 19163 162713 22147 165697
rect 22353 162713 25337 165697
rect 25543 162713 28527 165697
rect 28733 162713 31717 165697
rect 31923 162713 34907 165697
rect 35113 162713 38097 165697
rect 38303 162713 41287 165697
rect 41493 162713 44477 165697
rect 44683 162713 47667 165697
rect 47873 162713 50857 165697
rect 51063 162713 54047 165697
rect 54253 162713 57237 165697
rect 57443 162713 60427 165697
rect 60633 162713 63617 165697
rect 63823 162713 66807 165697
rect 67013 162713 69997 165697
rect 70203 162713 73187 165697
rect 73393 162713 76377 165697
rect 76583 162713 79567 165697
rect 79773 162713 82757 165697
rect 82963 162713 85947 165697
rect 86153 162713 89137 165697
rect 89343 162713 92327 165697
rect 92533 162713 95517 165697
rect 95723 162713 98707 165697
rect 98913 162713 101897 165697
rect 102103 162713 105087 165697
rect 105293 162713 108277 165697
rect 108483 162713 111467 165697
rect 111673 162713 114657 165697
rect 114863 162713 117847 165697
rect 118053 162713 121037 165697
rect 121243 162713 124227 165697
rect 124433 162713 127417 165697
rect 127623 162713 130607 165697
rect 130813 162713 133797 165697
rect 134003 162713 136987 165697
rect 23 159523 3007 162507
rect 3213 159523 6197 162507
rect 6403 159523 9387 162507
rect 9593 159523 12577 162507
rect 12783 159523 15767 162507
rect 15973 159523 18957 162507
rect 19163 159523 22147 162507
rect 22353 159523 25337 162507
rect 25543 159523 28527 162507
rect 28733 159523 31717 162507
rect 31923 159523 34907 162507
rect 35113 159523 38097 162507
rect 38303 159523 41287 162507
rect 41493 159523 44477 162507
rect 44683 159523 47667 162507
rect 47873 159523 50857 162507
rect 51063 159523 54047 162507
rect 54253 159523 57237 162507
rect 57443 159523 60427 162507
rect 60633 159523 63617 162507
rect 63823 159523 66807 162507
rect 67013 159523 69997 162507
rect 70203 159523 73187 162507
rect 73393 159523 76377 162507
rect 76583 159523 79567 162507
rect 79773 159523 82757 162507
rect 82963 159523 85947 162507
rect 86153 159523 89137 162507
rect 89343 159523 92327 162507
rect 92533 159523 95517 162507
rect 95723 159523 98707 162507
rect 98913 159523 101897 162507
rect 102103 159523 105087 162507
rect 105293 159523 108277 162507
rect 108483 159523 111467 162507
rect 111673 159523 114657 162507
rect 114863 159523 117847 162507
rect 118053 159523 121037 162507
rect 121243 159523 124227 162507
rect 124433 159523 127417 162507
rect 127623 159523 130607 162507
rect 130813 159523 133797 162507
rect 134003 159523 136987 162507
rect 23 156333 3007 159317
rect 3213 156333 6197 159317
rect 6403 156333 9387 159317
rect 9593 156333 12577 159317
rect 12783 156333 15767 159317
rect 15973 156333 18957 159317
rect 19163 156333 22147 159317
rect 22353 156333 25337 159317
rect 25543 156333 28527 159317
rect 28733 156333 31717 159317
rect 31923 156333 34907 159317
rect 35113 156333 38097 159317
rect 38303 156333 41287 159317
rect 41493 156333 44477 159317
rect 44683 156333 47667 159317
rect 47873 156333 50857 159317
rect 51063 156333 54047 159317
rect 54253 156333 57237 159317
rect 57443 156333 60427 159317
rect 60633 156333 63617 159317
rect 63823 156333 66807 159317
rect 67013 156333 69997 159317
rect 70203 156333 73187 159317
rect 73393 156333 76377 159317
rect 76583 156333 79567 159317
rect 79773 156333 82757 159317
rect 82963 156333 85947 159317
rect 86153 156333 89137 159317
rect 89343 156333 92327 159317
rect 92533 156333 95517 159317
rect 95723 156333 98707 159317
rect 98913 156333 101897 159317
rect 102103 156333 105087 159317
rect 105293 156333 108277 159317
rect 108483 156333 111467 159317
rect 111673 156333 114657 159317
rect 114863 156333 117847 159317
rect 118053 156333 121037 159317
rect 121243 156333 124227 159317
rect 124433 156333 127417 159317
rect 127623 156333 130607 159317
rect 130813 156333 133797 159317
rect 134003 156333 136987 159317
rect 23 153143 3007 156127
rect 3213 153143 6197 156127
rect 6403 153143 9387 156127
rect 9593 153143 12577 156127
rect 12783 153143 15767 156127
rect 15973 153143 18957 156127
rect 19163 153143 22147 156127
rect 22353 153143 25337 156127
rect 25543 153143 28527 156127
rect 28733 153143 31717 156127
rect 31923 153143 34907 156127
rect 35113 153143 38097 156127
rect 38303 153143 41287 156127
rect 41493 153143 44477 156127
rect 44683 153143 47667 156127
rect 47873 153143 50857 156127
rect 51063 153143 54047 156127
rect 54253 153143 57237 156127
rect 57443 153143 60427 156127
rect 60633 153143 63617 156127
rect 63823 153143 66807 156127
rect 67013 153143 69997 156127
rect 70203 153143 73187 156127
rect 73393 153143 76377 156127
rect 76583 153143 79567 156127
rect 79773 153143 82757 156127
rect 82963 153143 85947 156127
rect 86153 153143 89137 156127
rect 89343 153143 92327 156127
rect 92533 153143 95517 156127
rect 95723 153143 98707 156127
rect 98913 153143 101897 156127
rect 102103 153143 105087 156127
rect 105293 153143 108277 156127
rect 108483 153143 111467 156127
rect 111673 153143 114657 156127
rect 114863 153143 117847 156127
rect 118053 153143 121037 156127
rect 121243 153143 124227 156127
rect 124433 153143 127417 156127
rect 127623 153143 130607 156127
rect 130813 153143 133797 156127
rect 134003 153143 136987 156127
rect 23 149953 3007 152937
rect 3213 149953 6197 152937
rect 6403 149953 9387 152937
rect 9593 149953 12577 152937
rect 12783 149953 15767 152937
rect 15973 149953 18957 152937
rect 19163 149953 22147 152937
rect 22353 149953 25337 152937
rect 25543 149953 28527 152937
rect 28733 149953 31717 152937
rect 31923 149953 34907 152937
rect 35113 149953 38097 152937
rect 38303 149953 41287 152937
rect 41493 149953 44477 152937
rect 44683 149953 47667 152937
rect 47873 149953 50857 152937
rect 51063 149953 54047 152937
rect 54253 149953 57237 152937
rect 57443 149953 60427 152937
rect 60633 149953 63617 152937
rect 63823 149953 66807 152937
rect 67013 149953 69997 152937
rect 70203 149953 73187 152937
rect 73393 149953 76377 152937
rect 76583 149953 79567 152937
rect 79773 149953 82757 152937
rect 82963 149953 85947 152937
rect 86153 149953 89137 152937
rect 89343 149953 92327 152937
rect 92533 149953 95517 152937
rect 95723 149953 98707 152937
rect 98913 149953 101897 152937
rect 102103 149953 105087 152937
rect 105293 149953 108277 152937
rect 108483 149953 111467 152937
rect 111673 149953 114657 152937
rect 114863 149953 117847 152937
rect 118053 149953 121037 152937
rect 121243 149953 124227 152937
rect 124433 149953 127417 152937
rect 127623 149953 130607 152937
rect 130813 149953 133797 152937
rect 134003 149953 136987 152937
rect 23 146763 3007 149747
rect 3213 146763 6197 149747
rect 6403 146763 9387 149747
rect 9593 146763 12577 149747
rect 12783 146763 15767 149747
rect 15973 146763 18957 149747
rect 19163 146763 22147 149747
rect 22353 146763 25337 149747
rect 25543 146763 28527 149747
rect 28733 146763 31717 149747
rect 31923 146763 34907 149747
rect 35113 146763 38097 149747
rect 38303 146763 41287 149747
rect 41493 146763 44477 149747
rect 44683 146763 47667 149747
rect 47873 146763 50857 149747
rect 51063 146763 54047 149747
rect 54253 146763 57237 149747
rect 57443 146763 60427 149747
rect 60633 146763 63617 149747
rect 63823 146763 66807 149747
rect 67013 146763 69997 149747
rect 70203 146763 73187 149747
rect 73393 146763 76377 149747
rect 76583 146763 79567 149747
rect 79773 146763 82757 149747
rect 82963 146763 85947 149747
rect 86153 146763 89137 149747
rect 89343 146763 92327 149747
rect 92533 146763 95517 149747
rect 95723 146763 98707 149747
rect 98913 146763 101897 149747
rect 102103 146763 105087 149747
rect 105293 146763 108277 149747
rect 108483 146763 111467 149747
rect 111673 146763 114657 149747
rect 114863 146763 117847 149747
rect 118053 146763 121037 149747
rect 121243 146763 124227 149747
rect 124433 146763 127417 149747
rect 127623 146763 130607 149747
rect 130813 146763 133797 149747
rect 134003 146763 136987 149747
rect 23 143573 3007 146557
rect 3213 143573 6197 146557
rect 6403 143573 9387 146557
rect 9593 143573 12577 146557
rect 12783 143573 15767 146557
rect 15973 143573 18957 146557
rect 19163 143573 22147 146557
rect 22353 143573 25337 146557
rect 25543 143573 28527 146557
rect 28733 143573 31717 146557
rect 31923 143573 34907 146557
rect 35113 143573 38097 146557
rect 38303 143573 41287 146557
rect 41493 143573 44477 146557
rect 44683 143573 47667 146557
rect 47873 143573 50857 146557
rect 51063 143573 54047 146557
rect 54253 143573 57237 146557
rect 57443 143573 60427 146557
rect 60633 143573 63617 146557
rect 63823 143573 66807 146557
rect 67013 143573 69997 146557
rect 70203 143573 73187 146557
rect 73393 143573 76377 146557
rect 76583 143573 79567 146557
rect 79773 143573 82757 146557
rect 82963 143573 85947 146557
rect 86153 143573 89137 146557
rect 89343 143573 92327 146557
rect 92533 143573 95517 146557
rect 95723 143573 98707 146557
rect 98913 143573 101897 146557
rect 102103 143573 105087 146557
rect 105293 143573 108277 146557
rect 108483 143573 111467 146557
rect 111673 143573 114657 146557
rect 114863 143573 117847 146557
rect 118053 143573 121037 146557
rect 121243 143573 124227 146557
rect 124433 143573 127417 146557
rect 127623 143573 130607 146557
rect 130813 143573 133797 146557
rect 134003 143573 136987 146557
rect 23 140383 3007 143367
rect 3213 140383 6197 143367
rect 6403 140383 9387 143367
rect 9593 140383 12577 143367
rect 12783 140383 15767 143367
rect 15973 140383 18957 143367
rect 19163 140383 22147 143367
rect 22353 140383 25337 143367
rect 25543 140383 28527 143367
rect 28733 140383 31717 143367
rect 31923 140383 34907 143367
rect 35113 140383 38097 143367
rect 38303 140383 41287 143367
rect 41493 140383 44477 143367
rect 44683 140383 47667 143367
rect 47873 140383 50857 143367
rect 51063 140383 54047 143367
rect 54253 140383 57237 143367
rect 57443 140383 60427 143367
rect 60633 140383 63617 143367
rect 63823 140383 66807 143367
rect 67013 140383 69997 143367
rect 70203 140383 73187 143367
rect 73393 140383 76377 143367
rect 76583 140383 79567 143367
rect 79773 140383 82757 143367
rect 82963 140383 85947 143367
rect 86153 140383 89137 143367
rect 89343 140383 92327 143367
rect 92533 140383 95517 143367
rect 95723 140383 98707 143367
rect 98913 140383 101897 143367
rect 102103 140383 105087 143367
rect 105293 140383 108277 143367
rect 108483 140383 111467 143367
rect 111673 140383 114657 143367
rect 114863 140383 117847 143367
rect 118053 140383 121037 143367
rect 121243 140383 124227 143367
rect 124433 140383 127417 143367
rect 127623 140383 130607 143367
rect 130813 140383 133797 143367
rect 134003 140383 136987 143367
rect 9593 137193 12577 140177
rect 12783 137193 15767 140177
rect 15973 137193 18957 140177
rect 19163 137193 22147 140177
rect 22353 137193 25337 140177
rect 25543 137193 28527 140177
rect 28733 137193 31717 140177
rect 31923 137193 34907 140177
rect 35113 137193 38097 140177
rect 38303 137193 41287 140177
rect 41493 137193 44477 140177
rect 44683 137193 47667 140177
rect 47873 137193 50857 140177
rect 51063 137193 54047 140177
rect 54253 137193 57237 140177
rect 57443 137193 60427 140177
rect 60633 137193 63617 140177
rect 63823 137193 66807 140177
rect 67013 137193 69997 140177
rect 70203 137193 73187 140177
rect 73393 137193 76377 140177
rect 76583 137193 79567 140177
rect 79773 137193 82757 140177
rect 82963 137193 85947 140177
rect 86153 137193 89137 140177
rect 89343 137193 92327 140177
rect 92533 137193 95517 140177
rect 95723 137193 98707 140177
rect 98913 137193 101897 140177
rect 102103 137193 105087 140177
rect 105293 137193 108277 140177
rect 108483 137193 111467 140177
rect 111673 137193 114657 140177
rect 114863 137193 117847 140177
rect 118053 137193 121037 140177
rect 121243 137193 124227 140177
rect 124433 137193 127417 140177
rect 127623 137193 130607 140177
rect 130813 137193 133797 140177
rect 134003 137193 136987 140177
rect 9593 134003 12577 136987
rect 12783 134003 15767 136987
rect 15973 134003 18957 136987
rect 19163 134003 22147 136987
rect 22353 134003 25337 136987
rect 25543 134003 28527 136987
rect 28733 134003 31717 136987
rect 31923 134003 34907 136987
rect 35113 134003 38097 136987
rect 38303 134003 41287 136987
rect 41493 134003 44477 136987
rect 44683 134003 47667 136987
rect 47873 134003 50857 136987
rect 51063 134003 54047 136987
rect 54253 134003 57237 136987
rect 57443 134003 60427 136987
rect 60633 134003 63617 136987
rect 63823 134003 66807 136987
rect 67013 134003 69997 136987
rect 70203 134003 73187 136987
rect 73393 134003 76377 136987
rect 76583 134003 79567 136987
rect 79773 134003 82757 136987
rect 82963 134003 85947 136987
rect 86153 134003 89137 136987
rect 89343 134003 92327 136987
rect 92533 134003 95517 136987
rect 95723 134003 98707 136987
rect 98913 134003 101897 136987
rect 102103 134003 105087 136987
rect 105293 134003 108277 136987
rect 108483 134003 111467 136987
rect 111673 134003 114657 136987
rect 114863 134003 117847 136987
rect 118053 134003 121037 136987
rect 121243 134003 124227 136987
rect 124433 134003 127417 136987
rect 127623 134003 130607 136987
rect 130813 134003 133797 136987
rect 134003 134003 136987 136987
rect 9593 130813 12577 133797
rect 12783 130813 15767 133797
rect 15973 130813 18957 133797
rect 19163 130813 22147 133797
rect 22353 130813 25337 133797
rect 25543 130813 28527 133797
rect 28733 130813 31717 133797
rect 31923 130813 34907 133797
rect 35113 130813 38097 133797
rect 38303 130813 41287 133797
rect 41493 130813 44477 133797
rect 44683 130813 47667 133797
rect 47873 130813 50857 133797
rect 51063 130813 54047 133797
rect 54253 130813 57237 133797
rect 57443 130813 60427 133797
rect 60633 130813 63617 133797
rect 63823 130813 66807 133797
rect 67013 130813 69997 133797
rect 70203 130813 73187 133797
rect 73393 130813 76377 133797
rect 76583 130813 79567 133797
rect 79773 130813 82757 133797
rect 82963 130813 85947 133797
rect 86153 130813 89137 133797
rect 89343 130813 92327 133797
rect 92533 130813 95517 133797
rect 95723 130813 98707 133797
rect 98913 130813 101897 133797
rect 102103 130813 105087 133797
rect 105293 130813 108277 133797
rect 108483 130813 111467 133797
rect 111673 130813 114657 133797
rect 114863 130813 117847 133797
rect 118053 130813 121037 133797
rect 121243 130813 124227 133797
rect 124433 130813 127417 133797
rect 127623 130813 130607 133797
rect 130813 130813 133797 133797
rect 134003 130813 136987 133797
rect 9593 127623 12577 130607
rect 12783 127623 15767 130607
rect 15973 127623 18957 130607
rect 19163 127623 22147 130607
rect 22353 127623 25337 130607
rect 25543 127623 28527 130607
rect 28733 127623 31717 130607
rect 31923 127623 34907 130607
rect 35113 127623 38097 130607
rect 38303 127623 41287 130607
rect 41493 127623 44477 130607
rect 44683 127623 47667 130607
rect 47873 127623 50857 130607
rect 51063 127623 54047 130607
rect 54253 127623 57237 130607
rect 57443 127623 60427 130607
rect 60633 127623 63617 130607
rect 63823 127623 66807 130607
rect 67013 127623 69997 130607
rect 70203 127623 73187 130607
rect 73393 127623 76377 130607
rect 76583 127623 79567 130607
rect 79773 127623 82757 130607
rect 82963 127623 85947 130607
rect 86153 127623 89137 130607
rect 89343 127623 92327 130607
rect 92533 127623 95517 130607
rect 95723 127623 98707 130607
rect 98913 127623 101897 130607
rect 102103 127623 105087 130607
rect 105293 127623 108277 130607
rect 108483 127623 111467 130607
rect 111673 127623 114657 130607
rect 114863 127623 117847 130607
rect 118053 127623 121037 130607
rect 121243 127623 124227 130607
rect 124433 127623 127417 130607
rect 127623 127623 130607 130607
rect 130813 127623 133797 130607
rect 134003 127623 136987 130607
rect 9593 124433 12577 127417
rect 12783 124433 15767 127417
rect 15973 124433 18957 127417
rect 19163 124433 22147 127417
rect 22353 124433 25337 127417
rect 25543 124433 28527 127417
rect 28733 124433 31717 127417
rect 31923 124433 34907 127417
rect 35113 124433 38097 127417
rect 38303 124433 41287 127417
rect 41493 124433 44477 127417
rect 44683 124433 47667 127417
rect 47873 124433 50857 127417
rect 51063 124433 54047 127417
rect 54253 124433 57237 127417
rect 57443 124433 60427 127417
rect 60633 124433 63617 127417
rect 63823 124433 66807 127417
rect 67013 124433 69997 127417
rect 70203 124433 73187 127417
rect 73393 124433 76377 127417
rect 76583 124433 79567 127417
rect 79773 124433 82757 127417
rect 82963 124433 85947 127417
rect 86153 124433 89137 127417
rect 89343 124433 92327 127417
rect 92533 124433 95517 127417
rect 95723 124433 98707 127417
rect 98913 124433 101897 127417
rect 102103 124433 105087 127417
rect 105293 124433 108277 127417
rect 108483 124433 111467 127417
rect 111673 124433 114657 127417
rect 114863 124433 117847 127417
rect 118053 124433 121037 127417
rect 121243 124433 124227 127417
rect 124433 124433 127417 127417
rect 127623 124433 130607 127417
rect 130813 124433 133797 127417
rect 134003 124433 136987 127417
rect 9593 121243 12577 124227
rect 12783 121243 15767 124227
rect 15973 121243 18957 124227
rect 19163 121243 22147 124227
rect 22353 121243 25337 124227
rect 25543 121243 28527 124227
rect 28733 121243 31717 124227
rect 31923 121243 34907 124227
rect 35113 121243 38097 124227
rect 38303 121243 41287 124227
rect 41493 121243 44477 124227
rect 44683 121243 47667 124227
rect 47873 121243 50857 124227
rect 51063 121243 54047 124227
rect 54253 121243 57237 124227
rect 57443 121243 60427 124227
rect 60633 121243 63617 124227
rect 63823 121243 66807 124227
rect 67013 121243 69997 124227
rect 70203 121243 73187 124227
rect 73393 121243 76377 124227
rect 76583 121243 79567 124227
rect 79773 121243 82757 124227
rect 82963 121243 85947 124227
rect 86153 121243 89137 124227
rect 89343 121243 92327 124227
rect 92533 121243 95517 124227
rect 95723 121243 98707 124227
rect 98913 121243 101897 124227
rect 102103 121243 105087 124227
rect 105293 121243 108277 124227
rect 108483 121243 111467 124227
rect 111673 121243 114657 124227
rect 114863 121243 117847 124227
rect 118053 121243 121037 124227
rect 121243 121243 124227 124227
rect 124433 121243 127417 124227
rect 127623 121243 130607 124227
rect 130813 121243 133797 124227
rect 134003 121243 136987 124227
rect 23 118053 3007 121037
rect 3213 118053 6197 121037
rect 6403 118053 9387 121037
rect 9593 118053 12577 121037
rect 12783 118053 15767 121037
rect 15973 118053 18957 121037
rect 19163 118053 22147 121037
rect 22353 118053 25337 121037
rect 25543 118053 28527 121037
rect 28733 118053 31717 121037
rect 31923 118053 34907 121037
rect 35113 118053 38097 121037
rect 38303 118053 41287 121037
rect 41493 118053 44477 121037
rect 44683 118053 47667 121037
rect 47873 118053 50857 121037
rect 51063 118053 54047 121037
rect 54253 118053 57237 121037
rect 57443 118053 60427 121037
rect 60633 118053 63617 121037
rect 63823 118053 66807 121037
rect 67013 118053 69997 121037
rect 70203 118053 73187 121037
rect 73393 118053 76377 121037
rect 76583 118053 79567 121037
rect 79773 118053 82757 121037
rect 82963 118053 85947 121037
rect 86153 118053 89137 121037
rect 89343 118053 92327 121037
rect 92533 118053 95517 121037
rect 95723 118053 98707 121037
rect 98913 118053 101897 121037
rect 102103 118053 105087 121037
rect 105293 118053 108277 121037
rect 108483 118053 111467 121037
rect 111673 118053 114657 121037
rect 114863 118053 117847 121037
rect 118053 118053 121037 121037
rect 121243 118053 124227 121037
rect 124433 118053 127417 121037
rect 127623 118053 130607 121037
rect 130813 118053 133797 121037
rect 134003 118053 136987 121037
rect 23 114863 3007 117847
rect 3213 114863 6197 117847
rect 6403 114863 9387 117847
rect 9593 114863 12577 117847
rect 12783 114863 15767 117847
rect 15973 114863 18957 117847
rect 19163 114863 22147 117847
rect 22353 114863 25337 117847
rect 25543 114863 28527 117847
rect 28733 114863 31717 117847
rect 31923 114863 34907 117847
rect 35113 114863 38097 117847
rect 38303 114863 41287 117847
rect 41493 114863 44477 117847
rect 44683 114863 47667 117847
rect 47873 114863 50857 117847
rect 51063 114863 54047 117847
rect 54253 114863 57237 117847
rect 57443 114863 60427 117847
rect 60633 114863 63617 117847
rect 63823 114863 66807 117847
rect 67013 114863 69997 117847
rect 70203 114863 73187 117847
rect 73393 114863 76377 117847
rect 76583 114863 79567 117847
rect 79773 114863 82757 117847
rect 82963 114863 85947 117847
rect 86153 114863 89137 117847
rect 89343 114863 92327 117847
rect 92533 114863 95517 117847
rect 95723 114863 98707 117847
rect 98913 114863 101897 117847
rect 102103 114863 105087 117847
rect 105293 114863 108277 117847
rect 108483 114863 111467 117847
rect 111673 114863 114657 117847
rect 114863 114863 117847 117847
rect 118053 114863 121037 117847
rect 121243 114863 124227 117847
rect 124433 114863 127417 117847
rect 127623 114863 130607 117847
rect 130813 114863 133797 117847
rect 134003 114863 136987 117847
rect 23 111673 3007 114657
rect 3213 111673 6197 114657
rect 6403 111673 9387 114657
rect 9593 111673 12577 114657
rect 12783 111673 15767 114657
rect 15973 111673 18957 114657
rect 19163 111673 22147 114657
rect 22353 111673 25337 114657
rect 25543 111673 28527 114657
rect 28733 111673 31717 114657
rect 31923 111673 34907 114657
rect 35113 111673 38097 114657
rect 38303 111673 41287 114657
rect 41493 111673 44477 114657
rect 44683 111673 47667 114657
rect 47873 111673 50857 114657
rect 51063 111673 54047 114657
rect 54253 111673 57237 114657
rect 57443 111673 60427 114657
rect 60633 111673 63617 114657
rect 63823 111673 66807 114657
rect 67013 111673 69997 114657
rect 70203 111673 73187 114657
rect 73393 111673 76377 114657
rect 76583 111673 79567 114657
rect 79773 111673 82757 114657
rect 82963 111673 85947 114657
rect 86153 111673 89137 114657
rect 89343 111673 92327 114657
rect 92533 111673 95517 114657
rect 95723 111673 98707 114657
rect 98913 111673 101897 114657
rect 102103 111673 105087 114657
rect 105293 111673 108277 114657
rect 108483 111673 111467 114657
rect 111673 111673 114657 114657
rect 114863 111673 117847 114657
rect 118053 111673 121037 114657
rect 121243 111673 124227 114657
rect 124433 111673 127417 114657
rect 127623 111673 130607 114657
rect 130813 111673 133797 114657
rect 134003 111673 136987 114657
rect 23 108483 3007 111467
rect 3213 108483 6197 111467
rect 6403 108483 9387 111467
rect 9593 108483 12577 111467
rect 12783 108483 15767 111467
rect 15973 108483 18957 111467
rect 19163 108483 22147 111467
rect 22353 108483 25337 111467
rect 25543 108483 28527 111467
rect 28733 108483 31717 111467
rect 31923 108483 34907 111467
rect 35113 108483 38097 111467
rect 38303 108483 41287 111467
rect 41493 108483 44477 111467
rect 44683 108483 47667 111467
rect 47873 108483 50857 111467
rect 51063 108483 54047 111467
rect 54253 108483 57237 111467
rect 57443 108483 60427 111467
rect 60633 108483 63617 111467
rect 63823 108483 66807 111467
rect 67013 108483 69997 111467
rect 70203 108483 73187 111467
rect 73393 108483 76377 111467
rect 76583 108483 79567 111467
rect 79773 108483 82757 111467
rect 82963 108483 85947 111467
rect 86153 108483 89137 111467
rect 89343 108483 92327 111467
rect 92533 108483 95517 111467
rect 95723 108483 98707 111467
rect 98913 108483 101897 111467
rect 102103 108483 105087 111467
rect 105293 108483 108277 111467
rect 108483 108483 111467 111467
rect 111673 108483 114657 111467
rect 114863 108483 117847 111467
rect 118053 108483 121037 111467
rect 121243 108483 124227 111467
rect 124433 108483 127417 111467
rect 127623 108483 130607 111467
rect 130813 108483 133797 111467
rect 134003 108483 136987 111467
rect 23 105293 3007 108277
rect 3213 105293 6197 108277
rect 6403 105293 9387 108277
rect 9593 105293 12577 108277
rect 12783 105293 15767 108277
rect 15973 105293 18957 108277
rect 19163 105293 22147 108277
rect 22353 105293 25337 108277
rect 25543 105293 28527 108277
rect 28733 105293 31717 108277
rect 31923 105293 34907 108277
rect 35113 105293 38097 108277
rect 38303 105293 41287 108277
rect 41493 105293 44477 108277
rect 44683 105293 47667 108277
rect 47873 105293 50857 108277
rect 51063 105293 54047 108277
rect 54253 105293 57237 108277
rect 57443 105293 60427 108277
rect 60633 105293 63617 108277
rect 63823 105293 66807 108277
rect 67013 105293 69997 108277
rect 70203 105293 73187 108277
rect 73393 105293 76377 108277
rect 76583 105293 79567 108277
rect 79773 105293 82757 108277
rect 82963 105293 85947 108277
rect 86153 105293 89137 108277
rect 89343 105293 92327 108277
rect 92533 105293 95517 108277
rect 95723 105293 98707 108277
rect 98913 105293 101897 108277
rect 102103 105293 105087 108277
rect 105293 105293 108277 108277
rect 108483 105293 111467 108277
rect 111673 105293 114657 108277
rect 114863 105293 117847 108277
rect 118053 105293 121037 108277
rect 121243 105293 124227 108277
rect 124433 105293 127417 108277
rect 127623 105293 130607 108277
rect 130813 105293 133797 108277
rect 134003 105293 136987 108277
rect 23 102103 3007 105087
rect 3213 102103 6197 105087
rect 6403 102103 9387 105087
rect 9593 102103 12577 105087
rect 12783 102103 15767 105087
rect 15973 102103 18957 105087
rect 19163 102103 22147 105087
rect 22353 102103 25337 105087
rect 25543 102103 28527 105087
rect 28733 102103 31717 105087
rect 31923 102103 34907 105087
rect 35113 102103 38097 105087
rect 38303 102103 41287 105087
rect 41493 102103 44477 105087
rect 44683 102103 47667 105087
rect 47873 102103 50857 105087
rect 51063 102103 54047 105087
rect 54253 102103 57237 105087
rect 57443 102103 60427 105087
rect 60633 102103 63617 105087
rect 63823 102103 66807 105087
rect 67013 102103 69997 105087
rect 70203 102103 73187 105087
rect 73393 102103 76377 105087
rect 76583 102103 79567 105087
rect 79773 102103 82757 105087
rect 82963 102103 85947 105087
rect 86153 102103 89137 105087
rect 89343 102103 92327 105087
rect 92533 102103 95517 105087
rect 95723 102103 98707 105087
rect 98913 102103 101897 105087
rect 102103 102103 105087 105087
rect 105293 102103 108277 105087
rect 108483 102103 111467 105087
rect 111673 102103 114657 105087
rect 114863 102103 117847 105087
rect 118053 102103 121037 105087
rect 121243 102103 124227 105087
rect 124433 102103 127417 105087
rect 127623 102103 130607 105087
rect 130813 102103 133797 105087
rect 134003 102103 136987 105087
rect 23 98913 3007 101897
rect 3213 98913 6197 101897
rect 6403 98913 9387 101897
rect 9593 98913 12577 101897
rect 12783 98913 15767 101897
rect 15973 98913 18957 101897
rect 19163 98913 22147 101897
rect 22353 98913 25337 101897
rect 25543 98913 28527 101897
rect 28733 98913 31717 101897
rect 31923 98913 34907 101897
rect 35113 98913 38097 101897
rect 38303 98913 41287 101897
rect 41493 98913 44477 101897
rect 44683 98913 47667 101897
rect 47873 98913 50857 101897
rect 51063 98913 54047 101897
rect 54253 98913 57237 101897
rect 57443 98913 60427 101897
rect 60633 98913 63617 101897
rect 63823 98913 66807 101897
rect 67013 98913 69997 101897
rect 70203 98913 73187 101897
rect 73393 98913 76377 101897
rect 76583 98913 79567 101897
rect 79773 98913 82757 101897
rect 82963 98913 85947 101897
rect 86153 98913 89137 101897
rect 89343 98913 92327 101897
rect 92533 98913 95517 101897
rect 95723 98913 98707 101897
rect 98913 98913 101897 101897
rect 102103 98913 105087 101897
rect 105293 98913 108277 101897
rect 108483 98913 111467 101897
rect 111673 98913 114657 101897
rect 114863 98913 117847 101897
rect 118053 98913 121037 101897
rect 121243 98913 124227 101897
rect 124433 98913 127417 101897
rect 127623 98913 130607 101897
rect 130813 98913 133797 101897
rect 134003 98913 136987 101897
rect 9593 95723 12577 98707
rect 12783 95723 15767 98707
rect 15973 95723 18957 98707
rect 19163 95723 22147 98707
rect 22353 95723 25337 98707
rect 25543 95723 28527 98707
rect 28733 95723 31717 98707
rect 31923 95723 34907 98707
rect 35113 95723 38097 98707
rect 38303 95723 41287 98707
rect 41493 95723 44477 98707
rect 44683 95723 47667 98707
rect 47873 95723 50857 98707
rect 51063 95723 54047 98707
rect 54253 95723 57237 98707
rect 57443 95723 60427 98707
rect 60633 95723 63617 98707
rect 63823 95723 66807 98707
rect 67013 95723 69997 98707
rect 70203 95723 73187 98707
rect 73393 95723 76377 98707
rect 76583 95723 79567 98707
rect 79773 95723 82757 98707
rect 82963 95723 85947 98707
rect 86153 95723 89137 98707
rect 89343 95723 92327 98707
rect 92533 95723 95517 98707
rect 95723 95723 98707 98707
rect 98913 95723 101897 98707
rect 102103 95723 105087 98707
rect 105293 95723 108277 98707
rect 108483 95723 111467 98707
rect 111673 95723 114657 98707
rect 114863 95723 117847 98707
rect 118053 95723 121037 98707
rect 121243 95723 124227 98707
rect 124433 95723 127417 98707
rect 127623 95723 130607 98707
rect 130813 95723 133797 98707
rect 134003 95723 136987 98707
rect 9593 92533 12577 95517
rect 12783 92533 15767 95517
rect 15973 92533 18957 95517
rect 19163 92533 22147 95517
rect 22353 92533 25337 95517
rect 25543 92533 28527 95517
rect 28733 92533 31717 95517
rect 31923 92533 34907 95517
rect 35113 92533 38097 95517
rect 38303 92533 41287 95517
rect 41493 92533 44477 95517
rect 44683 92533 47667 95517
rect 47873 92533 50857 95517
rect 51063 92533 54047 95517
rect 54253 92533 57237 95517
rect 57443 92533 60427 95517
rect 60633 92533 63617 95517
rect 63823 92533 66807 95517
rect 67013 92533 69997 95517
rect 70203 92533 73187 95517
rect 73393 92533 76377 95517
rect 76583 92533 79567 95517
rect 79773 92533 82757 95517
rect 82963 92533 85947 95517
rect 86153 92533 89137 95517
rect 89343 92533 92327 95517
rect 92533 92533 95517 95517
rect 95723 92533 98707 95517
rect 98913 92533 101897 95517
rect 102103 92533 105087 95517
rect 105293 92533 108277 95517
rect 108483 92533 111467 95517
rect 111673 92533 114657 95517
rect 114863 92533 117847 95517
rect 118053 92533 121037 95517
rect 121243 92533 124227 95517
rect 124433 92533 127417 95517
rect 127623 92533 130607 95517
rect 130813 92533 133797 95517
rect 134003 92533 136987 95517
rect 9593 89343 12577 92327
rect 12783 89343 15767 92327
rect 15973 89343 18957 92327
rect 19163 89343 22147 92327
rect 22353 89343 25337 92327
rect 25543 89343 28527 92327
rect 28733 89343 31717 92327
rect 31923 89343 34907 92327
rect 35113 89343 38097 92327
rect 38303 89343 41287 92327
rect 41493 89343 44477 92327
rect 44683 89343 47667 92327
rect 47873 89343 50857 92327
rect 51063 89343 54047 92327
rect 54253 89343 57237 92327
rect 57443 89343 60427 92327
rect 60633 89343 63617 92327
rect 63823 89343 66807 92327
rect 67013 89343 69997 92327
rect 70203 89343 73187 92327
rect 73393 89343 76377 92327
rect 76583 89343 79567 92327
rect 79773 89343 82757 92327
rect 82963 89343 85947 92327
rect 86153 89343 89137 92327
rect 89343 89343 92327 92327
rect 92533 89343 95517 92327
rect 95723 89343 98707 92327
rect 98913 89343 101897 92327
rect 102103 89343 105087 92327
rect 105293 89343 108277 92327
rect 108483 89343 111467 92327
rect 111673 89343 114657 92327
rect 114863 89343 117847 92327
rect 118053 89343 121037 92327
rect 121243 89343 124227 92327
rect 124433 89343 127417 92327
rect 127623 89343 130607 92327
rect 130813 89343 133797 92327
rect 134003 89343 136987 92327
rect 9593 86153 12577 89137
rect 12783 86153 15767 89137
rect 15973 86153 18957 89137
rect 19163 86153 22147 89137
rect 22353 86153 25337 89137
rect 25543 86153 28527 89137
rect 28733 86153 31717 89137
rect 31923 86153 34907 89137
rect 35113 86153 38097 89137
rect 38303 86153 41287 89137
rect 41493 86153 44477 89137
rect 44683 86153 47667 89137
rect 47873 86153 50857 89137
rect 51063 86153 54047 89137
rect 54253 86153 57237 89137
rect 57443 86153 60427 89137
rect 60633 86153 63617 89137
rect 63823 86153 66807 89137
rect 67013 86153 69997 89137
rect 70203 86153 73187 89137
rect 73393 86153 76377 89137
rect 76583 86153 79567 89137
rect 79773 86153 82757 89137
rect 82963 86153 85947 89137
rect 86153 86153 89137 89137
rect 89343 86153 92327 89137
rect 92533 86153 95517 89137
rect 95723 86153 98707 89137
rect 98913 86153 101897 89137
rect 102103 86153 105087 89137
rect 105293 86153 108277 89137
rect 108483 86153 111467 89137
rect 111673 86153 114657 89137
rect 114863 86153 117847 89137
rect 118053 86153 121037 89137
rect 121243 86153 124227 89137
rect 124433 86153 127417 89137
rect 127623 86153 130607 89137
rect 130813 86153 133797 89137
rect 134003 86153 136987 89137
rect 9593 82963 12577 85947
rect 12783 82963 15767 85947
rect 15973 82963 18957 85947
rect 19163 82963 22147 85947
rect 22353 82963 25337 85947
rect 25543 82963 28527 85947
rect 28733 82963 31717 85947
rect 31923 82963 34907 85947
rect 35113 82963 38097 85947
rect 38303 82963 41287 85947
rect 41493 82963 44477 85947
rect 44683 82963 47667 85947
rect 47873 82963 50857 85947
rect 51063 82963 54047 85947
rect 54253 82963 57237 85947
rect 57443 82963 60427 85947
rect 60633 82963 63617 85947
rect 63823 82963 66807 85947
rect 67013 82963 69997 85947
rect 70203 82963 73187 85947
rect 73393 82963 76377 85947
rect 76583 82963 79567 85947
rect 79773 82963 82757 85947
rect 82963 82963 85947 85947
rect 86153 82963 89137 85947
rect 89343 82963 92327 85947
rect 92533 82963 95517 85947
rect 95723 82963 98707 85947
rect 98913 82963 101897 85947
rect 102103 82963 105087 85947
rect 105293 82963 108277 85947
rect 108483 82963 111467 85947
rect 111673 82963 114657 85947
rect 114863 82963 117847 85947
rect 118053 82963 121037 85947
rect 121243 82963 124227 85947
rect 124433 82963 127417 85947
rect 127623 82963 130607 85947
rect 130813 82963 133797 85947
rect 134003 82963 136987 85947
rect 9593 79773 12577 82757
rect 12783 79773 15767 82757
rect 15973 79773 18957 82757
rect 19163 79773 22147 82757
rect 22353 79773 25337 82757
rect 25543 79773 28527 82757
rect 28733 79773 31717 82757
rect 31923 79773 34907 82757
rect 35113 79773 38097 82757
rect 38303 79773 41287 82757
rect 41493 79773 44477 82757
rect 44683 79773 47667 82757
rect 47873 79773 50857 82757
rect 51063 79773 54047 82757
rect 54253 79773 57237 82757
rect 57443 79773 60427 82757
rect 60633 79773 63617 82757
rect 63823 79773 66807 82757
rect 67013 79773 69997 82757
rect 70203 79773 73187 82757
rect 73393 79773 76377 82757
rect 76583 79773 79567 82757
rect 79773 79773 82757 82757
rect 82963 79773 85947 82757
rect 86153 79773 89137 82757
rect 89343 79773 92327 82757
rect 92533 79773 95517 82757
rect 95723 79773 98707 82757
rect 98913 79773 101897 82757
rect 102103 79773 105087 82757
rect 105293 79773 108277 82757
rect 108483 79773 111467 82757
rect 111673 79773 114657 82757
rect 114863 79773 117847 82757
rect 118053 79773 121037 82757
rect 121243 79773 124227 82757
rect 124433 79773 127417 82757
rect 127623 79773 130607 82757
rect 130813 79773 133797 82757
rect 134003 79773 136987 82757
rect 23 76583 3007 79567
rect 3213 76583 6197 79567
rect 6403 76583 9387 79567
rect 9593 76583 12577 79567
rect 12783 76583 15767 79567
rect 15973 76583 18957 79567
rect 19163 76583 22147 79567
rect 22353 76583 25337 79567
rect 25543 76583 28527 79567
rect 28733 76583 31717 79567
rect 31923 76583 34907 79567
rect 35113 76583 38097 79567
rect 38303 76583 41287 79567
rect 41493 76583 44477 79567
rect 44683 76583 47667 79567
rect 47873 76583 50857 79567
rect 51063 76583 54047 79567
rect 54253 76583 57237 79567
rect 57443 76583 60427 79567
rect 60633 76583 63617 79567
rect 63823 76583 66807 79567
rect 67013 76583 69997 79567
rect 70203 76583 73187 79567
rect 73393 76583 76377 79567
rect 76583 76583 79567 79567
rect 79773 76583 82757 79567
rect 82963 76583 85947 79567
rect 86153 76583 89137 79567
rect 89343 76583 92327 79567
rect 92533 76583 95517 79567
rect 95723 76583 98707 79567
rect 98913 76583 101897 79567
rect 102103 76583 105087 79567
rect 105293 76583 108277 79567
rect 108483 76583 111467 79567
rect 111673 76583 114657 79567
rect 114863 76583 117847 79567
rect 118053 76583 121037 79567
rect 121243 76583 124227 79567
rect 124433 76583 127417 79567
rect 127623 76583 130607 79567
rect 130813 76583 133797 79567
rect 134003 76583 136987 79567
rect 23 73393 3007 76377
rect 3213 73393 6197 76377
rect 6403 73393 9387 76377
rect 9593 73393 12577 76377
rect 12783 73393 15767 76377
rect 15973 73393 18957 76377
rect 19163 73393 22147 76377
rect 22353 73393 25337 76377
rect 25543 73393 28527 76377
rect 28733 73393 31717 76377
rect 31923 73393 34907 76377
rect 35113 73393 38097 76377
rect 38303 73393 41287 76377
rect 41493 73393 44477 76377
rect 44683 73393 47667 76377
rect 47873 73393 50857 76377
rect 51063 73393 54047 76377
rect 54253 73393 57237 76377
rect 57443 73393 60427 76377
rect 60633 73393 63617 76377
rect 63823 73393 66807 76377
rect 67013 73393 69997 76377
rect 70203 73393 73187 76377
rect 73393 73393 76377 76377
rect 76583 73393 79567 76377
rect 79773 73393 82757 76377
rect 82963 73393 85947 76377
rect 86153 73393 89137 76377
rect 89343 73393 92327 76377
rect 92533 73393 95517 76377
rect 95723 73393 98707 76377
rect 98913 73393 101897 76377
rect 102103 73393 105087 76377
rect 105293 73393 108277 76377
rect 108483 73393 111467 76377
rect 111673 73393 114657 76377
rect 114863 73393 117847 76377
rect 118053 73393 121037 76377
rect 121243 73393 124227 76377
rect 124433 73393 127417 76377
rect 127623 73393 130607 76377
rect 130813 73393 133797 76377
rect 134003 73393 136987 76377
rect 23 70203 3007 73187
rect 3213 70203 6197 73187
rect 6403 70203 9387 73187
rect 9593 70203 12577 73187
rect 12783 70203 15767 73187
rect 15973 70203 18957 73187
rect 19163 70203 22147 73187
rect 22353 70203 25337 73187
rect 25543 70203 28527 73187
rect 28733 70203 31717 73187
rect 31923 70203 34907 73187
rect 35113 70203 38097 73187
rect 38303 70203 41287 73187
rect 41493 70203 44477 73187
rect 44683 70203 47667 73187
rect 47873 70203 50857 73187
rect 51063 70203 54047 73187
rect 54253 70203 57237 73187
rect 57443 70203 60427 73187
rect 60633 70203 63617 73187
rect 63823 70203 66807 73187
rect 67013 70203 69997 73187
rect 70203 70203 73187 73187
rect 73393 70203 76377 73187
rect 76583 70203 79567 73187
rect 79773 70203 82757 73187
rect 82963 70203 85947 73187
rect 86153 70203 89137 73187
rect 89343 70203 92327 73187
rect 92533 70203 95517 73187
rect 95723 70203 98707 73187
rect 98913 70203 101897 73187
rect 102103 70203 105087 73187
rect 105293 70203 108277 73187
rect 108483 70203 111467 73187
rect 111673 70203 114657 73187
rect 114863 70203 117847 73187
rect 118053 70203 121037 73187
rect 121243 70203 124227 73187
rect 124433 70203 127417 73187
rect 127623 70203 130607 73187
rect 130813 70203 133797 73187
rect 134003 70203 136987 73187
rect 23 67013 3007 69997
rect 3213 67013 6197 69997
rect 6403 67013 9387 69997
rect 9593 67013 12577 69997
rect 12783 67013 15767 69997
rect 15973 67013 18957 69997
rect 19163 67013 22147 69997
rect 22353 67013 25337 69997
rect 25543 67013 28527 69997
rect 28733 67013 31717 69997
rect 31923 67013 34907 69997
rect 35113 67013 38097 69997
rect 38303 67013 41287 69997
rect 41493 67013 44477 69997
rect 44683 67013 47667 69997
rect 47873 67013 50857 69997
rect 51063 67013 54047 69997
rect 54253 67013 57237 69997
rect 57443 67013 60427 69997
rect 60633 67013 63617 69997
rect 63823 67013 66807 69997
rect 67013 67013 69997 69997
rect 70203 67013 73187 69997
rect 73393 67013 76377 69997
rect 76583 67013 79567 69997
rect 79773 67013 82757 69997
rect 82963 67013 85947 69997
rect 86153 67013 89137 69997
rect 89343 67013 92327 69997
rect 92533 67013 95517 69997
rect 95723 67013 98707 69997
rect 98913 67013 101897 69997
rect 102103 67013 105087 69997
rect 105293 67013 108277 69997
rect 108483 67013 111467 69997
rect 111673 67013 114657 69997
rect 114863 67013 117847 69997
rect 118053 67013 121037 69997
rect 121243 67013 124227 69997
rect 124433 67013 127417 69997
rect 127623 67013 130607 69997
rect 130813 67013 133797 69997
rect 134003 67013 136987 69997
rect 23 63823 3007 66807
rect 3213 63823 6197 66807
rect 6403 63823 9387 66807
rect 9593 63823 12577 66807
rect 12783 63823 15767 66807
rect 15973 63823 18957 66807
rect 19163 63823 22147 66807
rect 22353 63823 25337 66807
rect 25543 63823 28527 66807
rect 28733 63823 31717 66807
rect 31923 63823 34907 66807
rect 35113 63823 38097 66807
rect 38303 63823 41287 66807
rect 41493 63823 44477 66807
rect 44683 63823 47667 66807
rect 47873 63823 50857 66807
rect 51063 63823 54047 66807
rect 54253 63823 57237 66807
rect 57443 63823 60427 66807
rect 60633 63823 63617 66807
rect 63823 63823 66807 66807
rect 67013 63823 69997 66807
rect 70203 63823 73187 66807
rect 73393 63823 76377 66807
rect 76583 63823 79567 66807
rect 79773 63823 82757 66807
rect 82963 63823 85947 66807
rect 86153 63823 89137 66807
rect 89343 63823 92327 66807
rect 92533 63823 95517 66807
rect 95723 63823 98707 66807
rect 98913 63823 101897 66807
rect 102103 63823 105087 66807
rect 105293 63823 108277 66807
rect 108483 63823 111467 66807
rect 111673 63823 114657 66807
rect 114863 63823 117847 66807
rect 118053 63823 121037 66807
rect 121243 63823 124227 66807
rect 124433 63823 127417 66807
rect 127623 63823 130607 66807
rect 130813 63823 133797 66807
rect 134003 63823 136987 66807
rect 23 60633 3007 63617
rect 3213 60633 6197 63617
rect 6403 60633 9387 63617
rect 9593 60633 12577 63617
rect 12783 60633 15767 63617
rect 15973 60633 18957 63617
rect 19163 60633 22147 63617
rect 22353 60633 25337 63617
rect 25543 60633 28527 63617
rect 28733 60633 31717 63617
rect 31923 60633 34907 63617
rect 35113 60633 38097 63617
rect 38303 60633 41287 63617
rect 41493 60633 44477 63617
rect 44683 60633 47667 63617
rect 47873 60633 50857 63617
rect 51063 60633 54047 63617
rect 54253 60633 57237 63617
rect 57443 60633 60427 63617
rect 60633 60633 63617 63617
rect 63823 60633 66807 63617
rect 67013 60633 69997 63617
rect 70203 60633 73187 63617
rect 73393 60633 76377 63617
rect 76583 60633 79567 63617
rect 79773 60633 82757 63617
rect 82963 60633 85947 63617
rect 86153 60633 89137 63617
rect 89343 60633 92327 63617
rect 92533 60633 95517 63617
rect 95723 60633 98707 63617
rect 98913 60633 101897 63617
rect 102103 60633 105087 63617
rect 105293 60633 108277 63617
rect 108483 60633 111467 63617
rect 111673 60633 114657 63617
rect 114863 60633 117847 63617
rect 118053 60633 121037 63617
rect 121243 60633 124227 63617
rect 124433 60633 127417 63617
rect 127623 60633 130607 63617
rect 130813 60633 133797 63617
rect 134003 60633 136987 63617
rect 23 57443 3007 60427
rect 3213 57443 6197 60427
rect 6403 57443 9387 60427
rect 9593 57443 12577 60427
rect 12783 57443 15767 60427
rect 15973 57443 18957 60427
rect 19163 57443 22147 60427
rect 22353 57443 25337 60427
rect 25543 57443 28527 60427
rect 28733 57443 31717 60427
rect 31923 57443 34907 60427
rect 35113 57443 38097 60427
rect 38303 57443 41287 60427
rect 41493 57443 44477 60427
rect 44683 57443 47667 60427
rect 47873 57443 50857 60427
rect 51063 57443 54047 60427
rect 54253 57443 57237 60427
rect 57443 57443 60427 60427
rect 60633 57443 63617 60427
rect 63823 57443 66807 60427
rect 67013 57443 69997 60427
rect 70203 57443 73187 60427
rect 73393 57443 76377 60427
rect 76583 57443 79567 60427
rect 79773 57443 82757 60427
rect 82963 57443 85947 60427
rect 86153 57443 89137 60427
rect 89343 57443 92327 60427
rect 92533 57443 95517 60427
rect 95723 57443 98707 60427
rect 98913 57443 101897 60427
rect 102103 57443 105087 60427
rect 105293 57443 108277 60427
rect 108483 57443 111467 60427
rect 111673 57443 114657 60427
rect 114863 57443 117847 60427
rect 118053 57443 121037 60427
rect 121243 57443 124227 60427
rect 124433 57443 127417 60427
rect 127623 57443 130607 60427
rect 130813 57443 133797 60427
rect 134003 57443 136987 60427
rect 23 54253 3007 57237
rect 3213 54253 6197 57237
rect 6403 54253 9387 57237
rect 9593 54253 12577 57237
rect 12783 54253 15767 57237
rect 15973 54253 18957 57237
rect 19163 54253 22147 57237
rect 22353 54253 25337 57237
rect 25543 54253 28527 57237
rect 28733 54253 31717 57237
rect 31923 54253 34907 57237
rect 35113 54253 38097 57237
rect 38303 54253 41287 57237
rect 41493 54253 44477 57237
rect 44683 54253 47667 57237
rect 47873 54253 50857 57237
rect 51063 54253 54047 57237
rect 54253 54253 57237 57237
rect 57443 54253 60427 57237
rect 60633 54253 63617 57237
rect 63823 54253 66807 57237
rect 67013 54253 69997 57237
rect 70203 54253 73187 57237
rect 73393 54253 76377 57237
rect 76583 54253 79567 57237
rect 79773 54253 82757 57237
rect 82963 54253 85947 57237
rect 86153 54253 89137 57237
rect 89343 54253 92327 57237
rect 92533 54253 95517 57237
rect 95723 54253 98707 57237
rect 98913 54253 101897 57237
rect 102103 54253 105087 57237
rect 105293 54253 108277 57237
rect 108483 54253 111467 57237
rect 111673 54253 114657 57237
rect 114863 54253 117847 57237
rect 118053 54253 121037 57237
rect 121243 54253 124227 57237
rect 124433 54253 127417 57237
rect 127623 54253 130607 57237
rect 130813 54253 133797 57237
rect 134003 54253 136987 57237
rect 23 51063 3007 54047
rect 3213 51063 6197 54047
rect 6403 51063 9387 54047
rect 9593 51063 12577 54047
rect 12783 51063 15767 54047
rect 15973 51063 18957 54047
rect 19163 51063 22147 54047
rect 22353 51063 25337 54047
rect 25543 51063 28527 54047
rect 28733 51063 31717 54047
rect 31923 51063 34907 54047
rect 35113 51063 38097 54047
rect 38303 51063 41287 54047
rect 41493 51063 44477 54047
rect 44683 51063 47667 54047
rect 47873 51063 50857 54047
rect 51063 51063 54047 54047
rect 54253 51063 57237 54047
rect 57443 51063 60427 54047
rect 60633 51063 63617 54047
rect 63823 51063 66807 54047
rect 67013 51063 69997 54047
rect 70203 51063 73187 54047
rect 73393 51063 76377 54047
rect 76583 51063 79567 54047
rect 79773 51063 82757 54047
rect 82963 51063 85947 54047
rect 86153 51063 89137 54047
rect 89343 51063 92327 54047
rect 92533 51063 95517 54047
rect 95723 51063 98707 54047
rect 98913 51063 101897 54047
rect 102103 51063 105087 54047
rect 105293 51063 108277 54047
rect 108483 51063 111467 54047
rect 111673 51063 114657 54047
rect 114863 51063 117847 54047
rect 118053 51063 121037 54047
rect 121243 51063 124227 54047
rect 124433 51063 127417 54047
rect 127623 51063 130607 54047
rect 130813 51063 133797 54047
rect 134003 51063 136987 54047
rect 23 47873 3007 50857
rect 3213 47873 6197 50857
rect 6403 47873 9387 50857
rect 9593 47873 12577 50857
rect 12783 47873 15767 50857
rect 15973 47873 18957 50857
rect 19163 47873 22147 50857
rect 22353 47873 25337 50857
rect 25543 47873 28527 50857
rect 28733 47873 31717 50857
rect 31923 47873 34907 50857
rect 35113 47873 38097 50857
rect 38303 47873 41287 50857
rect 41493 47873 44477 50857
rect 44683 47873 47667 50857
rect 47873 47873 50857 50857
rect 51063 47873 54047 50857
rect 54253 47873 57237 50857
rect 57443 47873 60427 50857
rect 60633 47873 63617 50857
rect 63823 47873 66807 50857
rect 67013 47873 69997 50857
rect 70203 47873 73187 50857
rect 73393 47873 76377 50857
rect 76583 47873 79567 50857
rect 79773 47873 82757 50857
rect 82963 47873 85947 50857
rect 86153 47873 89137 50857
rect 89343 47873 92327 50857
rect 92533 47873 95517 50857
rect 95723 47873 98707 50857
rect 98913 47873 101897 50857
rect 102103 47873 105087 50857
rect 105293 47873 108277 50857
rect 108483 47873 111467 50857
rect 111673 47873 114657 50857
rect 114863 47873 117847 50857
rect 118053 47873 121037 50857
rect 121243 47873 124227 50857
rect 124433 47873 127417 50857
rect 127623 47873 130607 50857
rect 130813 47873 133797 50857
rect 134003 47873 136987 50857
rect 23 44683 3007 47667
rect 3213 44683 6197 47667
rect 6403 44683 9387 47667
rect 9593 44683 12577 47667
rect 12783 44683 15767 47667
rect 15973 44683 18957 47667
rect 19163 44683 22147 47667
rect 22353 44683 25337 47667
rect 25543 44683 28527 47667
rect 28733 44683 31717 47667
rect 31923 44683 34907 47667
rect 35113 44683 38097 47667
rect 38303 44683 41287 47667
rect 41493 44683 44477 47667
rect 44683 44683 47667 47667
rect 47873 44683 50857 47667
rect 51063 44683 54047 47667
rect 54253 44683 57237 47667
rect 57443 44683 60427 47667
rect 60633 44683 63617 47667
rect 63823 44683 66807 47667
rect 67013 44683 69997 47667
rect 70203 44683 73187 47667
rect 73393 44683 76377 47667
rect 76583 44683 79567 47667
rect 79773 44683 82757 47667
rect 82963 44683 85947 47667
rect 86153 44683 89137 47667
rect 89343 44683 92327 47667
rect 92533 44683 95517 47667
rect 95723 44683 98707 47667
rect 98913 44683 101897 47667
rect 102103 44683 105087 47667
rect 105293 44683 108277 47667
rect 108483 44683 111467 47667
rect 111673 44683 114657 47667
rect 114863 44683 117847 47667
rect 118053 44683 121037 47667
rect 121243 44683 124227 47667
rect 124433 44683 127417 47667
rect 127623 44683 130607 47667
rect 130813 44683 133797 47667
rect 134003 44683 136987 47667
rect 23 41493 3007 44477
rect 3213 41493 6197 44477
rect 6403 41493 9387 44477
rect 9593 41493 12577 44477
rect 12783 41493 15767 44477
rect 15973 41493 18957 44477
rect 19163 41493 22147 44477
rect 22353 41493 25337 44477
rect 25543 41493 28527 44477
rect 28733 41493 31717 44477
rect 31923 41493 34907 44477
rect 35113 41493 38097 44477
rect 38303 41493 41287 44477
rect 41493 41493 44477 44477
rect 44683 41493 47667 44477
rect 47873 41493 50857 44477
rect 51063 41493 54047 44477
rect 54253 41493 57237 44477
rect 57443 41493 60427 44477
rect 60633 41493 63617 44477
rect 63823 41493 66807 44477
rect 67013 41493 69997 44477
rect 70203 41493 73187 44477
rect 73393 41493 76377 44477
rect 76583 41493 79567 44477
rect 79773 41493 82757 44477
rect 82963 41493 85947 44477
rect 86153 41493 89137 44477
rect 89343 41493 92327 44477
rect 92533 41493 95517 44477
rect 95723 41493 98707 44477
rect 98913 41493 101897 44477
rect 102103 41493 105087 44477
rect 105293 41493 108277 44477
rect 108483 41493 111467 44477
rect 111673 41493 114657 44477
rect 114863 41493 117847 44477
rect 118053 41493 121037 44477
rect 121243 41493 124227 44477
rect 124433 41493 127417 44477
rect 127623 41493 130607 44477
rect 130813 41493 133797 44477
rect 134003 41493 136987 44477
rect 23 38303 3007 41287
rect 3213 38303 6197 41287
rect 6403 38303 9387 41287
rect 9593 38303 12577 41287
rect 12783 38303 15767 41287
rect 15973 38303 18957 41287
rect 19163 38303 22147 41287
rect 22353 38303 25337 41287
rect 25543 38303 28527 41287
rect 28733 38303 31717 41287
rect 31923 38303 34907 41287
rect 35113 38303 38097 41287
rect 38303 38303 41287 41287
rect 41493 38303 44477 41287
rect 44683 38303 47667 41287
rect 47873 38303 50857 41287
rect 51063 38303 54047 41287
rect 54253 38303 57237 41287
rect 57443 38303 60427 41287
rect 60633 38303 63617 41287
rect 63823 38303 66807 41287
rect 67013 38303 69997 41287
rect 70203 38303 73187 41287
rect 73393 38303 76377 41287
rect 76583 38303 79567 41287
rect 79773 38303 82757 41287
rect 82963 38303 85947 41287
rect 86153 38303 89137 41287
rect 89343 38303 92327 41287
rect 92533 38303 95517 41287
rect 95723 38303 98707 41287
rect 98913 38303 101897 41287
rect 102103 38303 105087 41287
rect 105293 38303 108277 41287
rect 108483 38303 111467 41287
rect 111673 38303 114657 41287
rect 114863 38303 117847 41287
rect 118053 38303 121037 41287
rect 121243 38303 124227 41287
rect 124433 38303 127417 41287
rect 127623 38303 130607 41287
rect 130813 38303 133797 41287
rect 134003 38303 136987 41287
rect 23 35113 3007 38097
rect 3213 35113 6197 38097
rect 6403 35113 9387 38097
rect 9593 35113 12577 38097
rect 12783 35113 15767 38097
rect 15973 35113 18957 38097
rect 19163 35113 22147 38097
rect 22353 35113 25337 38097
rect 25543 35113 28527 38097
rect 28733 35113 31717 38097
rect 31923 35113 34907 38097
rect 35113 35113 38097 38097
rect 38303 35113 41287 38097
rect 41493 35113 44477 38097
rect 44683 35113 47667 38097
rect 47873 35113 50857 38097
rect 51063 35113 54047 38097
rect 54253 35113 57237 38097
rect 57443 35113 60427 38097
rect 60633 35113 63617 38097
rect 63823 35113 66807 38097
rect 67013 35113 69997 38097
rect 70203 35113 73187 38097
rect 73393 35113 76377 38097
rect 76583 35113 79567 38097
rect 79773 35113 82757 38097
rect 82963 35113 85947 38097
rect 86153 35113 89137 38097
rect 89343 35113 92327 38097
rect 92533 35113 95517 38097
rect 95723 35113 98707 38097
rect 98913 35113 101897 38097
rect 102103 35113 105087 38097
rect 105293 35113 108277 38097
rect 108483 35113 111467 38097
rect 111673 35113 114657 38097
rect 114863 35113 117847 38097
rect 118053 35113 121037 38097
rect 121243 35113 124227 38097
rect 124433 35113 127417 38097
rect 127623 35113 130607 38097
rect 130813 35113 133797 38097
rect 134003 35113 136987 38097
rect 23 31923 3007 34907
rect 3213 31923 6197 34907
rect 6403 31923 9387 34907
rect 9593 31923 12577 34907
rect 12783 31923 15767 34907
rect 15973 31923 18957 34907
rect 19163 31923 22147 34907
rect 22353 31923 25337 34907
rect 25543 31923 28527 34907
rect 28733 31923 31717 34907
rect 31923 31923 34907 34907
rect 35113 31923 38097 34907
rect 38303 31923 41287 34907
rect 41493 31923 44477 34907
rect 44683 31923 47667 34907
rect 47873 31923 50857 34907
rect 51063 31923 54047 34907
rect 54253 31923 57237 34907
rect 57443 31923 60427 34907
rect 60633 31923 63617 34907
rect 63823 31923 66807 34907
rect 67013 31923 69997 34907
rect 70203 31923 73187 34907
rect 73393 31923 76377 34907
rect 76583 31923 79567 34907
rect 79773 31923 82757 34907
rect 82963 31923 85947 34907
rect 86153 31923 89137 34907
rect 89343 31923 92327 34907
rect 92533 31923 95517 34907
rect 95723 31923 98707 34907
rect 98913 31923 101897 34907
rect 102103 31923 105087 34907
rect 105293 31923 108277 34907
rect 108483 31923 111467 34907
rect 111673 31923 114657 34907
rect 114863 31923 117847 34907
rect 118053 31923 121037 34907
rect 121243 31923 124227 34907
rect 124433 31923 127417 34907
rect 127623 31923 130607 34907
rect 130813 31923 133797 34907
rect 134003 31923 136987 34907
rect 23 28733 3007 31717
rect 3213 28733 6197 31717
rect 6403 28733 9387 31717
rect 9593 28733 12577 31717
rect 12783 28733 15767 31717
rect 15973 28733 18957 31717
rect 19163 28733 22147 31717
rect 22353 28733 25337 31717
rect 25543 28733 28527 31717
rect 28733 28733 31717 31717
rect 31923 28733 34907 31717
rect 35113 28733 38097 31717
rect 38303 28733 41287 31717
rect 41493 28733 44477 31717
rect 44683 28733 47667 31717
rect 47873 28733 50857 31717
rect 51063 28733 54047 31717
rect 54253 28733 57237 31717
rect 57443 28733 60427 31717
rect 60633 28733 63617 31717
rect 63823 28733 66807 31717
rect 67013 28733 69997 31717
rect 70203 28733 73187 31717
rect 73393 28733 76377 31717
rect 76583 28733 79567 31717
rect 79773 28733 82757 31717
rect 82963 28733 85947 31717
rect 86153 28733 89137 31717
rect 89343 28733 92327 31717
rect 92533 28733 95517 31717
rect 95723 28733 98707 31717
rect 98913 28733 101897 31717
rect 102103 28733 105087 31717
rect 105293 28733 108277 31717
rect 108483 28733 111467 31717
rect 111673 28733 114657 31717
rect 114863 28733 117847 31717
rect 118053 28733 121037 31717
rect 121243 28733 124227 31717
rect 124433 28733 127417 31717
rect 127623 28733 130607 31717
rect 130813 28733 133797 31717
rect 134003 28733 136987 31717
rect 23 25543 3007 28527
rect 3213 25543 6197 28527
rect 6403 25543 9387 28527
rect 9593 25543 12577 28527
rect 12783 25543 15767 28527
rect 15973 25543 18957 28527
rect 19163 25543 22147 28527
rect 22353 25543 25337 28527
rect 25543 25543 28527 28527
rect 28733 25543 31717 28527
rect 31923 25543 34907 28527
rect 35113 25543 38097 28527
rect 38303 25543 41287 28527
rect 41493 25543 44477 28527
rect 44683 25543 47667 28527
rect 47873 25543 50857 28527
rect 51063 25543 54047 28527
rect 54253 25543 57237 28527
rect 57443 25543 60427 28527
rect 60633 25543 63617 28527
rect 63823 25543 66807 28527
rect 67013 25543 69997 28527
rect 70203 25543 73187 28527
rect 73393 25543 76377 28527
rect 76583 25543 79567 28527
rect 79773 25543 82757 28527
rect 82963 25543 85947 28527
rect 86153 25543 89137 28527
rect 89343 25543 92327 28527
rect 92533 25543 95517 28527
rect 95723 25543 98707 28527
rect 98913 25543 101897 28527
rect 102103 25543 105087 28527
rect 105293 25543 108277 28527
rect 108483 25543 111467 28527
rect 111673 25543 114657 28527
rect 114863 25543 117847 28527
rect 118053 25543 121037 28527
rect 121243 25543 124227 28527
rect 124433 25543 127417 28527
rect 127623 25543 130607 28527
rect 130813 25543 133797 28527
rect 134003 25543 136987 28527
rect 23 22353 3007 25337
rect 3213 22353 6197 25337
rect 6403 22353 9387 25337
rect 9593 22353 12577 25337
rect 12783 22353 15767 25337
rect 15973 22353 18957 25337
rect 19163 22353 22147 25337
rect 22353 22353 25337 25337
rect 25543 22353 28527 25337
rect 28733 22353 31717 25337
rect 31923 22353 34907 25337
rect 35113 22353 38097 25337
rect 38303 22353 41287 25337
rect 41493 22353 44477 25337
rect 44683 22353 47667 25337
rect 47873 22353 50857 25337
rect 51063 22353 54047 25337
rect 54253 22353 57237 25337
rect 57443 22353 60427 25337
rect 60633 22353 63617 25337
rect 63823 22353 66807 25337
rect 67013 22353 69997 25337
rect 70203 22353 73187 25337
rect 73393 22353 76377 25337
rect 76583 22353 79567 25337
rect 79773 22353 82757 25337
rect 82963 22353 85947 25337
rect 86153 22353 89137 25337
rect 89343 22353 92327 25337
rect 92533 22353 95517 25337
rect 95723 22353 98707 25337
rect 98913 22353 101897 25337
rect 102103 22353 105087 25337
rect 105293 22353 108277 25337
rect 108483 22353 111467 25337
rect 111673 22353 114657 25337
rect 114863 22353 117847 25337
rect 118053 22353 121037 25337
rect 121243 22353 124227 25337
rect 124433 22353 127417 25337
rect 127623 22353 130607 25337
rect 130813 22353 133797 25337
rect 134003 22353 136987 25337
rect 23 19163 3007 22147
rect 3213 19163 6197 22147
rect 6403 19163 9387 22147
rect 9593 19163 12577 22147
rect 12783 19163 15767 22147
rect 15973 19163 18957 22147
rect 19163 19163 22147 22147
rect 22353 19163 25337 22147
rect 25543 19163 28527 22147
rect 28733 19163 31717 22147
rect 31923 19163 34907 22147
rect 35113 19163 38097 22147
rect 38303 19163 41287 22147
rect 41493 19163 44477 22147
rect 44683 19163 47667 22147
rect 47873 19163 50857 22147
rect 51063 19163 54047 22147
rect 54253 19163 57237 22147
rect 57443 19163 60427 22147
rect 60633 19163 63617 22147
rect 63823 19163 66807 22147
rect 67013 19163 69997 22147
rect 70203 19163 73187 22147
rect 73393 19163 76377 22147
rect 76583 19163 79567 22147
rect 79773 19163 82757 22147
rect 82963 19163 85947 22147
rect 86153 19163 89137 22147
rect 89343 19163 92327 22147
rect 92533 19163 95517 22147
rect 95723 19163 98707 22147
rect 98913 19163 101897 22147
rect 102103 19163 105087 22147
rect 105293 19163 108277 22147
rect 108483 19163 111467 22147
rect 111673 19163 114657 22147
rect 114863 19163 117847 22147
rect 118053 19163 121037 22147
rect 121243 19163 124227 22147
rect 124433 19163 127417 22147
rect 127623 19163 130607 22147
rect 130813 19163 133797 22147
rect 134003 19163 136987 22147
rect 23 15973 3007 18957
rect 3213 15973 6197 18957
rect 6403 15973 9387 18957
rect 9593 15973 12577 18957
rect 12783 15973 15767 18957
rect 15973 15973 18957 18957
rect 19163 15973 22147 18957
rect 22353 15973 25337 18957
rect 25543 15973 28527 18957
rect 28733 15973 31717 18957
rect 31923 15973 34907 18957
rect 35113 15973 38097 18957
rect 38303 15973 41287 18957
rect 41493 15973 44477 18957
rect 44683 15973 47667 18957
rect 47873 15973 50857 18957
rect 51063 15973 54047 18957
rect 54253 15973 57237 18957
rect 57443 15973 60427 18957
rect 60633 15973 63617 18957
rect 63823 15973 66807 18957
rect 67013 15973 69997 18957
rect 70203 15973 73187 18957
rect 73393 15973 76377 18957
rect 76583 15973 79567 18957
rect 79773 15973 82757 18957
rect 82963 15973 85947 18957
rect 86153 15973 89137 18957
rect 89343 15973 92327 18957
rect 92533 15973 95517 18957
rect 95723 15973 98707 18957
rect 98913 15973 101897 18957
rect 102103 15973 105087 18957
rect 105293 15973 108277 18957
rect 108483 15973 111467 18957
rect 111673 15973 114657 18957
rect 114863 15973 117847 18957
rect 118053 15973 121037 18957
rect 121243 15973 124227 18957
rect 124433 15973 127417 18957
rect 127623 15973 130607 18957
rect 130813 15973 133797 18957
rect 134003 15973 136987 18957
rect 23 12783 3007 15767
rect 3213 12783 6197 15767
rect 6403 12783 9387 15767
rect 9593 12783 12577 15767
rect 12783 12783 15767 15767
rect 15973 12783 18957 15767
rect 19163 12783 22147 15767
rect 22353 12783 25337 15767
rect 25543 12783 28527 15767
rect 28733 12783 31717 15767
rect 31923 12783 34907 15767
rect 35113 12783 38097 15767
rect 38303 12783 41287 15767
rect 41493 12783 44477 15767
rect 44683 12783 47667 15767
rect 47873 12783 50857 15767
rect 51063 12783 54047 15767
rect 54253 12783 57237 15767
rect 57443 12783 60427 15767
rect 60633 12783 63617 15767
rect 63823 12783 66807 15767
rect 67013 12783 69997 15767
rect 70203 12783 73187 15767
rect 73393 12783 76377 15767
rect 76583 12783 79567 15767
rect 79773 12783 82757 15767
rect 82963 12783 85947 15767
rect 86153 12783 89137 15767
rect 89343 12783 92327 15767
rect 92533 12783 95517 15767
rect 95723 12783 98707 15767
rect 98913 12783 101897 15767
rect 102103 12783 105087 15767
rect 105293 12783 108277 15767
rect 108483 12783 111467 15767
rect 111673 12783 114657 15767
rect 114863 12783 117847 15767
rect 118053 12783 121037 15767
rect 121243 12783 124227 15767
rect 124433 12783 127417 15767
rect 127623 12783 130607 15767
rect 130813 12783 133797 15767
rect 134003 12783 136987 15767
rect 23 9593 3007 12577
rect 3213 9593 6197 12577
rect 6403 9593 9387 12577
rect 9593 9593 12577 12577
rect 12783 9593 15767 12577
rect 15973 9593 18957 12577
rect 19163 9593 22147 12577
rect 22353 9593 25337 12577
rect 25543 9593 28527 12577
rect 28733 9593 31717 12577
rect 31923 9593 34907 12577
rect 35113 9593 38097 12577
rect 38303 9593 41287 12577
rect 41493 9593 44477 12577
rect 44683 9593 47667 12577
rect 47873 9593 50857 12577
rect 51063 9593 54047 12577
rect 54253 9593 57237 12577
rect 57443 9593 60427 12577
rect 60633 9593 63617 12577
rect 63823 9593 66807 12577
rect 67013 9593 69997 12577
rect 70203 9593 73187 12577
rect 73393 9593 76377 12577
rect 76583 9593 79567 12577
rect 79773 9593 82757 12577
rect 82963 9593 85947 12577
rect 86153 9593 89137 12577
rect 89343 9593 92327 12577
rect 92533 9593 95517 12577
rect 95723 9593 98707 12577
rect 98913 9593 101897 12577
rect 102103 9593 105087 12577
rect 105293 9593 108277 12577
rect 108483 9593 111467 12577
rect 111673 9593 114657 12577
rect 114863 9593 117847 12577
rect 118053 9593 121037 12577
rect 121243 9593 124227 12577
rect 124433 9593 127417 12577
rect 127623 9593 130607 12577
rect 130813 9593 133797 12577
rect 134003 9593 136987 12577
rect 23 6403 3007 9387
rect 3213 6403 6197 9387
rect 6403 6403 9387 9387
rect 9593 6403 12577 9387
rect 12783 6403 15767 9387
rect 15973 6403 18957 9387
rect 19163 6403 22147 9387
rect 22353 6403 25337 9387
rect 25543 6403 28527 9387
rect 28733 6403 31717 9387
rect 31923 6403 34907 9387
rect 35113 6403 38097 9387
rect 38303 6403 41287 9387
rect 41493 6403 44477 9387
rect 44683 6403 47667 9387
rect 47873 6403 50857 9387
rect 51063 6403 54047 9387
rect 54253 6403 57237 9387
rect 57443 6403 60427 9387
rect 60633 6403 63617 9387
rect 63823 6403 66807 9387
rect 67013 6403 69997 9387
rect 70203 6403 73187 9387
rect 73393 6403 76377 9387
rect 76583 6403 79567 9387
rect 79773 6403 82757 9387
rect 82963 6403 85947 9387
rect 86153 6403 89137 9387
rect 89343 6403 92327 9387
rect 92533 6403 95517 9387
rect 95723 6403 98707 9387
rect 98913 6403 101897 9387
rect 102103 6403 105087 9387
rect 105293 6403 108277 9387
rect 108483 6403 111467 9387
rect 111673 6403 114657 9387
rect 114863 6403 117847 9387
rect 118053 6403 121037 9387
rect 121243 6403 124227 9387
rect 124433 6403 127417 9387
rect 127623 6403 130607 9387
rect 130813 6403 133797 9387
rect 134003 6403 136987 9387
rect 23 3213 3007 6197
rect 3213 3213 6197 6197
rect 6403 3213 9387 6197
rect 9593 3213 12577 6197
rect 12783 3213 15767 6197
rect 15973 3213 18957 6197
rect 19163 3213 22147 6197
rect 22353 3213 25337 6197
rect 25543 3213 28527 6197
rect 28733 3213 31717 6197
rect 31923 3213 34907 6197
rect 35113 3213 38097 6197
rect 38303 3213 41287 6197
rect 41493 3213 44477 6197
rect 44683 3213 47667 6197
rect 47873 3213 50857 6197
rect 51063 3213 54047 6197
rect 54253 3213 57237 6197
rect 57443 3213 60427 6197
rect 60633 3213 63617 6197
rect 63823 3213 66807 6197
rect 67013 3213 69997 6197
rect 70203 3213 73187 6197
rect 73393 3213 76377 6197
rect 76583 3213 79567 6197
rect 79773 3213 82757 6197
rect 82963 3213 85947 6197
rect 86153 3213 89137 6197
rect 89343 3213 92327 6197
rect 92533 3213 95517 6197
rect 95723 3213 98707 6197
rect 98913 3213 101897 6197
rect 102103 3213 105087 6197
rect 105293 3213 108277 6197
rect 108483 3213 111467 6197
rect 111673 3213 114657 6197
rect 114863 3213 117847 6197
rect 118053 3213 121037 6197
rect 121243 3213 124227 6197
rect 124433 3213 127417 6197
rect 127623 3213 130607 6197
rect 130813 3213 133797 6197
rect 134003 3213 136987 6197
rect 23 23 3007 3007
rect 3213 23 6197 3007
rect 6403 23 9387 3007
rect 9593 23 12577 3007
rect 12783 23 15767 3007
rect 15973 23 18957 3007
rect 19163 23 22147 3007
rect 22353 23 25337 3007
rect 25543 23 28527 3007
rect 28733 23 31717 3007
rect 31923 23 34907 3007
rect 35113 23 38097 3007
rect 38303 23 41287 3007
rect 41493 23 44477 3007
rect 44683 23 47667 3007
rect 47873 23 50857 3007
rect 51063 23 54047 3007
rect 54253 23 57237 3007
rect 57443 23 60427 3007
rect 60633 23 63617 3007
rect 63823 23 66807 3007
rect 67013 23 69997 3007
rect 70203 23 73187 3007
rect 73393 23 76377 3007
rect 76583 23 79567 3007
rect 79773 23 82757 3007
rect 82963 23 85947 3007
rect 86153 23 89137 3007
rect 89343 23 92327 3007
rect 92533 23 95517 3007
rect 95723 23 98707 3007
rect 98913 23 101897 3007
rect 102103 23 105087 3007
rect 105293 23 108277 3007
rect 108483 23 111467 3007
rect 111673 23 114657 3007
rect 114863 23 117847 3007
rect 118053 23 121037 3007
rect 121243 23 124227 3007
rect 124433 23 127417 3007
rect 127623 23 130607 3007
rect 130813 23 133797 3007
rect 134003 23 136987 3007
<< metal5 >>
rect 1000 166980 68990 167000
rect 1000 166020 1020 166980
rect 68970 166020 68990 166980
rect 1000 165880 68990 166020
rect 71180 166980 135980 168000
rect 71180 166020 71200 166980
rect 135960 166020 135980 166980
rect 71180 166000 135980 166020
rect 1000 165720 2000 165880
rect 4190 165720 5190 165880
rect 7380 165720 8380 165880
rect 10570 165720 11570 165880
rect 13760 165720 14760 165880
rect 16950 165720 17950 165880
rect 20140 165720 21140 165880
rect 23330 165720 24330 165880
rect 26520 165720 27520 165880
rect 29710 165720 30710 165880
rect 32900 165720 33900 165880
rect 36090 165720 37090 165880
rect 39280 165720 40280 165880
rect 42470 165720 43470 165880
rect 45660 165720 46660 165880
rect 48850 165720 49850 165880
rect 52040 165720 53040 165880
rect 55230 165720 56230 165880
rect 58420 165720 59420 165880
rect 61610 165720 62610 165880
rect 64800 165720 65800 165880
rect 67990 165720 68990 165880
rect 71180 165720 72180 165800
rect 74370 165720 75370 165800
rect 77560 165720 78560 165800
rect 80750 165720 81750 165800
rect 83940 165720 84940 165800
rect 87130 165720 88130 165800
rect 90320 165720 91320 165800
rect 93510 165720 94510 165800
rect 96700 165720 97700 165800
rect 99890 165720 100890 165800
rect 103080 165720 104080 165800
rect 106270 165720 107270 165800
rect 109460 165720 110460 165800
rect 112650 165720 113650 165800
rect 115840 165720 116840 165800
rect 119030 165720 120030 165800
rect 122220 165720 123220 165800
rect 125410 165720 126410 165800
rect 128600 165720 129600 165800
rect 131790 165720 132790 165800
rect 134980 165720 135980 165800
rect 0 165697 3030 165720
rect 0 162713 23 165697
rect 3007 164690 3030 165697
rect 3190 165697 6220 165720
rect 3190 164690 3213 165697
rect 3007 163690 3213 164690
rect 3007 162713 3030 163690
rect 0 162690 3030 162713
rect 3190 162713 3213 163690
rect 6197 164690 6220 165697
rect 6380 165697 9410 165720
rect 6380 164690 6403 165697
rect 6197 163690 6403 164690
rect 6197 162713 6220 163690
rect 3190 162690 6220 162713
rect 6380 162713 6403 163690
rect 9387 164690 9410 165697
rect 9570 165697 12600 165720
rect 9570 164690 9593 165697
rect 9387 163690 9593 164690
rect 9387 162713 9410 163690
rect 6380 162690 9410 162713
rect 9570 162713 9593 163690
rect 12577 164690 12600 165697
rect 12760 165697 15790 165720
rect 12760 164690 12783 165697
rect 12577 163690 12783 164690
rect 12577 162713 12600 163690
rect 9570 162690 12600 162713
rect 12760 162713 12783 163690
rect 15767 164690 15790 165697
rect 15950 165697 18980 165720
rect 15950 164690 15973 165697
rect 15767 163690 15973 164690
rect 15767 162713 15790 163690
rect 12760 162690 15790 162713
rect 15950 162713 15973 163690
rect 18957 164690 18980 165697
rect 19140 165697 22170 165720
rect 19140 164690 19163 165697
rect 18957 163690 19163 164690
rect 18957 162713 18980 163690
rect 15950 162690 18980 162713
rect 19140 162713 19163 163690
rect 22147 164690 22170 165697
rect 22330 165697 25360 165720
rect 22330 164690 22353 165697
rect 22147 163690 22353 164690
rect 22147 162713 22170 163690
rect 19140 162690 22170 162713
rect 22330 162713 22353 163690
rect 25337 164690 25360 165697
rect 25520 165697 28550 165720
rect 25520 164690 25543 165697
rect 25337 163690 25543 164690
rect 25337 162713 25360 163690
rect 22330 162690 25360 162713
rect 25520 162713 25543 163690
rect 28527 164690 28550 165697
rect 28710 165697 31740 165720
rect 28710 164690 28733 165697
rect 28527 163690 28733 164690
rect 28527 162713 28550 163690
rect 25520 162690 28550 162713
rect 28710 162713 28733 163690
rect 31717 164690 31740 165697
rect 31900 165697 34930 165720
rect 31900 164690 31923 165697
rect 31717 163690 31923 164690
rect 31717 162713 31740 163690
rect 28710 162690 31740 162713
rect 31900 162713 31923 163690
rect 34907 164690 34930 165697
rect 35090 165697 38120 165720
rect 35090 164690 35113 165697
rect 34907 163690 35113 164690
rect 34907 162713 34930 163690
rect 31900 162690 34930 162713
rect 35090 162713 35113 163690
rect 38097 164690 38120 165697
rect 38280 165697 41310 165720
rect 38280 164690 38303 165697
rect 38097 163690 38303 164690
rect 38097 162713 38120 163690
rect 35090 162690 38120 162713
rect 38280 162713 38303 163690
rect 41287 164690 41310 165697
rect 41470 165697 44500 165720
rect 41470 164690 41493 165697
rect 41287 163690 41493 164690
rect 41287 162713 41310 163690
rect 38280 162690 41310 162713
rect 41470 162713 41493 163690
rect 44477 164690 44500 165697
rect 44660 165697 47690 165720
rect 44660 164690 44683 165697
rect 44477 163690 44683 164690
rect 44477 162713 44500 163690
rect 41470 162690 44500 162713
rect 44660 162713 44683 163690
rect 47667 164690 47690 165697
rect 47850 165697 50880 165720
rect 47850 164690 47873 165697
rect 47667 163690 47873 164690
rect 47667 162713 47690 163690
rect 44660 162690 47690 162713
rect 47850 162713 47873 163690
rect 50857 164690 50880 165697
rect 51040 165697 54070 165720
rect 51040 164690 51063 165697
rect 50857 163690 51063 164690
rect 50857 162713 50880 163690
rect 47850 162690 50880 162713
rect 51040 162713 51063 163690
rect 54047 164690 54070 165697
rect 54230 165697 57260 165720
rect 54230 164690 54253 165697
rect 54047 163690 54253 164690
rect 54047 162713 54070 163690
rect 51040 162690 54070 162713
rect 54230 162713 54253 163690
rect 57237 164690 57260 165697
rect 57420 165697 60450 165720
rect 57420 164690 57443 165697
rect 57237 163690 57443 164690
rect 57237 162713 57260 163690
rect 54230 162690 57260 162713
rect 57420 162713 57443 163690
rect 60427 164690 60450 165697
rect 60610 165697 63640 165720
rect 60610 164690 60633 165697
rect 60427 163690 60633 164690
rect 60427 162713 60450 163690
rect 57420 162690 60450 162713
rect 60610 162713 60633 163690
rect 63617 164690 63640 165697
rect 63800 165697 66830 165720
rect 63800 164690 63823 165697
rect 63617 163690 63823 164690
rect 63617 162713 63640 163690
rect 60610 162690 63640 162713
rect 63800 162713 63823 163690
rect 66807 164690 66830 165697
rect 66990 165697 70020 165720
rect 66990 164690 67013 165697
rect 66807 163690 67013 164690
rect 66807 162713 66830 163690
rect 63800 162690 66830 162713
rect 66990 162713 67013 163690
rect 69997 164690 70020 165697
rect 70180 165697 73210 165720
rect 70180 164690 70203 165697
rect 69997 163690 70203 164690
rect 69997 162713 70020 163690
rect 66990 162690 70020 162713
rect 70180 162713 70203 163690
rect 73187 164690 73210 165697
rect 73370 165697 76400 165720
rect 73370 164690 73393 165697
rect 73187 163690 73393 164690
rect 73187 162713 73210 163690
rect 70180 162690 73210 162713
rect 73370 162713 73393 163690
rect 76377 164690 76400 165697
rect 76560 165697 79590 165720
rect 76560 164690 76583 165697
rect 76377 163690 76583 164690
rect 76377 162713 76400 163690
rect 73370 162690 76400 162713
rect 76560 162713 76583 163690
rect 79567 164690 79590 165697
rect 79750 165697 82780 165720
rect 79750 164690 79773 165697
rect 79567 163690 79773 164690
rect 79567 162713 79590 163690
rect 76560 162690 79590 162713
rect 79750 162713 79773 163690
rect 82757 164690 82780 165697
rect 82940 165697 85970 165720
rect 82940 164690 82963 165697
rect 82757 163690 82963 164690
rect 82757 162713 82780 163690
rect 79750 162690 82780 162713
rect 82940 162713 82963 163690
rect 85947 164690 85970 165697
rect 86130 165697 89160 165720
rect 86130 164690 86153 165697
rect 85947 163690 86153 164690
rect 85947 162713 85970 163690
rect 82940 162690 85970 162713
rect 86130 162713 86153 163690
rect 89137 164690 89160 165697
rect 89320 165697 92350 165720
rect 89320 164690 89343 165697
rect 89137 163690 89343 164690
rect 89137 162713 89160 163690
rect 86130 162690 89160 162713
rect 89320 162713 89343 163690
rect 92327 164690 92350 165697
rect 92510 165697 95540 165720
rect 92510 164690 92533 165697
rect 92327 163690 92533 164690
rect 92327 162713 92350 163690
rect 89320 162690 92350 162713
rect 92510 162713 92533 163690
rect 95517 164690 95540 165697
rect 95700 165697 98730 165720
rect 95700 164690 95723 165697
rect 95517 163690 95723 164690
rect 95517 162713 95540 163690
rect 92510 162690 95540 162713
rect 95700 162713 95723 163690
rect 98707 164690 98730 165697
rect 98890 165697 101920 165720
rect 98890 164690 98913 165697
rect 98707 163690 98913 164690
rect 98707 162713 98730 163690
rect 95700 162690 98730 162713
rect 98890 162713 98913 163690
rect 101897 164690 101920 165697
rect 102080 165697 105110 165720
rect 102080 164690 102103 165697
rect 101897 163690 102103 164690
rect 101897 162713 101920 163690
rect 98890 162690 101920 162713
rect 102080 162713 102103 163690
rect 105087 164690 105110 165697
rect 105270 165697 108300 165720
rect 105270 164690 105293 165697
rect 105087 163690 105293 164690
rect 105087 162713 105110 163690
rect 102080 162690 105110 162713
rect 105270 162713 105293 163690
rect 108277 164690 108300 165697
rect 108460 165697 111490 165720
rect 108460 164690 108483 165697
rect 108277 163690 108483 164690
rect 108277 162713 108300 163690
rect 105270 162690 108300 162713
rect 108460 162713 108483 163690
rect 111467 164690 111490 165697
rect 111650 165697 114680 165720
rect 111650 164690 111673 165697
rect 111467 163690 111673 164690
rect 111467 162713 111490 163690
rect 108460 162690 111490 162713
rect 111650 162713 111673 163690
rect 114657 164690 114680 165697
rect 114840 165697 117870 165720
rect 114840 164690 114863 165697
rect 114657 163690 114863 164690
rect 114657 162713 114680 163690
rect 111650 162690 114680 162713
rect 114840 162713 114863 163690
rect 117847 164690 117870 165697
rect 118030 165697 121060 165720
rect 118030 164690 118053 165697
rect 117847 163690 118053 164690
rect 117847 162713 117870 163690
rect 114840 162690 117870 162713
rect 118030 162713 118053 163690
rect 121037 164690 121060 165697
rect 121220 165697 124250 165720
rect 121220 164690 121243 165697
rect 121037 163690 121243 164690
rect 121037 162713 121060 163690
rect 118030 162690 121060 162713
rect 121220 162713 121243 163690
rect 124227 164690 124250 165697
rect 124410 165697 127440 165720
rect 124410 164690 124433 165697
rect 124227 163690 124433 164690
rect 124227 162713 124250 163690
rect 121220 162690 124250 162713
rect 124410 162713 124433 163690
rect 127417 164690 127440 165697
rect 127600 165697 130630 165720
rect 127600 164690 127623 165697
rect 127417 163690 127623 164690
rect 127417 162713 127440 163690
rect 124410 162690 127440 162713
rect 127600 162713 127623 163690
rect 130607 164690 130630 165697
rect 130790 165697 133820 165720
rect 130790 164690 130813 165697
rect 130607 163690 130813 164690
rect 130607 162713 130630 163690
rect 127600 162690 130630 162713
rect 130790 162713 130813 163690
rect 133797 164690 133820 165697
rect 133980 165697 137010 165720
rect 133980 164690 134003 165697
rect 133797 163690 134003 164690
rect 133797 162713 133820 163690
rect 130790 162690 133820 162713
rect 133980 162713 134003 163690
rect 136987 164690 137010 165697
rect 136987 163690 137170 164690
rect 136987 162713 137010 163690
rect 133980 162690 137010 162713
rect 1000 162530 2000 162690
rect 4190 162530 5190 162690
rect 7380 162530 8380 162690
rect 10570 162530 11570 162690
rect 13760 162530 14760 162690
rect 16950 162530 17950 162690
rect 20140 162530 21140 162690
rect 23330 162530 24330 162690
rect 26520 162530 27520 162690
rect 29710 162530 30710 162690
rect 32900 162530 33900 162690
rect 36090 162530 37090 162690
rect 39280 162530 40280 162690
rect 42470 162530 43470 162690
rect 45660 162530 46660 162690
rect 48850 162530 49850 162690
rect 52040 162530 53040 162690
rect 55230 162530 56230 162690
rect 58420 162530 59420 162690
rect 61610 162530 62610 162690
rect 64800 162530 65800 162690
rect 67990 162530 68990 162690
rect 71180 162530 72180 162690
rect 74370 162530 75370 162690
rect 77560 162530 78560 162690
rect 80750 162530 81750 162690
rect 83940 162530 84940 162690
rect 87130 162530 88130 162690
rect 90320 162530 91320 162690
rect 93510 162530 94510 162690
rect 96700 162530 97700 162690
rect 99890 162530 100890 162690
rect 103080 162530 104080 162690
rect 106270 162530 107270 162690
rect 109460 162530 110460 162690
rect 112650 162530 113650 162690
rect 115840 162530 116840 162690
rect 119030 162530 120030 162690
rect 122220 162530 123220 162690
rect 125410 162530 126410 162690
rect 128600 162530 129600 162690
rect 131790 162530 132790 162690
rect 134980 162530 135980 162690
rect 0 162507 3030 162530
rect 0 159523 23 162507
rect 3007 161500 3030 162507
rect 3190 162507 6220 162530
rect 3190 161500 3213 162507
rect 3007 160500 3213 161500
rect 3007 159523 3030 160500
rect 0 159500 3030 159523
rect 3190 159523 3213 160500
rect 6197 161500 6220 162507
rect 6380 162507 9410 162530
rect 6380 161500 6403 162507
rect 6197 160500 6403 161500
rect 6197 159523 6220 160500
rect 3190 159500 6220 159523
rect 6380 159523 6403 160500
rect 9387 161500 9410 162507
rect 9570 162507 12600 162530
rect 9570 161500 9593 162507
rect 9387 160500 9593 161500
rect 9387 159523 9410 160500
rect 6380 159500 9410 159523
rect 9570 159523 9593 160500
rect 12577 161500 12600 162507
rect 12760 162507 15790 162530
rect 12760 161500 12783 162507
rect 12577 160500 12783 161500
rect 12577 159523 12600 160500
rect 9570 159500 12600 159523
rect 12760 159523 12783 160500
rect 15767 161500 15790 162507
rect 15950 162507 18980 162530
rect 15950 161500 15973 162507
rect 15767 160500 15973 161500
rect 15767 159523 15790 160500
rect 12760 159500 15790 159523
rect 15950 159523 15973 160500
rect 18957 161500 18980 162507
rect 19140 162507 22170 162530
rect 19140 161500 19163 162507
rect 18957 160500 19163 161500
rect 18957 159523 18980 160500
rect 15950 159500 18980 159523
rect 19140 159523 19163 160500
rect 22147 161500 22170 162507
rect 22330 162507 25360 162530
rect 22330 161500 22353 162507
rect 22147 160500 22353 161500
rect 22147 159523 22170 160500
rect 19140 159500 22170 159523
rect 22330 159523 22353 160500
rect 25337 161500 25360 162507
rect 25520 162507 28550 162530
rect 25520 161500 25543 162507
rect 25337 160500 25543 161500
rect 25337 159523 25360 160500
rect 22330 159500 25360 159523
rect 25520 159523 25543 160500
rect 28527 161500 28550 162507
rect 28710 162507 31740 162530
rect 28710 161500 28733 162507
rect 28527 160500 28733 161500
rect 28527 159523 28550 160500
rect 25520 159500 28550 159523
rect 28710 159523 28733 160500
rect 31717 161500 31740 162507
rect 31900 162507 34930 162530
rect 31900 161500 31923 162507
rect 31717 160500 31923 161500
rect 31717 159523 31740 160500
rect 28710 159500 31740 159523
rect 31900 159523 31923 160500
rect 34907 161500 34930 162507
rect 35090 162507 38120 162530
rect 35090 161500 35113 162507
rect 34907 160500 35113 161500
rect 34907 159523 34930 160500
rect 31900 159500 34930 159523
rect 35090 159523 35113 160500
rect 38097 161500 38120 162507
rect 38280 162507 41310 162530
rect 38280 161500 38303 162507
rect 38097 160500 38303 161500
rect 38097 159523 38120 160500
rect 35090 159500 38120 159523
rect 38280 159523 38303 160500
rect 41287 161500 41310 162507
rect 41470 162507 44500 162530
rect 41470 161500 41493 162507
rect 41287 160500 41493 161500
rect 41287 159523 41310 160500
rect 38280 159500 41310 159523
rect 41470 159523 41493 160500
rect 44477 161500 44500 162507
rect 44660 162507 47690 162530
rect 44660 161500 44683 162507
rect 44477 160500 44683 161500
rect 44477 159523 44500 160500
rect 41470 159500 44500 159523
rect 44660 159523 44683 160500
rect 47667 161500 47690 162507
rect 47850 162507 50880 162530
rect 47850 161500 47873 162507
rect 47667 160500 47873 161500
rect 47667 159523 47690 160500
rect 44660 159500 47690 159523
rect 47850 159523 47873 160500
rect 50857 161500 50880 162507
rect 51040 162507 54070 162530
rect 51040 161500 51063 162507
rect 50857 160500 51063 161500
rect 50857 159523 50880 160500
rect 47850 159500 50880 159523
rect 51040 159523 51063 160500
rect 54047 161500 54070 162507
rect 54230 162507 57260 162530
rect 54230 161500 54253 162507
rect 54047 160500 54253 161500
rect 54047 159523 54070 160500
rect 51040 159500 54070 159523
rect 54230 159523 54253 160500
rect 57237 161500 57260 162507
rect 57420 162507 60450 162530
rect 57420 161500 57443 162507
rect 57237 160500 57443 161500
rect 57237 159523 57260 160500
rect 54230 159500 57260 159523
rect 57420 159523 57443 160500
rect 60427 161500 60450 162507
rect 60610 162507 63640 162530
rect 60610 161500 60633 162507
rect 60427 160500 60633 161500
rect 60427 159523 60450 160500
rect 57420 159500 60450 159523
rect 60610 159523 60633 160500
rect 63617 161500 63640 162507
rect 63800 162507 66830 162530
rect 63800 161500 63823 162507
rect 63617 160500 63823 161500
rect 63617 159523 63640 160500
rect 60610 159500 63640 159523
rect 63800 159523 63823 160500
rect 66807 161500 66830 162507
rect 66990 162507 70020 162530
rect 66990 161500 67013 162507
rect 66807 160500 67013 161500
rect 66807 159523 66830 160500
rect 63800 159500 66830 159523
rect 66990 159523 67013 160500
rect 69997 161500 70020 162507
rect 70180 162507 73210 162530
rect 70180 161500 70203 162507
rect 69997 160500 70203 161500
rect 69997 159523 70020 160500
rect 66990 159500 70020 159523
rect 70180 159523 70203 160500
rect 73187 161500 73210 162507
rect 73370 162507 76400 162530
rect 73370 161500 73393 162507
rect 73187 160500 73393 161500
rect 73187 159523 73210 160500
rect 70180 159500 73210 159523
rect 73370 159523 73393 160500
rect 76377 161500 76400 162507
rect 76560 162507 79590 162530
rect 76560 161500 76583 162507
rect 76377 160500 76583 161500
rect 76377 159523 76400 160500
rect 73370 159500 76400 159523
rect 76560 159523 76583 160500
rect 79567 161500 79590 162507
rect 79750 162507 82780 162530
rect 79750 161500 79773 162507
rect 79567 160500 79773 161500
rect 79567 159523 79590 160500
rect 76560 159500 79590 159523
rect 79750 159523 79773 160500
rect 82757 161500 82780 162507
rect 82940 162507 85970 162530
rect 82940 161500 82963 162507
rect 82757 160500 82963 161500
rect 82757 159523 82780 160500
rect 79750 159500 82780 159523
rect 82940 159523 82963 160500
rect 85947 161500 85970 162507
rect 86130 162507 89160 162530
rect 86130 161500 86153 162507
rect 85947 160500 86153 161500
rect 85947 159523 85970 160500
rect 82940 159500 85970 159523
rect 86130 159523 86153 160500
rect 89137 161500 89160 162507
rect 89320 162507 92350 162530
rect 89320 161500 89343 162507
rect 89137 160500 89343 161500
rect 89137 159523 89160 160500
rect 86130 159500 89160 159523
rect 89320 159523 89343 160500
rect 92327 161500 92350 162507
rect 92510 162507 95540 162530
rect 92510 161500 92533 162507
rect 92327 160500 92533 161500
rect 92327 159523 92350 160500
rect 89320 159500 92350 159523
rect 92510 159523 92533 160500
rect 95517 161500 95540 162507
rect 95700 162507 98730 162530
rect 95700 161500 95723 162507
rect 95517 160500 95723 161500
rect 95517 159523 95540 160500
rect 92510 159500 95540 159523
rect 95700 159523 95723 160500
rect 98707 161500 98730 162507
rect 98890 162507 101920 162530
rect 98890 161500 98913 162507
rect 98707 160500 98913 161500
rect 98707 159523 98730 160500
rect 95700 159500 98730 159523
rect 98890 159523 98913 160500
rect 101897 161500 101920 162507
rect 102080 162507 105110 162530
rect 102080 161500 102103 162507
rect 101897 160500 102103 161500
rect 101897 159523 101920 160500
rect 98890 159500 101920 159523
rect 102080 159523 102103 160500
rect 105087 161500 105110 162507
rect 105270 162507 108300 162530
rect 105270 161500 105293 162507
rect 105087 160500 105293 161500
rect 105087 159523 105110 160500
rect 102080 159500 105110 159523
rect 105270 159523 105293 160500
rect 108277 161500 108300 162507
rect 108460 162507 111490 162530
rect 108460 161500 108483 162507
rect 108277 160500 108483 161500
rect 108277 159523 108300 160500
rect 105270 159500 108300 159523
rect 108460 159523 108483 160500
rect 111467 161500 111490 162507
rect 111650 162507 114680 162530
rect 111650 161500 111673 162507
rect 111467 160500 111673 161500
rect 111467 159523 111490 160500
rect 108460 159500 111490 159523
rect 111650 159523 111673 160500
rect 114657 161500 114680 162507
rect 114840 162507 117870 162530
rect 114840 161500 114863 162507
rect 114657 160500 114863 161500
rect 114657 159523 114680 160500
rect 111650 159500 114680 159523
rect 114840 159523 114863 160500
rect 117847 161500 117870 162507
rect 118030 162507 121060 162530
rect 118030 161500 118053 162507
rect 117847 160500 118053 161500
rect 117847 159523 117870 160500
rect 114840 159500 117870 159523
rect 118030 159523 118053 160500
rect 121037 161500 121060 162507
rect 121220 162507 124250 162530
rect 121220 161500 121243 162507
rect 121037 160500 121243 161500
rect 121037 159523 121060 160500
rect 118030 159500 121060 159523
rect 121220 159523 121243 160500
rect 124227 161500 124250 162507
rect 124410 162507 127440 162530
rect 124410 161500 124433 162507
rect 124227 160500 124433 161500
rect 124227 159523 124250 160500
rect 121220 159500 124250 159523
rect 124410 159523 124433 160500
rect 127417 161500 127440 162507
rect 127600 162507 130630 162530
rect 127600 161500 127623 162507
rect 127417 160500 127623 161500
rect 127417 159523 127440 160500
rect 124410 159500 127440 159523
rect 127600 159523 127623 160500
rect 130607 161500 130630 162507
rect 130790 162507 133820 162530
rect 130790 161500 130813 162507
rect 130607 160500 130813 161500
rect 130607 159523 130630 160500
rect 127600 159500 130630 159523
rect 130790 159523 130813 160500
rect 133797 161500 133820 162507
rect 133980 162507 137010 162530
rect 133980 161500 134003 162507
rect 133797 160500 134003 161500
rect 133797 159523 133820 160500
rect 130790 159500 133820 159523
rect 133980 159523 134003 160500
rect 136987 161500 137010 162507
rect 136987 160500 137170 161500
rect 136987 159523 137010 160500
rect 133980 159500 137010 159523
rect 1000 159340 2000 159500
rect 4190 159340 5190 159500
rect 7380 159340 8380 159500
rect 10570 159340 11570 159500
rect 13760 159340 14760 159500
rect 16950 159340 17950 159500
rect 20140 159340 21140 159500
rect 23330 159340 24330 159500
rect 26520 159340 27520 159500
rect 29710 159340 30710 159500
rect 32900 159340 33900 159500
rect 36090 159340 37090 159500
rect 39280 159340 40280 159500
rect 42470 159340 43470 159500
rect 45660 159340 46660 159500
rect 48850 159340 49850 159500
rect 52040 159340 53040 159500
rect 55230 159340 56230 159500
rect 58420 159340 59420 159500
rect 61610 159340 62610 159500
rect 64800 159340 65800 159500
rect 67990 159340 68990 159500
rect 71180 159340 72180 159500
rect 74370 159340 75370 159500
rect 77560 159340 78560 159500
rect 80750 159340 81750 159500
rect 83940 159340 84940 159500
rect 87130 159340 88130 159500
rect 90320 159340 91320 159500
rect 93510 159340 94510 159500
rect 96700 159340 97700 159500
rect 99890 159340 100890 159500
rect 103080 159340 104080 159500
rect 106270 159340 107270 159500
rect 109460 159340 110460 159500
rect 112650 159340 113650 159500
rect 115840 159340 116840 159500
rect 119030 159340 120030 159500
rect 122220 159340 123220 159500
rect 125410 159340 126410 159500
rect 128600 159340 129600 159500
rect 131790 159340 132790 159500
rect 134980 159340 135980 159500
rect 0 159317 3030 159340
rect 0 156333 23 159317
rect 3007 158310 3030 159317
rect 3190 159317 6220 159340
rect 3190 158310 3213 159317
rect 3007 157310 3213 158310
rect 3007 156333 3030 157310
rect 0 156310 3030 156333
rect 3190 156333 3213 157310
rect 6197 158310 6220 159317
rect 6380 159317 9410 159340
rect 6380 158310 6403 159317
rect 6197 157310 6403 158310
rect 6197 156333 6220 157310
rect 3190 156310 6220 156333
rect 6380 156333 6403 157310
rect 9387 158310 9410 159317
rect 9570 159317 12600 159340
rect 9570 158310 9593 159317
rect 9387 157310 9593 158310
rect 9387 156333 9410 157310
rect 6380 156310 9410 156333
rect 9570 156333 9593 157310
rect 12577 158310 12600 159317
rect 12760 159317 15790 159340
rect 12760 158310 12783 159317
rect 12577 157310 12783 158310
rect 12577 156333 12600 157310
rect 9570 156310 12600 156333
rect 12760 156333 12783 157310
rect 15767 158310 15790 159317
rect 15950 159317 18980 159340
rect 15950 158310 15973 159317
rect 15767 157310 15973 158310
rect 15767 156333 15790 157310
rect 12760 156310 15790 156333
rect 15950 156333 15973 157310
rect 18957 158310 18980 159317
rect 19140 159317 22170 159340
rect 19140 158310 19163 159317
rect 18957 157310 19163 158310
rect 18957 156333 18980 157310
rect 15950 156310 18980 156333
rect 19140 156333 19163 157310
rect 22147 158310 22170 159317
rect 22330 159317 25360 159340
rect 22330 158310 22353 159317
rect 22147 157310 22353 158310
rect 22147 156333 22170 157310
rect 19140 156310 22170 156333
rect 22330 156333 22353 157310
rect 25337 158310 25360 159317
rect 25520 159317 28550 159340
rect 25520 158310 25543 159317
rect 25337 157310 25543 158310
rect 25337 156333 25360 157310
rect 22330 156310 25360 156333
rect 25520 156333 25543 157310
rect 28527 158310 28550 159317
rect 28710 159317 31740 159340
rect 28710 158310 28733 159317
rect 28527 157310 28733 158310
rect 28527 156333 28550 157310
rect 25520 156310 28550 156333
rect 28710 156333 28733 157310
rect 31717 158310 31740 159317
rect 31900 159317 34930 159340
rect 31900 158310 31923 159317
rect 31717 157310 31923 158310
rect 31717 156333 31740 157310
rect 28710 156310 31740 156333
rect 31900 156333 31923 157310
rect 34907 158310 34930 159317
rect 35090 159317 38120 159340
rect 35090 158310 35113 159317
rect 34907 157310 35113 158310
rect 34907 156333 34930 157310
rect 31900 156310 34930 156333
rect 35090 156333 35113 157310
rect 38097 158310 38120 159317
rect 38280 159317 41310 159340
rect 38280 158310 38303 159317
rect 38097 157310 38303 158310
rect 38097 156333 38120 157310
rect 35090 156310 38120 156333
rect 38280 156333 38303 157310
rect 41287 158310 41310 159317
rect 41470 159317 44500 159340
rect 41470 158310 41493 159317
rect 41287 157310 41493 158310
rect 41287 156333 41310 157310
rect 38280 156310 41310 156333
rect 41470 156333 41493 157310
rect 44477 158310 44500 159317
rect 44660 159317 47690 159340
rect 44660 158310 44683 159317
rect 44477 157310 44683 158310
rect 44477 156333 44500 157310
rect 41470 156310 44500 156333
rect 44660 156333 44683 157310
rect 47667 158310 47690 159317
rect 47850 159317 50880 159340
rect 47850 158310 47873 159317
rect 47667 157310 47873 158310
rect 47667 156333 47690 157310
rect 44660 156310 47690 156333
rect 47850 156333 47873 157310
rect 50857 158310 50880 159317
rect 51040 159317 54070 159340
rect 51040 158310 51063 159317
rect 50857 157310 51063 158310
rect 50857 156333 50880 157310
rect 47850 156310 50880 156333
rect 51040 156333 51063 157310
rect 54047 158310 54070 159317
rect 54230 159317 57260 159340
rect 54230 158310 54253 159317
rect 54047 157310 54253 158310
rect 54047 156333 54070 157310
rect 51040 156310 54070 156333
rect 54230 156333 54253 157310
rect 57237 158310 57260 159317
rect 57420 159317 60450 159340
rect 57420 158310 57443 159317
rect 57237 157310 57443 158310
rect 57237 156333 57260 157310
rect 54230 156310 57260 156333
rect 57420 156333 57443 157310
rect 60427 158310 60450 159317
rect 60610 159317 63640 159340
rect 60610 158310 60633 159317
rect 60427 157310 60633 158310
rect 60427 156333 60450 157310
rect 57420 156310 60450 156333
rect 60610 156333 60633 157310
rect 63617 158310 63640 159317
rect 63800 159317 66830 159340
rect 63800 158310 63823 159317
rect 63617 157310 63823 158310
rect 63617 156333 63640 157310
rect 60610 156310 63640 156333
rect 63800 156333 63823 157310
rect 66807 158310 66830 159317
rect 66990 159317 70020 159340
rect 66990 158310 67013 159317
rect 66807 157310 67013 158310
rect 66807 156333 66830 157310
rect 63800 156310 66830 156333
rect 66990 156333 67013 157310
rect 69997 158310 70020 159317
rect 70180 159317 73210 159340
rect 70180 158310 70203 159317
rect 69997 157310 70203 158310
rect 69997 156333 70020 157310
rect 66990 156310 70020 156333
rect 70180 156333 70203 157310
rect 73187 158310 73210 159317
rect 73370 159317 76400 159340
rect 73370 158310 73393 159317
rect 73187 157310 73393 158310
rect 73187 156333 73210 157310
rect 70180 156310 73210 156333
rect 73370 156333 73393 157310
rect 76377 158310 76400 159317
rect 76560 159317 79590 159340
rect 76560 158310 76583 159317
rect 76377 157310 76583 158310
rect 76377 156333 76400 157310
rect 73370 156310 76400 156333
rect 76560 156333 76583 157310
rect 79567 158310 79590 159317
rect 79750 159317 82780 159340
rect 79750 158310 79773 159317
rect 79567 157310 79773 158310
rect 79567 156333 79590 157310
rect 76560 156310 79590 156333
rect 79750 156333 79773 157310
rect 82757 158310 82780 159317
rect 82940 159317 85970 159340
rect 82940 158310 82963 159317
rect 82757 157310 82963 158310
rect 82757 156333 82780 157310
rect 79750 156310 82780 156333
rect 82940 156333 82963 157310
rect 85947 158310 85970 159317
rect 86130 159317 89160 159340
rect 86130 158310 86153 159317
rect 85947 157310 86153 158310
rect 85947 156333 85970 157310
rect 82940 156310 85970 156333
rect 86130 156333 86153 157310
rect 89137 158310 89160 159317
rect 89320 159317 92350 159340
rect 89320 158310 89343 159317
rect 89137 157310 89343 158310
rect 89137 156333 89160 157310
rect 86130 156310 89160 156333
rect 89320 156333 89343 157310
rect 92327 158310 92350 159317
rect 92510 159317 95540 159340
rect 92510 158310 92533 159317
rect 92327 157310 92533 158310
rect 92327 156333 92350 157310
rect 89320 156310 92350 156333
rect 92510 156333 92533 157310
rect 95517 158310 95540 159317
rect 95700 159317 98730 159340
rect 95700 158310 95723 159317
rect 95517 157310 95723 158310
rect 95517 156333 95540 157310
rect 92510 156310 95540 156333
rect 95700 156333 95723 157310
rect 98707 158310 98730 159317
rect 98890 159317 101920 159340
rect 98890 158310 98913 159317
rect 98707 157310 98913 158310
rect 98707 156333 98730 157310
rect 95700 156310 98730 156333
rect 98890 156333 98913 157310
rect 101897 158310 101920 159317
rect 102080 159317 105110 159340
rect 102080 158310 102103 159317
rect 101897 157310 102103 158310
rect 101897 156333 101920 157310
rect 98890 156310 101920 156333
rect 102080 156333 102103 157310
rect 105087 158310 105110 159317
rect 105270 159317 108300 159340
rect 105270 158310 105293 159317
rect 105087 157310 105293 158310
rect 105087 156333 105110 157310
rect 102080 156310 105110 156333
rect 105270 156333 105293 157310
rect 108277 158310 108300 159317
rect 108460 159317 111490 159340
rect 108460 158310 108483 159317
rect 108277 157310 108483 158310
rect 108277 156333 108300 157310
rect 105270 156310 108300 156333
rect 108460 156333 108483 157310
rect 111467 158310 111490 159317
rect 111650 159317 114680 159340
rect 111650 158310 111673 159317
rect 111467 157310 111673 158310
rect 111467 156333 111490 157310
rect 108460 156310 111490 156333
rect 111650 156333 111673 157310
rect 114657 158310 114680 159317
rect 114840 159317 117870 159340
rect 114840 158310 114863 159317
rect 114657 157310 114863 158310
rect 114657 156333 114680 157310
rect 111650 156310 114680 156333
rect 114840 156333 114863 157310
rect 117847 158310 117870 159317
rect 118030 159317 121060 159340
rect 118030 158310 118053 159317
rect 117847 157310 118053 158310
rect 117847 156333 117870 157310
rect 114840 156310 117870 156333
rect 118030 156333 118053 157310
rect 121037 158310 121060 159317
rect 121220 159317 124250 159340
rect 121220 158310 121243 159317
rect 121037 157310 121243 158310
rect 121037 156333 121060 157310
rect 118030 156310 121060 156333
rect 121220 156333 121243 157310
rect 124227 158310 124250 159317
rect 124410 159317 127440 159340
rect 124410 158310 124433 159317
rect 124227 157310 124433 158310
rect 124227 156333 124250 157310
rect 121220 156310 124250 156333
rect 124410 156333 124433 157310
rect 127417 158310 127440 159317
rect 127600 159317 130630 159340
rect 127600 158310 127623 159317
rect 127417 157310 127623 158310
rect 127417 156333 127440 157310
rect 124410 156310 127440 156333
rect 127600 156333 127623 157310
rect 130607 158310 130630 159317
rect 130790 159317 133820 159340
rect 130790 158310 130813 159317
rect 130607 157310 130813 158310
rect 130607 156333 130630 157310
rect 127600 156310 130630 156333
rect 130790 156333 130813 157310
rect 133797 158310 133820 159317
rect 133980 159317 137010 159340
rect 133980 158310 134003 159317
rect 133797 157310 134003 158310
rect 133797 156333 133820 157310
rect 130790 156310 133820 156333
rect 133980 156333 134003 157310
rect 136987 158310 137010 159317
rect 136987 157310 137170 158310
rect 136987 156333 137010 157310
rect 133980 156310 137010 156333
rect 1000 156150 2000 156310
rect 4190 156150 5190 156310
rect 7380 156150 8380 156310
rect 10570 156150 11570 156310
rect 13760 156150 14760 156310
rect 16950 156150 17950 156310
rect 20140 156150 21140 156310
rect 23330 156150 24330 156310
rect 26520 156150 27520 156310
rect 29710 156150 30710 156310
rect 32900 156150 33900 156310
rect 36090 156150 37090 156310
rect 39280 156150 40280 156310
rect 42470 156150 43470 156310
rect 45660 156150 46660 156310
rect 48850 156150 49850 156310
rect 52040 156150 53040 156310
rect 55230 156150 56230 156310
rect 58420 156150 59420 156310
rect 61610 156150 62610 156310
rect 64800 156150 65800 156310
rect 67990 156150 68990 156310
rect 71180 156150 72180 156310
rect 74370 156150 75370 156310
rect 77560 156150 78560 156310
rect 80750 156150 81750 156310
rect 83940 156150 84940 156310
rect 87130 156150 88130 156310
rect 90320 156150 91320 156310
rect 93510 156150 94510 156310
rect 96700 156150 97700 156310
rect 99890 156150 100890 156310
rect 103080 156150 104080 156310
rect 106270 156150 107270 156310
rect 109460 156150 110460 156310
rect 112650 156150 113650 156310
rect 115840 156150 116840 156310
rect 119030 156150 120030 156310
rect 122220 156150 123220 156310
rect 125410 156150 126410 156310
rect 128600 156150 129600 156310
rect 131790 156150 132790 156310
rect 134980 156150 135980 156310
rect 0 156127 3030 156150
rect 0 153143 23 156127
rect 3007 155120 3030 156127
rect 3190 156127 6220 156150
rect 3190 155120 3213 156127
rect 3007 154120 3213 155120
rect 3007 153143 3030 154120
rect 0 153120 3030 153143
rect 3190 153143 3213 154120
rect 6197 155120 6220 156127
rect 6380 156127 9410 156150
rect 6380 155120 6403 156127
rect 6197 154120 6403 155120
rect 6197 153143 6220 154120
rect 3190 153120 6220 153143
rect 6380 153143 6403 154120
rect 9387 155120 9410 156127
rect 9570 156127 12600 156150
rect 9570 155120 9593 156127
rect 9387 154120 9593 155120
rect 9387 153143 9410 154120
rect 6380 153120 9410 153143
rect 9570 153143 9593 154120
rect 12577 155120 12600 156127
rect 12760 156127 15790 156150
rect 12760 155120 12783 156127
rect 12577 154120 12783 155120
rect 12577 153143 12600 154120
rect 9570 153120 12600 153143
rect 12760 153143 12783 154120
rect 15767 155120 15790 156127
rect 15950 156127 18980 156150
rect 15950 155120 15973 156127
rect 15767 154120 15973 155120
rect 15767 153143 15790 154120
rect 12760 153120 15790 153143
rect 15950 153143 15973 154120
rect 18957 155120 18980 156127
rect 19140 156127 22170 156150
rect 19140 155120 19163 156127
rect 18957 154120 19163 155120
rect 18957 153143 18980 154120
rect 15950 153120 18980 153143
rect 19140 153143 19163 154120
rect 22147 155120 22170 156127
rect 22330 156127 25360 156150
rect 22330 155120 22353 156127
rect 22147 154120 22353 155120
rect 22147 153143 22170 154120
rect 19140 153120 22170 153143
rect 22330 153143 22353 154120
rect 25337 155120 25360 156127
rect 25520 156127 28550 156150
rect 25520 155120 25543 156127
rect 25337 154120 25543 155120
rect 25337 153143 25360 154120
rect 22330 153120 25360 153143
rect 25520 153143 25543 154120
rect 28527 155120 28550 156127
rect 28710 156127 31740 156150
rect 28710 155120 28733 156127
rect 28527 154120 28733 155120
rect 28527 153143 28550 154120
rect 25520 153120 28550 153143
rect 28710 153143 28733 154120
rect 31717 155120 31740 156127
rect 31900 156127 34930 156150
rect 31900 155120 31923 156127
rect 31717 154120 31923 155120
rect 31717 153143 31740 154120
rect 28710 153120 31740 153143
rect 31900 153143 31923 154120
rect 34907 155120 34930 156127
rect 35090 156127 38120 156150
rect 35090 155120 35113 156127
rect 34907 154120 35113 155120
rect 34907 153143 34930 154120
rect 31900 153120 34930 153143
rect 35090 153143 35113 154120
rect 38097 155120 38120 156127
rect 38280 156127 41310 156150
rect 38280 155120 38303 156127
rect 38097 154120 38303 155120
rect 38097 153143 38120 154120
rect 35090 153120 38120 153143
rect 38280 153143 38303 154120
rect 41287 155120 41310 156127
rect 41470 156127 44500 156150
rect 41470 155120 41493 156127
rect 41287 154120 41493 155120
rect 41287 153143 41310 154120
rect 38280 153120 41310 153143
rect 41470 153143 41493 154120
rect 44477 155120 44500 156127
rect 44660 156127 47690 156150
rect 44660 155120 44683 156127
rect 44477 154120 44683 155120
rect 44477 153143 44500 154120
rect 41470 153120 44500 153143
rect 44660 153143 44683 154120
rect 47667 155120 47690 156127
rect 47850 156127 50880 156150
rect 47850 155120 47873 156127
rect 47667 154120 47873 155120
rect 47667 153143 47690 154120
rect 44660 153120 47690 153143
rect 47850 153143 47873 154120
rect 50857 155120 50880 156127
rect 51040 156127 54070 156150
rect 51040 155120 51063 156127
rect 50857 154120 51063 155120
rect 50857 153143 50880 154120
rect 47850 153120 50880 153143
rect 51040 153143 51063 154120
rect 54047 155120 54070 156127
rect 54230 156127 57260 156150
rect 54230 155120 54253 156127
rect 54047 154120 54253 155120
rect 54047 153143 54070 154120
rect 51040 153120 54070 153143
rect 54230 153143 54253 154120
rect 57237 155120 57260 156127
rect 57420 156127 60450 156150
rect 57420 155120 57443 156127
rect 57237 154120 57443 155120
rect 57237 153143 57260 154120
rect 54230 153120 57260 153143
rect 57420 153143 57443 154120
rect 60427 155120 60450 156127
rect 60610 156127 63640 156150
rect 60610 155120 60633 156127
rect 60427 154120 60633 155120
rect 60427 153143 60450 154120
rect 57420 153120 60450 153143
rect 60610 153143 60633 154120
rect 63617 155120 63640 156127
rect 63800 156127 66830 156150
rect 63800 155120 63823 156127
rect 63617 154120 63823 155120
rect 63617 153143 63640 154120
rect 60610 153120 63640 153143
rect 63800 153143 63823 154120
rect 66807 155120 66830 156127
rect 66990 156127 70020 156150
rect 66990 155120 67013 156127
rect 66807 154120 67013 155120
rect 66807 153143 66830 154120
rect 63800 153120 66830 153143
rect 66990 153143 67013 154120
rect 69997 155120 70020 156127
rect 70180 156127 73210 156150
rect 70180 155120 70203 156127
rect 69997 154120 70203 155120
rect 69997 153143 70020 154120
rect 66990 153120 70020 153143
rect 70180 153143 70203 154120
rect 73187 155120 73210 156127
rect 73370 156127 76400 156150
rect 73370 155120 73393 156127
rect 73187 154120 73393 155120
rect 73187 153143 73210 154120
rect 70180 153120 73210 153143
rect 73370 153143 73393 154120
rect 76377 155120 76400 156127
rect 76560 156127 79590 156150
rect 76560 155120 76583 156127
rect 76377 154120 76583 155120
rect 76377 153143 76400 154120
rect 73370 153120 76400 153143
rect 76560 153143 76583 154120
rect 79567 155120 79590 156127
rect 79750 156127 82780 156150
rect 79750 155120 79773 156127
rect 79567 154120 79773 155120
rect 79567 153143 79590 154120
rect 76560 153120 79590 153143
rect 79750 153143 79773 154120
rect 82757 155120 82780 156127
rect 82940 156127 85970 156150
rect 82940 155120 82963 156127
rect 82757 154120 82963 155120
rect 82757 153143 82780 154120
rect 79750 153120 82780 153143
rect 82940 153143 82963 154120
rect 85947 155120 85970 156127
rect 86130 156127 89160 156150
rect 86130 155120 86153 156127
rect 85947 154120 86153 155120
rect 85947 153143 85970 154120
rect 82940 153120 85970 153143
rect 86130 153143 86153 154120
rect 89137 155120 89160 156127
rect 89320 156127 92350 156150
rect 89320 155120 89343 156127
rect 89137 154120 89343 155120
rect 89137 153143 89160 154120
rect 86130 153120 89160 153143
rect 89320 153143 89343 154120
rect 92327 155120 92350 156127
rect 92510 156127 95540 156150
rect 92510 155120 92533 156127
rect 92327 154120 92533 155120
rect 92327 153143 92350 154120
rect 89320 153120 92350 153143
rect 92510 153143 92533 154120
rect 95517 155120 95540 156127
rect 95700 156127 98730 156150
rect 95700 155120 95723 156127
rect 95517 154120 95723 155120
rect 95517 153143 95540 154120
rect 92510 153120 95540 153143
rect 95700 153143 95723 154120
rect 98707 155120 98730 156127
rect 98890 156127 101920 156150
rect 98890 155120 98913 156127
rect 98707 154120 98913 155120
rect 98707 153143 98730 154120
rect 95700 153120 98730 153143
rect 98890 153143 98913 154120
rect 101897 155120 101920 156127
rect 102080 156127 105110 156150
rect 102080 155120 102103 156127
rect 101897 154120 102103 155120
rect 101897 153143 101920 154120
rect 98890 153120 101920 153143
rect 102080 153143 102103 154120
rect 105087 155120 105110 156127
rect 105270 156127 108300 156150
rect 105270 155120 105293 156127
rect 105087 154120 105293 155120
rect 105087 153143 105110 154120
rect 102080 153120 105110 153143
rect 105270 153143 105293 154120
rect 108277 155120 108300 156127
rect 108460 156127 111490 156150
rect 108460 155120 108483 156127
rect 108277 154120 108483 155120
rect 108277 153143 108300 154120
rect 105270 153120 108300 153143
rect 108460 153143 108483 154120
rect 111467 155120 111490 156127
rect 111650 156127 114680 156150
rect 111650 155120 111673 156127
rect 111467 154120 111673 155120
rect 111467 153143 111490 154120
rect 108460 153120 111490 153143
rect 111650 153143 111673 154120
rect 114657 155120 114680 156127
rect 114840 156127 117870 156150
rect 114840 155120 114863 156127
rect 114657 154120 114863 155120
rect 114657 153143 114680 154120
rect 111650 153120 114680 153143
rect 114840 153143 114863 154120
rect 117847 155120 117870 156127
rect 118030 156127 121060 156150
rect 118030 155120 118053 156127
rect 117847 154120 118053 155120
rect 117847 153143 117870 154120
rect 114840 153120 117870 153143
rect 118030 153143 118053 154120
rect 121037 155120 121060 156127
rect 121220 156127 124250 156150
rect 121220 155120 121243 156127
rect 121037 154120 121243 155120
rect 121037 153143 121060 154120
rect 118030 153120 121060 153143
rect 121220 153143 121243 154120
rect 124227 155120 124250 156127
rect 124410 156127 127440 156150
rect 124410 155120 124433 156127
rect 124227 154120 124433 155120
rect 124227 153143 124250 154120
rect 121220 153120 124250 153143
rect 124410 153143 124433 154120
rect 127417 155120 127440 156127
rect 127600 156127 130630 156150
rect 127600 155120 127623 156127
rect 127417 154120 127623 155120
rect 127417 153143 127440 154120
rect 124410 153120 127440 153143
rect 127600 153143 127623 154120
rect 130607 155120 130630 156127
rect 130790 156127 133820 156150
rect 130790 155120 130813 156127
rect 130607 154120 130813 155120
rect 130607 153143 130630 154120
rect 127600 153120 130630 153143
rect 130790 153143 130813 154120
rect 133797 155120 133820 156127
rect 133980 156127 137010 156150
rect 133980 155120 134003 156127
rect 133797 154120 134003 155120
rect 133797 153143 133820 154120
rect 130790 153120 133820 153143
rect 133980 153143 134003 154120
rect 136987 155120 137010 156127
rect 136987 154120 137170 155120
rect 136987 153143 137010 154120
rect 133980 153120 137010 153143
rect 1000 152960 2000 153120
rect 4190 152960 5190 153120
rect 7380 152960 8380 153120
rect 10570 152960 11570 153120
rect 13760 152960 14760 153120
rect 16950 152960 17950 153120
rect 20140 152960 21140 153120
rect 23330 152960 24330 153120
rect 26520 152960 27520 153120
rect 29710 152960 30710 153120
rect 32900 152960 33900 153120
rect 36090 152960 37090 153120
rect 39280 152960 40280 153120
rect 42470 152960 43470 153120
rect 45660 152960 46660 153120
rect 48850 152960 49850 153120
rect 52040 152960 53040 153120
rect 55230 152960 56230 153120
rect 58420 152960 59420 153120
rect 61610 152960 62610 153120
rect 64800 152960 65800 153120
rect 67990 152960 68990 153120
rect 71180 152960 72180 153120
rect 74370 152960 75370 153120
rect 77560 152960 78560 153120
rect 80750 152960 81750 153120
rect 83940 152960 84940 153120
rect 87130 152960 88130 153120
rect 90320 152960 91320 153120
rect 93510 152960 94510 153120
rect 96700 152960 97700 153120
rect 99890 152960 100890 153120
rect 103080 152960 104080 153120
rect 106270 152960 107270 153120
rect 109460 152960 110460 153120
rect 112650 152960 113650 153120
rect 115840 152960 116840 153120
rect 119030 152960 120030 153120
rect 122220 152960 123220 153120
rect 125410 152960 126410 153120
rect 128600 152960 129600 153120
rect 131790 152960 132790 153120
rect 134980 152960 135980 153120
rect 0 152937 3030 152960
rect 0 149953 23 152937
rect 3007 151930 3030 152937
rect 3190 152937 6220 152960
rect 3190 151930 3213 152937
rect 3007 150930 3213 151930
rect 3007 149953 3030 150930
rect 0 149930 3030 149953
rect 3190 149953 3213 150930
rect 6197 151930 6220 152937
rect 6380 152937 9410 152960
rect 6380 151930 6403 152937
rect 6197 150930 6403 151930
rect 6197 149953 6220 150930
rect 3190 149930 6220 149953
rect 6380 149953 6403 150930
rect 9387 151930 9410 152937
rect 9570 152937 12600 152960
rect 9570 151930 9593 152937
rect 9387 150930 9593 151930
rect 9387 149953 9410 150930
rect 6380 149930 9410 149953
rect 9570 149953 9593 150930
rect 12577 151930 12600 152937
rect 12760 152937 15790 152960
rect 12760 151930 12783 152937
rect 12577 150930 12783 151930
rect 12577 149953 12600 150930
rect 9570 149930 12600 149953
rect 12760 149953 12783 150930
rect 15767 151930 15790 152937
rect 15950 152937 18980 152960
rect 15950 151930 15973 152937
rect 15767 150930 15973 151930
rect 15767 149953 15790 150930
rect 12760 149930 15790 149953
rect 15950 149953 15973 150930
rect 18957 151930 18980 152937
rect 19140 152937 22170 152960
rect 19140 151930 19163 152937
rect 18957 150930 19163 151930
rect 18957 149953 18980 150930
rect 15950 149930 18980 149953
rect 19140 149953 19163 150930
rect 22147 151930 22170 152937
rect 22330 152937 25360 152960
rect 22330 151930 22353 152937
rect 22147 150930 22353 151930
rect 22147 149953 22170 150930
rect 19140 149930 22170 149953
rect 22330 149953 22353 150930
rect 25337 151930 25360 152937
rect 25520 152937 28550 152960
rect 25520 151930 25543 152937
rect 25337 150930 25543 151930
rect 25337 149953 25360 150930
rect 22330 149930 25360 149953
rect 25520 149953 25543 150930
rect 28527 151930 28550 152937
rect 28710 152937 31740 152960
rect 28710 151930 28733 152937
rect 28527 150930 28733 151930
rect 28527 149953 28550 150930
rect 25520 149930 28550 149953
rect 28710 149953 28733 150930
rect 31717 151930 31740 152937
rect 31900 152937 34930 152960
rect 31900 151930 31923 152937
rect 31717 150930 31923 151930
rect 31717 149953 31740 150930
rect 28710 149930 31740 149953
rect 31900 149953 31923 150930
rect 34907 151930 34930 152937
rect 35090 152937 38120 152960
rect 35090 151930 35113 152937
rect 34907 150930 35113 151930
rect 34907 149953 34930 150930
rect 31900 149930 34930 149953
rect 35090 149953 35113 150930
rect 38097 151930 38120 152937
rect 38280 152937 41310 152960
rect 38280 151930 38303 152937
rect 38097 150930 38303 151930
rect 38097 149953 38120 150930
rect 35090 149930 38120 149953
rect 38280 149953 38303 150930
rect 41287 151930 41310 152937
rect 41470 152937 44500 152960
rect 41470 151930 41493 152937
rect 41287 150930 41493 151930
rect 41287 149953 41310 150930
rect 38280 149930 41310 149953
rect 41470 149953 41493 150930
rect 44477 151930 44500 152937
rect 44660 152937 47690 152960
rect 44660 151930 44683 152937
rect 44477 150930 44683 151930
rect 44477 149953 44500 150930
rect 41470 149930 44500 149953
rect 44660 149953 44683 150930
rect 47667 151930 47690 152937
rect 47850 152937 50880 152960
rect 47850 151930 47873 152937
rect 47667 150930 47873 151930
rect 47667 149953 47690 150930
rect 44660 149930 47690 149953
rect 47850 149953 47873 150930
rect 50857 151930 50880 152937
rect 51040 152937 54070 152960
rect 51040 151930 51063 152937
rect 50857 150930 51063 151930
rect 50857 149953 50880 150930
rect 47850 149930 50880 149953
rect 51040 149953 51063 150930
rect 54047 151930 54070 152937
rect 54230 152937 57260 152960
rect 54230 151930 54253 152937
rect 54047 150930 54253 151930
rect 54047 149953 54070 150930
rect 51040 149930 54070 149953
rect 54230 149953 54253 150930
rect 57237 151930 57260 152937
rect 57420 152937 60450 152960
rect 57420 151930 57443 152937
rect 57237 150930 57443 151930
rect 57237 149953 57260 150930
rect 54230 149930 57260 149953
rect 57420 149953 57443 150930
rect 60427 151930 60450 152937
rect 60610 152937 63640 152960
rect 60610 151930 60633 152937
rect 60427 150930 60633 151930
rect 60427 149953 60450 150930
rect 57420 149930 60450 149953
rect 60610 149953 60633 150930
rect 63617 151930 63640 152937
rect 63800 152937 66830 152960
rect 63800 151930 63823 152937
rect 63617 150930 63823 151930
rect 63617 149953 63640 150930
rect 60610 149930 63640 149953
rect 63800 149953 63823 150930
rect 66807 151930 66830 152937
rect 66990 152937 70020 152960
rect 66990 151930 67013 152937
rect 66807 150930 67013 151930
rect 66807 149953 66830 150930
rect 63800 149930 66830 149953
rect 66990 149953 67013 150930
rect 69997 151930 70020 152937
rect 70180 152937 73210 152960
rect 70180 151930 70203 152937
rect 69997 150930 70203 151930
rect 69997 149953 70020 150930
rect 66990 149930 70020 149953
rect 70180 149953 70203 150930
rect 73187 151930 73210 152937
rect 73370 152937 76400 152960
rect 73370 151930 73393 152937
rect 73187 150930 73393 151930
rect 73187 149953 73210 150930
rect 70180 149930 73210 149953
rect 73370 149953 73393 150930
rect 76377 151930 76400 152937
rect 76560 152937 79590 152960
rect 76560 151930 76583 152937
rect 76377 150930 76583 151930
rect 76377 149953 76400 150930
rect 73370 149930 76400 149953
rect 76560 149953 76583 150930
rect 79567 151930 79590 152937
rect 79750 152937 82780 152960
rect 79750 151930 79773 152937
rect 79567 150930 79773 151930
rect 79567 149953 79590 150930
rect 76560 149930 79590 149953
rect 79750 149953 79773 150930
rect 82757 151930 82780 152937
rect 82940 152937 85970 152960
rect 82940 151930 82963 152937
rect 82757 150930 82963 151930
rect 82757 149953 82780 150930
rect 79750 149930 82780 149953
rect 82940 149953 82963 150930
rect 85947 151930 85970 152937
rect 86130 152937 89160 152960
rect 86130 151930 86153 152937
rect 85947 150930 86153 151930
rect 85947 149953 85970 150930
rect 82940 149930 85970 149953
rect 86130 149953 86153 150930
rect 89137 151930 89160 152937
rect 89320 152937 92350 152960
rect 89320 151930 89343 152937
rect 89137 150930 89343 151930
rect 89137 149953 89160 150930
rect 86130 149930 89160 149953
rect 89320 149953 89343 150930
rect 92327 151930 92350 152937
rect 92510 152937 95540 152960
rect 92510 151930 92533 152937
rect 92327 150930 92533 151930
rect 92327 149953 92350 150930
rect 89320 149930 92350 149953
rect 92510 149953 92533 150930
rect 95517 151930 95540 152937
rect 95700 152937 98730 152960
rect 95700 151930 95723 152937
rect 95517 150930 95723 151930
rect 95517 149953 95540 150930
rect 92510 149930 95540 149953
rect 95700 149953 95723 150930
rect 98707 151930 98730 152937
rect 98890 152937 101920 152960
rect 98890 151930 98913 152937
rect 98707 150930 98913 151930
rect 98707 149953 98730 150930
rect 95700 149930 98730 149953
rect 98890 149953 98913 150930
rect 101897 151930 101920 152937
rect 102080 152937 105110 152960
rect 102080 151930 102103 152937
rect 101897 150930 102103 151930
rect 101897 149953 101920 150930
rect 98890 149930 101920 149953
rect 102080 149953 102103 150930
rect 105087 151930 105110 152937
rect 105270 152937 108300 152960
rect 105270 151930 105293 152937
rect 105087 150930 105293 151930
rect 105087 149953 105110 150930
rect 102080 149930 105110 149953
rect 105270 149953 105293 150930
rect 108277 151930 108300 152937
rect 108460 152937 111490 152960
rect 108460 151930 108483 152937
rect 108277 150930 108483 151930
rect 108277 149953 108300 150930
rect 105270 149930 108300 149953
rect 108460 149953 108483 150930
rect 111467 151930 111490 152937
rect 111650 152937 114680 152960
rect 111650 151930 111673 152937
rect 111467 150930 111673 151930
rect 111467 149953 111490 150930
rect 108460 149930 111490 149953
rect 111650 149953 111673 150930
rect 114657 151930 114680 152937
rect 114840 152937 117870 152960
rect 114840 151930 114863 152937
rect 114657 150930 114863 151930
rect 114657 149953 114680 150930
rect 111650 149930 114680 149953
rect 114840 149953 114863 150930
rect 117847 151930 117870 152937
rect 118030 152937 121060 152960
rect 118030 151930 118053 152937
rect 117847 150930 118053 151930
rect 117847 149953 117870 150930
rect 114840 149930 117870 149953
rect 118030 149953 118053 150930
rect 121037 151930 121060 152937
rect 121220 152937 124250 152960
rect 121220 151930 121243 152937
rect 121037 150930 121243 151930
rect 121037 149953 121060 150930
rect 118030 149930 121060 149953
rect 121220 149953 121243 150930
rect 124227 151930 124250 152937
rect 124410 152937 127440 152960
rect 124410 151930 124433 152937
rect 124227 150930 124433 151930
rect 124227 149953 124250 150930
rect 121220 149930 124250 149953
rect 124410 149953 124433 150930
rect 127417 151930 127440 152937
rect 127600 152937 130630 152960
rect 127600 151930 127623 152937
rect 127417 150930 127623 151930
rect 127417 149953 127440 150930
rect 124410 149930 127440 149953
rect 127600 149953 127623 150930
rect 130607 151930 130630 152937
rect 130790 152937 133820 152960
rect 130790 151930 130813 152937
rect 130607 150930 130813 151930
rect 130607 149953 130630 150930
rect 127600 149930 130630 149953
rect 130790 149953 130813 150930
rect 133797 151930 133820 152937
rect 133980 152937 137010 152960
rect 133980 151930 134003 152937
rect 133797 150930 134003 151930
rect 133797 149953 133820 150930
rect 130790 149930 133820 149953
rect 133980 149953 134003 150930
rect 136987 151930 137010 152937
rect 136987 150930 137170 151930
rect 136987 149953 137010 150930
rect 133980 149930 137010 149953
rect 1000 149770 2000 149930
rect 4190 149770 5190 149930
rect 7380 149770 8380 149930
rect 10570 149770 11570 149930
rect 13760 149770 14760 149930
rect 16950 149770 17950 149930
rect 20140 149770 21140 149930
rect 23330 149770 24330 149930
rect 26520 149770 27520 149930
rect 29710 149770 30710 149930
rect 32900 149770 33900 149930
rect 36090 149770 37090 149930
rect 39280 149770 40280 149930
rect 42470 149770 43470 149930
rect 45660 149770 46660 149930
rect 48850 149770 49850 149930
rect 52040 149770 53040 149930
rect 55230 149770 56230 149930
rect 58420 149770 59420 149930
rect 61610 149770 62610 149930
rect 64800 149770 65800 149930
rect 67990 149770 68990 149930
rect 71180 149770 72180 149930
rect 74370 149770 75370 149930
rect 77560 149770 78560 149930
rect 80750 149770 81750 149930
rect 83940 149770 84940 149930
rect 87130 149770 88130 149930
rect 90320 149770 91320 149930
rect 93510 149770 94510 149930
rect 96700 149770 97700 149930
rect 99890 149770 100890 149930
rect 103080 149770 104080 149930
rect 106270 149770 107270 149930
rect 109460 149770 110460 149930
rect 112650 149770 113650 149930
rect 115840 149770 116840 149930
rect 119030 149770 120030 149930
rect 122220 149770 123220 149930
rect 125410 149770 126410 149930
rect 128600 149770 129600 149930
rect 131790 149770 132790 149930
rect 134980 149770 135980 149930
rect 0 149747 3030 149770
rect 0 146763 23 149747
rect 3007 148740 3030 149747
rect 3190 149747 6220 149770
rect 3190 148740 3213 149747
rect 3007 147740 3213 148740
rect 3007 146763 3030 147740
rect 0 146740 3030 146763
rect 3190 146763 3213 147740
rect 6197 148740 6220 149747
rect 6380 149747 9410 149770
rect 6380 148740 6403 149747
rect 6197 147740 6403 148740
rect 6197 146763 6220 147740
rect 3190 146740 6220 146763
rect 6380 146763 6403 147740
rect 9387 148740 9410 149747
rect 9570 149747 12600 149770
rect 9570 148740 9593 149747
rect 9387 147740 9593 148740
rect 9387 146763 9410 147740
rect 6380 146740 9410 146763
rect 9570 146763 9593 147740
rect 12577 148740 12600 149747
rect 12760 149747 15790 149770
rect 12760 148740 12783 149747
rect 12577 147740 12783 148740
rect 12577 146763 12600 147740
rect 9570 146740 12600 146763
rect 12760 146763 12783 147740
rect 15767 148740 15790 149747
rect 15950 149747 18980 149770
rect 15950 148740 15973 149747
rect 15767 147740 15973 148740
rect 15767 146763 15790 147740
rect 12760 146740 15790 146763
rect 15950 146763 15973 147740
rect 18957 148740 18980 149747
rect 19140 149747 22170 149770
rect 19140 148740 19163 149747
rect 18957 147740 19163 148740
rect 18957 146763 18980 147740
rect 15950 146740 18980 146763
rect 19140 146763 19163 147740
rect 22147 148740 22170 149747
rect 22330 149747 25360 149770
rect 22330 148740 22353 149747
rect 22147 147740 22353 148740
rect 22147 146763 22170 147740
rect 19140 146740 22170 146763
rect 22330 146763 22353 147740
rect 25337 148740 25360 149747
rect 25520 149747 28550 149770
rect 25520 148740 25543 149747
rect 25337 147740 25543 148740
rect 25337 146763 25360 147740
rect 22330 146740 25360 146763
rect 25520 146763 25543 147740
rect 28527 148740 28550 149747
rect 28710 149747 31740 149770
rect 28710 148740 28733 149747
rect 28527 147740 28733 148740
rect 28527 146763 28550 147740
rect 25520 146740 28550 146763
rect 28710 146763 28733 147740
rect 31717 148740 31740 149747
rect 31900 149747 34930 149770
rect 31900 148740 31923 149747
rect 31717 147740 31923 148740
rect 31717 146763 31740 147740
rect 28710 146740 31740 146763
rect 31900 146763 31923 147740
rect 34907 148740 34930 149747
rect 35090 149747 38120 149770
rect 35090 148740 35113 149747
rect 34907 147740 35113 148740
rect 34907 146763 34930 147740
rect 31900 146740 34930 146763
rect 35090 146763 35113 147740
rect 38097 148740 38120 149747
rect 38280 149747 41310 149770
rect 38280 148740 38303 149747
rect 38097 147740 38303 148740
rect 38097 146763 38120 147740
rect 35090 146740 38120 146763
rect 38280 146763 38303 147740
rect 41287 148740 41310 149747
rect 41470 149747 44500 149770
rect 41470 148740 41493 149747
rect 41287 147740 41493 148740
rect 41287 146763 41310 147740
rect 38280 146740 41310 146763
rect 41470 146763 41493 147740
rect 44477 148740 44500 149747
rect 44660 149747 47690 149770
rect 44660 148740 44683 149747
rect 44477 147740 44683 148740
rect 44477 146763 44500 147740
rect 41470 146740 44500 146763
rect 44660 146763 44683 147740
rect 47667 148740 47690 149747
rect 47850 149747 50880 149770
rect 47850 148740 47873 149747
rect 47667 147740 47873 148740
rect 47667 146763 47690 147740
rect 44660 146740 47690 146763
rect 47850 146763 47873 147740
rect 50857 148740 50880 149747
rect 51040 149747 54070 149770
rect 51040 148740 51063 149747
rect 50857 147740 51063 148740
rect 50857 146763 50880 147740
rect 47850 146740 50880 146763
rect 51040 146763 51063 147740
rect 54047 148740 54070 149747
rect 54230 149747 57260 149770
rect 54230 148740 54253 149747
rect 54047 147740 54253 148740
rect 54047 146763 54070 147740
rect 51040 146740 54070 146763
rect 54230 146763 54253 147740
rect 57237 148740 57260 149747
rect 57420 149747 60450 149770
rect 57420 148740 57443 149747
rect 57237 147740 57443 148740
rect 57237 146763 57260 147740
rect 54230 146740 57260 146763
rect 57420 146763 57443 147740
rect 60427 148740 60450 149747
rect 60610 149747 63640 149770
rect 60610 148740 60633 149747
rect 60427 147740 60633 148740
rect 60427 146763 60450 147740
rect 57420 146740 60450 146763
rect 60610 146763 60633 147740
rect 63617 148740 63640 149747
rect 63800 149747 66830 149770
rect 63800 148740 63823 149747
rect 63617 147740 63823 148740
rect 63617 146763 63640 147740
rect 60610 146740 63640 146763
rect 63800 146763 63823 147740
rect 66807 148740 66830 149747
rect 66990 149747 70020 149770
rect 66990 148740 67013 149747
rect 66807 147740 67013 148740
rect 66807 146763 66830 147740
rect 63800 146740 66830 146763
rect 66990 146763 67013 147740
rect 69997 148740 70020 149747
rect 70180 149747 73210 149770
rect 70180 148740 70203 149747
rect 69997 147740 70203 148740
rect 69997 146763 70020 147740
rect 66990 146740 70020 146763
rect 70180 146763 70203 147740
rect 73187 148740 73210 149747
rect 73370 149747 76400 149770
rect 73370 148740 73393 149747
rect 73187 147740 73393 148740
rect 73187 146763 73210 147740
rect 70180 146740 73210 146763
rect 73370 146763 73393 147740
rect 76377 148740 76400 149747
rect 76560 149747 79590 149770
rect 76560 148740 76583 149747
rect 76377 147740 76583 148740
rect 76377 146763 76400 147740
rect 73370 146740 76400 146763
rect 76560 146763 76583 147740
rect 79567 148740 79590 149747
rect 79750 149747 82780 149770
rect 79750 148740 79773 149747
rect 79567 147740 79773 148740
rect 79567 146763 79590 147740
rect 76560 146740 79590 146763
rect 79750 146763 79773 147740
rect 82757 148740 82780 149747
rect 82940 149747 85970 149770
rect 82940 148740 82963 149747
rect 82757 147740 82963 148740
rect 82757 146763 82780 147740
rect 79750 146740 82780 146763
rect 82940 146763 82963 147740
rect 85947 148740 85970 149747
rect 86130 149747 89160 149770
rect 86130 148740 86153 149747
rect 85947 147740 86153 148740
rect 85947 146763 85970 147740
rect 82940 146740 85970 146763
rect 86130 146763 86153 147740
rect 89137 148740 89160 149747
rect 89320 149747 92350 149770
rect 89320 148740 89343 149747
rect 89137 147740 89343 148740
rect 89137 146763 89160 147740
rect 86130 146740 89160 146763
rect 89320 146763 89343 147740
rect 92327 148740 92350 149747
rect 92510 149747 95540 149770
rect 92510 148740 92533 149747
rect 92327 147740 92533 148740
rect 92327 146763 92350 147740
rect 89320 146740 92350 146763
rect 92510 146763 92533 147740
rect 95517 148740 95540 149747
rect 95700 149747 98730 149770
rect 95700 148740 95723 149747
rect 95517 147740 95723 148740
rect 95517 146763 95540 147740
rect 92510 146740 95540 146763
rect 95700 146763 95723 147740
rect 98707 148740 98730 149747
rect 98890 149747 101920 149770
rect 98890 148740 98913 149747
rect 98707 147740 98913 148740
rect 98707 146763 98730 147740
rect 95700 146740 98730 146763
rect 98890 146763 98913 147740
rect 101897 148740 101920 149747
rect 102080 149747 105110 149770
rect 102080 148740 102103 149747
rect 101897 147740 102103 148740
rect 101897 146763 101920 147740
rect 98890 146740 101920 146763
rect 102080 146763 102103 147740
rect 105087 148740 105110 149747
rect 105270 149747 108300 149770
rect 105270 148740 105293 149747
rect 105087 147740 105293 148740
rect 105087 146763 105110 147740
rect 102080 146740 105110 146763
rect 105270 146763 105293 147740
rect 108277 148740 108300 149747
rect 108460 149747 111490 149770
rect 108460 148740 108483 149747
rect 108277 147740 108483 148740
rect 108277 146763 108300 147740
rect 105270 146740 108300 146763
rect 108460 146763 108483 147740
rect 111467 148740 111490 149747
rect 111650 149747 114680 149770
rect 111650 148740 111673 149747
rect 111467 147740 111673 148740
rect 111467 146763 111490 147740
rect 108460 146740 111490 146763
rect 111650 146763 111673 147740
rect 114657 148740 114680 149747
rect 114840 149747 117870 149770
rect 114840 148740 114863 149747
rect 114657 147740 114863 148740
rect 114657 146763 114680 147740
rect 111650 146740 114680 146763
rect 114840 146763 114863 147740
rect 117847 148740 117870 149747
rect 118030 149747 121060 149770
rect 118030 148740 118053 149747
rect 117847 147740 118053 148740
rect 117847 146763 117870 147740
rect 114840 146740 117870 146763
rect 118030 146763 118053 147740
rect 121037 148740 121060 149747
rect 121220 149747 124250 149770
rect 121220 148740 121243 149747
rect 121037 147740 121243 148740
rect 121037 146763 121060 147740
rect 118030 146740 121060 146763
rect 121220 146763 121243 147740
rect 124227 148740 124250 149747
rect 124410 149747 127440 149770
rect 124410 148740 124433 149747
rect 124227 147740 124433 148740
rect 124227 146763 124250 147740
rect 121220 146740 124250 146763
rect 124410 146763 124433 147740
rect 127417 148740 127440 149747
rect 127600 149747 130630 149770
rect 127600 148740 127623 149747
rect 127417 147740 127623 148740
rect 127417 146763 127440 147740
rect 124410 146740 127440 146763
rect 127600 146763 127623 147740
rect 130607 148740 130630 149747
rect 130790 149747 133820 149770
rect 130790 148740 130813 149747
rect 130607 147740 130813 148740
rect 130607 146763 130630 147740
rect 127600 146740 130630 146763
rect 130790 146763 130813 147740
rect 133797 148740 133820 149747
rect 133980 149747 137010 149770
rect 133980 148740 134003 149747
rect 133797 147740 134003 148740
rect 133797 146763 133820 147740
rect 130790 146740 133820 146763
rect 133980 146763 134003 147740
rect 136987 148740 137010 149747
rect 136987 147740 137170 148740
rect 136987 146763 137010 147740
rect 133980 146740 137010 146763
rect 1000 146580 2000 146740
rect 4190 146580 5190 146740
rect 7380 146580 8380 146740
rect 10570 146580 11570 146740
rect 13760 146580 14760 146740
rect 16950 146580 17950 146740
rect 20140 146580 21140 146740
rect 23330 146580 24330 146740
rect 26520 146580 27520 146740
rect 29710 146580 30710 146740
rect 32900 146580 33900 146740
rect 36090 146580 37090 146740
rect 39280 146580 40280 146740
rect 42470 146580 43470 146740
rect 45660 146580 46660 146740
rect 48850 146580 49850 146740
rect 52040 146580 53040 146740
rect 55230 146580 56230 146740
rect 58420 146580 59420 146740
rect 61610 146580 62610 146740
rect 64800 146580 65800 146740
rect 67990 146580 68990 146740
rect 71180 146580 72180 146740
rect 74370 146580 75370 146740
rect 77560 146580 78560 146740
rect 80750 146580 81750 146740
rect 83940 146580 84940 146740
rect 87130 146580 88130 146740
rect 90320 146580 91320 146740
rect 93510 146580 94510 146740
rect 96700 146580 97700 146740
rect 99890 146580 100890 146740
rect 103080 146580 104080 146740
rect 106270 146580 107270 146740
rect 109460 146580 110460 146740
rect 112650 146580 113650 146740
rect 115840 146580 116840 146740
rect 119030 146580 120030 146740
rect 122220 146580 123220 146740
rect 125410 146580 126410 146740
rect 128600 146580 129600 146740
rect 131790 146580 132790 146740
rect 134980 146580 135980 146740
rect 0 146557 3030 146580
rect 0 143573 23 146557
rect 3007 145550 3030 146557
rect 3190 146557 6220 146580
rect 3190 145550 3213 146557
rect 3007 144550 3213 145550
rect 3007 143573 3030 144550
rect 0 143550 3030 143573
rect 3190 143573 3213 144550
rect 6197 145550 6220 146557
rect 6380 146557 9410 146580
rect 6380 145550 6403 146557
rect 6197 144550 6403 145550
rect 6197 143573 6220 144550
rect 3190 143550 6220 143573
rect 6380 143573 6403 144550
rect 9387 145550 9410 146557
rect 9570 146557 12600 146580
rect 9570 145550 9593 146557
rect 9387 144550 9593 145550
rect 9387 143573 9410 144550
rect 6380 143550 9410 143573
rect 9570 143573 9593 144550
rect 12577 145550 12600 146557
rect 12760 146557 15790 146580
rect 12760 145550 12783 146557
rect 12577 144550 12783 145550
rect 12577 143573 12600 144550
rect 9570 143550 12600 143573
rect 12760 143573 12783 144550
rect 15767 145550 15790 146557
rect 15950 146557 18980 146580
rect 15950 145550 15973 146557
rect 15767 144550 15973 145550
rect 15767 143573 15790 144550
rect 12760 143550 15790 143573
rect 15950 143573 15973 144550
rect 18957 145550 18980 146557
rect 19140 146557 22170 146580
rect 19140 145550 19163 146557
rect 18957 144550 19163 145550
rect 18957 143573 18980 144550
rect 15950 143550 18980 143573
rect 19140 143573 19163 144550
rect 22147 145550 22170 146557
rect 22330 146557 25360 146580
rect 22330 145550 22353 146557
rect 22147 144550 22353 145550
rect 22147 143573 22170 144550
rect 19140 143550 22170 143573
rect 22330 143573 22353 144550
rect 25337 145550 25360 146557
rect 25520 146557 28550 146580
rect 25520 145550 25543 146557
rect 25337 144550 25543 145550
rect 25337 143573 25360 144550
rect 22330 143550 25360 143573
rect 25520 143573 25543 144550
rect 28527 145550 28550 146557
rect 28710 146557 31740 146580
rect 28710 145550 28733 146557
rect 28527 144550 28733 145550
rect 28527 143573 28550 144550
rect 25520 143550 28550 143573
rect 28710 143573 28733 144550
rect 31717 145550 31740 146557
rect 31900 146557 34930 146580
rect 31900 145550 31923 146557
rect 31717 144550 31923 145550
rect 31717 143573 31740 144550
rect 28710 143550 31740 143573
rect 31900 143573 31923 144550
rect 34907 145550 34930 146557
rect 35090 146557 38120 146580
rect 35090 145550 35113 146557
rect 34907 144550 35113 145550
rect 34907 143573 34930 144550
rect 31900 143550 34930 143573
rect 35090 143573 35113 144550
rect 38097 145550 38120 146557
rect 38280 146557 41310 146580
rect 38280 145550 38303 146557
rect 38097 144550 38303 145550
rect 38097 143573 38120 144550
rect 35090 143550 38120 143573
rect 38280 143573 38303 144550
rect 41287 145550 41310 146557
rect 41470 146557 44500 146580
rect 41470 145550 41493 146557
rect 41287 144550 41493 145550
rect 41287 143573 41310 144550
rect 38280 143550 41310 143573
rect 41470 143573 41493 144550
rect 44477 145550 44500 146557
rect 44660 146557 47690 146580
rect 44660 145550 44683 146557
rect 44477 144550 44683 145550
rect 44477 143573 44500 144550
rect 41470 143550 44500 143573
rect 44660 143573 44683 144550
rect 47667 145550 47690 146557
rect 47850 146557 50880 146580
rect 47850 145550 47873 146557
rect 47667 144550 47873 145550
rect 47667 143573 47690 144550
rect 44660 143550 47690 143573
rect 47850 143573 47873 144550
rect 50857 145550 50880 146557
rect 51040 146557 54070 146580
rect 51040 145550 51063 146557
rect 50857 144550 51063 145550
rect 50857 143573 50880 144550
rect 47850 143550 50880 143573
rect 51040 143573 51063 144550
rect 54047 145550 54070 146557
rect 54230 146557 57260 146580
rect 54230 145550 54253 146557
rect 54047 144550 54253 145550
rect 54047 143573 54070 144550
rect 51040 143550 54070 143573
rect 54230 143573 54253 144550
rect 57237 145550 57260 146557
rect 57420 146557 60450 146580
rect 57420 145550 57443 146557
rect 57237 144550 57443 145550
rect 57237 143573 57260 144550
rect 54230 143550 57260 143573
rect 57420 143573 57443 144550
rect 60427 145550 60450 146557
rect 60610 146557 63640 146580
rect 60610 145550 60633 146557
rect 60427 144550 60633 145550
rect 60427 143573 60450 144550
rect 57420 143550 60450 143573
rect 60610 143573 60633 144550
rect 63617 145550 63640 146557
rect 63800 146557 66830 146580
rect 63800 145550 63823 146557
rect 63617 144550 63823 145550
rect 63617 143573 63640 144550
rect 60610 143550 63640 143573
rect 63800 143573 63823 144550
rect 66807 145550 66830 146557
rect 66990 146557 70020 146580
rect 66990 145550 67013 146557
rect 66807 144550 67013 145550
rect 66807 143573 66830 144550
rect 63800 143550 66830 143573
rect 66990 143573 67013 144550
rect 69997 145550 70020 146557
rect 70180 146557 73210 146580
rect 70180 145550 70203 146557
rect 69997 144550 70203 145550
rect 69997 143573 70020 144550
rect 66990 143550 70020 143573
rect 70180 143573 70203 144550
rect 73187 145550 73210 146557
rect 73370 146557 76400 146580
rect 73370 145550 73393 146557
rect 73187 144550 73393 145550
rect 73187 143573 73210 144550
rect 70180 143550 73210 143573
rect 73370 143573 73393 144550
rect 76377 145550 76400 146557
rect 76560 146557 79590 146580
rect 76560 145550 76583 146557
rect 76377 144550 76583 145550
rect 76377 143573 76400 144550
rect 73370 143550 76400 143573
rect 76560 143573 76583 144550
rect 79567 145550 79590 146557
rect 79750 146557 82780 146580
rect 79750 145550 79773 146557
rect 79567 144550 79773 145550
rect 79567 143573 79590 144550
rect 76560 143550 79590 143573
rect 79750 143573 79773 144550
rect 82757 145550 82780 146557
rect 82940 146557 85970 146580
rect 82940 145550 82963 146557
rect 82757 144550 82963 145550
rect 82757 143573 82780 144550
rect 79750 143550 82780 143573
rect 82940 143573 82963 144550
rect 85947 145550 85970 146557
rect 86130 146557 89160 146580
rect 86130 145550 86153 146557
rect 85947 144550 86153 145550
rect 85947 143573 85970 144550
rect 82940 143550 85970 143573
rect 86130 143573 86153 144550
rect 89137 145550 89160 146557
rect 89320 146557 92350 146580
rect 89320 145550 89343 146557
rect 89137 144550 89343 145550
rect 89137 143573 89160 144550
rect 86130 143550 89160 143573
rect 89320 143573 89343 144550
rect 92327 145550 92350 146557
rect 92510 146557 95540 146580
rect 92510 145550 92533 146557
rect 92327 144550 92533 145550
rect 92327 143573 92350 144550
rect 89320 143550 92350 143573
rect 92510 143573 92533 144550
rect 95517 145550 95540 146557
rect 95700 146557 98730 146580
rect 95700 145550 95723 146557
rect 95517 144550 95723 145550
rect 95517 143573 95540 144550
rect 92510 143550 95540 143573
rect 95700 143573 95723 144550
rect 98707 145550 98730 146557
rect 98890 146557 101920 146580
rect 98890 145550 98913 146557
rect 98707 144550 98913 145550
rect 98707 143573 98730 144550
rect 95700 143550 98730 143573
rect 98890 143573 98913 144550
rect 101897 145550 101920 146557
rect 102080 146557 105110 146580
rect 102080 145550 102103 146557
rect 101897 144550 102103 145550
rect 101897 143573 101920 144550
rect 98890 143550 101920 143573
rect 102080 143573 102103 144550
rect 105087 145550 105110 146557
rect 105270 146557 108300 146580
rect 105270 145550 105293 146557
rect 105087 144550 105293 145550
rect 105087 143573 105110 144550
rect 102080 143550 105110 143573
rect 105270 143573 105293 144550
rect 108277 145550 108300 146557
rect 108460 146557 111490 146580
rect 108460 145550 108483 146557
rect 108277 144550 108483 145550
rect 108277 143573 108300 144550
rect 105270 143550 108300 143573
rect 108460 143573 108483 144550
rect 111467 145550 111490 146557
rect 111650 146557 114680 146580
rect 111650 145550 111673 146557
rect 111467 144550 111673 145550
rect 111467 143573 111490 144550
rect 108460 143550 111490 143573
rect 111650 143573 111673 144550
rect 114657 145550 114680 146557
rect 114840 146557 117870 146580
rect 114840 145550 114863 146557
rect 114657 144550 114863 145550
rect 114657 143573 114680 144550
rect 111650 143550 114680 143573
rect 114840 143573 114863 144550
rect 117847 145550 117870 146557
rect 118030 146557 121060 146580
rect 118030 145550 118053 146557
rect 117847 144550 118053 145550
rect 117847 143573 117870 144550
rect 114840 143550 117870 143573
rect 118030 143573 118053 144550
rect 121037 145550 121060 146557
rect 121220 146557 124250 146580
rect 121220 145550 121243 146557
rect 121037 144550 121243 145550
rect 121037 143573 121060 144550
rect 118030 143550 121060 143573
rect 121220 143573 121243 144550
rect 124227 145550 124250 146557
rect 124410 146557 127440 146580
rect 124410 145550 124433 146557
rect 124227 144550 124433 145550
rect 124227 143573 124250 144550
rect 121220 143550 124250 143573
rect 124410 143573 124433 144550
rect 127417 145550 127440 146557
rect 127600 146557 130630 146580
rect 127600 145550 127623 146557
rect 127417 144550 127623 145550
rect 127417 143573 127440 144550
rect 124410 143550 127440 143573
rect 127600 143573 127623 144550
rect 130607 145550 130630 146557
rect 130790 146557 133820 146580
rect 130790 145550 130813 146557
rect 130607 144550 130813 145550
rect 130607 143573 130630 144550
rect 127600 143550 130630 143573
rect 130790 143573 130813 144550
rect 133797 145550 133820 146557
rect 133980 146557 137010 146580
rect 133980 145550 134003 146557
rect 133797 144550 134003 145550
rect 133797 143573 133820 144550
rect 130790 143550 133820 143573
rect 133980 143573 134003 144550
rect 136987 145550 137010 146557
rect 136987 144550 137170 145550
rect 136987 143573 137010 144550
rect 133980 143550 137010 143573
rect 1000 143390 2000 143550
rect 4190 143390 5190 143550
rect 7380 143390 8380 143550
rect 10570 143390 11570 143550
rect 13760 143390 14760 143550
rect 16950 143390 17950 143550
rect 20140 143390 21140 143550
rect 23330 143390 24330 143550
rect 26520 143390 27520 143550
rect 29710 143390 30710 143550
rect 32900 143390 33900 143550
rect 36090 143390 37090 143550
rect 39280 143390 40280 143550
rect 42470 143390 43470 143550
rect 45660 143390 46660 143550
rect 48850 143390 49850 143550
rect 52040 143390 53040 143550
rect 55230 143390 56230 143550
rect 58420 143390 59420 143550
rect 61610 143390 62610 143550
rect 64800 143390 65800 143550
rect 67990 143390 68990 143550
rect 71180 143390 72180 143550
rect 74370 143390 75370 143550
rect 77560 143390 78560 143550
rect 80750 143390 81750 143550
rect 83940 143390 84940 143550
rect 87130 143390 88130 143550
rect 90320 143390 91320 143550
rect 93510 143390 94510 143550
rect 96700 143390 97700 143550
rect 99890 143390 100890 143550
rect 103080 143390 104080 143550
rect 106270 143390 107270 143550
rect 109460 143390 110460 143550
rect 112650 143390 113650 143550
rect 115840 143390 116840 143550
rect 119030 143390 120030 143550
rect 122220 143390 123220 143550
rect 125410 143390 126410 143550
rect 128600 143390 129600 143550
rect 131790 143390 132790 143550
rect 134980 143390 135980 143550
rect 0 143367 3030 143390
rect 0 140383 23 143367
rect 3007 142360 3030 143367
rect 3190 143367 6220 143390
rect 3190 142360 3213 143367
rect 3007 141360 3213 142360
rect 3007 140383 3030 141360
rect 0 140360 3030 140383
rect 3190 140383 3213 141360
rect 6197 142360 6220 143367
rect 6380 143367 9410 143390
rect 6380 142360 6403 143367
rect 6197 141360 6403 142360
rect 6197 140383 6220 141360
rect 3190 140360 6220 140383
rect 6380 140383 6403 141360
rect 9387 142360 9410 143367
rect 9570 143367 12600 143390
rect 9570 142360 9593 143367
rect 9387 141360 9593 142360
rect 9387 140383 9410 141360
rect 6380 140360 9410 140383
rect 9570 140383 9593 141360
rect 12577 142360 12600 143367
rect 12760 143367 15790 143390
rect 12760 142360 12783 143367
rect 12577 141360 12783 142360
rect 12577 140383 12600 141360
rect 9570 140360 12600 140383
rect 12760 140383 12783 141360
rect 15767 142360 15790 143367
rect 15950 143367 18980 143390
rect 15950 142360 15973 143367
rect 15767 141360 15973 142360
rect 15767 140383 15790 141360
rect 12760 140360 15790 140383
rect 15950 140383 15973 141360
rect 18957 142360 18980 143367
rect 19140 143367 22170 143390
rect 19140 142360 19163 143367
rect 18957 141360 19163 142360
rect 18957 140383 18980 141360
rect 15950 140360 18980 140383
rect 19140 140383 19163 141360
rect 22147 142360 22170 143367
rect 22330 143367 25360 143390
rect 22330 142360 22353 143367
rect 22147 141360 22353 142360
rect 22147 140383 22170 141360
rect 19140 140360 22170 140383
rect 22330 140383 22353 141360
rect 25337 142360 25360 143367
rect 25520 143367 28550 143390
rect 25520 142360 25543 143367
rect 25337 141360 25543 142360
rect 25337 140383 25360 141360
rect 22330 140360 25360 140383
rect 25520 140383 25543 141360
rect 28527 142360 28550 143367
rect 28710 143367 31740 143390
rect 28710 142360 28733 143367
rect 28527 141360 28733 142360
rect 28527 140383 28550 141360
rect 25520 140360 28550 140383
rect 28710 140383 28733 141360
rect 31717 142360 31740 143367
rect 31900 143367 34930 143390
rect 31900 142360 31923 143367
rect 31717 141360 31923 142360
rect 31717 140383 31740 141360
rect 28710 140360 31740 140383
rect 31900 140383 31923 141360
rect 34907 142360 34930 143367
rect 35090 143367 38120 143390
rect 35090 142360 35113 143367
rect 34907 141360 35113 142360
rect 34907 140383 34930 141360
rect 31900 140360 34930 140383
rect 35090 140383 35113 141360
rect 38097 142360 38120 143367
rect 38280 143367 41310 143390
rect 38280 142360 38303 143367
rect 38097 141360 38303 142360
rect 38097 140383 38120 141360
rect 35090 140360 38120 140383
rect 38280 140383 38303 141360
rect 41287 142360 41310 143367
rect 41470 143367 44500 143390
rect 41470 142360 41493 143367
rect 41287 141360 41493 142360
rect 41287 140383 41310 141360
rect 38280 140360 41310 140383
rect 41470 140383 41493 141360
rect 44477 142360 44500 143367
rect 44660 143367 47690 143390
rect 44660 142360 44683 143367
rect 44477 141360 44683 142360
rect 44477 140383 44500 141360
rect 41470 140360 44500 140383
rect 44660 140383 44683 141360
rect 47667 142360 47690 143367
rect 47850 143367 50880 143390
rect 47850 142360 47873 143367
rect 47667 141360 47873 142360
rect 47667 140383 47690 141360
rect 44660 140360 47690 140383
rect 47850 140383 47873 141360
rect 50857 142360 50880 143367
rect 51040 143367 54070 143390
rect 51040 142360 51063 143367
rect 50857 141360 51063 142360
rect 50857 140383 50880 141360
rect 47850 140360 50880 140383
rect 51040 140383 51063 141360
rect 54047 142360 54070 143367
rect 54230 143367 57260 143390
rect 54230 142360 54253 143367
rect 54047 141360 54253 142360
rect 54047 140383 54070 141360
rect 51040 140360 54070 140383
rect 54230 140383 54253 141360
rect 57237 142360 57260 143367
rect 57420 143367 60450 143390
rect 57420 142360 57443 143367
rect 57237 141360 57443 142360
rect 57237 140383 57260 141360
rect 54230 140360 57260 140383
rect 57420 140383 57443 141360
rect 60427 142360 60450 143367
rect 60610 143367 63640 143390
rect 60610 142360 60633 143367
rect 60427 141360 60633 142360
rect 60427 140383 60450 141360
rect 57420 140360 60450 140383
rect 60610 140383 60633 141360
rect 63617 142360 63640 143367
rect 63800 143367 66830 143390
rect 63800 142360 63823 143367
rect 63617 141360 63823 142360
rect 63617 140383 63640 141360
rect 60610 140360 63640 140383
rect 63800 140383 63823 141360
rect 66807 142360 66830 143367
rect 66990 143367 70020 143390
rect 66990 142360 67013 143367
rect 66807 141360 67013 142360
rect 66807 140383 66830 141360
rect 63800 140360 66830 140383
rect 66990 140383 67013 141360
rect 69997 142360 70020 143367
rect 70180 143367 73210 143390
rect 70180 142360 70203 143367
rect 69997 141360 70203 142360
rect 69997 140383 70020 141360
rect 66990 140360 70020 140383
rect 70180 140383 70203 141360
rect 73187 142360 73210 143367
rect 73370 143367 76400 143390
rect 73370 142360 73393 143367
rect 73187 141360 73393 142360
rect 73187 140383 73210 141360
rect 70180 140360 73210 140383
rect 73370 140383 73393 141360
rect 76377 142360 76400 143367
rect 76560 143367 79590 143390
rect 76560 142360 76583 143367
rect 76377 141360 76583 142360
rect 76377 140383 76400 141360
rect 73370 140360 76400 140383
rect 76560 140383 76583 141360
rect 79567 142360 79590 143367
rect 79750 143367 82780 143390
rect 79750 142360 79773 143367
rect 79567 141360 79773 142360
rect 79567 140383 79590 141360
rect 76560 140360 79590 140383
rect 79750 140383 79773 141360
rect 82757 142360 82780 143367
rect 82940 143367 85970 143390
rect 82940 142360 82963 143367
rect 82757 141360 82963 142360
rect 82757 140383 82780 141360
rect 79750 140360 82780 140383
rect 82940 140383 82963 141360
rect 85947 142360 85970 143367
rect 86130 143367 89160 143390
rect 86130 142360 86153 143367
rect 85947 141360 86153 142360
rect 85947 140383 85970 141360
rect 82940 140360 85970 140383
rect 86130 140383 86153 141360
rect 89137 142360 89160 143367
rect 89320 143367 92350 143390
rect 89320 142360 89343 143367
rect 89137 141360 89343 142360
rect 89137 140383 89160 141360
rect 86130 140360 89160 140383
rect 89320 140383 89343 141360
rect 92327 142360 92350 143367
rect 92510 143367 95540 143390
rect 92510 142360 92533 143367
rect 92327 141360 92533 142360
rect 92327 140383 92350 141360
rect 89320 140360 92350 140383
rect 92510 140383 92533 141360
rect 95517 142360 95540 143367
rect 95700 143367 98730 143390
rect 95700 142360 95723 143367
rect 95517 141360 95723 142360
rect 95517 140383 95540 141360
rect 92510 140360 95540 140383
rect 95700 140383 95723 141360
rect 98707 142360 98730 143367
rect 98890 143367 101920 143390
rect 98890 142360 98913 143367
rect 98707 141360 98913 142360
rect 98707 140383 98730 141360
rect 95700 140360 98730 140383
rect 98890 140383 98913 141360
rect 101897 142360 101920 143367
rect 102080 143367 105110 143390
rect 102080 142360 102103 143367
rect 101897 141360 102103 142360
rect 101897 140383 101920 141360
rect 98890 140360 101920 140383
rect 102080 140383 102103 141360
rect 105087 142360 105110 143367
rect 105270 143367 108300 143390
rect 105270 142360 105293 143367
rect 105087 141360 105293 142360
rect 105087 140383 105110 141360
rect 102080 140360 105110 140383
rect 105270 140383 105293 141360
rect 108277 142360 108300 143367
rect 108460 143367 111490 143390
rect 108460 142360 108483 143367
rect 108277 141360 108483 142360
rect 108277 140383 108300 141360
rect 105270 140360 108300 140383
rect 108460 140383 108483 141360
rect 111467 142360 111490 143367
rect 111650 143367 114680 143390
rect 111650 142360 111673 143367
rect 111467 141360 111673 142360
rect 111467 140383 111490 141360
rect 108460 140360 111490 140383
rect 111650 140383 111673 141360
rect 114657 142360 114680 143367
rect 114840 143367 117870 143390
rect 114840 142360 114863 143367
rect 114657 141360 114863 142360
rect 114657 140383 114680 141360
rect 111650 140360 114680 140383
rect 114840 140383 114863 141360
rect 117847 142360 117870 143367
rect 118030 143367 121060 143390
rect 118030 142360 118053 143367
rect 117847 141360 118053 142360
rect 117847 140383 117870 141360
rect 114840 140360 117870 140383
rect 118030 140383 118053 141360
rect 121037 142360 121060 143367
rect 121220 143367 124250 143390
rect 121220 142360 121243 143367
rect 121037 141360 121243 142360
rect 121037 140383 121060 141360
rect 118030 140360 121060 140383
rect 121220 140383 121243 141360
rect 124227 142360 124250 143367
rect 124410 143367 127440 143390
rect 124410 142360 124433 143367
rect 124227 141360 124433 142360
rect 124227 140383 124250 141360
rect 121220 140360 124250 140383
rect 124410 140383 124433 141360
rect 127417 142360 127440 143367
rect 127600 143367 130630 143390
rect 127600 142360 127623 143367
rect 127417 141360 127623 142360
rect 127417 140383 127440 141360
rect 124410 140360 127440 140383
rect 127600 140383 127623 141360
rect 130607 142360 130630 143367
rect 130790 143367 133820 143390
rect 130790 142360 130813 143367
rect 130607 141360 130813 142360
rect 130607 140383 130630 141360
rect 127600 140360 130630 140383
rect 130790 140383 130813 141360
rect 133797 142360 133820 143367
rect 133980 143367 137010 143390
rect 133980 142360 134003 143367
rect 133797 141360 134003 142360
rect 133797 140383 133820 141360
rect 130790 140360 133820 140383
rect 133980 140383 134003 141360
rect 136987 142360 137010 143367
rect 136987 141360 137170 142360
rect 136987 140383 137010 141360
rect 133980 140360 137010 140383
rect 1000 140200 2000 140360
rect 4190 140200 5190 140360
rect 7380 140200 8380 140360
rect 10570 140200 11570 140360
rect 13760 140200 14760 140360
rect 16950 140200 17950 140360
rect 20140 140200 21140 140360
rect 23330 140200 24330 140360
rect 26520 140200 27520 140360
rect 29710 140200 30710 140360
rect 32900 140200 33900 140360
rect 36090 140200 37090 140360
rect 39280 140200 40280 140360
rect 42470 140200 43470 140360
rect 45660 140200 46660 140360
rect 48850 140200 49850 140360
rect 52040 140200 53040 140360
rect 55230 140200 56230 140360
rect 58420 140200 59420 140360
rect 61610 140200 62610 140360
rect 64800 140200 65800 140360
rect 67990 140200 68990 140360
rect 71180 140200 72180 140360
rect 74370 140200 75370 140360
rect 77560 140200 78560 140360
rect 80750 140200 81750 140360
rect 83940 140200 84940 140360
rect 87130 140200 88130 140360
rect 90320 140200 91320 140360
rect 93510 140200 94510 140360
rect 96700 140200 97700 140360
rect 99890 140200 100890 140360
rect 103080 140200 104080 140360
rect 106270 140200 107270 140360
rect 109460 140200 110460 140360
rect 112650 140200 113650 140360
rect 115840 140200 116840 140360
rect 119030 140200 120030 140360
rect 122220 140200 123220 140360
rect 125410 140200 126410 140360
rect 128600 140200 129600 140360
rect 131790 140200 132790 140360
rect 134980 140200 135980 140360
rect 0 140160 3030 140200
rect 3190 140160 6220 140200
rect 6380 140160 9410 140200
rect 0 140110 9410 140160
rect 0 121310 50 140110
rect 9320 139170 9410 140110
rect 9570 140177 12600 140200
rect 9570 139170 9593 140177
rect 9320 138170 9593 139170
rect 9320 137170 9410 138170
rect 9570 137193 9593 138170
rect 12577 139170 12600 140177
rect 12760 140177 15790 140200
rect 12760 139170 12783 140177
rect 12577 138170 12783 139170
rect 12577 137193 12600 138170
rect 9570 137170 12600 137193
rect 12760 137193 12783 138170
rect 15767 139170 15790 140177
rect 15950 140177 18980 140200
rect 15950 139170 15973 140177
rect 15767 138170 15973 139170
rect 15767 137193 15790 138170
rect 12760 137170 15790 137193
rect 15950 137193 15973 138170
rect 18957 139170 18980 140177
rect 19140 140177 22170 140200
rect 19140 139170 19163 140177
rect 18957 138170 19163 139170
rect 18957 137193 18980 138170
rect 15950 137170 18980 137193
rect 19140 137193 19163 138170
rect 22147 139170 22170 140177
rect 22330 140177 25360 140200
rect 22330 139170 22353 140177
rect 22147 138170 22353 139170
rect 22147 137193 22170 138170
rect 19140 137170 22170 137193
rect 22330 137193 22353 138170
rect 25337 139170 25360 140177
rect 25520 140177 28550 140200
rect 25520 139170 25543 140177
rect 25337 138170 25543 139170
rect 25337 137193 25360 138170
rect 22330 137170 25360 137193
rect 25520 137193 25543 138170
rect 28527 139170 28550 140177
rect 28710 140177 31740 140200
rect 28710 139170 28733 140177
rect 28527 138170 28733 139170
rect 28527 137193 28550 138170
rect 25520 137170 28550 137193
rect 28710 137193 28733 138170
rect 31717 139170 31740 140177
rect 31900 140177 34930 140200
rect 31900 139170 31923 140177
rect 31717 138170 31923 139170
rect 31717 137193 31740 138170
rect 28710 137170 31740 137193
rect 31900 137193 31923 138170
rect 34907 139170 34930 140177
rect 35090 140177 38120 140200
rect 35090 139170 35113 140177
rect 34907 138170 35113 139170
rect 34907 137193 34930 138170
rect 31900 137170 34930 137193
rect 35090 137193 35113 138170
rect 38097 139170 38120 140177
rect 38280 140177 41310 140200
rect 38280 139170 38303 140177
rect 38097 138170 38303 139170
rect 38097 137193 38120 138170
rect 35090 137170 38120 137193
rect 38280 137193 38303 138170
rect 41287 139170 41310 140177
rect 41470 140177 44500 140200
rect 41470 139170 41493 140177
rect 41287 138170 41493 139170
rect 41287 137193 41310 138170
rect 38280 137170 41310 137193
rect 41470 137193 41493 138170
rect 44477 139170 44500 140177
rect 44660 140177 47690 140200
rect 44660 139170 44683 140177
rect 44477 138170 44683 139170
rect 44477 137193 44500 138170
rect 41470 137170 44500 137193
rect 44660 137193 44683 138170
rect 47667 139170 47690 140177
rect 47850 140177 50880 140200
rect 47850 139170 47873 140177
rect 47667 138170 47873 139170
rect 47667 137193 47690 138170
rect 44660 137170 47690 137193
rect 47850 137193 47873 138170
rect 50857 139170 50880 140177
rect 51040 140177 54070 140200
rect 51040 139170 51063 140177
rect 50857 138170 51063 139170
rect 50857 137193 50880 138170
rect 47850 137170 50880 137193
rect 51040 137193 51063 138170
rect 54047 139170 54070 140177
rect 54230 140177 57260 140200
rect 54230 139170 54253 140177
rect 54047 138170 54253 139170
rect 54047 137193 54070 138170
rect 51040 137170 54070 137193
rect 54230 137193 54253 138170
rect 57237 139170 57260 140177
rect 57420 140177 60450 140200
rect 57420 139170 57443 140177
rect 57237 138170 57443 139170
rect 57237 137193 57260 138170
rect 54230 137170 57260 137193
rect 57420 137193 57443 138170
rect 60427 139170 60450 140177
rect 60610 140177 63640 140200
rect 60610 139170 60633 140177
rect 60427 138170 60633 139170
rect 60427 137193 60450 138170
rect 57420 137170 60450 137193
rect 60610 137193 60633 138170
rect 63617 139170 63640 140177
rect 63800 140177 66830 140200
rect 63800 139170 63823 140177
rect 63617 138170 63823 139170
rect 63617 137193 63640 138170
rect 60610 137170 63640 137193
rect 63800 137193 63823 138170
rect 66807 139170 66830 140177
rect 66990 140177 70020 140200
rect 66990 139170 67013 140177
rect 66807 138170 67013 139170
rect 66807 137193 66830 138170
rect 63800 137170 66830 137193
rect 66990 137193 67013 138170
rect 69997 139170 70020 140177
rect 70180 140177 73210 140200
rect 70180 139170 70203 140177
rect 69997 138170 70203 139170
rect 69997 137193 70020 138170
rect 66990 137170 70020 137193
rect 70180 137193 70203 138170
rect 73187 139170 73210 140177
rect 73370 140177 76400 140200
rect 73370 139170 73393 140177
rect 73187 138170 73393 139170
rect 73187 137193 73210 138170
rect 70180 137170 73210 137193
rect 73370 137193 73393 138170
rect 76377 139170 76400 140177
rect 76560 140177 79590 140200
rect 76560 139170 76583 140177
rect 76377 138170 76583 139170
rect 76377 137193 76400 138170
rect 73370 137170 76400 137193
rect 76560 137193 76583 138170
rect 79567 139170 79590 140177
rect 79750 140177 82780 140200
rect 79750 139170 79773 140177
rect 79567 138170 79773 139170
rect 79567 137193 79590 138170
rect 76560 137170 79590 137193
rect 79750 137193 79773 138170
rect 82757 139170 82780 140177
rect 82940 140177 85970 140200
rect 82940 139170 82963 140177
rect 82757 138170 82963 139170
rect 82757 137193 82780 138170
rect 79750 137170 82780 137193
rect 82940 137193 82963 138170
rect 85947 139170 85970 140177
rect 86130 140177 89160 140200
rect 86130 139170 86153 140177
rect 85947 138170 86153 139170
rect 85947 137193 85970 138170
rect 82940 137170 85970 137193
rect 86130 137193 86153 138170
rect 89137 139170 89160 140177
rect 89320 140177 92350 140200
rect 89320 139170 89343 140177
rect 89137 138170 89343 139170
rect 89137 137193 89160 138170
rect 86130 137170 89160 137193
rect 89320 137193 89343 138170
rect 92327 139170 92350 140177
rect 92510 140177 95540 140200
rect 92510 139170 92533 140177
rect 92327 138170 92533 139170
rect 92327 137193 92350 138170
rect 89320 137170 92350 137193
rect 92510 137193 92533 138170
rect 95517 139170 95540 140177
rect 95700 140177 98730 140200
rect 95700 139170 95723 140177
rect 95517 138170 95723 139170
rect 95517 137193 95540 138170
rect 92510 137170 95540 137193
rect 95700 137193 95723 138170
rect 98707 139170 98730 140177
rect 98890 140177 101920 140200
rect 98890 139170 98913 140177
rect 98707 138170 98913 139170
rect 98707 137193 98730 138170
rect 95700 137170 98730 137193
rect 98890 137193 98913 138170
rect 101897 139170 101920 140177
rect 102080 140177 105110 140200
rect 102080 139170 102103 140177
rect 101897 138170 102103 139170
rect 101897 137193 101920 138170
rect 98890 137170 101920 137193
rect 102080 137193 102103 138170
rect 105087 139170 105110 140177
rect 105270 140177 108300 140200
rect 105270 139170 105293 140177
rect 105087 138170 105293 139170
rect 105087 137193 105110 138170
rect 102080 137170 105110 137193
rect 105270 137193 105293 138170
rect 108277 139170 108300 140177
rect 108460 140177 111490 140200
rect 108460 139170 108483 140177
rect 108277 138170 108483 139170
rect 108277 137193 108300 138170
rect 105270 137170 108300 137193
rect 108460 137193 108483 138170
rect 111467 139170 111490 140177
rect 111650 140177 114680 140200
rect 111650 139170 111673 140177
rect 111467 138170 111673 139170
rect 111467 137193 111490 138170
rect 108460 137170 111490 137193
rect 111650 137193 111673 138170
rect 114657 139170 114680 140177
rect 114840 140177 117870 140200
rect 114840 139170 114863 140177
rect 114657 138170 114863 139170
rect 114657 137193 114680 138170
rect 111650 137170 114680 137193
rect 114840 137193 114863 138170
rect 117847 139170 117870 140177
rect 118030 140177 121060 140200
rect 118030 139170 118053 140177
rect 117847 138170 118053 139170
rect 117847 137193 117870 138170
rect 114840 137170 117870 137193
rect 118030 137193 118053 138170
rect 121037 139170 121060 140177
rect 121220 140177 124250 140200
rect 121220 139170 121243 140177
rect 121037 138170 121243 139170
rect 121037 137193 121060 138170
rect 118030 137170 121060 137193
rect 121220 137193 121243 138170
rect 124227 139170 124250 140177
rect 124410 140177 127440 140200
rect 124410 139170 124433 140177
rect 124227 138170 124433 139170
rect 124227 137193 124250 138170
rect 121220 137170 124250 137193
rect 124410 137193 124433 138170
rect 127417 139170 127440 140177
rect 127600 140177 130630 140200
rect 127600 139170 127623 140177
rect 127417 138170 127623 139170
rect 127417 137193 127440 138170
rect 124410 137170 127440 137193
rect 127600 137193 127623 138170
rect 130607 139170 130630 140177
rect 130790 140177 133820 140200
rect 130790 139170 130813 140177
rect 130607 138170 130813 139170
rect 130607 137193 130630 138170
rect 127600 137170 130630 137193
rect 130790 137193 130813 138170
rect 133797 139170 133820 140177
rect 133980 140177 137010 140200
rect 133980 139170 134003 140177
rect 133797 138170 134003 139170
rect 133797 137193 133820 138170
rect 130790 137170 133820 137193
rect 133980 137193 134003 138170
rect 136987 139170 137010 140177
rect 136987 138170 137170 139170
rect 136987 137193 137010 138170
rect 133980 137170 137010 137193
rect 9320 137010 9370 137170
rect 10570 137010 11570 137170
rect 13760 137010 14760 137170
rect 16950 137010 17950 137170
rect 20140 137010 21140 137170
rect 23330 137010 24330 137170
rect 26520 137010 27520 137170
rect 29710 137010 30710 137170
rect 32900 137010 33900 137170
rect 36090 137010 37090 137170
rect 39280 137010 40280 137170
rect 42470 137010 43470 137170
rect 45660 137010 46660 137170
rect 48850 137010 49850 137170
rect 52040 137010 53040 137170
rect 55230 137010 56230 137170
rect 58420 137010 59420 137170
rect 61610 137010 62610 137170
rect 64800 137010 65800 137170
rect 67990 137010 68990 137170
rect 71180 137010 72180 137170
rect 74370 137010 75370 137170
rect 77560 137010 78560 137170
rect 80750 137010 81750 137170
rect 83940 137010 84940 137170
rect 87130 137010 88130 137170
rect 90320 137010 91320 137170
rect 93510 137010 94510 137170
rect 96700 137010 97700 137170
rect 99890 137010 100890 137170
rect 103080 137010 104080 137170
rect 106270 137010 107270 137170
rect 109460 137010 110460 137170
rect 112650 137010 113650 137170
rect 115840 137010 116840 137170
rect 119030 137010 120030 137170
rect 122220 137010 123220 137170
rect 125410 137010 126410 137170
rect 128600 137010 129600 137170
rect 131790 137010 132790 137170
rect 134980 137010 135980 137170
rect 9320 135980 9410 137010
rect 9570 136987 12600 137010
rect 9570 135980 9593 136987
rect 9320 134980 9593 135980
rect 9320 133980 9410 134980
rect 9570 134003 9593 134980
rect 12577 135980 12600 136987
rect 12760 136987 15790 137010
rect 12760 135980 12783 136987
rect 12577 134980 12783 135980
rect 12577 134003 12600 134980
rect 9570 133980 12600 134003
rect 12760 134003 12783 134980
rect 15767 135980 15790 136987
rect 15950 136987 18980 137010
rect 15950 135980 15973 136987
rect 15767 134980 15973 135980
rect 15767 134003 15790 134980
rect 12760 133980 15790 134003
rect 15950 134003 15973 134980
rect 18957 135980 18980 136987
rect 19140 136987 22170 137010
rect 19140 135980 19163 136987
rect 18957 134980 19163 135980
rect 18957 134003 18980 134980
rect 15950 133980 18980 134003
rect 19140 134003 19163 134980
rect 22147 135980 22170 136987
rect 22330 136987 25360 137010
rect 22330 135980 22353 136987
rect 22147 134980 22353 135980
rect 22147 134003 22170 134980
rect 19140 133980 22170 134003
rect 22330 134003 22353 134980
rect 25337 135980 25360 136987
rect 25520 136987 28550 137010
rect 25520 135980 25543 136987
rect 25337 134980 25543 135980
rect 25337 134003 25360 134980
rect 22330 133980 25360 134003
rect 25520 134003 25543 134980
rect 28527 135980 28550 136987
rect 28710 136987 31740 137010
rect 28710 135980 28733 136987
rect 28527 134980 28733 135980
rect 28527 134003 28550 134980
rect 25520 133980 28550 134003
rect 28710 134003 28733 134980
rect 31717 135980 31740 136987
rect 31900 136987 34930 137010
rect 31900 135980 31923 136987
rect 31717 134980 31923 135980
rect 31717 134003 31740 134980
rect 28710 133980 31740 134003
rect 31900 134003 31923 134980
rect 34907 135980 34930 136987
rect 35090 136987 38120 137010
rect 35090 135980 35113 136987
rect 34907 134980 35113 135980
rect 34907 134003 34930 134980
rect 31900 133980 34930 134003
rect 35090 134003 35113 134980
rect 38097 135980 38120 136987
rect 38280 136987 41310 137010
rect 38280 135980 38303 136987
rect 38097 134980 38303 135980
rect 38097 134003 38120 134980
rect 35090 133980 38120 134003
rect 38280 134003 38303 134980
rect 41287 135980 41310 136987
rect 41470 136987 44500 137010
rect 41470 135980 41493 136987
rect 41287 134980 41493 135980
rect 41287 134003 41310 134980
rect 38280 133980 41310 134003
rect 41470 134003 41493 134980
rect 44477 135980 44500 136987
rect 44660 136987 47690 137010
rect 44660 135980 44683 136987
rect 44477 134980 44683 135980
rect 44477 134003 44500 134980
rect 41470 133980 44500 134003
rect 44660 134003 44683 134980
rect 47667 135980 47690 136987
rect 47850 136987 50880 137010
rect 47850 135980 47873 136987
rect 47667 134980 47873 135980
rect 47667 134003 47690 134980
rect 44660 133980 47690 134003
rect 47850 134003 47873 134980
rect 50857 135980 50880 136987
rect 51040 136987 54070 137010
rect 51040 135980 51063 136987
rect 50857 134980 51063 135980
rect 50857 134003 50880 134980
rect 47850 133980 50880 134003
rect 51040 134003 51063 134980
rect 54047 135980 54070 136987
rect 54230 136987 57260 137010
rect 54230 135980 54253 136987
rect 54047 134980 54253 135980
rect 54047 134003 54070 134980
rect 51040 133980 54070 134003
rect 54230 134003 54253 134980
rect 57237 135980 57260 136987
rect 57420 136987 60450 137010
rect 57420 135980 57443 136987
rect 57237 134980 57443 135980
rect 57237 134003 57260 134980
rect 54230 133980 57260 134003
rect 57420 134003 57443 134980
rect 60427 135980 60450 136987
rect 60610 136987 63640 137010
rect 60610 135980 60633 136987
rect 60427 134980 60633 135980
rect 60427 134003 60450 134980
rect 57420 133980 60450 134003
rect 60610 134003 60633 134980
rect 63617 135980 63640 136987
rect 63800 136987 66830 137010
rect 63800 135980 63823 136987
rect 63617 134980 63823 135980
rect 63617 134003 63640 134980
rect 60610 133980 63640 134003
rect 63800 134003 63823 134980
rect 66807 135980 66830 136987
rect 66990 136987 70020 137010
rect 66990 135980 67013 136987
rect 66807 134980 67013 135980
rect 66807 134003 66830 134980
rect 63800 133980 66830 134003
rect 66990 134003 67013 134980
rect 69997 135980 70020 136987
rect 70180 136987 73210 137010
rect 70180 135980 70203 136987
rect 69997 134980 70203 135980
rect 69997 134003 70020 134980
rect 66990 133980 70020 134003
rect 70180 134003 70203 134980
rect 73187 135980 73210 136987
rect 73370 136987 76400 137010
rect 73370 135980 73393 136987
rect 73187 134980 73393 135980
rect 73187 134003 73210 134980
rect 70180 133980 73210 134003
rect 73370 134003 73393 134980
rect 76377 135980 76400 136987
rect 76560 136987 79590 137010
rect 76560 135980 76583 136987
rect 76377 134980 76583 135980
rect 76377 134003 76400 134980
rect 73370 133980 76400 134003
rect 76560 134003 76583 134980
rect 79567 135980 79590 136987
rect 79750 136987 82780 137010
rect 79750 135980 79773 136987
rect 79567 134980 79773 135980
rect 79567 134003 79590 134980
rect 76560 133980 79590 134003
rect 79750 134003 79773 134980
rect 82757 135980 82780 136987
rect 82940 136987 85970 137010
rect 82940 135980 82963 136987
rect 82757 134980 82963 135980
rect 82757 134003 82780 134980
rect 79750 133980 82780 134003
rect 82940 134003 82963 134980
rect 85947 135980 85970 136987
rect 86130 136987 89160 137010
rect 86130 135980 86153 136987
rect 85947 134980 86153 135980
rect 85947 134003 85970 134980
rect 82940 133980 85970 134003
rect 86130 134003 86153 134980
rect 89137 135980 89160 136987
rect 89320 136987 92350 137010
rect 89320 135980 89343 136987
rect 89137 134980 89343 135980
rect 89137 134003 89160 134980
rect 86130 133980 89160 134003
rect 89320 134003 89343 134980
rect 92327 135980 92350 136987
rect 92510 136987 95540 137010
rect 92510 135980 92533 136987
rect 92327 134980 92533 135980
rect 92327 134003 92350 134980
rect 89320 133980 92350 134003
rect 92510 134003 92533 134980
rect 95517 135980 95540 136987
rect 95700 136987 98730 137010
rect 95700 135980 95723 136987
rect 95517 134980 95723 135980
rect 95517 134003 95540 134980
rect 92510 133980 95540 134003
rect 95700 134003 95723 134980
rect 98707 135980 98730 136987
rect 98890 136987 101920 137010
rect 98890 135980 98913 136987
rect 98707 134980 98913 135980
rect 98707 134003 98730 134980
rect 95700 133980 98730 134003
rect 98890 134003 98913 134980
rect 101897 135980 101920 136987
rect 102080 136987 105110 137010
rect 102080 135980 102103 136987
rect 101897 134980 102103 135980
rect 101897 134003 101920 134980
rect 98890 133980 101920 134003
rect 102080 134003 102103 134980
rect 105087 135980 105110 136987
rect 105270 136987 108300 137010
rect 105270 135980 105293 136987
rect 105087 134980 105293 135980
rect 105087 134003 105110 134980
rect 102080 133980 105110 134003
rect 105270 134003 105293 134980
rect 108277 135980 108300 136987
rect 108460 136987 111490 137010
rect 108460 135980 108483 136987
rect 108277 134980 108483 135980
rect 108277 134003 108300 134980
rect 105270 133980 108300 134003
rect 108460 134003 108483 134980
rect 111467 135980 111490 136987
rect 111650 136987 114680 137010
rect 111650 135980 111673 136987
rect 111467 134980 111673 135980
rect 111467 134003 111490 134980
rect 108460 133980 111490 134003
rect 111650 134003 111673 134980
rect 114657 135980 114680 136987
rect 114840 136987 117870 137010
rect 114840 135980 114863 136987
rect 114657 134980 114863 135980
rect 114657 134003 114680 134980
rect 111650 133980 114680 134003
rect 114840 134003 114863 134980
rect 117847 135980 117870 136987
rect 118030 136987 121060 137010
rect 118030 135980 118053 136987
rect 117847 134980 118053 135980
rect 117847 134003 117870 134980
rect 114840 133980 117870 134003
rect 118030 134003 118053 134980
rect 121037 135980 121060 136987
rect 121220 136987 124250 137010
rect 121220 135980 121243 136987
rect 121037 134980 121243 135980
rect 121037 134003 121060 134980
rect 118030 133980 121060 134003
rect 121220 134003 121243 134980
rect 124227 135980 124250 136987
rect 124410 136987 127440 137010
rect 124410 135980 124433 136987
rect 124227 134980 124433 135980
rect 124227 134003 124250 134980
rect 121220 133980 124250 134003
rect 124410 134003 124433 134980
rect 127417 135980 127440 136987
rect 127600 136987 130630 137010
rect 127600 135980 127623 136987
rect 127417 134980 127623 135980
rect 127417 134003 127440 134980
rect 124410 133980 127440 134003
rect 127600 134003 127623 134980
rect 130607 135980 130630 136987
rect 130790 136987 133820 137010
rect 130790 135980 130813 136987
rect 130607 134980 130813 135980
rect 130607 134003 130630 134980
rect 127600 133980 130630 134003
rect 130790 134003 130813 134980
rect 133797 135980 133820 136987
rect 133980 136987 137010 137010
rect 133980 135980 134003 136987
rect 133797 134980 134003 135980
rect 133797 134003 133820 134980
rect 130790 133980 133820 134003
rect 133980 134003 134003 134980
rect 136987 135980 137010 136987
rect 136987 134980 137170 135980
rect 136987 134003 137010 134980
rect 133980 133980 137010 134003
rect 9320 133820 9370 133980
rect 10570 133820 11570 133980
rect 13760 133820 14760 133980
rect 16950 133820 17950 133980
rect 20140 133820 21140 133980
rect 23330 133820 24330 133980
rect 26520 133820 27520 133980
rect 29710 133820 30710 133980
rect 32900 133820 33900 133980
rect 36090 133820 37090 133980
rect 39280 133820 40280 133980
rect 42470 133820 43470 133980
rect 45660 133820 46660 133980
rect 48850 133820 49850 133980
rect 52040 133820 53040 133980
rect 55230 133820 56230 133980
rect 58420 133820 59420 133980
rect 61610 133820 62610 133980
rect 64800 133820 65800 133980
rect 67990 133820 68990 133980
rect 71180 133820 72180 133980
rect 74370 133820 75370 133980
rect 77560 133820 78560 133980
rect 80750 133820 81750 133980
rect 83940 133820 84940 133980
rect 87130 133820 88130 133980
rect 90320 133820 91320 133980
rect 93510 133820 94510 133980
rect 96700 133820 97700 133980
rect 99890 133820 100890 133980
rect 103080 133820 104080 133980
rect 106270 133820 107270 133980
rect 109460 133820 110460 133980
rect 112650 133820 113650 133980
rect 115840 133820 116840 133980
rect 119030 133820 120030 133980
rect 122220 133820 123220 133980
rect 125410 133820 126410 133980
rect 128600 133820 129600 133980
rect 131790 133820 132790 133980
rect 134980 133820 135980 133980
rect 9320 132790 9410 133820
rect 9570 133797 12600 133820
rect 9570 132790 9593 133797
rect 9320 131790 9593 132790
rect 9320 130790 9410 131790
rect 9570 130813 9593 131790
rect 12577 132790 12600 133797
rect 12760 133797 15790 133820
rect 12760 132790 12783 133797
rect 12577 131790 12783 132790
rect 12577 130813 12600 131790
rect 9570 130790 12600 130813
rect 12760 130813 12783 131790
rect 15767 132790 15790 133797
rect 15950 133797 18980 133820
rect 15950 132790 15973 133797
rect 15767 131790 15973 132790
rect 15767 130813 15790 131790
rect 12760 130790 15790 130813
rect 15950 130813 15973 131790
rect 18957 132790 18980 133797
rect 19140 133797 22170 133820
rect 19140 132790 19163 133797
rect 18957 131790 19163 132790
rect 18957 130813 18980 131790
rect 15950 130790 18980 130813
rect 19140 130813 19163 131790
rect 22147 132790 22170 133797
rect 22330 133797 25360 133820
rect 22330 132790 22353 133797
rect 22147 131790 22353 132790
rect 22147 130813 22170 131790
rect 19140 130790 22170 130813
rect 22330 130813 22353 131790
rect 25337 132790 25360 133797
rect 25520 133797 28550 133820
rect 25520 132790 25543 133797
rect 25337 131790 25543 132790
rect 25337 130813 25360 131790
rect 22330 130790 25360 130813
rect 25520 130813 25543 131790
rect 28527 132790 28550 133797
rect 28710 133797 31740 133820
rect 28710 132790 28733 133797
rect 28527 131790 28733 132790
rect 28527 130813 28550 131790
rect 25520 130790 28550 130813
rect 28710 130813 28733 131790
rect 31717 132790 31740 133797
rect 31900 133797 34930 133820
rect 31900 132790 31923 133797
rect 31717 131790 31923 132790
rect 31717 130813 31740 131790
rect 28710 130790 31740 130813
rect 31900 130813 31923 131790
rect 34907 132790 34930 133797
rect 35090 133797 38120 133820
rect 35090 132790 35113 133797
rect 34907 131790 35113 132790
rect 34907 130813 34930 131790
rect 31900 130790 34930 130813
rect 35090 130813 35113 131790
rect 38097 132790 38120 133797
rect 38280 133797 41310 133820
rect 38280 132790 38303 133797
rect 38097 131790 38303 132790
rect 38097 130813 38120 131790
rect 35090 130790 38120 130813
rect 38280 130813 38303 131790
rect 41287 132790 41310 133797
rect 41470 133797 44500 133820
rect 41470 132790 41493 133797
rect 41287 131790 41493 132790
rect 41287 130813 41310 131790
rect 38280 130790 41310 130813
rect 41470 130813 41493 131790
rect 44477 132790 44500 133797
rect 44660 133797 47690 133820
rect 44660 132790 44683 133797
rect 44477 131790 44683 132790
rect 44477 130813 44500 131790
rect 41470 130790 44500 130813
rect 44660 130813 44683 131790
rect 47667 132790 47690 133797
rect 47850 133797 50880 133820
rect 47850 132790 47873 133797
rect 47667 131790 47873 132790
rect 47667 130813 47690 131790
rect 44660 130790 47690 130813
rect 47850 130813 47873 131790
rect 50857 132790 50880 133797
rect 51040 133797 54070 133820
rect 51040 132790 51063 133797
rect 50857 131790 51063 132790
rect 50857 130813 50880 131790
rect 47850 130790 50880 130813
rect 51040 130813 51063 131790
rect 54047 132790 54070 133797
rect 54230 133797 57260 133820
rect 54230 132790 54253 133797
rect 54047 131790 54253 132790
rect 54047 130813 54070 131790
rect 51040 130790 54070 130813
rect 54230 130813 54253 131790
rect 57237 132790 57260 133797
rect 57420 133797 60450 133820
rect 57420 132790 57443 133797
rect 57237 131790 57443 132790
rect 57237 130813 57260 131790
rect 54230 130790 57260 130813
rect 57420 130813 57443 131790
rect 60427 132790 60450 133797
rect 60610 133797 63640 133820
rect 60610 132790 60633 133797
rect 60427 131790 60633 132790
rect 60427 130813 60450 131790
rect 57420 130790 60450 130813
rect 60610 130813 60633 131790
rect 63617 132790 63640 133797
rect 63800 133797 66830 133820
rect 63800 132790 63823 133797
rect 63617 131790 63823 132790
rect 63617 130813 63640 131790
rect 60610 130790 63640 130813
rect 63800 130813 63823 131790
rect 66807 132790 66830 133797
rect 66990 133797 70020 133820
rect 66990 132790 67013 133797
rect 66807 131790 67013 132790
rect 66807 130813 66830 131790
rect 63800 130790 66830 130813
rect 66990 130813 67013 131790
rect 69997 132790 70020 133797
rect 70180 133797 73210 133820
rect 70180 132790 70203 133797
rect 69997 131790 70203 132790
rect 69997 130813 70020 131790
rect 66990 130790 70020 130813
rect 70180 130813 70203 131790
rect 73187 132790 73210 133797
rect 73370 133797 76400 133820
rect 73370 132790 73393 133797
rect 73187 131790 73393 132790
rect 73187 130813 73210 131790
rect 70180 130790 73210 130813
rect 73370 130813 73393 131790
rect 76377 132790 76400 133797
rect 76560 133797 79590 133820
rect 76560 132790 76583 133797
rect 76377 131790 76583 132790
rect 76377 130813 76400 131790
rect 73370 130790 76400 130813
rect 76560 130813 76583 131790
rect 79567 132790 79590 133797
rect 79750 133797 82780 133820
rect 79750 132790 79773 133797
rect 79567 131790 79773 132790
rect 79567 130813 79590 131790
rect 76560 130790 79590 130813
rect 79750 130813 79773 131790
rect 82757 132790 82780 133797
rect 82940 133797 85970 133820
rect 82940 132790 82963 133797
rect 82757 131790 82963 132790
rect 82757 130813 82780 131790
rect 79750 130790 82780 130813
rect 82940 130813 82963 131790
rect 85947 132790 85970 133797
rect 86130 133797 89160 133820
rect 86130 132790 86153 133797
rect 85947 131790 86153 132790
rect 85947 130813 85970 131790
rect 82940 130790 85970 130813
rect 86130 130813 86153 131790
rect 89137 132790 89160 133797
rect 89320 133797 92350 133820
rect 89320 132790 89343 133797
rect 89137 131790 89343 132790
rect 89137 130813 89160 131790
rect 86130 130790 89160 130813
rect 89320 130813 89343 131790
rect 92327 132790 92350 133797
rect 92510 133797 95540 133820
rect 92510 132790 92533 133797
rect 92327 131790 92533 132790
rect 92327 130813 92350 131790
rect 89320 130790 92350 130813
rect 92510 130813 92533 131790
rect 95517 132790 95540 133797
rect 95700 133797 98730 133820
rect 95700 132790 95723 133797
rect 95517 131790 95723 132790
rect 95517 130813 95540 131790
rect 92510 130790 95540 130813
rect 95700 130813 95723 131790
rect 98707 132790 98730 133797
rect 98890 133797 101920 133820
rect 98890 132790 98913 133797
rect 98707 131790 98913 132790
rect 98707 130813 98730 131790
rect 95700 130790 98730 130813
rect 98890 130813 98913 131790
rect 101897 132790 101920 133797
rect 102080 133797 105110 133820
rect 102080 132790 102103 133797
rect 101897 131790 102103 132790
rect 101897 130813 101920 131790
rect 98890 130790 101920 130813
rect 102080 130813 102103 131790
rect 105087 132790 105110 133797
rect 105270 133797 108300 133820
rect 105270 132790 105293 133797
rect 105087 131790 105293 132790
rect 105087 130813 105110 131790
rect 102080 130790 105110 130813
rect 105270 130813 105293 131790
rect 108277 132790 108300 133797
rect 108460 133797 111490 133820
rect 108460 132790 108483 133797
rect 108277 131790 108483 132790
rect 108277 130813 108300 131790
rect 105270 130790 108300 130813
rect 108460 130813 108483 131790
rect 111467 132790 111490 133797
rect 111650 133797 114680 133820
rect 111650 132790 111673 133797
rect 111467 131790 111673 132790
rect 111467 130813 111490 131790
rect 108460 130790 111490 130813
rect 111650 130813 111673 131790
rect 114657 132790 114680 133797
rect 114840 133797 117870 133820
rect 114840 132790 114863 133797
rect 114657 131790 114863 132790
rect 114657 130813 114680 131790
rect 111650 130790 114680 130813
rect 114840 130813 114863 131790
rect 117847 132790 117870 133797
rect 118030 133797 121060 133820
rect 118030 132790 118053 133797
rect 117847 131790 118053 132790
rect 117847 130813 117870 131790
rect 114840 130790 117870 130813
rect 118030 130813 118053 131790
rect 121037 132790 121060 133797
rect 121220 133797 124250 133820
rect 121220 132790 121243 133797
rect 121037 131790 121243 132790
rect 121037 130813 121060 131790
rect 118030 130790 121060 130813
rect 121220 130813 121243 131790
rect 124227 132790 124250 133797
rect 124410 133797 127440 133820
rect 124410 132790 124433 133797
rect 124227 131790 124433 132790
rect 124227 130813 124250 131790
rect 121220 130790 124250 130813
rect 124410 130813 124433 131790
rect 127417 132790 127440 133797
rect 127600 133797 130630 133820
rect 127600 132790 127623 133797
rect 127417 131790 127623 132790
rect 127417 130813 127440 131790
rect 124410 130790 127440 130813
rect 127600 130813 127623 131790
rect 130607 132790 130630 133797
rect 130790 133797 133820 133820
rect 130790 132790 130813 133797
rect 130607 131790 130813 132790
rect 130607 130813 130630 131790
rect 127600 130790 130630 130813
rect 130790 130813 130813 131790
rect 133797 132790 133820 133797
rect 133980 133797 137010 133820
rect 133980 132790 134003 133797
rect 133797 131790 134003 132790
rect 133797 130813 133820 131790
rect 130790 130790 133820 130813
rect 133980 130813 134003 131790
rect 136987 132790 137010 133797
rect 136987 131790 137170 132790
rect 136987 130813 137010 131790
rect 133980 130790 137010 130813
rect 9320 130630 9370 130790
rect 10570 130630 11570 130790
rect 13760 130630 14760 130790
rect 16950 130630 17950 130790
rect 20140 130630 21140 130790
rect 23330 130630 24330 130790
rect 26520 130630 27520 130790
rect 29710 130630 30710 130790
rect 32900 130630 33900 130790
rect 36090 130630 37090 130790
rect 39280 130630 40280 130790
rect 42470 130630 43470 130790
rect 45660 130630 46660 130790
rect 48850 130630 49850 130790
rect 52040 130630 53040 130790
rect 55230 130630 56230 130790
rect 58420 130630 59420 130790
rect 61610 130630 62610 130790
rect 64800 130630 65800 130790
rect 67990 130630 68990 130790
rect 71180 130630 72180 130790
rect 74370 130630 75370 130790
rect 77560 130630 78560 130790
rect 80750 130630 81750 130790
rect 83940 130630 84940 130790
rect 87130 130630 88130 130790
rect 90320 130630 91320 130790
rect 93510 130630 94510 130790
rect 96700 130630 97700 130790
rect 99890 130630 100890 130790
rect 103080 130630 104080 130790
rect 106270 130630 107270 130790
rect 109460 130630 110460 130790
rect 112650 130630 113650 130790
rect 115840 130630 116840 130790
rect 119030 130630 120030 130790
rect 122220 130630 123220 130790
rect 125410 130630 126410 130790
rect 128600 130630 129600 130790
rect 131790 130630 132790 130790
rect 134980 130630 135980 130790
rect 9320 129600 9410 130630
rect 9570 130607 12600 130630
rect 9570 129600 9593 130607
rect 9320 128600 9593 129600
rect 9320 127600 9410 128600
rect 9570 127623 9593 128600
rect 12577 129600 12600 130607
rect 12760 130607 15790 130630
rect 12760 129600 12783 130607
rect 12577 128600 12783 129600
rect 12577 127623 12600 128600
rect 9570 127600 12600 127623
rect 12760 127623 12783 128600
rect 15767 129600 15790 130607
rect 15950 130607 18980 130630
rect 15950 129600 15973 130607
rect 15767 128600 15973 129600
rect 15767 127623 15790 128600
rect 12760 127600 15790 127623
rect 15950 127623 15973 128600
rect 18957 129600 18980 130607
rect 19140 130607 22170 130630
rect 19140 129600 19163 130607
rect 18957 128600 19163 129600
rect 18957 127623 18980 128600
rect 15950 127600 18980 127623
rect 19140 127623 19163 128600
rect 22147 129600 22170 130607
rect 22330 130607 25360 130630
rect 22330 129600 22353 130607
rect 22147 128600 22353 129600
rect 22147 127623 22170 128600
rect 19140 127600 22170 127623
rect 22330 127623 22353 128600
rect 25337 129600 25360 130607
rect 25520 130607 28550 130630
rect 25520 129600 25543 130607
rect 25337 128600 25543 129600
rect 25337 127623 25360 128600
rect 22330 127600 25360 127623
rect 25520 127623 25543 128600
rect 28527 129600 28550 130607
rect 28710 130607 31740 130630
rect 28710 129600 28733 130607
rect 28527 128600 28733 129600
rect 28527 127623 28550 128600
rect 25520 127600 28550 127623
rect 28710 127623 28733 128600
rect 31717 129600 31740 130607
rect 31900 130607 34930 130630
rect 31900 129600 31923 130607
rect 31717 128600 31923 129600
rect 31717 127623 31740 128600
rect 28710 127600 31740 127623
rect 31900 127623 31923 128600
rect 34907 129600 34930 130607
rect 35090 130607 38120 130630
rect 35090 129600 35113 130607
rect 34907 128600 35113 129600
rect 34907 127623 34930 128600
rect 31900 127600 34930 127623
rect 35090 127623 35113 128600
rect 38097 129600 38120 130607
rect 38280 130607 41310 130630
rect 38280 129600 38303 130607
rect 38097 128600 38303 129600
rect 38097 127623 38120 128600
rect 35090 127600 38120 127623
rect 38280 127623 38303 128600
rect 41287 129600 41310 130607
rect 41470 130607 44500 130630
rect 41470 129600 41493 130607
rect 41287 128600 41493 129600
rect 41287 127623 41310 128600
rect 38280 127600 41310 127623
rect 41470 127623 41493 128600
rect 44477 129600 44500 130607
rect 44660 130607 47690 130630
rect 44660 129600 44683 130607
rect 44477 128600 44683 129600
rect 44477 127623 44500 128600
rect 41470 127600 44500 127623
rect 44660 127623 44683 128600
rect 47667 129600 47690 130607
rect 47850 130607 50880 130630
rect 47850 129600 47873 130607
rect 47667 128600 47873 129600
rect 47667 127623 47690 128600
rect 44660 127600 47690 127623
rect 47850 127623 47873 128600
rect 50857 129600 50880 130607
rect 51040 130607 54070 130630
rect 51040 129600 51063 130607
rect 50857 128600 51063 129600
rect 50857 127623 50880 128600
rect 47850 127600 50880 127623
rect 51040 127623 51063 128600
rect 54047 129600 54070 130607
rect 54230 130607 57260 130630
rect 54230 129600 54253 130607
rect 54047 128600 54253 129600
rect 54047 127623 54070 128600
rect 51040 127600 54070 127623
rect 54230 127623 54253 128600
rect 57237 129600 57260 130607
rect 57420 130607 60450 130630
rect 57420 129600 57443 130607
rect 57237 128600 57443 129600
rect 57237 127623 57260 128600
rect 54230 127600 57260 127623
rect 57420 127623 57443 128600
rect 60427 129600 60450 130607
rect 60610 130607 63640 130630
rect 60610 129600 60633 130607
rect 60427 128600 60633 129600
rect 60427 127623 60450 128600
rect 57420 127600 60450 127623
rect 60610 127623 60633 128600
rect 63617 129600 63640 130607
rect 63800 130607 66830 130630
rect 63800 129600 63823 130607
rect 63617 128600 63823 129600
rect 63617 127623 63640 128600
rect 60610 127600 63640 127623
rect 63800 127623 63823 128600
rect 66807 129600 66830 130607
rect 66990 130607 70020 130630
rect 66990 129600 67013 130607
rect 66807 128600 67013 129600
rect 66807 127623 66830 128600
rect 63800 127600 66830 127623
rect 66990 127623 67013 128600
rect 69997 129600 70020 130607
rect 70180 130607 73210 130630
rect 70180 129600 70203 130607
rect 69997 128600 70203 129600
rect 69997 127623 70020 128600
rect 66990 127600 70020 127623
rect 70180 127623 70203 128600
rect 73187 129600 73210 130607
rect 73370 130607 76400 130630
rect 73370 129600 73393 130607
rect 73187 128600 73393 129600
rect 73187 127623 73210 128600
rect 70180 127600 73210 127623
rect 73370 127623 73393 128600
rect 76377 129600 76400 130607
rect 76560 130607 79590 130630
rect 76560 129600 76583 130607
rect 76377 128600 76583 129600
rect 76377 127623 76400 128600
rect 73370 127600 76400 127623
rect 76560 127623 76583 128600
rect 79567 129600 79590 130607
rect 79750 130607 82780 130630
rect 79750 129600 79773 130607
rect 79567 128600 79773 129600
rect 79567 127623 79590 128600
rect 76560 127600 79590 127623
rect 79750 127623 79773 128600
rect 82757 129600 82780 130607
rect 82940 130607 85970 130630
rect 82940 129600 82963 130607
rect 82757 128600 82963 129600
rect 82757 127623 82780 128600
rect 79750 127600 82780 127623
rect 82940 127623 82963 128600
rect 85947 129600 85970 130607
rect 86130 130607 89160 130630
rect 86130 129600 86153 130607
rect 85947 128600 86153 129600
rect 85947 127623 85970 128600
rect 82940 127600 85970 127623
rect 86130 127623 86153 128600
rect 89137 129600 89160 130607
rect 89320 130607 92350 130630
rect 89320 129600 89343 130607
rect 89137 128600 89343 129600
rect 89137 127623 89160 128600
rect 86130 127600 89160 127623
rect 89320 127623 89343 128600
rect 92327 129600 92350 130607
rect 92510 130607 95540 130630
rect 92510 129600 92533 130607
rect 92327 128600 92533 129600
rect 92327 127623 92350 128600
rect 89320 127600 92350 127623
rect 92510 127623 92533 128600
rect 95517 129600 95540 130607
rect 95700 130607 98730 130630
rect 95700 129600 95723 130607
rect 95517 128600 95723 129600
rect 95517 127623 95540 128600
rect 92510 127600 95540 127623
rect 95700 127623 95723 128600
rect 98707 129600 98730 130607
rect 98890 130607 101920 130630
rect 98890 129600 98913 130607
rect 98707 128600 98913 129600
rect 98707 127623 98730 128600
rect 95700 127600 98730 127623
rect 98890 127623 98913 128600
rect 101897 129600 101920 130607
rect 102080 130607 105110 130630
rect 102080 129600 102103 130607
rect 101897 128600 102103 129600
rect 101897 127623 101920 128600
rect 98890 127600 101920 127623
rect 102080 127623 102103 128600
rect 105087 129600 105110 130607
rect 105270 130607 108300 130630
rect 105270 129600 105293 130607
rect 105087 128600 105293 129600
rect 105087 127623 105110 128600
rect 102080 127600 105110 127623
rect 105270 127623 105293 128600
rect 108277 129600 108300 130607
rect 108460 130607 111490 130630
rect 108460 129600 108483 130607
rect 108277 128600 108483 129600
rect 108277 127623 108300 128600
rect 105270 127600 108300 127623
rect 108460 127623 108483 128600
rect 111467 129600 111490 130607
rect 111650 130607 114680 130630
rect 111650 129600 111673 130607
rect 111467 128600 111673 129600
rect 111467 127623 111490 128600
rect 108460 127600 111490 127623
rect 111650 127623 111673 128600
rect 114657 129600 114680 130607
rect 114840 130607 117870 130630
rect 114840 129600 114863 130607
rect 114657 128600 114863 129600
rect 114657 127623 114680 128600
rect 111650 127600 114680 127623
rect 114840 127623 114863 128600
rect 117847 129600 117870 130607
rect 118030 130607 121060 130630
rect 118030 129600 118053 130607
rect 117847 128600 118053 129600
rect 117847 127623 117870 128600
rect 114840 127600 117870 127623
rect 118030 127623 118053 128600
rect 121037 129600 121060 130607
rect 121220 130607 124250 130630
rect 121220 129600 121243 130607
rect 121037 128600 121243 129600
rect 121037 127623 121060 128600
rect 118030 127600 121060 127623
rect 121220 127623 121243 128600
rect 124227 129600 124250 130607
rect 124410 130607 127440 130630
rect 124410 129600 124433 130607
rect 124227 128600 124433 129600
rect 124227 127623 124250 128600
rect 121220 127600 124250 127623
rect 124410 127623 124433 128600
rect 127417 129600 127440 130607
rect 127600 130607 130630 130630
rect 127600 129600 127623 130607
rect 127417 128600 127623 129600
rect 127417 127623 127440 128600
rect 124410 127600 127440 127623
rect 127600 127623 127623 128600
rect 130607 129600 130630 130607
rect 130790 130607 133820 130630
rect 130790 129600 130813 130607
rect 130607 128600 130813 129600
rect 130607 127623 130630 128600
rect 127600 127600 130630 127623
rect 130790 127623 130813 128600
rect 133797 129600 133820 130607
rect 133980 130607 137010 130630
rect 133980 129600 134003 130607
rect 133797 128600 134003 129600
rect 133797 127623 133820 128600
rect 130790 127600 133820 127623
rect 133980 127623 134003 128600
rect 136987 129600 137010 130607
rect 136987 128600 137170 129600
rect 136987 127623 137010 128600
rect 133980 127600 137010 127623
rect 9320 127440 9370 127600
rect 10570 127440 11570 127600
rect 13760 127440 14760 127600
rect 16950 127440 17950 127600
rect 20140 127440 21140 127600
rect 23330 127440 24330 127600
rect 26520 127440 27520 127600
rect 29710 127440 30710 127600
rect 32900 127440 33900 127600
rect 36090 127440 37090 127600
rect 39280 127440 40280 127600
rect 42470 127440 43470 127600
rect 45660 127440 46660 127600
rect 48850 127440 49850 127600
rect 52040 127440 53040 127600
rect 55230 127440 56230 127600
rect 58420 127440 59420 127600
rect 61610 127440 62610 127600
rect 64800 127440 65800 127600
rect 67990 127440 68990 127600
rect 71180 127440 72180 127600
rect 74370 127440 75370 127600
rect 77560 127440 78560 127600
rect 80750 127440 81750 127600
rect 83940 127440 84940 127600
rect 87130 127440 88130 127600
rect 90320 127440 91320 127600
rect 93510 127440 94510 127600
rect 96700 127440 97700 127600
rect 99890 127440 100890 127600
rect 103080 127440 104080 127600
rect 106270 127440 107270 127600
rect 109460 127440 110460 127600
rect 112650 127440 113650 127600
rect 115840 127440 116840 127600
rect 119030 127440 120030 127600
rect 122220 127440 123220 127600
rect 125410 127440 126410 127600
rect 128600 127440 129600 127600
rect 131790 127440 132790 127600
rect 134980 127440 135980 127600
rect 9320 126410 9410 127440
rect 9570 127417 12600 127440
rect 9570 126410 9593 127417
rect 9320 125410 9593 126410
rect 9320 124410 9410 125410
rect 9570 124433 9593 125410
rect 12577 126410 12600 127417
rect 12760 127417 15790 127440
rect 12760 126410 12783 127417
rect 12577 125410 12783 126410
rect 12577 124433 12600 125410
rect 9570 124410 12600 124433
rect 12760 124433 12783 125410
rect 15767 126410 15790 127417
rect 15950 127417 18980 127440
rect 15950 126410 15973 127417
rect 15767 125410 15973 126410
rect 15767 124433 15790 125410
rect 12760 124410 15790 124433
rect 15950 124433 15973 125410
rect 18957 126410 18980 127417
rect 19140 127417 22170 127440
rect 19140 126410 19163 127417
rect 18957 125410 19163 126410
rect 18957 124433 18980 125410
rect 15950 124410 18980 124433
rect 19140 124433 19163 125410
rect 22147 126410 22170 127417
rect 22330 127417 25360 127440
rect 22330 126410 22353 127417
rect 22147 125410 22353 126410
rect 22147 124433 22170 125410
rect 19140 124410 22170 124433
rect 22330 124433 22353 125410
rect 25337 126410 25360 127417
rect 25520 127417 28550 127440
rect 25520 126410 25543 127417
rect 25337 125410 25543 126410
rect 25337 124433 25360 125410
rect 22330 124410 25360 124433
rect 25520 124433 25543 125410
rect 28527 126410 28550 127417
rect 28710 127417 31740 127440
rect 28710 126410 28733 127417
rect 28527 125410 28733 126410
rect 28527 124433 28550 125410
rect 25520 124410 28550 124433
rect 28710 124433 28733 125410
rect 31717 126410 31740 127417
rect 31900 127417 34930 127440
rect 31900 126410 31923 127417
rect 31717 125410 31923 126410
rect 31717 124433 31740 125410
rect 28710 124410 31740 124433
rect 31900 124433 31923 125410
rect 34907 126410 34930 127417
rect 35090 127417 38120 127440
rect 35090 126410 35113 127417
rect 34907 125410 35113 126410
rect 34907 124433 34930 125410
rect 31900 124410 34930 124433
rect 35090 124433 35113 125410
rect 38097 126410 38120 127417
rect 38280 127417 41310 127440
rect 38280 126410 38303 127417
rect 38097 125410 38303 126410
rect 38097 124433 38120 125410
rect 35090 124410 38120 124433
rect 38280 124433 38303 125410
rect 41287 126410 41310 127417
rect 41470 127417 44500 127440
rect 41470 126410 41493 127417
rect 41287 125410 41493 126410
rect 41287 124433 41310 125410
rect 38280 124410 41310 124433
rect 41470 124433 41493 125410
rect 44477 126410 44500 127417
rect 44660 127417 47690 127440
rect 44660 126410 44683 127417
rect 44477 125410 44683 126410
rect 44477 124433 44500 125410
rect 41470 124410 44500 124433
rect 44660 124433 44683 125410
rect 47667 126410 47690 127417
rect 47850 127417 50880 127440
rect 47850 126410 47873 127417
rect 47667 125410 47873 126410
rect 47667 124433 47690 125410
rect 44660 124410 47690 124433
rect 47850 124433 47873 125410
rect 50857 126410 50880 127417
rect 51040 127417 54070 127440
rect 51040 126410 51063 127417
rect 50857 125410 51063 126410
rect 50857 124433 50880 125410
rect 47850 124410 50880 124433
rect 51040 124433 51063 125410
rect 54047 126410 54070 127417
rect 54230 127417 57260 127440
rect 54230 126410 54253 127417
rect 54047 125410 54253 126410
rect 54047 124433 54070 125410
rect 51040 124410 54070 124433
rect 54230 124433 54253 125410
rect 57237 126410 57260 127417
rect 57420 127417 60450 127440
rect 57420 126410 57443 127417
rect 57237 125410 57443 126410
rect 57237 124433 57260 125410
rect 54230 124410 57260 124433
rect 57420 124433 57443 125410
rect 60427 126410 60450 127417
rect 60610 127417 63640 127440
rect 60610 126410 60633 127417
rect 60427 125410 60633 126410
rect 60427 124433 60450 125410
rect 57420 124410 60450 124433
rect 60610 124433 60633 125410
rect 63617 126410 63640 127417
rect 63800 127417 66830 127440
rect 63800 126410 63823 127417
rect 63617 125410 63823 126410
rect 63617 124433 63640 125410
rect 60610 124410 63640 124433
rect 63800 124433 63823 125410
rect 66807 126410 66830 127417
rect 66990 127417 70020 127440
rect 66990 126410 67013 127417
rect 66807 125410 67013 126410
rect 66807 124433 66830 125410
rect 63800 124410 66830 124433
rect 66990 124433 67013 125410
rect 69997 126410 70020 127417
rect 70180 127417 73210 127440
rect 70180 126410 70203 127417
rect 69997 125410 70203 126410
rect 69997 124433 70020 125410
rect 66990 124410 70020 124433
rect 70180 124433 70203 125410
rect 73187 126410 73210 127417
rect 73370 127417 76400 127440
rect 73370 126410 73393 127417
rect 73187 125410 73393 126410
rect 73187 124433 73210 125410
rect 70180 124410 73210 124433
rect 73370 124433 73393 125410
rect 76377 126410 76400 127417
rect 76560 127417 79590 127440
rect 76560 126410 76583 127417
rect 76377 125410 76583 126410
rect 76377 124433 76400 125410
rect 73370 124410 76400 124433
rect 76560 124433 76583 125410
rect 79567 126410 79590 127417
rect 79750 127417 82780 127440
rect 79750 126410 79773 127417
rect 79567 125410 79773 126410
rect 79567 124433 79590 125410
rect 76560 124410 79590 124433
rect 79750 124433 79773 125410
rect 82757 126410 82780 127417
rect 82940 127417 85970 127440
rect 82940 126410 82963 127417
rect 82757 125410 82963 126410
rect 82757 124433 82780 125410
rect 79750 124410 82780 124433
rect 82940 124433 82963 125410
rect 85947 126410 85970 127417
rect 86130 127417 89160 127440
rect 86130 126410 86153 127417
rect 85947 125410 86153 126410
rect 85947 124433 85970 125410
rect 82940 124410 85970 124433
rect 86130 124433 86153 125410
rect 89137 126410 89160 127417
rect 89320 127417 92350 127440
rect 89320 126410 89343 127417
rect 89137 125410 89343 126410
rect 89137 124433 89160 125410
rect 86130 124410 89160 124433
rect 89320 124433 89343 125410
rect 92327 126410 92350 127417
rect 92510 127417 95540 127440
rect 92510 126410 92533 127417
rect 92327 125410 92533 126410
rect 92327 124433 92350 125410
rect 89320 124410 92350 124433
rect 92510 124433 92533 125410
rect 95517 126410 95540 127417
rect 95700 127417 98730 127440
rect 95700 126410 95723 127417
rect 95517 125410 95723 126410
rect 95517 124433 95540 125410
rect 92510 124410 95540 124433
rect 95700 124433 95723 125410
rect 98707 126410 98730 127417
rect 98890 127417 101920 127440
rect 98890 126410 98913 127417
rect 98707 125410 98913 126410
rect 98707 124433 98730 125410
rect 95700 124410 98730 124433
rect 98890 124433 98913 125410
rect 101897 126410 101920 127417
rect 102080 127417 105110 127440
rect 102080 126410 102103 127417
rect 101897 125410 102103 126410
rect 101897 124433 101920 125410
rect 98890 124410 101920 124433
rect 102080 124433 102103 125410
rect 105087 126410 105110 127417
rect 105270 127417 108300 127440
rect 105270 126410 105293 127417
rect 105087 125410 105293 126410
rect 105087 124433 105110 125410
rect 102080 124410 105110 124433
rect 105270 124433 105293 125410
rect 108277 126410 108300 127417
rect 108460 127417 111490 127440
rect 108460 126410 108483 127417
rect 108277 125410 108483 126410
rect 108277 124433 108300 125410
rect 105270 124410 108300 124433
rect 108460 124433 108483 125410
rect 111467 126410 111490 127417
rect 111650 127417 114680 127440
rect 111650 126410 111673 127417
rect 111467 125410 111673 126410
rect 111467 124433 111490 125410
rect 108460 124410 111490 124433
rect 111650 124433 111673 125410
rect 114657 126410 114680 127417
rect 114840 127417 117870 127440
rect 114840 126410 114863 127417
rect 114657 125410 114863 126410
rect 114657 124433 114680 125410
rect 111650 124410 114680 124433
rect 114840 124433 114863 125410
rect 117847 126410 117870 127417
rect 118030 127417 121060 127440
rect 118030 126410 118053 127417
rect 117847 125410 118053 126410
rect 117847 124433 117870 125410
rect 114840 124410 117870 124433
rect 118030 124433 118053 125410
rect 121037 126410 121060 127417
rect 121220 127417 124250 127440
rect 121220 126410 121243 127417
rect 121037 125410 121243 126410
rect 121037 124433 121060 125410
rect 118030 124410 121060 124433
rect 121220 124433 121243 125410
rect 124227 126410 124250 127417
rect 124410 127417 127440 127440
rect 124410 126410 124433 127417
rect 124227 125410 124433 126410
rect 124227 124433 124250 125410
rect 121220 124410 124250 124433
rect 124410 124433 124433 125410
rect 127417 126410 127440 127417
rect 127600 127417 130630 127440
rect 127600 126410 127623 127417
rect 127417 125410 127623 126410
rect 127417 124433 127440 125410
rect 124410 124410 127440 124433
rect 127600 124433 127623 125410
rect 130607 126410 130630 127417
rect 130790 127417 133820 127440
rect 130790 126410 130813 127417
rect 130607 125410 130813 126410
rect 130607 124433 130630 125410
rect 127600 124410 130630 124433
rect 130790 124433 130813 125410
rect 133797 126410 133820 127417
rect 133980 127417 137010 127440
rect 133980 126410 134003 127417
rect 133797 125410 134003 126410
rect 133797 124433 133820 125410
rect 130790 124410 133820 124433
rect 133980 124433 134003 125410
rect 136987 126410 137010 127417
rect 136987 125410 137170 126410
rect 136987 124433 137010 125410
rect 133980 124410 137010 124433
rect 9320 124250 9370 124410
rect 10570 124250 11570 124410
rect 13760 124250 14760 124410
rect 16950 124250 17950 124410
rect 20140 124250 21140 124410
rect 23330 124250 24330 124410
rect 26520 124250 27520 124410
rect 29710 124250 30710 124410
rect 32900 124250 33900 124410
rect 36090 124250 37090 124410
rect 39280 124250 40280 124410
rect 42470 124250 43470 124410
rect 45660 124250 46660 124410
rect 48850 124250 49850 124410
rect 52040 124250 53040 124410
rect 55230 124250 56230 124410
rect 58420 124250 59420 124410
rect 61610 124250 62610 124410
rect 64800 124250 65800 124410
rect 67990 124250 68990 124410
rect 71180 124250 72180 124410
rect 74370 124250 75370 124410
rect 77560 124250 78560 124410
rect 80750 124250 81750 124410
rect 83940 124250 84940 124410
rect 87130 124250 88130 124410
rect 90320 124250 91320 124410
rect 93510 124250 94510 124410
rect 96700 124250 97700 124410
rect 99890 124250 100890 124410
rect 103080 124250 104080 124410
rect 106270 124250 107270 124410
rect 109460 124250 110460 124410
rect 112650 124250 113650 124410
rect 115840 124250 116840 124410
rect 119030 124250 120030 124410
rect 122220 124250 123220 124410
rect 125410 124250 126410 124410
rect 128600 124250 129600 124410
rect 131790 124250 132790 124410
rect 134980 124250 135980 124410
rect 9320 123220 9410 124250
rect 9570 124227 12600 124250
rect 9570 123220 9593 124227
rect 9320 122220 9593 123220
rect 9320 121310 9410 122220
rect 0 121260 9410 121310
rect 0 121220 3030 121260
rect 3190 121220 6220 121260
rect 6380 121220 9410 121260
rect 9570 121243 9593 122220
rect 12577 123220 12600 124227
rect 12760 124227 15790 124250
rect 12760 123220 12783 124227
rect 12577 122220 12783 123220
rect 12577 121243 12600 122220
rect 9570 121220 12600 121243
rect 12760 121243 12783 122220
rect 15767 123220 15790 124227
rect 15950 124227 18980 124250
rect 15950 123220 15973 124227
rect 15767 122220 15973 123220
rect 15767 121243 15790 122220
rect 12760 121220 15790 121243
rect 15950 121243 15973 122220
rect 18957 123220 18980 124227
rect 19140 124227 22170 124250
rect 19140 123220 19163 124227
rect 18957 122220 19163 123220
rect 18957 121243 18980 122220
rect 15950 121220 18980 121243
rect 19140 121243 19163 122220
rect 22147 123220 22170 124227
rect 22330 124227 25360 124250
rect 22330 123220 22353 124227
rect 22147 122220 22353 123220
rect 22147 121243 22170 122220
rect 19140 121220 22170 121243
rect 22330 121243 22353 122220
rect 25337 123220 25360 124227
rect 25520 124227 28550 124250
rect 25520 123220 25543 124227
rect 25337 122220 25543 123220
rect 25337 121243 25360 122220
rect 22330 121220 25360 121243
rect 25520 121243 25543 122220
rect 28527 123220 28550 124227
rect 28710 124227 31740 124250
rect 28710 123220 28733 124227
rect 28527 122220 28733 123220
rect 28527 121243 28550 122220
rect 25520 121220 28550 121243
rect 28710 121243 28733 122220
rect 31717 123220 31740 124227
rect 31900 124227 34930 124250
rect 31900 123220 31923 124227
rect 31717 122220 31923 123220
rect 31717 121243 31740 122220
rect 28710 121220 31740 121243
rect 31900 121243 31923 122220
rect 34907 123220 34930 124227
rect 35090 124227 38120 124250
rect 35090 123220 35113 124227
rect 34907 122220 35113 123220
rect 34907 121243 34930 122220
rect 31900 121220 34930 121243
rect 35090 121243 35113 122220
rect 38097 123220 38120 124227
rect 38280 124227 41310 124250
rect 38280 123220 38303 124227
rect 38097 122220 38303 123220
rect 38097 121243 38120 122220
rect 35090 121220 38120 121243
rect 38280 121243 38303 122220
rect 41287 123220 41310 124227
rect 41470 124227 44500 124250
rect 41470 123220 41493 124227
rect 41287 122220 41493 123220
rect 41287 121243 41310 122220
rect 38280 121220 41310 121243
rect 41470 121243 41493 122220
rect 44477 123220 44500 124227
rect 44660 124227 47690 124250
rect 44660 123220 44683 124227
rect 44477 122220 44683 123220
rect 44477 121243 44500 122220
rect 41470 121220 44500 121243
rect 44660 121243 44683 122220
rect 47667 123220 47690 124227
rect 47850 124227 50880 124250
rect 47850 123220 47873 124227
rect 47667 122220 47873 123220
rect 47667 121243 47690 122220
rect 44660 121220 47690 121243
rect 47850 121243 47873 122220
rect 50857 123220 50880 124227
rect 51040 124227 54070 124250
rect 51040 123220 51063 124227
rect 50857 122220 51063 123220
rect 50857 121243 50880 122220
rect 47850 121220 50880 121243
rect 51040 121243 51063 122220
rect 54047 123220 54070 124227
rect 54230 124227 57260 124250
rect 54230 123220 54253 124227
rect 54047 122220 54253 123220
rect 54047 121243 54070 122220
rect 51040 121220 54070 121243
rect 54230 121243 54253 122220
rect 57237 123220 57260 124227
rect 57420 124227 60450 124250
rect 57420 123220 57443 124227
rect 57237 122220 57443 123220
rect 57237 121243 57260 122220
rect 54230 121220 57260 121243
rect 57420 121243 57443 122220
rect 60427 123220 60450 124227
rect 60610 124227 63640 124250
rect 60610 123220 60633 124227
rect 60427 122220 60633 123220
rect 60427 121243 60450 122220
rect 57420 121220 60450 121243
rect 60610 121243 60633 122220
rect 63617 123220 63640 124227
rect 63800 124227 66830 124250
rect 63800 123220 63823 124227
rect 63617 122220 63823 123220
rect 63617 121243 63640 122220
rect 60610 121220 63640 121243
rect 63800 121243 63823 122220
rect 66807 123220 66830 124227
rect 66990 124227 70020 124250
rect 66990 123220 67013 124227
rect 66807 122220 67013 123220
rect 66807 121243 66830 122220
rect 63800 121220 66830 121243
rect 66990 121243 67013 122220
rect 69997 123220 70020 124227
rect 70180 124227 73210 124250
rect 70180 123220 70203 124227
rect 69997 122220 70203 123220
rect 69997 121243 70020 122220
rect 66990 121220 70020 121243
rect 70180 121243 70203 122220
rect 73187 123220 73210 124227
rect 73370 124227 76400 124250
rect 73370 123220 73393 124227
rect 73187 122220 73393 123220
rect 73187 121243 73210 122220
rect 70180 121220 73210 121243
rect 73370 121243 73393 122220
rect 76377 123220 76400 124227
rect 76560 124227 79590 124250
rect 76560 123220 76583 124227
rect 76377 122220 76583 123220
rect 76377 121243 76400 122220
rect 73370 121220 76400 121243
rect 76560 121243 76583 122220
rect 79567 123220 79590 124227
rect 79750 124227 82780 124250
rect 79750 123220 79773 124227
rect 79567 122220 79773 123220
rect 79567 121243 79590 122220
rect 76560 121220 79590 121243
rect 79750 121243 79773 122220
rect 82757 123220 82780 124227
rect 82940 124227 85970 124250
rect 82940 123220 82963 124227
rect 82757 122220 82963 123220
rect 82757 121243 82780 122220
rect 79750 121220 82780 121243
rect 82940 121243 82963 122220
rect 85947 123220 85970 124227
rect 86130 124227 89160 124250
rect 86130 123220 86153 124227
rect 85947 122220 86153 123220
rect 85947 121243 85970 122220
rect 82940 121220 85970 121243
rect 86130 121243 86153 122220
rect 89137 123220 89160 124227
rect 89320 124227 92350 124250
rect 89320 123220 89343 124227
rect 89137 122220 89343 123220
rect 89137 121243 89160 122220
rect 86130 121220 89160 121243
rect 89320 121243 89343 122220
rect 92327 123220 92350 124227
rect 92510 124227 95540 124250
rect 92510 123220 92533 124227
rect 92327 122220 92533 123220
rect 92327 121243 92350 122220
rect 89320 121220 92350 121243
rect 92510 121243 92533 122220
rect 95517 123220 95540 124227
rect 95700 124227 98730 124250
rect 95700 123220 95723 124227
rect 95517 122220 95723 123220
rect 95517 121243 95540 122220
rect 92510 121220 95540 121243
rect 95700 121243 95723 122220
rect 98707 123220 98730 124227
rect 98890 124227 101920 124250
rect 98890 123220 98913 124227
rect 98707 122220 98913 123220
rect 98707 121243 98730 122220
rect 95700 121220 98730 121243
rect 98890 121243 98913 122220
rect 101897 123220 101920 124227
rect 102080 124227 105110 124250
rect 102080 123220 102103 124227
rect 101897 122220 102103 123220
rect 101897 121243 101920 122220
rect 98890 121220 101920 121243
rect 102080 121243 102103 122220
rect 105087 123220 105110 124227
rect 105270 124227 108300 124250
rect 105270 123220 105293 124227
rect 105087 122220 105293 123220
rect 105087 121243 105110 122220
rect 102080 121220 105110 121243
rect 105270 121243 105293 122220
rect 108277 123220 108300 124227
rect 108460 124227 111490 124250
rect 108460 123220 108483 124227
rect 108277 122220 108483 123220
rect 108277 121243 108300 122220
rect 105270 121220 108300 121243
rect 108460 121243 108483 122220
rect 111467 123220 111490 124227
rect 111650 124227 114680 124250
rect 111650 123220 111673 124227
rect 111467 122220 111673 123220
rect 111467 121243 111490 122220
rect 108460 121220 111490 121243
rect 111650 121243 111673 122220
rect 114657 123220 114680 124227
rect 114840 124227 117870 124250
rect 114840 123220 114863 124227
rect 114657 122220 114863 123220
rect 114657 121243 114680 122220
rect 111650 121220 114680 121243
rect 114840 121243 114863 122220
rect 117847 123220 117870 124227
rect 118030 124227 121060 124250
rect 118030 123220 118053 124227
rect 117847 122220 118053 123220
rect 117847 121243 117870 122220
rect 114840 121220 117870 121243
rect 118030 121243 118053 122220
rect 121037 123220 121060 124227
rect 121220 124227 124250 124250
rect 121220 123220 121243 124227
rect 121037 122220 121243 123220
rect 121037 121243 121060 122220
rect 118030 121220 121060 121243
rect 121220 121243 121243 122220
rect 124227 123220 124250 124227
rect 124410 124227 127440 124250
rect 124410 123220 124433 124227
rect 124227 122220 124433 123220
rect 124227 121243 124250 122220
rect 121220 121220 124250 121243
rect 124410 121243 124433 122220
rect 127417 123220 127440 124227
rect 127600 124227 130630 124250
rect 127600 123220 127623 124227
rect 127417 122220 127623 123220
rect 127417 121243 127440 122220
rect 124410 121220 127440 121243
rect 127600 121243 127623 122220
rect 130607 123220 130630 124227
rect 130790 124227 133820 124250
rect 130790 123220 130813 124227
rect 130607 122220 130813 123220
rect 130607 121243 130630 122220
rect 127600 121220 130630 121243
rect 130790 121243 130813 122220
rect 133797 123220 133820 124227
rect 133980 124227 137010 124250
rect 133980 123220 134003 124227
rect 133797 122220 134003 123220
rect 133797 121243 133820 122220
rect 130790 121220 133820 121243
rect 133980 121243 134003 122220
rect 136987 123220 137010 124227
rect 136987 122220 137170 123220
rect 136987 121243 137010 122220
rect 133980 121220 137010 121243
rect 1000 121060 2000 121220
rect 4190 121060 5190 121220
rect 7380 121060 8380 121220
rect 10570 121060 11570 121220
rect 13760 121060 14760 121220
rect 16950 121060 17950 121220
rect 20140 121060 21140 121220
rect 23330 121060 24330 121220
rect 26520 121060 27520 121220
rect 29710 121060 30710 121220
rect 32900 121060 33900 121220
rect 36090 121060 37090 121220
rect 39280 121060 40280 121220
rect 42470 121060 43470 121220
rect 45660 121060 46660 121220
rect 48850 121060 49850 121220
rect 52040 121060 53040 121220
rect 55230 121060 56230 121220
rect 58420 121060 59420 121220
rect 61610 121060 62610 121220
rect 64800 121060 65800 121220
rect 67990 121060 68990 121220
rect 71180 121060 72180 121220
rect 74370 121060 75370 121220
rect 77560 121060 78560 121220
rect 80750 121060 81750 121220
rect 83940 121060 84940 121220
rect 87130 121060 88130 121220
rect 90320 121060 91320 121220
rect 93510 121060 94510 121220
rect 96700 121060 97700 121220
rect 99890 121060 100890 121220
rect 103080 121060 104080 121220
rect 106270 121060 107270 121220
rect 109460 121060 110460 121220
rect 112650 121060 113650 121220
rect 115840 121060 116840 121220
rect 119030 121060 120030 121220
rect 122220 121060 123220 121220
rect 125410 121060 126410 121220
rect 128600 121060 129600 121220
rect 131790 121060 132790 121220
rect 134980 121060 135980 121220
rect 0 121037 3030 121060
rect 0 118053 23 121037
rect 3007 120030 3030 121037
rect 3190 121037 6220 121060
rect 3190 120030 3213 121037
rect 3007 119030 3213 120030
rect 3007 118053 3030 119030
rect 0 118030 3030 118053
rect 3190 118053 3213 119030
rect 6197 120030 6220 121037
rect 6380 121037 9410 121060
rect 6380 120030 6403 121037
rect 6197 119030 6403 120030
rect 6197 118053 6220 119030
rect 3190 118030 6220 118053
rect 6380 118053 6403 119030
rect 9387 120030 9410 121037
rect 9570 121037 12600 121060
rect 9570 120030 9593 121037
rect 9387 119030 9593 120030
rect 9387 118053 9410 119030
rect 6380 118030 9410 118053
rect 9570 118053 9593 119030
rect 12577 120030 12600 121037
rect 12760 121037 15790 121060
rect 12760 120030 12783 121037
rect 12577 119030 12783 120030
rect 12577 118053 12600 119030
rect 9570 118030 12600 118053
rect 12760 118053 12783 119030
rect 15767 120030 15790 121037
rect 15950 121037 18980 121060
rect 15950 120030 15973 121037
rect 15767 119030 15973 120030
rect 15767 118053 15790 119030
rect 12760 118030 15790 118053
rect 15950 118053 15973 119030
rect 18957 120030 18980 121037
rect 19140 121037 22170 121060
rect 19140 120030 19163 121037
rect 18957 119030 19163 120030
rect 18957 118053 18980 119030
rect 15950 118030 18980 118053
rect 19140 118053 19163 119030
rect 22147 120030 22170 121037
rect 22330 121037 25360 121060
rect 22330 120030 22353 121037
rect 22147 119030 22353 120030
rect 22147 118053 22170 119030
rect 19140 118030 22170 118053
rect 22330 118053 22353 119030
rect 25337 120030 25360 121037
rect 25520 121037 28550 121060
rect 25520 120030 25543 121037
rect 25337 119030 25543 120030
rect 25337 118053 25360 119030
rect 22330 118030 25360 118053
rect 25520 118053 25543 119030
rect 28527 120030 28550 121037
rect 28710 121037 31740 121060
rect 28710 120030 28733 121037
rect 28527 119030 28733 120030
rect 28527 118053 28550 119030
rect 25520 118030 28550 118053
rect 28710 118053 28733 119030
rect 31717 120030 31740 121037
rect 31900 121037 34930 121060
rect 31900 120030 31923 121037
rect 31717 119030 31923 120030
rect 31717 118053 31740 119030
rect 28710 118030 31740 118053
rect 31900 118053 31923 119030
rect 34907 120030 34930 121037
rect 35090 121037 38120 121060
rect 35090 120030 35113 121037
rect 34907 119030 35113 120030
rect 34907 118053 34930 119030
rect 31900 118030 34930 118053
rect 35090 118053 35113 119030
rect 38097 120030 38120 121037
rect 38280 121037 41310 121060
rect 38280 120030 38303 121037
rect 38097 119030 38303 120030
rect 38097 118053 38120 119030
rect 35090 118030 38120 118053
rect 38280 118053 38303 119030
rect 41287 120030 41310 121037
rect 41470 121037 44500 121060
rect 41470 120030 41493 121037
rect 41287 119030 41493 120030
rect 41287 118053 41310 119030
rect 38280 118030 41310 118053
rect 41470 118053 41493 119030
rect 44477 120030 44500 121037
rect 44660 121037 47690 121060
rect 44660 120030 44683 121037
rect 44477 119030 44683 120030
rect 44477 118053 44500 119030
rect 41470 118030 44500 118053
rect 44660 118053 44683 119030
rect 47667 120030 47690 121037
rect 47850 121037 50880 121060
rect 47850 120030 47873 121037
rect 47667 119030 47873 120030
rect 47667 118053 47690 119030
rect 44660 118030 47690 118053
rect 47850 118053 47873 119030
rect 50857 120030 50880 121037
rect 51040 121037 54070 121060
rect 51040 120030 51063 121037
rect 50857 119030 51063 120030
rect 50857 118053 50880 119030
rect 47850 118030 50880 118053
rect 51040 118053 51063 119030
rect 54047 120030 54070 121037
rect 54230 121037 57260 121060
rect 54230 120030 54253 121037
rect 54047 119030 54253 120030
rect 54047 118053 54070 119030
rect 51040 118030 54070 118053
rect 54230 118053 54253 119030
rect 57237 120030 57260 121037
rect 57420 121037 60450 121060
rect 57420 120030 57443 121037
rect 57237 119030 57443 120030
rect 57237 118053 57260 119030
rect 54230 118030 57260 118053
rect 57420 118053 57443 119030
rect 60427 120030 60450 121037
rect 60610 121037 63640 121060
rect 60610 120030 60633 121037
rect 60427 119030 60633 120030
rect 60427 118053 60450 119030
rect 57420 118030 60450 118053
rect 60610 118053 60633 119030
rect 63617 120030 63640 121037
rect 63800 121037 66830 121060
rect 63800 120030 63823 121037
rect 63617 119030 63823 120030
rect 63617 118053 63640 119030
rect 60610 118030 63640 118053
rect 63800 118053 63823 119030
rect 66807 120030 66830 121037
rect 66990 121037 70020 121060
rect 66990 120030 67013 121037
rect 66807 119030 67013 120030
rect 66807 118053 66830 119030
rect 63800 118030 66830 118053
rect 66990 118053 67013 119030
rect 69997 120030 70020 121037
rect 70180 121037 73210 121060
rect 70180 120030 70203 121037
rect 69997 119030 70203 120030
rect 69997 118053 70020 119030
rect 66990 118030 70020 118053
rect 70180 118053 70203 119030
rect 73187 120030 73210 121037
rect 73370 121037 76400 121060
rect 73370 120030 73393 121037
rect 73187 119030 73393 120030
rect 73187 118053 73210 119030
rect 70180 118030 73210 118053
rect 73370 118053 73393 119030
rect 76377 120030 76400 121037
rect 76560 121037 79590 121060
rect 76560 120030 76583 121037
rect 76377 119030 76583 120030
rect 76377 118053 76400 119030
rect 73370 118030 76400 118053
rect 76560 118053 76583 119030
rect 79567 120030 79590 121037
rect 79750 121037 82780 121060
rect 79750 120030 79773 121037
rect 79567 119030 79773 120030
rect 79567 118053 79590 119030
rect 76560 118030 79590 118053
rect 79750 118053 79773 119030
rect 82757 120030 82780 121037
rect 82940 121037 85970 121060
rect 82940 120030 82963 121037
rect 82757 119030 82963 120030
rect 82757 118053 82780 119030
rect 79750 118030 82780 118053
rect 82940 118053 82963 119030
rect 85947 120030 85970 121037
rect 86130 121037 89160 121060
rect 86130 120030 86153 121037
rect 85947 119030 86153 120030
rect 85947 118053 85970 119030
rect 82940 118030 85970 118053
rect 86130 118053 86153 119030
rect 89137 120030 89160 121037
rect 89320 121037 92350 121060
rect 89320 120030 89343 121037
rect 89137 119030 89343 120030
rect 89137 118053 89160 119030
rect 86130 118030 89160 118053
rect 89320 118053 89343 119030
rect 92327 120030 92350 121037
rect 92510 121037 95540 121060
rect 92510 120030 92533 121037
rect 92327 119030 92533 120030
rect 92327 118053 92350 119030
rect 89320 118030 92350 118053
rect 92510 118053 92533 119030
rect 95517 120030 95540 121037
rect 95700 121037 98730 121060
rect 95700 120030 95723 121037
rect 95517 119030 95723 120030
rect 95517 118053 95540 119030
rect 92510 118030 95540 118053
rect 95700 118053 95723 119030
rect 98707 120030 98730 121037
rect 98890 121037 101920 121060
rect 98890 120030 98913 121037
rect 98707 119030 98913 120030
rect 98707 118053 98730 119030
rect 95700 118030 98730 118053
rect 98890 118053 98913 119030
rect 101897 120030 101920 121037
rect 102080 121037 105110 121060
rect 102080 120030 102103 121037
rect 101897 119030 102103 120030
rect 101897 118053 101920 119030
rect 98890 118030 101920 118053
rect 102080 118053 102103 119030
rect 105087 120030 105110 121037
rect 105270 121037 108300 121060
rect 105270 120030 105293 121037
rect 105087 119030 105293 120030
rect 105087 118053 105110 119030
rect 102080 118030 105110 118053
rect 105270 118053 105293 119030
rect 108277 120030 108300 121037
rect 108460 121037 111490 121060
rect 108460 120030 108483 121037
rect 108277 119030 108483 120030
rect 108277 118053 108300 119030
rect 105270 118030 108300 118053
rect 108460 118053 108483 119030
rect 111467 120030 111490 121037
rect 111650 121037 114680 121060
rect 111650 120030 111673 121037
rect 111467 119030 111673 120030
rect 111467 118053 111490 119030
rect 108460 118030 111490 118053
rect 111650 118053 111673 119030
rect 114657 120030 114680 121037
rect 114840 121037 117870 121060
rect 114840 120030 114863 121037
rect 114657 119030 114863 120030
rect 114657 118053 114680 119030
rect 111650 118030 114680 118053
rect 114840 118053 114863 119030
rect 117847 120030 117870 121037
rect 118030 121037 121060 121060
rect 118030 120030 118053 121037
rect 117847 119030 118053 120030
rect 117847 118053 117870 119030
rect 114840 118030 117870 118053
rect 118030 118053 118053 119030
rect 121037 120030 121060 121037
rect 121220 121037 124250 121060
rect 121220 120030 121243 121037
rect 121037 119030 121243 120030
rect 121037 118053 121060 119030
rect 118030 118030 121060 118053
rect 121220 118053 121243 119030
rect 124227 120030 124250 121037
rect 124410 121037 127440 121060
rect 124410 120030 124433 121037
rect 124227 119030 124433 120030
rect 124227 118053 124250 119030
rect 121220 118030 124250 118053
rect 124410 118053 124433 119030
rect 127417 120030 127440 121037
rect 127600 121037 130630 121060
rect 127600 120030 127623 121037
rect 127417 119030 127623 120030
rect 127417 118053 127440 119030
rect 124410 118030 127440 118053
rect 127600 118053 127623 119030
rect 130607 120030 130630 121037
rect 130790 121037 133820 121060
rect 130790 120030 130813 121037
rect 130607 119030 130813 120030
rect 130607 118053 130630 119030
rect 127600 118030 130630 118053
rect 130790 118053 130813 119030
rect 133797 120030 133820 121037
rect 133980 121037 137010 121060
rect 133980 120030 134003 121037
rect 133797 119030 134003 120030
rect 133797 118053 133820 119030
rect 130790 118030 133820 118053
rect 133980 118053 134003 119030
rect 136987 120030 137010 121037
rect 136987 119030 137170 120030
rect 136987 118053 137010 119030
rect 133980 118030 137010 118053
rect 1000 117870 2000 118030
rect 4190 117870 5190 118030
rect 7380 117870 8380 118030
rect 10570 117870 11570 118030
rect 13760 117870 14760 118030
rect 16950 117870 17950 118030
rect 20140 117870 21140 118030
rect 23330 117870 24330 118030
rect 26520 117870 27520 118030
rect 29710 117870 30710 118030
rect 32900 117870 33900 118030
rect 36090 117870 37090 118030
rect 39280 117870 40280 118030
rect 42470 117870 43470 118030
rect 45660 117870 46660 118030
rect 48850 117870 49850 118030
rect 52040 117870 53040 118030
rect 55230 117870 56230 118030
rect 58420 117870 59420 118030
rect 61610 117870 62610 118030
rect 64800 117870 65800 118030
rect 67990 117870 68990 118030
rect 71180 117870 72180 118030
rect 74370 117870 75370 118030
rect 77560 117870 78560 118030
rect 80750 117870 81750 118030
rect 83940 117870 84940 118030
rect 87130 117870 88130 118030
rect 90320 117870 91320 118030
rect 93510 117870 94510 118030
rect 96700 117870 97700 118030
rect 99890 117870 100890 118030
rect 103080 117870 104080 118030
rect 106270 117870 107270 118030
rect 109460 117870 110460 118030
rect 112650 117870 113650 118030
rect 115840 117870 116840 118030
rect 119030 117870 120030 118030
rect 122220 117870 123220 118030
rect 125410 117870 126410 118030
rect 128600 117870 129600 118030
rect 131790 117870 132790 118030
rect 134980 117870 135980 118030
rect 0 117847 3030 117870
rect 0 114863 23 117847
rect 3007 116840 3030 117847
rect 3190 117847 6220 117870
rect 3190 116840 3213 117847
rect 3007 115840 3213 116840
rect 3007 114863 3030 115840
rect 0 114840 3030 114863
rect 3190 114863 3213 115840
rect 6197 116840 6220 117847
rect 6380 117847 9410 117870
rect 6380 116840 6403 117847
rect 6197 115840 6403 116840
rect 6197 114863 6220 115840
rect 3190 114840 6220 114863
rect 6380 114863 6403 115840
rect 9387 116840 9410 117847
rect 9570 117847 12600 117870
rect 9570 116840 9593 117847
rect 9387 115840 9593 116840
rect 9387 114863 9410 115840
rect 6380 114840 9410 114863
rect 9570 114863 9593 115840
rect 12577 116840 12600 117847
rect 12760 117847 15790 117870
rect 12760 116840 12783 117847
rect 12577 115840 12783 116840
rect 12577 114863 12600 115840
rect 9570 114840 12600 114863
rect 12760 114863 12783 115840
rect 15767 116840 15790 117847
rect 15950 117847 18980 117870
rect 15950 116840 15973 117847
rect 15767 115840 15973 116840
rect 15767 114863 15790 115840
rect 12760 114840 15790 114863
rect 15950 114863 15973 115840
rect 18957 116840 18980 117847
rect 19140 117847 22170 117870
rect 19140 116840 19163 117847
rect 18957 115840 19163 116840
rect 18957 114863 18980 115840
rect 15950 114840 18980 114863
rect 19140 114863 19163 115840
rect 22147 116840 22170 117847
rect 22330 117847 25360 117870
rect 22330 116840 22353 117847
rect 22147 115840 22353 116840
rect 22147 114863 22170 115840
rect 19140 114840 22170 114863
rect 22330 114863 22353 115840
rect 25337 116840 25360 117847
rect 25520 117847 28550 117870
rect 25520 116840 25543 117847
rect 25337 115840 25543 116840
rect 25337 114863 25360 115840
rect 22330 114840 25360 114863
rect 25520 114863 25543 115840
rect 28527 116840 28550 117847
rect 28710 117847 31740 117870
rect 28710 116840 28733 117847
rect 28527 115840 28733 116840
rect 28527 114863 28550 115840
rect 25520 114840 28550 114863
rect 28710 114863 28733 115840
rect 31717 116840 31740 117847
rect 31900 117847 34930 117870
rect 31900 116840 31923 117847
rect 31717 115840 31923 116840
rect 31717 114863 31740 115840
rect 28710 114840 31740 114863
rect 31900 114863 31923 115840
rect 34907 116840 34930 117847
rect 35090 117847 38120 117870
rect 35090 116840 35113 117847
rect 34907 115840 35113 116840
rect 34907 114863 34930 115840
rect 31900 114840 34930 114863
rect 35090 114863 35113 115840
rect 38097 116840 38120 117847
rect 38280 117847 41310 117870
rect 38280 116840 38303 117847
rect 38097 115840 38303 116840
rect 38097 114863 38120 115840
rect 35090 114840 38120 114863
rect 38280 114863 38303 115840
rect 41287 116840 41310 117847
rect 41470 117847 44500 117870
rect 41470 116840 41493 117847
rect 41287 115840 41493 116840
rect 41287 114863 41310 115840
rect 38280 114840 41310 114863
rect 41470 114863 41493 115840
rect 44477 116840 44500 117847
rect 44660 117847 47690 117870
rect 44660 116840 44683 117847
rect 44477 115840 44683 116840
rect 44477 114863 44500 115840
rect 41470 114840 44500 114863
rect 44660 114863 44683 115840
rect 47667 116840 47690 117847
rect 47850 117847 50880 117870
rect 47850 116840 47873 117847
rect 47667 115840 47873 116840
rect 47667 114863 47690 115840
rect 44660 114840 47690 114863
rect 47850 114863 47873 115840
rect 50857 116840 50880 117847
rect 51040 117847 54070 117870
rect 51040 116840 51063 117847
rect 50857 115840 51063 116840
rect 50857 114863 50880 115840
rect 47850 114840 50880 114863
rect 51040 114863 51063 115840
rect 54047 116840 54070 117847
rect 54230 117847 57260 117870
rect 54230 116840 54253 117847
rect 54047 115840 54253 116840
rect 54047 114863 54070 115840
rect 51040 114840 54070 114863
rect 54230 114863 54253 115840
rect 57237 116840 57260 117847
rect 57420 117847 60450 117870
rect 57420 116840 57443 117847
rect 57237 115840 57443 116840
rect 57237 114863 57260 115840
rect 54230 114840 57260 114863
rect 57420 114863 57443 115840
rect 60427 116840 60450 117847
rect 60610 117847 63640 117870
rect 60610 116840 60633 117847
rect 60427 115840 60633 116840
rect 60427 114863 60450 115840
rect 57420 114840 60450 114863
rect 60610 114863 60633 115840
rect 63617 116840 63640 117847
rect 63800 117847 66830 117870
rect 63800 116840 63823 117847
rect 63617 115840 63823 116840
rect 63617 114863 63640 115840
rect 60610 114840 63640 114863
rect 63800 114863 63823 115840
rect 66807 116840 66830 117847
rect 66990 117847 70020 117870
rect 66990 116840 67013 117847
rect 66807 115840 67013 116840
rect 66807 114863 66830 115840
rect 63800 114840 66830 114863
rect 66990 114863 67013 115840
rect 69997 116840 70020 117847
rect 70180 117847 73210 117870
rect 70180 116840 70203 117847
rect 69997 115840 70203 116840
rect 69997 114863 70020 115840
rect 66990 114840 70020 114863
rect 70180 114863 70203 115840
rect 73187 116840 73210 117847
rect 73370 117847 76400 117870
rect 73370 116840 73393 117847
rect 73187 115840 73393 116840
rect 73187 114863 73210 115840
rect 70180 114840 73210 114863
rect 73370 114863 73393 115840
rect 76377 116840 76400 117847
rect 76560 117847 79590 117870
rect 76560 116840 76583 117847
rect 76377 115840 76583 116840
rect 76377 114863 76400 115840
rect 73370 114840 76400 114863
rect 76560 114863 76583 115840
rect 79567 116840 79590 117847
rect 79750 117847 82780 117870
rect 79750 116840 79773 117847
rect 79567 115840 79773 116840
rect 79567 114863 79590 115840
rect 76560 114840 79590 114863
rect 79750 114863 79773 115840
rect 82757 116840 82780 117847
rect 82940 117847 85970 117870
rect 82940 116840 82963 117847
rect 82757 115840 82963 116840
rect 82757 114863 82780 115840
rect 79750 114840 82780 114863
rect 82940 114863 82963 115840
rect 85947 116840 85970 117847
rect 86130 117847 89160 117870
rect 86130 116840 86153 117847
rect 85947 115840 86153 116840
rect 85947 114863 85970 115840
rect 82940 114840 85970 114863
rect 86130 114863 86153 115840
rect 89137 116840 89160 117847
rect 89320 117847 92350 117870
rect 89320 116840 89343 117847
rect 89137 115840 89343 116840
rect 89137 114863 89160 115840
rect 86130 114840 89160 114863
rect 89320 114863 89343 115840
rect 92327 116840 92350 117847
rect 92510 117847 95540 117870
rect 92510 116840 92533 117847
rect 92327 115840 92533 116840
rect 92327 114863 92350 115840
rect 89320 114840 92350 114863
rect 92510 114863 92533 115840
rect 95517 116840 95540 117847
rect 95700 117847 98730 117870
rect 95700 116840 95723 117847
rect 95517 115840 95723 116840
rect 95517 114863 95540 115840
rect 92510 114840 95540 114863
rect 95700 114863 95723 115840
rect 98707 116840 98730 117847
rect 98890 117847 101920 117870
rect 98890 116840 98913 117847
rect 98707 115840 98913 116840
rect 98707 114863 98730 115840
rect 95700 114840 98730 114863
rect 98890 114863 98913 115840
rect 101897 116840 101920 117847
rect 102080 117847 105110 117870
rect 102080 116840 102103 117847
rect 101897 115840 102103 116840
rect 101897 114863 101920 115840
rect 98890 114840 101920 114863
rect 102080 114863 102103 115840
rect 105087 116840 105110 117847
rect 105270 117847 108300 117870
rect 105270 116840 105293 117847
rect 105087 115840 105293 116840
rect 105087 114863 105110 115840
rect 102080 114840 105110 114863
rect 105270 114863 105293 115840
rect 108277 116840 108300 117847
rect 108460 117847 111490 117870
rect 108460 116840 108483 117847
rect 108277 115840 108483 116840
rect 108277 114863 108300 115840
rect 105270 114840 108300 114863
rect 108460 114863 108483 115840
rect 111467 116840 111490 117847
rect 111650 117847 114680 117870
rect 111650 116840 111673 117847
rect 111467 115840 111673 116840
rect 111467 114863 111490 115840
rect 108460 114840 111490 114863
rect 111650 114863 111673 115840
rect 114657 116840 114680 117847
rect 114840 117847 117870 117870
rect 114840 116840 114863 117847
rect 114657 115840 114863 116840
rect 114657 114863 114680 115840
rect 111650 114840 114680 114863
rect 114840 114863 114863 115840
rect 117847 116840 117870 117847
rect 118030 117847 121060 117870
rect 118030 116840 118053 117847
rect 117847 115840 118053 116840
rect 117847 114863 117870 115840
rect 114840 114840 117870 114863
rect 118030 114863 118053 115840
rect 121037 116840 121060 117847
rect 121220 117847 124250 117870
rect 121220 116840 121243 117847
rect 121037 115840 121243 116840
rect 121037 114863 121060 115840
rect 118030 114840 121060 114863
rect 121220 114863 121243 115840
rect 124227 116840 124250 117847
rect 124410 117847 127440 117870
rect 124410 116840 124433 117847
rect 124227 115840 124433 116840
rect 124227 114863 124250 115840
rect 121220 114840 124250 114863
rect 124410 114863 124433 115840
rect 127417 116840 127440 117847
rect 127600 117847 130630 117870
rect 127600 116840 127623 117847
rect 127417 115840 127623 116840
rect 127417 114863 127440 115840
rect 124410 114840 127440 114863
rect 127600 114863 127623 115840
rect 130607 116840 130630 117847
rect 130790 117847 133820 117870
rect 130790 116840 130813 117847
rect 130607 115840 130813 116840
rect 130607 114863 130630 115840
rect 127600 114840 130630 114863
rect 130790 114863 130813 115840
rect 133797 116840 133820 117847
rect 133980 117847 137010 117870
rect 133980 116840 134003 117847
rect 133797 115840 134003 116840
rect 133797 114863 133820 115840
rect 130790 114840 133820 114863
rect 133980 114863 134003 115840
rect 136987 116840 137010 117847
rect 136987 115840 137170 116840
rect 136987 114863 137010 115840
rect 133980 114840 137010 114863
rect 1000 114680 2000 114840
rect 4190 114680 5190 114840
rect 7380 114680 8380 114840
rect 10570 114680 11570 114840
rect 13760 114680 14760 114840
rect 16950 114680 17950 114840
rect 20140 114680 21140 114840
rect 23330 114680 24330 114840
rect 26520 114680 27520 114840
rect 29710 114680 30710 114840
rect 32900 114680 33900 114840
rect 36090 114680 37090 114840
rect 39280 114680 40280 114840
rect 42470 114680 43470 114840
rect 45660 114680 46660 114840
rect 48850 114680 49850 114840
rect 52040 114680 53040 114840
rect 55230 114680 56230 114840
rect 58420 114680 59420 114840
rect 61610 114680 62610 114840
rect 64800 114680 65800 114840
rect 67990 114680 68990 114840
rect 71180 114680 72180 114840
rect 74370 114680 75370 114840
rect 77560 114680 78560 114840
rect 80750 114680 81750 114840
rect 83940 114680 84940 114840
rect 87130 114680 88130 114840
rect 90320 114680 91320 114840
rect 93510 114680 94510 114840
rect 96700 114680 97700 114840
rect 99890 114680 100890 114840
rect 103080 114680 104080 114840
rect 106270 114680 107270 114840
rect 109460 114680 110460 114840
rect 112650 114680 113650 114840
rect 115840 114680 116840 114840
rect 119030 114680 120030 114840
rect 122220 114680 123220 114840
rect 125410 114680 126410 114840
rect 128600 114680 129600 114840
rect 131790 114680 132790 114840
rect 134980 114680 135980 114840
rect 0 114657 3030 114680
rect 0 111673 23 114657
rect 3007 113650 3030 114657
rect 3190 114657 6220 114680
rect 3190 113650 3213 114657
rect 3007 112650 3213 113650
rect 3007 111673 3030 112650
rect 0 111650 3030 111673
rect 3190 111673 3213 112650
rect 6197 113650 6220 114657
rect 6380 114657 9410 114680
rect 6380 113650 6403 114657
rect 6197 112650 6403 113650
rect 6197 111673 6220 112650
rect 3190 111650 6220 111673
rect 6380 111673 6403 112650
rect 9387 113650 9410 114657
rect 9570 114657 12600 114680
rect 9570 113650 9593 114657
rect 9387 112650 9593 113650
rect 9387 111673 9410 112650
rect 6380 111650 9410 111673
rect 9570 111673 9593 112650
rect 12577 113650 12600 114657
rect 12760 114657 15790 114680
rect 12760 113650 12783 114657
rect 12577 112650 12783 113650
rect 12577 111673 12600 112650
rect 9570 111650 12600 111673
rect 12760 111673 12783 112650
rect 15767 113650 15790 114657
rect 15950 114657 18980 114680
rect 15950 113650 15973 114657
rect 15767 112650 15973 113650
rect 15767 111673 15790 112650
rect 12760 111650 15790 111673
rect 15950 111673 15973 112650
rect 18957 113650 18980 114657
rect 19140 114657 22170 114680
rect 19140 113650 19163 114657
rect 18957 112650 19163 113650
rect 18957 111673 18980 112650
rect 15950 111650 18980 111673
rect 19140 111673 19163 112650
rect 22147 113650 22170 114657
rect 22330 114657 25360 114680
rect 22330 113650 22353 114657
rect 22147 112650 22353 113650
rect 22147 111673 22170 112650
rect 19140 111650 22170 111673
rect 22330 111673 22353 112650
rect 25337 113650 25360 114657
rect 25520 114657 28550 114680
rect 25520 113650 25543 114657
rect 25337 112650 25543 113650
rect 25337 111673 25360 112650
rect 22330 111650 25360 111673
rect 25520 111673 25543 112650
rect 28527 113650 28550 114657
rect 28710 114657 31740 114680
rect 28710 113650 28733 114657
rect 28527 112650 28733 113650
rect 28527 111673 28550 112650
rect 25520 111650 28550 111673
rect 28710 111673 28733 112650
rect 31717 113650 31740 114657
rect 31900 114657 34930 114680
rect 31900 113650 31923 114657
rect 31717 112650 31923 113650
rect 31717 111673 31740 112650
rect 28710 111650 31740 111673
rect 31900 111673 31923 112650
rect 34907 113650 34930 114657
rect 35090 114657 38120 114680
rect 35090 113650 35113 114657
rect 34907 112650 35113 113650
rect 34907 111673 34930 112650
rect 31900 111650 34930 111673
rect 35090 111673 35113 112650
rect 38097 113650 38120 114657
rect 38280 114657 41310 114680
rect 38280 113650 38303 114657
rect 38097 112650 38303 113650
rect 38097 111673 38120 112650
rect 35090 111650 38120 111673
rect 38280 111673 38303 112650
rect 41287 113650 41310 114657
rect 41470 114657 44500 114680
rect 41470 113650 41493 114657
rect 41287 112650 41493 113650
rect 41287 111673 41310 112650
rect 38280 111650 41310 111673
rect 41470 111673 41493 112650
rect 44477 113650 44500 114657
rect 44660 114657 47690 114680
rect 44660 113650 44683 114657
rect 44477 112650 44683 113650
rect 44477 111673 44500 112650
rect 41470 111650 44500 111673
rect 44660 111673 44683 112650
rect 47667 113650 47690 114657
rect 47850 114657 50880 114680
rect 47850 113650 47873 114657
rect 47667 112650 47873 113650
rect 47667 111673 47690 112650
rect 44660 111650 47690 111673
rect 47850 111673 47873 112650
rect 50857 113650 50880 114657
rect 51040 114657 54070 114680
rect 51040 113650 51063 114657
rect 50857 112650 51063 113650
rect 50857 111673 50880 112650
rect 47850 111650 50880 111673
rect 51040 111673 51063 112650
rect 54047 113650 54070 114657
rect 54230 114657 57260 114680
rect 54230 113650 54253 114657
rect 54047 112650 54253 113650
rect 54047 111673 54070 112650
rect 51040 111650 54070 111673
rect 54230 111673 54253 112650
rect 57237 113650 57260 114657
rect 57420 114657 60450 114680
rect 57420 113650 57443 114657
rect 57237 112650 57443 113650
rect 57237 111673 57260 112650
rect 54230 111650 57260 111673
rect 57420 111673 57443 112650
rect 60427 113650 60450 114657
rect 60610 114657 63640 114680
rect 60610 113650 60633 114657
rect 60427 112650 60633 113650
rect 60427 111673 60450 112650
rect 57420 111650 60450 111673
rect 60610 111673 60633 112650
rect 63617 113650 63640 114657
rect 63800 114657 66830 114680
rect 63800 113650 63823 114657
rect 63617 112650 63823 113650
rect 63617 111673 63640 112650
rect 60610 111650 63640 111673
rect 63800 111673 63823 112650
rect 66807 113650 66830 114657
rect 66990 114657 70020 114680
rect 66990 113650 67013 114657
rect 66807 112650 67013 113650
rect 66807 111673 66830 112650
rect 63800 111650 66830 111673
rect 66990 111673 67013 112650
rect 69997 113650 70020 114657
rect 70180 114657 73210 114680
rect 70180 113650 70203 114657
rect 69997 112650 70203 113650
rect 69997 111673 70020 112650
rect 66990 111650 70020 111673
rect 70180 111673 70203 112650
rect 73187 113650 73210 114657
rect 73370 114657 76400 114680
rect 73370 113650 73393 114657
rect 73187 112650 73393 113650
rect 73187 111673 73210 112650
rect 70180 111650 73210 111673
rect 73370 111673 73393 112650
rect 76377 113650 76400 114657
rect 76560 114657 79590 114680
rect 76560 113650 76583 114657
rect 76377 112650 76583 113650
rect 76377 111673 76400 112650
rect 73370 111650 76400 111673
rect 76560 111673 76583 112650
rect 79567 113650 79590 114657
rect 79750 114657 82780 114680
rect 79750 113650 79773 114657
rect 79567 112650 79773 113650
rect 79567 111673 79590 112650
rect 76560 111650 79590 111673
rect 79750 111673 79773 112650
rect 82757 113650 82780 114657
rect 82940 114657 85970 114680
rect 82940 113650 82963 114657
rect 82757 112650 82963 113650
rect 82757 111673 82780 112650
rect 79750 111650 82780 111673
rect 82940 111673 82963 112650
rect 85947 113650 85970 114657
rect 86130 114657 89160 114680
rect 86130 113650 86153 114657
rect 85947 112650 86153 113650
rect 85947 111673 85970 112650
rect 82940 111650 85970 111673
rect 86130 111673 86153 112650
rect 89137 113650 89160 114657
rect 89320 114657 92350 114680
rect 89320 113650 89343 114657
rect 89137 112650 89343 113650
rect 89137 111673 89160 112650
rect 86130 111650 89160 111673
rect 89320 111673 89343 112650
rect 92327 113650 92350 114657
rect 92510 114657 95540 114680
rect 92510 113650 92533 114657
rect 92327 112650 92533 113650
rect 92327 111673 92350 112650
rect 89320 111650 92350 111673
rect 92510 111673 92533 112650
rect 95517 113650 95540 114657
rect 95700 114657 98730 114680
rect 95700 113650 95723 114657
rect 95517 112650 95723 113650
rect 95517 111673 95540 112650
rect 92510 111650 95540 111673
rect 95700 111673 95723 112650
rect 98707 113650 98730 114657
rect 98890 114657 101920 114680
rect 98890 113650 98913 114657
rect 98707 112650 98913 113650
rect 98707 111673 98730 112650
rect 95700 111650 98730 111673
rect 98890 111673 98913 112650
rect 101897 113650 101920 114657
rect 102080 114657 105110 114680
rect 102080 113650 102103 114657
rect 101897 112650 102103 113650
rect 101897 111673 101920 112650
rect 98890 111650 101920 111673
rect 102080 111673 102103 112650
rect 105087 113650 105110 114657
rect 105270 114657 108300 114680
rect 105270 113650 105293 114657
rect 105087 112650 105293 113650
rect 105087 111673 105110 112650
rect 102080 111650 105110 111673
rect 105270 111673 105293 112650
rect 108277 113650 108300 114657
rect 108460 114657 111490 114680
rect 108460 113650 108483 114657
rect 108277 112650 108483 113650
rect 108277 111673 108300 112650
rect 105270 111650 108300 111673
rect 108460 111673 108483 112650
rect 111467 113650 111490 114657
rect 111650 114657 114680 114680
rect 111650 113650 111673 114657
rect 111467 112650 111673 113650
rect 111467 111673 111490 112650
rect 108460 111650 111490 111673
rect 111650 111673 111673 112650
rect 114657 113650 114680 114657
rect 114840 114657 117870 114680
rect 114840 113650 114863 114657
rect 114657 112650 114863 113650
rect 114657 111673 114680 112650
rect 111650 111650 114680 111673
rect 114840 111673 114863 112650
rect 117847 113650 117870 114657
rect 118030 114657 121060 114680
rect 118030 113650 118053 114657
rect 117847 112650 118053 113650
rect 117847 111673 117870 112650
rect 114840 111650 117870 111673
rect 118030 111673 118053 112650
rect 121037 113650 121060 114657
rect 121220 114657 124250 114680
rect 121220 113650 121243 114657
rect 121037 112650 121243 113650
rect 121037 111673 121060 112650
rect 118030 111650 121060 111673
rect 121220 111673 121243 112650
rect 124227 113650 124250 114657
rect 124410 114657 127440 114680
rect 124410 113650 124433 114657
rect 124227 112650 124433 113650
rect 124227 111673 124250 112650
rect 121220 111650 124250 111673
rect 124410 111673 124433 112650
rect 127417 113650 127440 114657
rect 127600 114657 130630 114680
rect 127600 113650 127623 114657
rect 127417 112650 127623 113650
rect 127417 111673 127440 112650
rect 124410 111650 127440 111673
rect 127600 111673 127623 112650
rect 130607 113650 130630 114657
rect 130790 114657 133820 114680
rect 130790 113650 130813 114657
rect 130607 112650 130813 113650
rect 130607 111673 130630 112650
rect 127600 111650 130630 111673
rect 130790 111673 130813 112650
rect 133797 113650 133820 114657
rect 133980 114657 137010 114680
rect 133980 113650 134003 114657
rect 133797 112650 134003 113650
rect 133797 111673 133820 112650
rect 130790 111650 133820 111673
rect 133980 111673 134003 112650
rect 136987 113650 137010 114657
rect 136987 112650 137170 113650
rect 136987 111673 137010 112650
rect 133980 111650 137010 111673
rect 1000 111490 2000 111650
rect 4190 111490 5190 111650
rect 7380 111490 8380 111650
rect 10570 111490 11570 111650
rect 13760 111490 14760 111650
rect 16950 111490 17950 111650
rect 20140 111490 21140 111650
rect 23330 111490 24330 111650
rect 26520 111490 27520 111650
rect 29710 111490 30710 111650
rect 32900 111490 33900 111650
rect 36090 111490 37090 111650
rect 39280 111490 40280 111650
rect 42470 111490 43470 111650
rect 45660 111490 46660 111650
rect 48850 111490 49850 111650
rect 52040 111490 53040 111650
rect 55230 111490 56230 111650
rect 58420 111490 59420 111650
rect 61610 111490 62610 111650
rect 64800 111490 65800 111650
rect 67990 111490 68990 111650
rect 71180 111490 72180 111650
rect 74370 111490 75370 111650
rect 77560 111490 78560 111650
rect 80750 111490 81750 111650
rect 83940 111490 84940 111650
rect 87130 111490 88130 111650
rect 90320 111490 91320 111650
rect 93510 111490 94510 111650
rect 96700 111490 97700 111650
rect 99890 111490 100890 111650
rect 103080 111490 104080 111650
rect 106270 111490 107270 111650
rect 109460 111490 110460 111650
rect 112650 111490 113650 111650
rect 115840 111490 116840 111650
rect 119030 111490 120030 111650
rect 122220 111490 123220 111650
rect 125410 111490 126410 111650
rect 128600 111490 129600 111650
rect 131790 111490 132790 111650
rect 134980 111490 135980 111650
rect 0 111467 3030 111490
rect 0 108483 23 111467
rect 3007 110460 3030 111467
rect 3190 111467 6220 111490
rect 3190 110460 3213 111467
rect 3007 109460 3213 110460
rect 3007 108483 3030 109460
rect 0 108460 3030 108483
rect 3190 108483 3213 109460
rect 6197 110460 6220 111467
rect 6380 111467 9410 111490
rect 6380 110460 6403 111467
rect 6197 109460 6403 110460
rect 6197 108483 6220 109460
rect 3190 108460 6220 108483
rect 6380 108483 6403 109460
rect 9387 110460 9410 111467
rect 9570 111467 12600 111490
rect 9570 110460 9593 111467
rect 9387 109460 9593 110460
rect 9387 108483 9410 109460
rect 6380 108460 9410 108483
rect 9570 108483 9593 109460
rect 12577 110460 12600 111467
rect 12760 111467 15790 111490
rect 12760 110460 12783 111467
rect 12577 109460 12783 110460
rect 12577 108483 12600 109460
rect 9570 108460 12600 108483
rect 12760 108483 12783 109460
rect 15767 110460 15790 111467
rect 15950 111467 18980 111490
rect 15950 110460 15973 111467
rect 15767 109460 15973 110460
rect 15767 108483 15790 109460
rect 12760 108460 15790 108483
rect 15950 108483 15973 109460
rect 18957 110460 18980 111467
rect 19140 111467 22170 111490
rect 19140 110460 19163 111467
rect 18957 109460 19163 110460
rect 18957 108483 18980 109460
rect 15950 108460 18980 108483
rect 19140 108483 19163 109460
rect 22147 110460 22170 111467
rect 22330 111467 25360 111490
rect 22330 110460 22353 111467
rect 22147 109460 22353 110460
rect 22147 108483 22170 109460
rect 19140 108460 22170 108483
rect 22330 108483 22353 109460
rect 25337 110460 25360 111467
rect 25520 111467 28550 111490
rect 25520 110460 25543 111467
rect 25337 109460 25543 110460
rect 25337 108483 25360 109460
rect 22330 108460 25360 108483
rect 25520 108483 25543 109460
rect 28527 110460 28550 111467
rect 28710 111467 31740 111490
rect 28710 110460 28733 111467
rect 28527 109460 28733 110460
rect 28527 108483 28550 109460
rect 25520 108460 28550 108483
rect 28710 108483 28733 109460
rect 31717 110460 31740 111467
rect 31900 111467 34930 111490
rect 31900 110460 31923 111467
rect 31717 109460 31923 110460
rect 31717 108483 31740 109460
rect 28710 108460 31740 108483
rect 31900 108483 31923 109460
rect 34907 110460 34930 111467
rect 35090 111467 38120 111490
rect 35090 110460 35113 111467
rect 34907 109460 35113 110460
rect 34907 108483 34930 109460
rect 31900 108460 34930 108483
rect 35090 108483 35113 109460
rect 38097 110460 38120 111467
rect 38280 111467 41310 111490
rect 38280 110460 38303 111467
rect 38097 109460 38303 110460
rect 38097 108483 38120 109460
rect 35090 108460 38120 108483
rect 38280 108483 38303 109460
rect 41287 110460 41310 111467
rect 41470 111467 44500 111490
rect 41470 110460 41493 111467
rect 41287 109460 41493 110460
rect 41287 108483 41310 109460
rect 38280 108460 41310 108483
rect 41470 108483 41493 109460
rect 44477 110460 44500 111467
rect 44660 111467 47690 111490
rect 44660 110460 44683 111467
rect 44477 109460 44683 110460
rect 44477 108483 44500 109460
rect 41470 108460 44500 108483
rect 44660 108483 44683 109460
rect 47667 110460 47690 111467
rect 47850 111467 50880 111490
rect 47850 110460 47873 111467
rect 47667 109460 47873 110460
rect 47667 108483 47690 109460
rect 44660 108460 47690 108483
rect 47850 108483 47873 109460
rect 50857 110460 50880 111467
rect 51040 111467 54070 111490
rect 51040 110460 51063 111467
rect 50857 109460 51063 110460
rect 50857 108483 50880 109460
rect 47850 108460 50880 108483
rect 51040 108483 51063 109460
rect 54047 110460 54070 111467
rect 54230 111467 57260 111490
rect 54230 110460 54253 111467
rect 54047 109460 54253 110460
rect 54047 108483 54070 109460
rect 51040 108460 54070 108483
rect 54230 108483 54253 109460
rect 57237 110460 57260 111467
rect 57420 111467 60450 111490
rect 57420 110460 57443 111467
rect 57237 109460 57443 110460
rect 57237 108483 57260 109460
rect 54230 108460 57260 108483
rect 57420 108483 57443 109460
rect 60427 110460 60450 111467
rect 60610 111467 63640 111490
rect 60610 110460 60633 111467
rect 60427 109460 60633 110460
rect 60427 108483 60450 109460
rect 57420 108460 60450 108483
rect 60610 108483 60633 109460
rect 63617 110460 63640 111467
rect 63800 111467 66830 111490
rect 63800 110460 63823 111467
rect 63617 109460 63823 110460
rect 63617 108483 63640 109460
rect 60610 108460 63640 108483
rect 63800 108483 63823 109460
rect 66807 110460 66830 111467
rect 66990 111467 70020 111490
rect 66990 110460 67013 111467
rect 66807 109460 67013 110460
rect 66807 108483 66830 109460
rect 63800 108460 66830 108483
rect 66990 108483 67013 109460
rect 69997 110460 70020 111467
rect 70180 111467 73210 111490
rect 70180 110460 70203 111467
rect 69997 109460 70203 110460
rect 69997 108483 70020 109460
rect 66990 108460 70020 108483
rect 70180 108483 70203 109460
rect 73187 110460 73210 111467
rect 73370 111467 76400 111490
rect 73370 110460 73393 111467
rect 73187 109460 73393 110460
rect 73187 108483 73210 109460
rect 70180 108460 73210 108483
rect 73370 108483 73393 109460
rect 76377 110460 76400 111467
rect 76560 111467 79590 111490
rect 76560 110460 76583 111467
rect 76377 109460 76583 110460
rect 76377 108483 76400 109460
rect 73370 108460 76400 108483
rect 76560 108483 76583 109460
rect 79567 110460 79590 111467
rect 79750 111467 82780 111490
rect 79750 110460 79773 111467
rect 79567 109460 79773 110460
rect 79567 108483 79590 109460
rect 76560 108460 79590 108483
rect 79750 108483 79773 109460
rect 82757 110460 82780 111467
rect 82940 111467 85970 111490
rect 82940 110460 82963 111467
rect 82757 109460 82963 110460
rect 82757 108483 82780 109460
rect 79750 108460 82780 108483
rect 82940 108483 82963 109460
rect 85947 110460 85970 111467
rect 86130 111467 89160 111490
rect 86130 110460 86153 111467
rect 85947 109460 86153 110460
rect 85947 108483 85970 109460
rect 82940 108460 85970 108483
rect 86130 108483 86153 109460
rect 89137 110460 89160 111467
rect 89320 111467 92350 111490
rect 89320 110460 89343 111467
rect 89137 109460 89343 110460
rect 89137 108483 89160 109460
rect 86130 108460 89160 108483
rect 89320 108483 89343 109460
rect 92327 110460 92350 111467
rect 92510 111467 95540 111490
rect 92510 110460 92533 111467
rect 92327 109460 92533 110460
rect 92327 108483 92350 109460
rect 89320 108460 92350 108483
rect 92510 108483 92533 109460
rect 95517 110460 95540 111467
rect 95700 111467 98730 111490
rect 95700 110460 95723 111467
rect 95517 109460 95723 110460
rect 95517 108483 95540 109460
rect 92510 108460 95540 108483
rect 95700 108483 95723 109460
rect 98707 110460 98730 111467
rect 98890 111467 101920 111490
rect 98890 110460 98913 111467
rect 98707 109460 98913 110460
rect 98707 108483 98730 109460
rect 95700 108460 98730 108483
rect 98890 108483 98913 109460
rect 101897 110460 101920 111467
rect 102080 111467 105110 111490
rect 102080 110460 102103 111467
rect 101897 109460 102103 110460
rect 101897 108483 101920 109460
rect 98890 108460 101920 108483
rect 102080 108483 102103 109460
rect 105087 110460 105110 111467
rect 105270 111467 108300 111490
rect 105270 110460 105293 111467
rect 105087 109460 105293 110460
rect 105087 108483 105110 109460
rect 102080 108460 105110 108483
rect 105270 108483 105293 109460
rect 108277 110460 108300 111467
rect 108460 111467 111490 111490
rect 108460 110460 108483 111467
rect 108277 109460 108483 110460
rect 108277 108483 108300 109460
rect 105270 108460 108300 108483
rect 108460 108483 108483 109460
rect 111467 110460 111490 111467
rect 111650 111467 114680 111490
rect 111650 110460 111673 111467
rect 111467 109460 111673 110460
rect 111467 108483 111490 109460
rect 108460 108460 111490 108483
rect 111650 108483 111673 109460
rect 114657 110460 114680 111467
rect 114840 111467 117870 111490
rect 114840 110460 114863 111467
rect 114657 109460 114863 110460
rect 114657 108483 114680 109460
rect 111650 108460 114680 108483
rect 114840 108483 114863 109460
rect 117847 110460 117870 111467
rect 118030 111467 121060 111490
rect 118030 110460 118053 111467
rect 117847 109460 118053 110460
rect 117847 108483 117870 109460
rect 114840 108460 117870 108483
rect 118030 108483 118053 109460
rect 121037 110460 121060 111467
rect 121220 111467 124250 111490
rect 121220 110460 121243 111467
rect 121037 109460 121243 110460
rect 121037 108483 121060 109460
rect 118030 108460 121060 108483
rect 121220 108483 121243 109460
rect 124227 110460 124250 111467
rect 124410 111467 127440 111490
rect 124410 110460 124433 111467
rect 124227 109460 124433 110460
rect 124227 108483 124250 109460
rect 121220 108460 124250 108483
rect 124410 108483 124433 109460
rect 127417 110460 127440 111467
rect 127600 111467 130630 111490
rect 127600 110460 127623 111467
rect 127417 109460 127623 110460
rect 127417 108483 127440 109460
rect 124410 108460 127440 108483
rect 127600 108483 127623 109460
rect 130607 110460 130630 111467
rect 130790 111467 133820 111490
rect 130790 110460 130813 111467
rect 130607 109460 130813 110460
rect 130607 108483 130630 109460
rect 127600 108460 130630 108483
rect 130790 108483 130813 109460
rect 133797 110460 133820 111467
rect 133980 111467 137010 111490
rect 133980 110460 134003 111467
rect 133797 109460 134003 110460
rect 133797 108483 133820 109460
rect 130790 108460 133820 108483
rect 133980 108483 134003 109460
rect 136987 110460 137010 111467
rect 136987 109460 137170 110460
rect 136987 108483 137010 109460
rect 133980 108460 137010 108483
rect 1000 108300 2000 108460
rect 4190 108300 5190 108460
rect 7380 108300 8380 108460
rect 10570 108300 11570 108460
rect 13760 108300 14760 108460
rect 16950 108300 17950 108460
rect 20140 108300 21140 108460
rect 23330 108300 24330 108460
rect 26520 108300 27520 108460
rect 29710 108300 30710 108460
rect 32900 108300 33900 108460
rect 36090 108300 37090 108460
rect 39280 108300 40280 108460
rect 42470 108300 43470 108460
rect 45660 108300 46660 108460
rect 48850 108300 49850 108460
rect 52040 108300 53040 108460
rect 55230 108300 56230 108460
rect 58420 108300 59420 108460
rect 61610 108300 62610 108460
rect 64800 108300 65800 108460
rect 67990 108300 68990 108460
rect 71180 108300 72180 108460
rect 74370 108300 75370 108460
rect 77560 108300 78560 108460
rect 80750 108300 81750 108460
rect 83940 108300 84940 108460
rect 87130 108300 88130 108460
rect 90320 108300 91320 108460
rect 93510 108300 94510 108460
rect 96700 108300 97700 108460
rect 99890 108300 100890 108460
rect 103080 108300 104080 108460
rect 106270 108300 107270 108460
rect 109460 108300 110460 108460
rect 112650 108300 113650 108460
rect 115840 108300 116840 108460
rect 119030 108300 120030 108460
rect 122220 108300 123220 108460
rect 125410 108300 126410 108460
rect 128600 108300 129600 108460
rect 131790 108300 132790 108460
rect 134980 108300 135980 108460
rect 0 108277 3030 108300
rect 0 105293 23 108277
rect 3007 107270 3030 108277
rect 3190 108277 6220 108300
rect 3190 107270 3213 108277
rect 3007 106270 3213 107270
rect 3007 105293 3030 106270
rect 0 105270 3030 105293
rect 3190 105293 3213 106270
rect 6197 107270 6220 108277
rect 6380 108277 9410 108300
rect 6380 107270 6403 108277
rect 6197 106270 6403 107270
rect 6197 105293 6220 106270
rect 3190 105270 6220 105293
rect 6380 105293 6403 106270
rect 9387 107270 9410 108277
rect 9570 108277 12600 108300
rect 9570 107270 9593 108277
rect 9387 106270 9593 107270
rect 9387 105293 9410 106270
rect 6380 105270 9410 105293
rect 9570 105293 9593 106270
rect 12577 107270 12600 108277
rect 12760 108277 15790 108300
rect 12760 107270 12783 108277
rect 12577 106270 12783 107270
rect 12577 105293 12600 106270
rect 9570 105270 12600 105293
rect 12760 105293 12783 106270
rect 15767 107270 15790 108277
rect 15950 108277 18980 108300
rect 15950 107270 15973 108277
rect 15767 106270 15973 107270
rect 15767 105293 15790 106270
rect 12760 105270 15790 105293
rect 15950 105293 15973 106270
rect 18957 107270 18980 108277
rect 19140 108277 22170 108300
rect 19140 107270 19163 108277
rect 18957 106270 19163 107270
rect 18957 105293 18980 106270
rect 15950 105270 18980 105293
rect 19140 105293 19163 106270
rect 22147 107270 22170 108277
rect 22330 108277 25360 108300
rect 22330 107270 22353 108277
rect 22147 106270 22353 107270
rect 22147 105293 22170 106270
rect 19140 105270 22170 105293
rect 22330 105293 22353 106270
rect 25337 107270 25360 108277
rect 25520 108277 28550 108300
rect 25520 107270 25543 108277
rect 25337 106270 25543 107270
rect 25337 105293 25360 106270
rect 22330 105270 25360 105293
rect 25520 105293 25543 106270
rect 28527 107270 28550 108277
rect 28710 108277 31740 108300
rect 28710 107270 28733 108277
rect 28527 106270 28733 107270
rect 28527 105293 28550 106270
rect 25520 105270 28550 105293
rect 28710 105293 28733 106270
rect 31717 107270 31740 108277
rect 31900 108277 34930 108300
rect 31900 107270 31923 108277
rect 31717 106270 31923 107270
rect 31717 105293 31740 106270
rect 28710 105270 31740 105293
rect 31900 105293 31923 106270
rect 34907 107270 34930 108277
rect 35090 108277 38120 108300
rect 35090 107270 35113 108277
rect 34907 106270 35113 107270
rect 34907 105293 34930 106270
rect 31900 105270 34930 105293
rect 35090 105293 35113 106270
rect 38097 107270 38120 108277
rect 38280 108277 41310 108300
rect 38280 107270 38303 108277
rect 38097 106270 38303 107270
rect 38097 105293 38120 106270
rect 35090 105270 38120 105293
rect 38280 105293 38303 106270
rect 41287 107270 41310 108277
rect 41470 108277 44500 108300
rect 41470 107270 41493 108277
rect 41287 106270 41493 107270
rect 41287 105293 41310 106270
rect 38280 105270 41310 105293
rect 41470 105293 41493 106270
rect 44477 107270 44500 108277
rect 44660 108277 47690 108300
rect 44660 107270 44683 108277
rect 44477 106270 44683 107270
rect 44477 105293 44500 106270
rect 41470 105270 44500 105293
rect 44660 105293 44683 106270
rect 47667 107270 47690 108277
rect 47850 108277 50880 108300
rect 47850 107270 47873 108277
rect 47667 106270 47873 107270
rect 47667 105293 47690 106270
rect 44660 105270 47690 105293
rect 47850 105293 47873 106270
rect 50857 107270 50880 108277
rect 51040 108277 54070 108300
rect 51040 107270 51063 108277
rect 50857 106270 51063 107270
rect 50857 105293 50880 106270
rect 47850 105270 50880 105293
rect 51040 105293 51063 106270
rect 54047 107270 54070 108277
rect 54230 108277 57260 108300
rect 54230 107270 54253 108277
rect 54047 106270 54253 107270
rect 54047 105293 54070 106270
rect 51040 105270 54070 105293
rect 54230 105293 54253 106270
rect 57237 107270 57260 108277
rect 57420 108277 60450 108300
rect 57420 107270 57443 108277
rect 57237 106270 57443 107270
rect 57237 105293 57260 106270
rect 54230 105270 57260 105293
rect 57420 105293 57443 106270
rect 60427 107270 60450 108277
rect 60610 108277 63640 108300
rect 60610 107270 60633 108277
rect 60427 106270 60633 107270
rect 60427 105293 60450 106270
rect 57420 105270 60450 105293
rect 60610 105293 60633 106270
rect 63617 107270 63640 108277
rect 63800 108277 66830 108300
rect 63800 107270 63823 108277
rect 63617 106270 63823 107270
rect 63617 105293 63640 106270
rect 60610 105270 63640 105293
rect 63800 105293 63823 106270
rect 66807 107270 66830 108277
rect 66990 108277 70020 108300
rect 66990 107270 67013 108277
rect 66807 106270 67013 107270
rect 66807 105293 66830 106270
rect 63800 105270 66830 105293
rect 66990 105293 67013 106270
rect 69997 107270 70020 108277
rect 70180 108277 73210 108300
rect 70180 107270 70203 108277
rect 69997 106270 70203 107270
rect 69997 105293 70020 106270
rect 66990 105270 70020 105293
rect 70180 105293 70203 106270
rect 73187 107270 73210 108277
rect 73370 108277 76400 108300
rect 73370 107270 73393 108277
rect 73187 106270 73393 107270
rect 73187 105293 73210 106270
rect 70180 105270 73210 105293
rect 73370 105293 73393 106270
rect 76377 107270 76400 108277
rect 76560 108277 79590 108300
rect 76560 107270 76583 108277
rect 76377 106270 76583 107270
rect 76377 105293 76400 106270
rect 73370 105270 76400 105293
rect 76560 105293 76583 106270
rect 79567 107270 79590 108277
rect 79750 108277 82780 108300
rect 79750 107270 79773 108277
rect 79567 106270 79773 107270
rect 79567 105293 79590 106270
rect 76560 105270 79590 105293
rect 79750 105293 79773 106270
rect 82757 107270 82780 108277
rect 82940 108277 85970 108300
rect 82940 107270 82963 108277
rect 82757 106270 82963 107270
rect 82757 105293 82780 106270
rect 79750 105270 82780 105293
rect 82940 105293 82963 106270
rect 85947 107270 85970 108277
rect 86130 108277 89160 108300
rect 86130 107270 86153 108277
rect 85947 106270 86153 107270
rect 85947 105293 85970 106270
rect 82940 105270 85970 105293
rect 86130 105293 86153 106270
rect 89137 107270 89160 108277
rect 89320 108277 92350 108300
rect 89320 107270 89343 108277
rect 89137 106270 89343 107270
rect 89137 105293 89160 106270
rect 86130 105270 89160 105293
rect 89320 105293 89343 106270
rect 92327 107270 92350 108277
rect 92510 108277 95540 108300
rect 92510 107270 92533 108277
rect 92327 106270 92533 107270
rect 92327 105293 92350 106270
rect 89320 105270 92350 105293
rect 92510 105293 92533 106270
rect 95517 107270 95540 108277
rect 95700 108277 98730 108300
rect 95700 107270 95723 108277
rect 95517 106270 95723 107270
rect 95517 105293 95540 106270
rect 92510 105270 95540 105293
rect 95700 105293 95723 106270
rect 98707 107270 98730 108277
rect 98890 108277 101920 108300
rect 98890 107270 98913 108277
rect 98707 106270 98913 107270
rect 98707 105293 98730 106270
rect 95700 105270 98730 105293
rect 98890 105293 98913 106270
rect 101897 107270 101920 108277
rect 102080 108277 105110 108300
rect 102080 107270 102103 108277
rect 101897 106270 102103 107270
rect 101897 105293 101920 106270
rect 98890 105270 101920 105293
rect 102080 105293 102103 106270
rect 105087 107270 105110 108277
rect 105270 108277 108300 108300
rect 105270 107270 105293 108277
rect 105087 106270 105293 107270
rect 105087 105293 105110 106270
rect 102080 105270 105110 105293
rect 105270 105293 105293 106270
rect 108277 107270 108300 108277
rect 108460 108277 111490 108300
rect 108460 107270 108483 108277
rect 108277 106270 108483 107270
rect 108277 105293 108300 106270
rect 105270 105270 108300 105293
rect 108460 105293 108483 106270
rect 111467 107270 111490 108277
rect 111650 108277 114680 108300
rect 111650 107270 111673 108277
rect 111467 106270 111673 107270
rect 111467 105293 111490 106270
rect 108460 105270 111490 105293
rect 111650 105293 111673 106270
rect 114657 107270 114680 108277
rect 114840 108277 117870 108300
rect 114840 107270 114863 108277
rect 114657 106270 114863 107270
rect 114657 105293 114680 106270
rect 111650 105270 114680 105293
rect 114840 105293 114863 106270
rect 117847 107270 117870 108277
rect 118030 108277 121060 108300
rect 118030 107270 118053 108277
rect 117847 106270 118053 107270
rect 117847 105293 117870 106270
rect 114840 105270 117870 105293
rect 118030 105293 118053 106270
rect 121037 107270 121060 108277
rect 121220 108277 124250 108300
rect 121220 107270 121243 108277
rect 121037 106270 121243 107270
rect 121037 105293 121060 106270
rect 118030 105270 121060 105293
rect 121220 105293 121243 106270
rect 124227 107270 124250 108277
rect 124410 108277 127440 108300
rect 124410 107270 124433 108277
rect 124227 106270 124433 107270
rect 124227 105293 124250 106270
rect 121220 105270 124250 105293
rect 124410 105293 124433 106270
rect 127417 107270 127440 108277
rect 127600 108277 130630 108300
rect 127600 107270 127623 108277
rect 127417 106270 127623 107270
rect 127417 105293 127440 106270
rect 124410 105270 127440 105293
rect 127600 105293 127623 106270
rect 130607 107270 130630 108277
rect 130790 108277 133820 108300
rect 130790 107270 130813 108277
rect 130607 106270 130813 107270
rect 130607 105293 130630 106270
rect 127600 105270 130630 105293
rect 130790 105293 130813 106270
rect 133797 107270 133820 108277
rect 133980 108277 137010 108300
rect 133980 107270 134003 108277
rect 133797 106270 134003 107270
rect 133797 105293 133820 106270
rect 130790 105270 133820 105293
rect 133980 105293 134003 106270
rect 136987 107270 137010 108277
rect 136987 106270 137170 107270
rect 136987 105293 137010 106270
rect 133980 105270 137010 105293
rect 1000 105110 2000 105270
rect 4190 105110 5190 105270
rect 7380 105110 8380 105270
rect 10570 105110 11570 105270
rect 13760 105110 14760 105270
rect 16950 105110 17950 105270
rect 20140 105110 21140 105270
rect 23330 105110 24330 105270
rect 26520 105110 27520 105270
rect 29710 105110 30710 105270
rect 32900 105110 33900 105270
rect 36090 105110 37090 105270
rect 39280 105110 40280 105270
rect 42470 105110 43470 105270
rect 45660 105110 46660 105270
rect 48850 105110 49850 105270
rect 52040 105110 53040 105270
rect 55230 105110 56230 105270
rect 58420 105110 59420 105270
rect 61610 105110 62610 105270
rect 64800 105110 65800 105270
rect 67990 105110 68990 105270
rect 71180 105110 72180 105270
rect 74370 105110 75370 105270
rect 77560 105110 78560 105270
rect 80750 105110 81750 105270
rect 83940 105110 84940 105270
rect 87130 105110 88130 105270
rect 90320 105110 91320 105270
rect 93510 105110 94510 105270
rect 96700 105110 97700 105270
rect 99890 105110 100890 105270
rect 103080 105110 104080 105270
rect 106270 105110 107270 105270
rect 109460 105110 110460 105270
rect 112650 105110 113650 105270
rect 115840 105110 116840 105270
rect 119030 105110 120030 105270
rect 122220 105110 123220 105270
rect 125410 105110 126410 105270
rect 128600 105110 129600 105270
rect 131790 105110 132790 105270
rect 134980 105110 135980 105270
rect 0 105087 3030 105110
rect 0 102103 23 105087
rect 3007 104080 3030 105087
rect 3190 105087 6220 105110
rect 3190 104080 3213 105087
rect 3007 103080 3213 104080
rect 3007 102103 3030 103080
rect 0 102080 3030 102103
rect 3190 102103 3213 103080
rect 6197 104080 6220 105087
rect 6380 105087 9410 105110
rect 6380 104080 6403 105087
rect 6197 103080 6403 104080
rect 6197 102103 6220 103080
rect 3190 102080 6220 102103
rect 6380 102103 6403 103080
rect 9387 104080 9410 105087
rect 9570 105087 12600 105110
rect 9570 104080 9593 105087
rect 9387 103080 9593 104080
rect 9387 102103 9410 103080
rect 6380 102080 9410 102103
rect 9570 102103 9593 103080
rect 12577 104080 12600 105087
rect 12760 105087 15790 105110
rect 12760 104080 12783 105087
rect 12577 103080 12783 104080
rect 12577 102103 12600 103080
rect 9570 102080 12600 102103
rect 12760 102103 12783 103080
rect 15767 104080 15790 105087
rect 15950 105087 18980 105110
rect 15950 104080 15973 105087
rect 15767 103080 15973 104080
rect 15767 102103 15790 103080
rect 12760 102080 15790 102103
rect 15950 102103 15973 103080
rect 18957 104080 18980 105087
rect 19140 105087 22170 105110
rect 19140 104080 19163 105087
rect 18957 103080 19163 104080
rect 18957 102103 18980 103080
rect 15950 102080 18980 102103
rect 19140 102103 19163 103080
rect 22147 104080 22170 105087
rect 22330 105087 25360 105110
rect 22330 104080 22353 105087
rect 22147 103080 22353 104080
rect 22147 102103 22170 103080
rect 19140 102080 22170 102103
rect 22330 102103 22353 103080
rect 25337 104080 25360 105087
rect 25520 105087 28550 105110
rect 25520 104080 25543 105087
rect 25337 103080 25543 104080
rect 25337 102103 25360 103080
rect 22330 102080 25360 102103
rect 25520 102103 25543 103080
rect 28527 104080 28550 105087
rect 28710 105087 31740 105110
rect 28710 104080 28733 105087
rect 28527 103080 28733 104080
rect 28527 102103 28550 103080
rect 25520 102080 28550 102103
rect 28710 102103 28733 103080
rect 31717 104080 31740 105087
rect 31900 105087 34930 105110
rect 31900 104080 31923 105087
rect 31717 103080 31923 104080
rect 31717 102103 31740 103080
rect 28710 102080 31740 102103
rect 31900 102103 31923 103080
rect 34907 104080 34930 105087
rect 35090 105087 38120 105110
rect 35090 104080 35113 105087
rect 34907 103080 35113 104080
rect 34907 102103 34930 103080
rect 31900 102080 34930 102103
rect 35090 102103 35113 103080
rect 38097 104080 38120 105087
rect 38280 105087 41310 105110
rect 38280 104080 38303 105087
rect 38097 103080 38303 104080
rect 38097 102103 38120 103080
rect 35090 102080 38120 102103
rect 38280 102103 38303 103080
rect 41287 104080 41310 105087
rect 41470 105087 44500 105110
rect 41470 104080 41493 105087
rect 41287 103080 41493 104080
rect 41287 102103 41310 103080
rect 38280 102080 41310 102103
rect 41470 102103 41493 103080
rect 44477 104080 44500 105087
rect 44660 105087 47690 105110
rect 44660 104080 44683 105087
rect 44477 103080 44683 104080
rect 44477 102103 44500 103080
rect 41470 102080 44500 102103
rect 44660 102103 44683 103080
rect 47667 104080 47690 105087
rect 47850 105087 50880 105110
rect 47850 104080 47873 105087
rect 47667 103080 47873 104080
rect 47667 102103 47690 103080
rect 44660 102080 47690 102103
rect 47850 102103 47873 103080
rect 50857 104080 50880 105087
rect 51040 105087 54070 105110
rect 51040 104080 51063 105087
rect 50857 103080 51063 104080
rect 50857 102103 50880 103080
rect 47850 102080 50880 102103
rect 51040 102103 51063 103080
rect 54047 104080 54070 105087
rect 54230 105087 57260 105110
rect 54230 104080 54253 105087
rect 54047 103080 54253 104080
rect 54047 102103 54070 103080
rect 51040 102080 54070 102103
rect 54230 102103 54253 103080
rect 57237 104080 57260 105087
rect 57420 105087 60450 105110
rect 57420 104080 57443 105087
rect 57237 103080 57443 104080
rect 57237 102103 57260 103080
rect 54230 102080 57260 102103
rect 57420 102103 57443 103080
rect 60427 104080 60450 105087
rect 60610 105087 63640 105110
rect 60610 104080 60633 105087
rect 60427 103080 60633 104080
rect 60427 102103 60450 103080
rect 57420 102080 60450 102103
rect 60610 102103 60633 103080
rect 63617 104080 63640 105087
rect 63800 105087 66830 105110
rect 63800 104080 63823 105087
rect 63617 103080 63823 104080
rect 63617 102103 63640 103080
rect 60610 102080 63640 102103
rect 63800 102103 63823 103080
rect 66807 104080 66830 105087
rect 66990 105087 70020 105110
rect 66990 104080 67013 105087
rect 66807 103080 67013 104080
rect 66807 102103 66830 103080
rect 63800 102080 66830 102103
rect 66990 102103 67013 103080
rect 69997 104080 70020 105087
rect 70180 105087 73210 105110
rect 70180 104080 70203 105087
rect 69997 103080 70203 104080
rect 69997 102103 70020 103080
rect 66990 102080 70020 102103
rect 70180 102103 70203 103080
rect 73187 104080 73210 105087
rect 73370 105087 76400 105110
rect 73370 104080 73393 105087
rect 73187 103080 73393 104080
rect 73187 102103 73210 103080
rect 70180 102080 73210 102103
rect 73370 102103 73393 103080
rect 76377 104080 76400 105087
rect 76560 105087 79590 105110
rect 76560 104080 76583 105087
rect 76377 103080 76583 104080
rect 76377 102103 76400 103080
rect 73370 102080 76400 102103
rect 76560 102103 76583 103080
rect 79567 104080 79590 105087
rect 79750 105087 82780 105110
rect 79750 104080 79773 105087
rect 79567 103080 79773 104080
rect 79567 102103 79590 103080
rect 76560 102080 79590 102103
rect 79750 102103 79773 103080
rect 82757 104080 82780 105087
rect 82940 105087 85970 105110
rect 82940 104080 82963 105087
rect 82757 103080 82963 104080
rect 82757 102103 82780 103080
rect 79750 102080 82780 102103
rect 82940 102103 82963 103080
rect 85947 104080 85970 105087
rect 86130 105087 89160 105110
rect 86130 104080 86153 105087
rect 85947 103080 86153 104080
rect 85947 102103 85970 103080
rect 82940 102080 85970 102103
rect 86130 102103 86153 103080
rect 89137 104080 89160 105087
rect 89320 105087 92350 105110
rect 89320 104080 89343 105087
rect 89137 103080 89343 104080
rect 89137 102103 89160 103080
rect 86130 102080 89160 102103
rect 89320 102103 89343 103080
rect 92327 104080 92350 105087
rect 92510 105087 95540 105110
rect 92510 104080 92533 105087
rect 92327 103080 92533 104080
rect 92327 102103 92350 103080
rect 89320 102080 92350 102103
rect 92510 102103 92533 103080
rect 95517 104080 95540 105087
rect 95700 105087 98730 105110
rect 95700 104080 95723 105087
rect 95517 103080 95723 104080
rect 95517 102103 95540 103080
rect 92510 102080 95540 102103
rect 95700 102103 95723 103080
rect 98707 104080 98730 105087
rect 98890 105087 101920 105110
rect 98890 104080 98913 105087
rect 98707 103080 98913 104080
rect 98707 102103 98730 103080
rect 95700 102080 98730 102103
rect 98890 102103 98913 103080
rect 101897 104080 101920 105087
rect 102080 105087 105110 105110
rect 102080 104080 102103 105087
rect 101897 103080 102103 104080
rect 101897 102103 101920 103080
rect 98890 102080 101920 102103
rect 102080 102103 102103 103080
rect 105087 104080 105110 105087
rect 105270 105087 108300 105110
rect 105270 104080 105293 105087
rect 105087 103080 105293 104080
rect 105087 102103 105110 103080
rect 102080 102080 105110 102103
rect 105270 102103 105293 103080
rect 108277 104080 108300 105087
rect 108460 105087 111490 105110
rect 108460 104080 108483 105087
rect 108277 103080 108483 104080
rect 108277 102103 108300 103080
rect 105270 102080 108300 102103
rect 108460 102103 108483 103080
rect 111467 104080 111490 105087
rect 111650 105087 114680 105110
rect 111650 104080 111673 105087
rect 111467 103080 111673 104080
rect 111467 102103 111490 103080
rect 108460 102080 111490 102103
rect 111650 102103 111673 103080
rect 114657 104080 114680 105087
rect 114840 105087 117870 105110
rect 114840 104080 114863 105087
rect 114657 103080 114863 104080
rect 114657 102103 114680 103080
rect 111650 102080 114680 102103
rect 114840 102103 114863 103080
rect 117847 104080 117870 105087
rect 118030 105087 121060 105110
rect 118030 104080 118053 105087
rect 117847 103080 118053 104080
rect 117847 102103 117870 103080
rect 114840 102080 117870 102103
rect 118030 102103 118053 103080
rect 121037 104080 121060 105087
rect 121220 105087 124250 105110
rect 121220 104080 121243 105087
rect 121037 103080 121243 104080
rect 121037 102103 121060 103080
rect 118030 102080 121060 102103
rect 121220 102103 121243 103080
rect 124227 104080 124250 105087
rect 124410 105087 127440 105110
rect 124410 104080 124433 105087
rect 124227 103080 124433 104080
rect 124227 102103 124250 103080
rect 121220 102080 124250 102103
rect 124410 102103 124433 103080
rect 127417 104080 127440 105087
rect 127600 105087 130630 105110
rect 127600 104080 127623 105087
rect 127417 103080 127623 104080
rect 127417 102103 127440 103080
rect 124410 102080 127440 102103
rect 127600 102103 127623 103080
rect 130607 104080 130630 105087
rect 130790 105087 133820 105110
rect 130790 104080 130813 105087
rect 130607 103080 130813 104080
rect 130607 102103 130630 103080
rect 127600 102080 130630 102103
rect 130790 102103 130813 103080
rect 133797 104080 133820 105087
rect 133980 105087 137010 105110
rect 133980 104080 134003 105087
rect 133797 103080 134003 104080
rect 133797 102103 133820 103080
rect 130790 102080 133820 102103
rect 133980 102103 134003 103080
rect 136987 104080 137010 105087
rect 136987 103080 137170 104080
rect 136987 102103 137010 103080
rect 133980 102080 137010 102103
rect 1000 101920 2000 102080
rect 4190 101920 5190 102080
rect 7380 101920 8380 102080
rect 10570 101920 11570 102080
rect 13760 101920 14760 102080
rect 16950 101920 17950 102080
rect 20140 101920 21140 102080
rect 23330 101920 24330 102080
rect 26520 101920 27520 102080
rect 29710 101920 30710 102080
rect 32900 101920 33900 102080
rect 36090 101920 37090 102080
rect 39280 101920 40280 102080
rect 42470 101920 43470 102080
rect 45660 101920 46660 102080
rect 48850 101920 49850 102080
rect 52040 101920 53040 102080
rect 55230 101920 56230 102080
rect 58420 101920 59420 102080
rect 61610 101920 62610 102080
rect 64800 101920 65800 102080
rect 67990 101920 68990 102080
rect 71180 101920 72180 102080
rect 74370 101920 75370 102080
rect 77560 101920 78560 102080
rect 80750 101920 81750 102080
rect 83940 101920 84940 102080
rect 87130 101920 88130 102080
rect 90320 101920 91320 102080
rect 93510 101920 94510 102080
rect 96700 101920 97700 102080
rect 99890 101920 100890 102080
rect 103080 101920 104080 102080
rect 106270 101920 107270 102080
rect 109460 101920 110460 102080
rect 112650 101920 113650 102080
rect 115840 101920 116840 102080
rect 119030 101920 120030 102080
rect 122220 101920 123220 102080
rect 125410 101920 126410 102080
rect 128600 101920 129600 102080
rect 131790 101920 132790 102080
rect 134980 101920 135980 102080
rect 0 101897 3030 101920
rect 0 98913 23 101897
rect 3007 100890 3030 101897
rect 3190 101897 6220 101920
rect 3190 100890 3213 101897
rect 3007 99890 3213 100890
rect 3007 98913 3030 99890
rect 0 98890 3030 98913
rect 3190 98913 3213 99890
rect 6197 100890 6220 101897
rect 6380 101897 9410 101920
rect 6380 100890 6403 101897
rect 6197 99890 6403 100890
rect 6197 98913 6220 99890
rect 3190 98890 6220 98913
rect 6380 98913 6403 99890
rect 9387 100890 9410 101897
rect 9570 101897 12600 101920
rect 9570 100890 9593 101897
rect 9387 99890 9593 100890
rect 9387 98913 9410 99890
rect 6380 98890 9410 98913
rect 9570 98913 9593 99890
rect 12577 100890 12600 101897
rect 12760 101897 15790 101920
rect 12760 100890 12783 101897
rect 12577 99890 12783 100890
rect 12577 98913 12600 99890
rect 9570 98890 12600 98913
rect 12760 98913 12783 99890
rect 15767 100890 15790 101897
rect 15950 101897 18980 101920
rect 15950 100890 15973 101897
rect 15767 99890 15973 100890
rect 15767 98913 15790 99890
rect 12760 98890 15790 98913
rect 15950 98913 15973 99890
rect 18957 100890 18980 101897
rect 19140 101897 22170 101920
rect 19140 100890 19163 101897
rect 18957 99890 19163 100890
rect 18957 98913 18980 99890
rect 15950 98890 18980 98913
rect 19140 98913 19163 99890
rect 22147 100890 22170 101897
rect 22330 101897 25360 101920
rect 22330 100890 22353 101897
rect 22147 99890 22353 100890
rect 22147 98913 22170 99890
rect 19140 98890 22170 98913
rect 22330 98913 22353 99890
rect 25337 100890 25360 101897
rect 25520 101897 28550 101920
rect 25520 100890 25543 101897
rect 25337 99890 25543 100890
rect 25337 98913 25360 99890
rect 22330 98890 25360 98913
rect 25520 98913 25543 99890
rect 28527 100890 28550 101897
rect 28710 101897 31740 101920
rect 28710 100890 28733 101897
rect 28527 99890 28733 100890
rect 28527 98913 28550 99890
rect 25520 98890 28550 98913
rect 28710 98913 28733 99890
rect 31717 100890 31740 101897
rect 31900 101897 34930 101920
rect 31900 100890 31923 101897
rect 31717 99890 31923 100890
rect 31717 98913 31740 99890
rect 28710 98890 31740 98913
rect 31900 98913 31923 99890
rect 34907 100890 34930 101897
rect 35090 101897 38120 101920
rect 35090 100890 35113 101897
rect 34907 99890 35113 100890
rect 34907 98913 34930 99890
rect 31900 98890 34930 98913
rect 35090 98913 35113 99890
rect 38097 100890 38120 101897
rect 38280 101897 41310 101920
rect 38280 100890 38303 101897
rect 38097 99890 38303 100890
rect 38097 98913 38120 99890
rect 35090 98890 38120 98913
rect 38280 98913 38303 99890
rect 41287 100890 41310 101897
rect 41470 101897 44500 101920
rect 41470 100890 41493 101897
rect 41287 99890 41493 100890
rect 41287 98913 41310 99890
rect 38280 98890 41310 98913
rect 41470 98913 41493 99890
rect 44477 100890 44500 101897
rect 44660 101897 47690 101920
rect 44660 100890 44683 101897
rect 44477 99890 44683 100890
rect 44477 98913 44500 99890
rect 41470 98890 44500 98913
rect 44660 98913 44683 99890
rect 47667 100890 47690 101897
rect 47850 101897 50880 101920
rect 47850 100890 47873 101897
rect 47667 99890 47873 100890
rect 47667 98913 47690 99890
rect 44660 98890 47690 98913
rect 47850 98913 47873 99890
rect 50857 100890 50880 101897
rect 51040 101897 54070 101920
rect 51040 100890 51063 101897
rect 50857 99890 51063 100890
rect 50857 98913 50880 99890
rect 47850 98890 50880 98913
rect 51040 98913 51063 99890
rect 54047 100890 54070 101897
rect 54230 101897 57260 101920
rect 54230 100890 54253 101897
rect 54047 99890 54253 100890
rect 54047 98913 54070 99890
rect 51040 98890 54070 98913
rect 54230 98913 54253 99890
rect 57237 100890 57260 101897
rect 57420 101897 60450 101920
rect 57420 100890 57443 101897
rect 57237 99890 57443 100890
rect 57237 98913 57260 99890
rect 54230 98890 57260 98913
rect 57420 98913 57443 99890
rect 60427 100890 60450 101897
rect 60610 101897 63640 101920
rect 60610 100890 60633 101897
rect 60427 99890 60633 100890
rect 60427 98913 60450 99890
rect 57420 98890 60450 98913
rect 60610 98913 60633 99890
rect 63617 100890 63640 101897
rect 63800 101897 66830 101920
rect 63800 100890 63823 101897
rect 63617 99890 63823 100890
rect 63617 98913 63640 99890
rect 60610 98890 63640 98913
rect 63800 98913 63823 99890
rect 66807 100890 66830 101897
rect 66990 101897 70020 101920
rect 66990 100890 67013 101897
rect 66807 99890 67013 100890
rect 66807 98913 66830 99890
rect 63800 98890 66830 98913
rect 66990 98913 67013 99890
rect 69997 100890 70020 101897
rect 70180 101897 73210 101920
rect 70180 100890 70203 101897
rect 69997 99890 70203 100890
rect 69997 98913 70020 99890
rect 66990 98890 70020 98913
rect 70180 98913 70203 99890
rect 73187 100890 73210 101897
rect 73370 101897 76400 101920
rect 73370 100890 73393 101897
rect 73187 99890 73393 100890
rect 73187 98913 73210 99890
rect 70180 98890 73210 98913
rect 73370 98913 73393 99890
rect 76377 100890 76400 101897
rect 76560 101897 79590 101920
rect 76560 100890 76583 101897
rect 76377 99890 76583 100890
rect 76377 98913 76400 99890
rect 73370 98890 76400 98913
rect 76560 98913 76583 99890
rect 79567 100890 79590 101897
rect 79750 101897 82780 101920
rect 79750 100890 79773 101897
rect 79567 99890 79773 100890
rect 79567 98913 79590 99890
rect 76560 98890 79590 98913
rect 79750 98913 79773 99890
rect 82757 100890 82780 101897
rect 82940 101897 85970 101920
rect 82940 100890 82963 101897
rect 82757 99890 82963 100890
rect 82757 98913 82780 99890
rect 79750 98890 82780 98913
rect 82940 98913 82963 99890
rect 85947 100890 85970 101897
rect 86130 101897 89160 101920
rect 86130 100890 86153 101897
rect 85947 99890 86153 100890
rect 85947 98913 85970 99890
rect 82940 98890 85970 98913
rect 86130 98913 86153 99890
rect 89137 100890 89160 101897
rect 89320 101897 92350 101920
rect 89320 100890 89343 101897
rect 89137 99890 89343 100890
rect 89137 98913 89160 99890
rect 86130 98890 89160 98913
rect 89320 98913 89343 99890
rect 92327 100890 92350 101897
rect 92510 101897 95540 101920
rect 92510 100890 92533 101897
rect 92327 99890 92533 100890
rect 92327 98913 92350 99890
rect 89320 98890 92350 98913
rect 92510 98913 92533 99890
rect 95517 100890 95540 101897
rect 95700 101897 98730 101920
rect 95700 100890 95723 101897
rect 95517 99890 95723 100890
rect 95517 98913 95540 99890
rect 92510 98890 95540 98913
rect 95700 98913 95723 99890
rect 98707 100890 98730 101897
rect 98890 101897 101920 101920
rect 98890 100890 98913 101897
rect 98707 99890 98913 100890
rect 98707 98913 98730 99890
rect 95700 98890 98730 98913
rect 98890 98913 98913 99890
rect 101897 100890 101920 101897
rect 102080 101897 105110 101920
rect 102080 100890 102103 101897
rect 101897 99890 102103 100890
rect 101897 98913 101920 99890
rect 98890 98890 101920 98913
rect 102080 98913 102103 99890
rect 105087 100890 105110 101897
rect 105270 101897 108300 101920
rect 105270 100890 105293 101897
rect 105087 99890 105293 100890
rect 105087 98913 105110 99890
rect 102080 98890 105110 98913
rect 105270 98913 105293 99890
rect 108277 100890 108300 101897
rect 108460 101897 111490 101920
rect 108460 100890 108483 101897
rect 108277 99890 108483 100890
rect 108277 98913 108300 99890
rect 105270 98890 108300 98913
rect 108460 98913 108483 99890
rect 111467 100890 111490 101897
rect 111650 101897 114680 101920
rect 111650 100890 111673 101897
rect 111467 99890 111673 100890
rect 111467 98913 111490 99890
rect 108460 98890 111490 98913
rect 111650 98913 111673 99890
rect 114657 100890 114680 101897
rect 114840 101897 117870 101920
rect 114840 100890 114863 101897
rect 114657 99890 114863 100890
rect 114657 98913 114680 99890
rect 111650 98890 114680 98913
rect 114840 98913 114863 99890
rect 117847 100890 117870 101897
rect 118030 101897 121060 101920
rect 118030 100890 118053 101897
rect 117847 99890 118053 100890
rect 117847 98913 117870 99890
rect 114840 98890 117870 98913
rect 118030 98913 118053 99890
rect 121037 100890 121060 101897
rect 121220 101897 124250 101920
rect 121220 100890 121243 101897
rect 121037 99890 121243 100890
rect 121037 98913 121060 99890
rect 118030 98890 121060 98913
rect 121220 98913 121243 99890
rect 124227 100890 124250 101897
rect 124410 101897 127440 101920
rect 124410 100890 124433 101897
rect 124227 99890 124433 100890
rect 124227 98913 124250 99890
rect 121220 98890 124250 98913
rect 124410 98913 124433 99890
rect 127417 100890 127440 101897
rect 127600 101897 130630 101920
rect 127600 100890 127623 101897
rect 127417 99890 127623 100890
rect 127417 98913 127440 99890
rect 124410 98890 127440 98913
rect 127600 98913 127623 99890
rect 130607 100890 130630 101897
rect 130790 101897 133820 101920
rect 130790 100890 130813 101897
rect 130607 99890 130813 100890
rect 130607 98913 130630 99890
rect 127600 98890 130630 98913
rect 130790 98913 130813 99890
rect 133797 100890 133820 101897
rect 133980 101897 137010 101920
rect 133980 100890 134003 101897
rect 133797 99890 134003 100890
rect 133797 98913 133820 99890
rect 130790 98890 133820 98913
rect 133980 98913 134003 99890
rect 136987 100890 137010 101897
rect 136987 99890 137170 100890
rect 136987 98913 137010 99890
rect 133980 98890 137010 98913
rect 1000 98889 2000 98890
rect 4190 98889 5190 98890
rect 7380 98889 8380 98890
rect 10570 98730 11570 98890
rect 13760 98730 14760 98890
rect 16950 98730 17950 98890
rect 20140 98730 21140 98890
rect 23330 98730 24330 98890
rect 26520 98730 27520 98890
rect 29710 98730 30710 98890
rect 32900 98730 33900 98890
rect 36090 98730 37090 98890
rect 39280 98730 40280 98890
rect 42470 98730 43470 98890
rect 45660 98730 46660 98890
rect 48850 98730 49850 98890
rect 52040 98730 53040 98890
rect 55230 98730 56230 98890
rect 58420 98730 59420 98890
rect 61610 98730 62610 98890
rect 64800 98730 65800 98890
rect 67990 98730 68990 98890
rect 71180 98730 72180 98890
rect 74370 98730 75370 98890
rect 77560 98730 78560 98890
rect 80750 98730 81750 98890
rect 83940 98730 84940 98890
rect 87130 98730 88130 98890
rect 90320 98730 91320 98890
rect 93510 98730 94510 98890
rect 96700 98730 97700 98890
rect 99890 98730 100890 98890
rect 103080 98730 104080 98890
rect 106270 98730 107270 98890
rect 109460 98730 110460 98890
rect 112650 98730 113650 98890
rect 115840 98730 116840 98890
rect 119030 98730 120030 98890
rect 122220 98730 123220 98890
rect 125410 98730 126410 98890
rect 128600 98730 129600 98890
rect 131790 98730 132790 98890
rect 134980 98730 135980 98890
rect 9570 98707 12600 98730
rect 0 98639 9370 98689
rect 0 79839 50 98639
rect 9320 79839 9370 98639
rect 9570 95723 9593 98707
rect 12577 97700 12600 98707
rect 12760 98707 15790 98730
rect 12760 97700 12783 98707
rect 12577 96700 12783 97700
rect 12577 95723 12600 96700
rect 9570 95700 12600 95723
rect 12760 95723 12783 96700
rect 15767 97700 15790 98707
rect 15950 98707 18980 98730
rect 15950 97700 15973 98707
rect 15767 96700 15973 97700
rect 15767 95723 15790 96700
rect 12760 95700 15790 95723
rect 15950 95723 15973 96700
rect 18957 97700 18980 98707
rect 19140 98707 22170 98730
rect 19140 97700 19163 98707
rect 18957 96700 19163 97700
rect 18957 95723 18980 96700
rect 15950 95700 18980 95723
rect 19140 95723 19163 96700
rect 22147 97700 22170 98707
rect 22330 98707 25360 98730
rect 22330 97700 22353 98707
rect 22147 96700 22353 97700
rect 22147 95723 22170 96700
rect 19140 95700 22170 95723
rect 22330 95723 22353 96700
rect 25337 97700 25360 98707
rect 25520 98707 28550 98730
rect 25520 97700 25543 98707
rect 25337 96700 25543 97700
rect 25337 95723 25360 96700
rect 22330 95700 25360 95723
rect 25520 95723 25543 96700
rect 28527 97700 28550 98707
rect 28710 98707 31740 98730
rect 28710 97700 28733 98707
rect 28527 96700 28733 97700
rect 28527 95723 28550 96700
rect 25520 95700 28550 95723
rect 28710 95723 28733 96700
rect 31717 97700 31740 98707
rect 31900 98707 34930 98730
rect 31900 97700 31923 98707
rect 31717 96700 31923 97700
rect 31717 95723 31740 96700
rect 28710 95700 31740 95723
rect 31900 95723 31923 96700
rect 34907 97700 34930 98707
rect 35090 98707 38120 98730
rect 35090 97700 35113 98707
rect 34907 96700 35113 97700
rect 34907 95723 34930 96700
rect 31900 95700 34930 95723
rect 35090 95723 35113 96700
rect 38097 97700 38120 98707
rect 38280 98707 41310 98730
rect 38280 97700 38303 98707
rect 38097 96700 38303 97700
rect 38097 95723 38120 96700
rect 35090 95700 38120 95723
rect 38280 95723 38303 96700
rect 41287 97700 41310 98707
rect 41470 98707 44500 98730
rect 41470 97700 41493 98707
rect 41287 96700 41493 97700
rect 41287 95723 41310 96700
rect 38280 95700 41310 95723
rect 41470 95723 41493 96700
rect 44477 97700 44500 98707
rect 44660 98707 47690 98730
rect 44660 97700 44683 98707
rect 44477 96700 44683 97700
rect 44477 95723 44500 96700
rect 41470 95700 44500 95723
rect 44660 95723 44683 96700
rect 47667 97700 47690 98707
rect 47850 98707 50880 98730
rect 47850 97700 47873 98707
rect 47667 96700 47873 97700
rect 47667 95723 47690 96700
rect 44660 95700 47690 95723
rect 47850 95723 47873 96700
rect 50857 97700 50880 98707
rect 51040 98707 54070 98730
rect 51040 97700 51063 98707
rect 50857 96700 51063 97700
rect 50857 95723 50880 96700
rect 47850 95700 50880 95723
rect 51040 95723 51063 96700
rect 54047 97700 54070 98707
rect 54230 98707 57260 98730
rect 54230 97700 54253 98707
rect 54047 96700 54253 97700
rect 54047 95723 54070 96700
rect 51040 95700 54070 95723
rect 54230 95723 54253 96700
rect 57237 97700 57260 98707
rect 57420 98707 60450 98730
rect 57420 97700 57443 98707
rect 57237 96700 57443 97700
rect 57237 95723 57260 96700
rect 54230 95700 57260 95723
rect 57420 95723 57443 96700
rect 60427 97700 60450 98707
rect 60610 98707 63640 98730
rect 60610 97700 60633 98707
rect 60427 96700 60633 97700
rect 60427 95723 60450 96700
rect 57420 95700 60450 95723
rect 60610 95723 60633 96700
rect 63617 97700 63640 98707
rect 63800 98707 66830 98730
rect 63800 97700 63823 98707
rect 63617 96700 63823 97700
rect 63617 95723 63640 96700
rect 60610 95700 63640 95723
rect 63800 95723 63823 96700
rect 66807 97700 66830 98707
rect 66990 98707 70020 98730
rect 66990 97700 67013 98707
rect 66807 96700 67013 97700
rect 66807 95723 66830 96700
rect 63800 95700 66830 95723
rect 66990 95723 67013 96700
rect 69997 97700 70020 98707
rect 70180 98707 73210 98730
rect 70180 97700 70203 98707
rect 69997 96700 70203 97700
rect 69997 95723 70020 96700
rect 66990 95700 70020 95723
rect 70180 95723 70203 96700
rect 73187 97700 73210 98707
rect 73370 98707 76400 98730
rect 73370 97700 73393 98707
rect 73187 96700 73393 97700
rect 73187 95723 73210 96700
rect 70180 95700 73210 95723
rect 73370 95723 73393 96700
rect 76377 97700 76400 98707
rect 76560 98707 79590 98730
rect 76560 97700 76583 98707
rect 76377 96700 76583 97700
rect 76377 95723 76400 96700
rect 73370 95700 76400 95723
rect 76560 95723 76583 96700
rect 79567 97700 79590 98707
rect 79750 98707 82780 98730
rect 79750 97700 79773 98707
rect 79567 96700 79773 97700
rect 79567 95723 79590 96700
rect 76560 95700 79590 95723
rect 79750 95723 79773 96700
rect 82757 97700 82780 98707
rect 82940 98707 85970 98730
rect 82940 97700 82963 98707
rect 82757 96700 82963 97700
rect 82757 95723 82780 96700
rect 79750 95700 82780 95723
rect 82940 95723 82963 96700
rect 85947 97700 85970 98707
rect 86130 98707 89160 98730
rect 86130 97700 86153 98707
rect 85947 96700 86153 97700
rect 85947 95723 85970 96700
rect 82940 95700 85970 95723
rect 86130 95723 86153 96700
rect 89137 97700 89160 98707
rect 89320 98707 92350 98730
rect 89320 97700 89343 98707
rect 89137 96700 89343 97700
rect 89137 95723 89160 96700
rect 86130 95700 89160 95723
rect 89320 95723 89343 96700
rect 92327 97700 92350 98707
rect 92510 98707 95540 98730
rect 92510 97700 92533 98707
rect 92327 96700 92533 97700
rect 92327 95723 92350 96700
rect 89320 95700 92350 95723
rect 92510 95723 92533 96700
rect 95517 97700 95540 98707
rect 95700 98707 98730 98730
rect 95700 97700 95723 98707
rect 95517 96700 95723 97700
rect 95517 95723 95540 96700
rect 92510 95700 95540 95723
rect 95700 95723 95723 96700
rect 98707 97700 98730 98707
rect 98890 98707 101920 98730
rect 98890 97700 98913 98707
rect 98707 96700 98913 97700
rect 98707 95723 98730 96700
rect 95700 95700 98730 95723
rect 98890 95723 98913 96700
rect 101897 97700 101920 98707
rect 102080 98707 105110 98730
rect 102080 97700 102103 98707
rect 101897 96700 102103 97700
rect 101897 95723 101920 96700
rect 98890 95700 101920 95723
rect 102080 95723 102103 96700
rect 105087 97700 105110 98707
rect 105270 98707 108300 98730
rect 105270 97700 105293 98707
rect 105087 96700 105293 97700
rect 105087 95723 105110 96700
rect 102080 95700 105110 95723
rect 105270 95723 105293 96700
rect 108277 97700 108300 98707
rect 108460 98707 111490 98730
rect 108460 97700 108483 98707
rect 108277 96700 108483 97700
rect 108277 95723 108300 96700
rect 105270 95700 108300 95723
rect 108460 95723 108483 96700
rect 111467 97700 111490 98707
rect 111650 98707 114680 98730
rect 111650 97700 111673 98707
rect 111467 96700 111673 97700
rect 111467 95723 111490 96700
rect 108460 95700 111490 95723
rect 111650 95723 111673 96700
rect 114657 97700 114680 98707
rect 114840 98707 117870 98730
rect 114840 97700 114863 98707
rect 114657 96700 114863 97700
rect 114657 95723 114680 96700
rect 111650 95700 114680 95723
rect 114840 95723 114863 96700
rect 117847 97700 117870 98707
rect 118030 98707 121060 98730
rect 118030 97700 118053 98707
rect 117847 96700 118053 97700
rect 117847 95723 117870 96700
rect 114840 95700 117870 95723
rect 118030 95723 118053 96700
rect 121037 97700 121060 98707
rect 121220 98707 124250 98730
rect 121220 97700 121243 98707
rect 121037 96700 121243 97700
rect 121037 95723 121060 96700
rect 118030 95700 121060 95723
rect 121220 95723 121243 96700
rect 124227 97700 124250 98707
rect 124410 98707 127440 98730
rect 124410 97700 124433 98707
rect 124227 96700 124433 97700
rect 124227 95723 124250 96700
rect 121220 95700 124250 95723
rect 124410 95723 124433 96700
rect 127417 97700 127440 98707
rect 127600 98707 130630 98730
rect 127600 97700 127623 98707
rect 127417 96700 127623 97700
rect 127417 95723 127440 96700
rect 124410 95700 127440 95723
rect 127600 95723 127623 96700
rect 130607 97700 130630 98707
rect 130790 98707 133820 98730
rect 130790 97700 130813 98707
rect 130607 96700 130813 97700
rect 130607 95723 130630 96700
rect 127600 95700 130630 95723
rect 130790 95723 130813 96700
rect 133797 97700 133820 98707
rect 133980 98707 137010 98730
rect 133980 97700 134003 98707
rect 133797 96700 134003 97700
rect 133797 95723 133820 96700
rect 130790 95700 133820 95723
rect 133980 95723 134003 96700
rect 136987 97700 137010 98707
rect 136987 96700 137170 97700
rect 136987 95723 137010 96700
rect 133980 95700 137010 95723
rect 10570 95540 11570 95700
rect 13760 95540 14760 95700
rect 16950 95540 17950 95700
rect 20140 95540 21140 95700
rect 23330 95540 24330 95700
rect 26520 95540 27520 95700
rect 29710 95540 30710 95700
rect 32900 95540 33900 95700
rect 36090 95540 37090 95700
rect 39280 95540 40280 95700
rect 42470 95540 43470 95700
rect 45660 95540 46660 95700
rect 48850 95540 49850 95700
rect 52040 95540 53040 95700
rect 55230 95540 56230 95700
rect 58420 95540 59420 95700
rect 61610 95540 62610 95700
rect 64800 95540 65800 95700
rect 67990 95540 68990 95700
rect 71180 95540 72180 95700
rect 74370 95540 75370 95700
rect 77560 95540 78560 95700
rect 80750 95540 81750 95700
rect 83940 95540 84940 95700
rect 87130 95540 88130 95700
rect 90320 95540 91320 95700
rect 93510 95540 94510 95700
rect 96700 95540 97700 95700
rect 99890 95540 100890 95700
rect 103080 95540 104080 95700
rect 106270 95540 107270 95700
rect 109460 95540 110460 95700
rect 112650 95540 113650 95700
rect 115840 95540 116840 95700
rect 119030 95540 120030 95700
rect 122220 95540 123220 95700
rect 125410 95540 126410 95700
rect 128600 95540 129600 95700
rect 131790 95540 132790 95700
rect 134980 95540 135980 95700
rect 9570 95517 12600 95540
rect 9570 92533 9593 95517
rect 12577 94510 12600 95517
rect 12760 95517 15790 95540
rect 12760 94510 12783 95517
rect 12577 93510 12783 94510
rect 12577 92533 12600 93510
rect 9570 92510 12600 92533
rect 12760 92533 12783 93510
rect 15767 94510 15790 95517
rect 15950 95517 18980 95540
rect 15950 94510 15973 95517
rect 15767 93510 15973 94510
rect 15767 92533 15790 93510
rect 12760 92510 15790 92533
rect 15950 92533 15973 93510
rect 18957 94510 18980 95517
rect 19140 95517 22170 95540
rect 19140 94510 19163 95517
rect 18957 93510 19163 94510
rect 18957 92533 18980 93510
rect 15950 92510 18980 92533
rect 19140 92533 19163 93510
rect 22147 94510 22170 95517
rect 22330 95517 25360 95540
rect 22330 94510 22353 95517
rect 22147 93510 22353 94510
rect 22147 92533 22170 93510
rect 19140 92510 22170 92533
rect 22330 92533 22353 93510
rect 25337 94510 25360 95517
rect 25520 95517 28550 95540
rect 25520 94510 25543 95517
rect 25337 93510 25543 94510
rect 25337 92533 25360 93510
rect 22330 92510 25360 92533
rect 25520 92533 25543 93510
rect 28527 94510 28550 95517
rect 28710 95517 31740 95540
rect 28710 94510 28733 95517
rect 28527 93510 28733 94510
rect 28527 92533 28550 93510
rect 25520 92510 28550 92533
rect 28710 92533 28733 93510
rect 31717 94510 31740 95517
rect 31900 95517 34930 95540
rect 31900 94510 31923 95517
rect 31717 93510 31923 94510
rect 31717 92533 31740 93510
rect 28710 92510 31740 92533
rect 31900 92533 31923 93510
rect 34907 94510 34930 95517
rect 35090 95517 38120 95540
rect 35090 94510 35113 95517
rect 34907 93510 35113 94510
rect 34907 92533 34930 93510
rect 31900 92510 34930 92533
rect 35090 92533 35113 93510
rect 38097 94510 38120 95517
rect 38280 95517 41310 95540
rect 38280 94510 38303 95517
rect 38097 93510 38303 94510
rect 38097 92533 38120 93510
rect 35090 92510 38120 92533
rect 38280 92533 38303 93510
rect 41287 94510 41310 95517
rect 41470 95517 44500 95540
rect 41470 94510 41493 95517
rect 41287 93510 41493 94510
rect 41287 92533 41310 93510
rect 38280 92510 41310 92533
rect 41470 92533 41493 93510
rect 44477 94510 44500 95517
rect 44660 95517 47690 95540
rect 44660 94510 44683 95517
rect 44477 93510 44683 94510
rect 44477 92533 44500 93510
rect 41470 92510 44500 92533
rect 44660 92533 44683 93510
rect 47667 94510 47690 95517
rect 47850 95517 50880 95540
rect 47850 94510 47873 95517
rect 47667 93510 47873 94510
rect 47667 92533 47690 93510
rect 44660 92510 47690 92533
rect 47850 92533 47873 93510
rect 50857 94510 50880 95517
rect 51040 95517 54070 95540
rect 51040 94510 51063 95517
rect 50857 93510 51063 94510
rect 50857 92533 50880 93510
rect 47850 92510 50880 92533
rect 51040 92533 51063 93510
rect 54047 94510 54070 95517
rect 54230 95517 57260 95540
rect 54230 94510 54253 95517
rect 54047 93510 54253 94510
rect 54047 92533 54070 93510
rect 51040 92510 54070 92533
rect 54230 92533 54253 93510
rect 57237 94510 57260 95517
rect 57420 95517 60450 95540
rect 57420 94510 57443 95517
rect 57237 93510 57443 94510
rect 57237 92533 57260 93510
rect 54230 92510 57260 92533
rect 57420 92533 57443 93510
rect 60427 94510 60450 95517
rect 60610 95517 63640 95540
rect 60610 94510 60633 95517
rect 60427 93510 60633 94510
rect 60427 92533 60450 93510
rect 57420 92510 60450 92533
rect 60610 92533 60633 93510
rect 63617 94510 63640 95517
rect 63800 95517 66830 95540
rect 63800 94510 63823 95517
rect 63617 93510 63823 94510
rect 63617 92533 63640 93510
rect 60610 92510 63640 92533
rect 63800 92533 63823 93510
rect 66807 94510 66830 95517
rect 66990 95517 70020 95540
rect 66990 94510 67013 95517
rect 66807 93510 67013 94510
rect 66807 92533 66830 93510
rect 63800 92510 66830 92533
rect 66990 92533 67013 93510
rect 69997 94510 70020 95517
rect 70180 95517 73210 95540
rect 70180 94510 70203 95517
rect 69997 93510 70203 94510
rect 69997 92533 70020 93510
rect 66990 92510 70020 92533
rect 70180 92533 70203 93510
rect 73187 94510 73210 95517
rect 73370 95517 76400 95540
rect 73370 94510 73393 95517
rect 73187 93510 73393 94510
rect 73187 92533 73210 93510
rect 70180 92510 73210 92533
rect 73370 92533 73393 93510
rect 76377 94510 76400 95517
rect 76560 95517 79590 95540
rect 76560 94510 76583 95517
rect 76377 93510 76583 94510
rect 76377 92533 76400 93510
rect 73370 92510 76400 92533
rect 76560 92533 76583 93510
rect 79567 94510 79590 95517
rect 79750 95517 82780 95540
rect 79750 94510 79773 95517
rect 79567 93510 79773 94510
rect 79567 92533 79590 93510
rect 76560 92510 79590 92533
rect 79750 92533 79773 93510
rect 82757 94510 82780 95517
rect 82940 95517 85970 95540
rect 82940 94510 82963 95517
rect 82757 93510 82963 94510
rect 82757 92533 82780 93510
rect 79750 92510 82780 92533
rect 82940 92533 82963 93510
rect 85947 94510 85970 95517
rect 86130 95517 89160 95540
rect 86130 94510 86153 95517
rect 85947 93510 86153 94510
rect 85947 92533 85970 93510
rect 82940 92510 85970 92533
rect 86130 92533 86153 93510
rect 89137 94510 89160 95517
rect 89320 95517 92350 95540
rect 89320 94510 89343 95517
rect 89137 93510 89343 94510
rect 89137 92533 89160 93510
rect 86130 92510 89160 92533
rect 89320 92533 89343 93510
rect 92327 94510 92350 95517
rect 92510 95517 95540 95540
rect 92510 94510 92533 95517
rect 92327 93510 92533 94510
rect 92327 92533 92350 93510
rect 89320 92510 92350 92533
rect 92510 92533 92533 93510
rect 95517 94510 95540 95517
rect 95700 95517 98730 95540
rect 95700 94510 95723 95517
rect 95517 93510 95723 94510
rect 95517 92533 95540 93510
rect 92510 92510 95540 92533
rect 95700 92533 95723 93510
rect 98707 94510 98730 95517
rect 98890 95517 101920 95540
rect 98890 94510 98913 95517
rect 98707 93510 98913 94510
rect 98707 92533 98730 93510
rect 95700 92510 98730 92533
rect 98890 92533 98913 93510
rect 101897 94510 101920 95517
rect 102080 95517 105110 95540
rect 102080 94510 102103 95517
rect 101897 93510 102103 94510
rect 101897 92533 101920 93510
rect 98890 92510 101920 92533
rect 102080 92533 102103 93510
rect 105087 94510 105110 95517
rect 105270 95517 108300 95540
rect 105270 94510 105293 95517
rect 105087 93510 105293 94510
rect 105087 92533 105110 93510
rect 102080 92510 105110 92533
rect 105270 92533 105293 93510
rect 108277 94510 108300 95517
rect 108460 95517 111490 95540
rect 108460 94510 108483 95517
rect 108277 93510 108483 94510
rect 108277 92533 108300 93510
rect 105270 92510 108300 92533
rect 108460 92533 108483 93510
rect 111467 94510 111490 95517
rect 111650 95517 114680 95540
rect 111650 94510 111673 95517
rect 111467 93510 111673 94510
rect 111467 92533 111490 93510
rect 108460 92510 111490 92533
rect 111650 92533 111673 93510
rect 114657 94510 114680 95517
rect 114840 95517 117870 95540
rect 114840 94510 114863 95517
rect 114657 93510 114863 94510
rect 114657 92533 114680 93510
rect 111650 92510 114680 92533
rect 114840 92533 114863 93510
rect 117847 94510 117870 95517
rect 118030 95517 121060 95540
rect 118030 94510 118053 95517
rect 117847 93510 118053 94510
rect 117847 92533 117870 93510
rect 114840 92510 117870 92533
rect 118030 92533 118053 93510
rect 121037 94510 121060 95517
rect 121220 95517 124250 95540
rect 121220 94510 121243 95517
rect 121037 93510 121243 94510
rect 121037 92533 121060 93510
rect 118030 92510 121060 92533
rect 121220 92533 121243 93510
rect 124227 94510 124250 95517
rect 124410 95517 127440 95540
rect 124410 94510 124433 95517
rect 124227 93510 124433 94510
rect 124227 92533 124250 93510
rect 121220 92510 124250 92533
rect 124410 92533 124433 93510
rect 127417 94510 127440 95517
rect 127600 95517 130630 95540
rect 127600 94510 127623 95517
rect 127417 93510 127623 94510
rect 127417 92533 127440 93510
rect 124410 92510 127440 92533
rect 127600 92533 127623 93510
rect 130607 94510 130630 95517
rect 130790 95517 133820 95540
rect 130790 94510 130813 95517
rect 130607 93510 130813 94510
rect 130607 92533 130630 93510
rect 127600 92510 130630 92533
rect 130790 92533 130813 93510
rect 133797 94510 133820 95517
rect 133980 95517 137010 95540
rect 133980 94510 134003 95517
rect 133797 93510 134003 94510
rect 133797 92533 133820 93510
rect 130790 92510 133820 92533
rect 133980 92533 134003 93510
rect 136987 94510 137010 95517
rect 136987 93510 137170 94510
rect 136987 92533 137010 93510
rect 133980 92510 137010 92533
rect 10570 92350 11570 92510
rect 13760 92350 14760 92510
rect 16950 92350 17950 92510
rect 20140 92350 21140 92510
rect 23330 92350 24330 92510
rect 26520 92350 27520 92510
rect 29710 92350 30710 92510
rect 32900 92350 33900 92510
rect 36090 92350 37090 92510
rect 39280 92350 40280 92510
rect 42470 92350 43470 92510
rect 45660 92350 46660 92510
rect 48850 92350 49850 92510
rect 52040 92350 53040 92510
rect 55230 92350 56230 92510
rect 58420 92350 59420 92510
rect 61610 92350 62610 92510
rect 64800 92350 65800 92510
rect 67990 92350 68990 92510
rect 71180 92350 72180 92510
rect 74370 92350 75370 92510
rect 77560 92350 78560 92510
rect 80750 92350 81750 92510
rect 83940 92350 84940 92510
rect 87130 92350 88130 92510
rect 90320 92350 91320 92510
rect 93510 92350 94510 92510
rect 96700 92350 97700 92510
rect 99890 92350 100890 92510
rect 103080 92350 104080 92510
rect 106270 92350 107270 92510
rect 109460 92350 110460 92510
rect 112650 92350 113650 92510
rect 115840 92350 116840 92510
rect 119030 92350 120030 92510
rect 122220 92350 123220 92510
rect 125410 92350 126410 92510
rect 128600 92350 129600 92510
rect 131790 92350 132790 92510
rect 134980 92350 135980 92510
rect 9570 92327 12600 92350
rect 9570 89343 9593 92327
rect 12577 91320 12600 92327
rect 12760 92327 15790 92350
rect 12760 91320 12783 92327
rect 12577 90320 12783 91320
rect 12577 89343 12600 90320
rect 9570 89320 12600 89343
rect 12760 89343 12783 90320
rect 15767 91320 15790 92327
rect 15950 92327 18980 92350
rect 15950 91320 15973 92327
rect 15767 90320 15973 91320
rect 15767 89343 15790 90320
rect 12760 89320 15790 89343
rect 15950 89343 15973 90320
rect 18957 91320 18980 92327
rect 19140 92327 22170 92350
rect 19140 91320 19163 92327
rect 18957 90320 19163 91320
rect 18957 89343 18980 90320
rect 15950 89320 18980 89343
rect 19140 89343 19163 90320
rect 22147 91320 22170 92327
rect 22330 92327 25360 92350
rect 22330 91320 22353 92327
rect 22147 90320 22353 91320
rect 22147 89343 22170 90320
rect 19140 89320 22170 89343
rect 22330 89343 22353 90320
rect 25337 91320 25360 92327
rect 25520 92327 28550 92350
rect 25520 91320 25543 92327
rect 25337 90320 25543 91320
rect 25337 89343 25360 90320
rect 22330 89320 25360 89343
rect 25520 89343 25543 90320
rect 28527 91320 28550 92327
rect 28710 92327 31740 92350
rect 28710 91320 28733 92327
rect 28527 90320 28733 91320
rect 28527 89343 28550 90320
rect 25520 89320 28550 89343
rect 28710 89343 28733 90320
rect 31717 91320 31740 92327
rect 31900 92327 34930 92350
rect 31900 91320 31923 92327
rect 31717 90320 31923 91320
rect 31717 89343 31740 90320
rect 28710 89320 31740 89343
rect 31900 89343 31923 90320
rect 34907 91320 34930 92327
rect 35090 92327 38120 92350
rect 35090 91320 35113 92327
rect 34907 90320 35113 91320
rect 34907 89343 34930 90320
rect 31900 89320 34930 89343
rect 35090 89343 35113 90320
rect 38097 91320 38120 92327
rect 38280 92327 41310 92350
rect 38280 91320 38303 92327
rect 38097 90320 38303 91320
rect 38097 89343 38120 90320
rect 35090 89320 38120 89343
rect 38280 89343 38303 90320
rect 41287 91320 41310 92327
rect 41470 92327 44500 92350
rect 41470 91320 41493 92327
rect 41287 90320 41493 91320
rect 41287 89343 41310 90320
rect 38280 89320 41310 89343
rect 41470 89343 41493 90320
rect 44477 91320 44500 92327
rect 44660 92327 47690 92350
rect 44660 91320 44683 92327
rect 44477 90320 44683 91320
rect 44477 89343 44500 90320
rect 41470 89320 44500 89343
rect 44660 89343 44683 90320
rect 47667 91320 47690 92327
rect 47850 92327 50880 92350
rect 47850 91320 47873 92327
rect 47667 90320 47873 91320
rect 47667 89343 47690 90320
rect 44660 89320 47690 89343
rect 47850 89343 47873 90320
rect 50857 91320 50880 92327
rect 51040 92327 54070 92350
rect 51040 91320 51063 92327
rect 50857 90320 51063 91320
rect 50857 89343 50880 90320
rect 47850 89320 50880 89343
rect 51040 89343 51063 90320
rect 54047 91320 54070 92327
rect 54230 92327 57260 92350
rect 54230 91320 54253 92327
rect 54047 90320 54253 91320
rect 54047 89343 54070 90320
rect 51040 89320 54070 89343
rect 54230 89343 54253 90320
rect 57237 91320 57260 92327
rect 57420 92327 60450 92350
rect 57420 91320 57443 92327
rect 57237 90320 57443 91320
rect 57237 89343 57260 90320
rect 54230 89320 57260 89343
rect 57420 89343 57443 90320
rect 60427 91320 60450 92327
rect 60610 92327 63640 92350
rect 60610 91320 60633 92327
rect 60427 90320 60633 91320
rect 60427 89343 60450 90320
rect 57420 89320 60450 89343
rect 60610 89343 60633 90320
rect 63617 91320 63640 92327
rect 63800 92327 66830 92350
rect 63800 91320 63823 92327
rect 63617 90320 63823 91320
rect 63617 89343 63640 90320
rect 60610 89320 63640 89343
rect 63800 89343 63823 90320
rect 66807 91320 66830 92327
rect 66990 92327 70020 92350
rect 66990 91320 67013 92327
rect 66807 90320 67013 91320
rect 66807 89343 66830 90320
rect 63800 89320 66830 89343
rect 66990 89343 67013 90320
rect 69997 91320 70020 92327
rect 70180 92327 73210 92350
rect 70180 91320 70203 92327
rect 69997 90320 70203 91320
rect 69997 89343 70020 90320
rect 66990 89320 70020 89343
rect 70180 89343 70203 90320
rect 73187 91320 73210 92327
rect 73370 92327 76400 92350
rect 73370 91320 73393 92327
rect 73187 90320 73393 91320
rect 73187 89343 73210 90320
rect 70180 89320 73210 89343
rect 73370 89343 73393 90320
rect 76377 91320 76400 92327
rect 76560 92327 79590 92350
rect 76560 91320 76583 92327
rect 76377 90320 76583 91320
rect 76377 89343 76400 90320
rect 73370 89320 76400 89343
rect 76560 89343 76583 90320
rect 79567 91320 79590 92327
rect 79750 92327 82780 92350
rect 79750 91320 79773 92327
rect 79567 90320 79773 91320
rect 79567 89343 79590 90320
rect 76560 89320 79590 89343
rect 79750 89343 79773 90320
rect 82757 91320 82780 92327
rect 82940 92327 85970 92350
rect 82940 91320 82963 92327
rect 82757 90320 82963 91320
rect 82757 89343 82780 90320
rect 79750 89320 82780 89343
rect 82940 89343 82963 90320
rect 85947 91320 85970 92327
rect 86130 92327 89160 92350
rect 86130 91320 86153 92327
rect 85947 90320 86153 91320
rect 85947 89343 85970 90320
rect 82940 89320 85970 89343
rect 86130 89343 86153 90320
rect 89137 91320 89160 92327
rect 89320 92327 92350 92350
rect 89320 91320 89343 92327
rect 89137 90320 89343 91320
rect 89137 89343 89160 90320
rect 86130 89320 89160 89343
rect 89320 89343 89343 90320
rect 92327 91320 92350 92327
rect 92510 92327 95540 92350
rect 92510 91320 92533 92327
rect 92327 90320 92533 91320
rect 92327 89343 92350 90320
rect 89320 89320 92350 89343
rect 92510 89343 92533 90320
rect 95517 91320 95540 92327
rect 95700 92327 98730 92350
rect 95700 91320 95723 92327
rect 95517 90320 95723 91320
rect 95517 89343 95540 90320
rect 92510 89320 95540 89343
rect 95700 89343 95723 90320
rect 98707 91320 98730 92327
rect 98890 92327 101920 92350
rect 98890 91320 98913 92327
rect 98707 90320 98913 91320
rect 98707 89343 98730 90320
rect 95700 89320 98730 89343
rect 98890 89343 98913 90320
rect 101897 91320 101920 92327
rect 102080 92327 105110 92350
rect 102080 91320 102103 92327
rect 101897 90320 102103 91320
rect 101897 89343 101920 90320
rect 98890 89320 101920 89343
rect 102080 89343 102103 90320
rect 105087 91320 105110 92327
rect 105270 92327 108300 92350
rect 105270 91320 105293 92327
rect 105087 90320 105293 91320
rect 105087 89343 105110 90320
rect 102080 89320 105110 89343
rect 105270 89343 105293 90320
rect 108277 91320 108300 92327
rect 108460 92327 111490 92350
rect 108460 91320 108483 92327
rect 108277 90320 108483 91320
rect 108277 89343 108300 90320
rect 105270 89320 108300 89343
rect 108460 89343 108483 90320
rect 111467 91320 111490 92327
rect 111650 92327 114680 92350
rect 111650 91320 111673 92327
rect 111467 90320 111673 91320
rect 111467 89343 111490 90320
rect 108460 89320 111490 89343
rect 111650 89343 111673 90320
rect 114657 91320 114680 92327
rect 114840 92327 117870 92350
rect 114840 91320 114863 92327
rect 114657 90320 114863 91320
rect 114657 89343 114680 90320
rect 111650 89320 114680 89343
rect 114840 89343 114863 90320
rect 117847 91320 117870 92327
rect 118030 92327 121060 92350
rect 118030 91320 118053 92327
rect 117847 90320 118053 91320
rect 117847 89343 117870 90320
rect 114840 89320 117870 89343
rect 118030 89343 118053 90320
rect 121037 91320 121060 92327
rect 121220 92327 124250 92350
rect 121220 91320 121243 92327
rect 121037 90320 121243 91320
rect 121037 89343 121060 90320
rect 118030 89320 121060 89343
rect 121220 89343 121243 90320
rect 124227 91320 124250 92327
rect 124410 92327 127440 92350
rect 124410 91320 124433 92327
rect 124227 90320 124433 91320
rect 124227 89343 124250 90320
rect 121220 89320 124250 89343
rect 124410 89343 124433 90320
rect 127417 91320 127440 92327
rect 127600 92327 130630 92350
rect 127600 91320 127623 92327
rect 127417 90320 127623 91320
rect 127417 89343 127440 90320
rect 124410 89320 127440 89343
rect 127600 89343 127623 90320
rect 130607 91320 130630 92327
rect 130790 92327 133820 92350
rect 130790 91320 130813 92327
rect 130607 90320 130813 91320
rect 130607 89343 130630 90320
rect 127600 89320 130630 89343
rect 130790 89343 130813 90320
rect 133797 91320 133820 92327
rect 133980 92327 137010 92350
rect 133980 91320 134003 92327
rect 133797 90320 134003 91320
rect 133797 89343 133820 90320
rect 130790 89320 133820 89343
rect 133980 89343 134003 90320
rect 136987 91320 137010 92327
rect 136987 90320 137170 91320
rect 136987 89343 137010 90320
rect 133980 89320 137010 89343
rect 10570 89160 11570 89320
rect 13760 89160 14760 89320
rect 16950 89160 17950 89320
rect 20140 89160 21140 89320
rect 23330 89160 24330 89320
rect 26520 89160 27520 89320
rect 29710 89160 30710 89320
rect 32900 89160 33900 89320
rect 36090 89160 37090 89320
rect 39280 89160 40280 89320
rect 42470 89160 43470 89320
rect 45660 89160 46660 89320
rect 48850 89160 49850 89320
rect 52040 89160 53040 89320
rect 55230 89160 56230 89320
rect 58420 89160 59420 89320
rect 61610 89160 62610 89320
rect 64800 89160 65800 89320
rect 67990 89160 68990 89320
rect 71180 89160 72180 89320
rect 74370 89160 75370 89320
rect 77560 89160 78560 89320
rect 80750 89160 81750 89320
rect 83940 89160 84940 89320
rect 87130 89160 88130 89320
rect 90320 89160 91320 89320
rect 93510 89160 94510 89320
rect 96700 89160 97700 89320
rect 99890 89160 100890 89320
rect 103080 89160 104080 89320
rect 106270 89160 107270 89320
rect 109460 89160 110460 89320
rect 112650 89160 113650 89320
rect 115840 89160 116840 89320
rect 119030 89160 120030 89320
rect 122220 89160 123220 89320
rect 125410 89160 126410 89320
rect 128600 89160 129600 89320
rect 131790 89160 132790 89320
rect 134980 89160 135980 89320
rect 9570 89137 12600 89160
rect 9570 86153 9593 89137
rect 12577 88130 12600 89137
rect 12760 89137 15790 89160
rect 12760 88130 12783 89137
rect 12577 87130 12783 88130
rect 12577 86153 12600 87130
rect 9570 86130 12600 86153
rect 12760 86153 12783 87130
rect 15767 88130 15790 89137
rect 15950 89137 18980 89160
rect 15950 88130 15973 89137
rect 15767 87130 15973 88130
rect 15767 86153 15790 87130
rect 12760 86130 15790 86153
rect 15950 86153 15973 87130
rect 18957 88130 18980 89137
rect 19140 89137 22170 89160
rect 19140 88130 19163 89137
rect 18957 87130 19163 88130
rect 18957 86153 18980 87130
rect 15950 86130 18980 86153
rect 19140 86153 19163 87130
rect 22147 88130 22170 89137
rect 22330 89137 25360 89160
rect 22330 88130 22353 89137
rect 22147 87130 22353 88130
rect 22147 86153 22170 87130
rect 19140 86130 22170 86153
rect 22330 86153 22353 87130
rect 25337 88130 25360 89137
rect 25520 89137 28550 89160
rect 25520 88130 25543 89137
rect 25337 87130 25543 88130
rect 25337 86153 25360 87130
rect 22330 86130 25360 86153
rect 25520 86153 25543 87130
rect 28527 88130 28550 89137
rect 28710 89137 31740 89160
rect 28710 88130 28733 89137
rect 28527 87130 28733 88130
rect 28527 86153 28550 87130
rect 25520 86130 28550 86153
rect 28710 86153 28733 87130
rect 31717 88130 31740 89137
rect 31900 89137 34930 89160
rect 31900 88130 31923 89137
rect 31717 87130 31923 88130
rect 31717 86153 31740 87130
rect 28710 86130 31740 86153
rect 31900 86153 31923 87130
rect 34907 88130 34930 89137
rect 35090 89137 38120 89160
rect 35090 88130 35113 89137
rect 34907 87130 35113 88130
rect 34907 86153 34930 87130
rect 31900 86130 34930 86153
rect 35090 86153 35113 87130
rect 38097 88130 38120 89137
rect 38280 89137 41310 89160
rect 38280 88130 38303 89137
rect 38097 87130 38303 88130
rect 38097 86153 38120 87130
rect 35090 86130 38120 86153
rect 38280 86153 38303 87130
rect 41287 88130 41310 89137
rect 41470 89137 44500 89160
rect 41470 88130 41493 89137
rect 41287 87130 41493 88130
rect 41287 86153 41310 87130
rect 38280 86130 41310 86153
rect 41470 86153 41493 87130
rect 44477 88130 44500 89137
rect 44660 89137 47690 89160
rect 44660 88130 44683 89137
rect 44477 87130 44683 88130
rect 44477 86153 44500 87130
rect 41470 86130 44500 86153
rect 44660 86153 44683 87130
rect 47667 88130 47690 89137
rect 47850 89137 50880 89160
rect 47850 88130 47873 89137
rect 47667 87130 47873 88130
rect 47667 86153 47690 87130
rect 44660 86130 47690 86153
rect 47850 86153 47873 87130
rect 50857 88130 50880 89137
rect 51040 89137 54070 89160
rect 51040 88130 51063 89137
rect 50857 87130 51063 88130
rect 50857 86153 50880 87130
rect 47850 86130 50880 86153
rect 51040 86153 51063 87130
rect 54047 88130 54070 89137
rect 54230 89137 57260 89160
rect 54230 88130 54253 89137
rect 54047 87130 54253 88130
rect 54047 86153 54070 87130
rect 51040 86130 54070 86153
rect 54230 86153 54253 87130
rect 57237 88130 57260 89137
rect 57420 89137 60450 89160
rect 57420 88130 57443 89137
rect 57237 87130 57443 88130
rect 57237 86153 57260 87130
rect 54230 86130 57260 86153
rect 57420 86153 57443 87130
rect 60427 88130 60450 89137
rect 60610 89137 63640 89160
rect 60610 88130 60633 89137
rect 60427 87130 60633 88130
rect 60427 86153 60450 87130
rect 57420 86130 60450 86153
rect 60610 86153 60633 87130
rect 63617 88130 63640 89137
rect 63800 89137 66830 89160
rect 63800 88130 63823 89137
rect 63617 87130 63823 88130
rect 63617 86153 63640 87130
rect 60610 86130 63640 86153
rect 63800 86153 63823 87130
rect 66807 88130 66830 89137
rect 66990 89137 70020 89160
rect 66990 88130 67013 89137
rect 66807 87130 67013 88130
rect 66807 86153 66830 87130
rect 63800 86130 66830 86153
rect 66990 86153 67013 87130
rect 69997 88130 70020 89137
rect 70180 89137 73210 89160
rect 70180 88130 70203 89137
rect 69997 87130 70203 88130
rect 69997 86153 70020 87130
rect 66990 86130 70020 86153
rect 70180 86153 70203 87130
rect 73187 88130 73210 89137
rect 73370 89137 76400 89160
rect 73370 88130 73393 89137
rect 73187 87130 73393 88130
rect 73187 86153 73210 87130
rect 70180 86130 73210 86153
rect 73370 86153 73393 87130
rect 76377 88130 76400 89137
rect 76560 89137 79590 89160
rect 76560 88130 76583 89137
rect 76377 87130 76583 88130
rect 76377 86153 76400 87130
rect 73370 86130 76400 86153
rect 76560 86153 76583 87130
rect 79567 88130 79590 89137
rect 79750 89137 82780 89160
rect 79750 88130 79773 89137
rect 79567 87130 79773 88130
rect 79567 86153 79590 87130
rect 76560 86130 79590 86153
rect 79750 86153 79773 87130
rect 82757 88130 82780 89137
rect 82940 89137 85970 89160
rect 82940 88130 82963 89137
rect 82757 87130 82963 88130
rect 82757 86153 82780 87130
rect 79750 86130 82780 86153
rect 82940 86153 82963 87130
rect 85947 88130 85970 89137
rect 86130 89137 89160 89160
rect 86130 88130 86153 89137
rect 85947 87130 86153 88130
rect 85947 86153 85970 87130
rect 82940 86130 85970 86153
rect 86130 86153 86153 87130
rect 89137 88130 89160 89137
rect 89320 89137 92350 89160
rect 89320 88130 89343 89137
rect 89137 87130 89343 88130
rect 89137 86153 89160 87130
rect 86130 86130 89160 86153
rect 89320 86153 89343 87130
rect 92327 88130 92350 89137
rect 92510 89137 95540 89160
rect 92510 88130 92533 89137
rect 92327 87130 92533 88130
rect 92327 86153 92350 87130
rect 89320 86130 92350 86153
rect 92510 86153 92533 87130
rect 95517 88130 95540 89137
rect 95700 89137 98730 89160
rect 95700 88130 95723 89137
rect 95517 87130 95723 88130
rect 95517 86153 95540 87130
rect 92510 86130 95540 86153
rect 95700 86153 95723 87130
rect 98707 88130 98730 89137
rect 98890 89137 101920 89160
rect 98890 88130 98913 89137
rect 98707 87130 98913 88130
rect 98707 86153 98730 87130
rect 95700 86130 98730 86153
rect 98890 86153 98913 87130
rect 101897 88130 101920 89137
rect 102080 89137 105110 89160
rect 102080 88130 102103 89137
rect 101897 87130 102103 88130
rect 101897 86153 101920 87130
rect 98890 86130 101920 86153
rect 102080 86153 102103 87130
rect 105087 88130 105110 89137
rect 105270 89137 108300 89160
rect 105270 88130 105293 89137
rect 105087 87130 105293 88130
rect 105087 86153 105110 87130
rect 102080 86130 105110 86153
rect 105270 86153 105293 87130
rect 108277 88130 108300 89137
rect 108460 89137 111490 89160
rect 108460 88130 108483 89137
rect 108277 87130 108483 88130
rect 108277 86153 108300 87130
rect 105270 86130 108300 86153
rect 108460 86153 108483 87130
rect 111467 88130 111490 89137
rect 111650 89137 114680 89160
rect 111650 88130 111673 89137
rect 111467 87130 111673 88130
rect 111467 86153 111490 87130
rect 108460 86130 111490 86153
rect 111650 86153 111673 87130
rect 114657 88130 114680 89137
rect 114840 89137 117870 89160
rect 114840 88130 114863 89137
rect 114657 87130 114863 88130
rect 114657 86153 114680 87130
rect 111650 86130 114680 86153
rect 114840 86153 114863 87130
rect 117847 88130 117870 89137
rect 118030 89137 121060 89160
rect 118030 88130 118053 89137
rect 117847 87130 118053 88130
rect 117847 86153 117870 87130
rect 114840 86130 117870 86153
rect 118030 86153 118053 87130
rect 121037 88130 121060 89137
rect 121220 89137 124250 89160
rect 121220 88130 121243 89137
rect 121037 87130 121243 88130
rect 121037 86153 121060 87130
rect 118030 86130 121060 86153
rect 121220 86153 121243 87130
rect 124227 88130 124250 89137
rect 124410 89137 127440 89160
rect 124410 88130 124433 89137
rect 124227 87130 124433 88130
rect 124227 86153 124250 87130
rect 121220 86130 124250 86153
rect 124410 86153 124433 87130
rect 127417 88130 127440 89137
rect 127600 89137 130630 89160
rect 127600 88130 127623 89137
rect 127417 87130 127623 88130
rect 127417 86153 127440 87130
rect 124410 86130 127440 86153
rect 127600 86153 127623 87130
rect 130607 88130 130630 89137
rect 130790 89137 133820 89160
rect 130790 88130 130813 89137
rect 130607 87130 130813 88130
rect 130607 86153 130630 87130
rect 127600 86130 130630 86153
rect 130790 86153 130813 87130
rect 133797 88130 133820 89137
rect 133980 89137 137010 89160
rect 133980 88130 134003 89137
rect 133797 87130 134003 88130
rect 133797 86153 133820 87130
rect 130790 86130 133820 86153
rect 133980 86153 134003 87130
rect 136987 88130 137010 89137
rect 136987 87130 137170 88130
rect 136987 86153 137010 87130
rect 133980 86130 137010 86153
rect 10570 85970 11570 86130
rect 13760 85970 14760 86130
rect 16950 85970 17950 86130
rect 20140 85970 21140 86130
rect 23330 85970 24330 86130
rect 26520 85970 27520 86130
rect 29710 85970 30710 86130
rect 32900 85970 33900 86130
rect 36090 85970 37090 86130
rect 39280 85970 40280 86130
rect 42470 85970 43470 86130
rect 45660 85970 46660 86130
rect 48850 85970 49850 86130
rect 52040 85970 53040 86130
rect 55230 85970 56230 86130
rect 58420 85970 59420 86130
rect 61610 85970 62610 86130
rect 64800 85970 65800 86130
rect 67990 85970 68990 86130
rect 71180 85970 72180 86130
rect 74370 85970 75370 86130
rect 77560 85970 78560 86130
rect 80750 85970 81750 86130
rect 83940 85970 84940 86130
rect 87130 85970 88130 86130
rect 90320 85970 91320 86130
rect 93510 85970 94510 86130
rect 96700 85970 97700 86130
rect 99890 85970 100890 86130
rect 103080 85970 104080 86130
rect 106270 85970 107270 86130
rect 109460 85970 110460 86130
rect 112650 85970 113650 86130
rect 115840 85970 116840 86130
rect 119030 85970 120030 86130
rect 122220 85970 123220 86130
rect 125410 85970 126410 86130
rect 128600 85970 129600 86130
rect 131790 85970 132790 86130
rect 134980 85970 135980 86130
rect 9570 85947 12600 85970
rect 9570 82963 9593 85947
rect 12577 84940 12600 85947
rect 12760 85947 15790 85970
rect 12760 84940 12783 85947
rect 12577 83940 12783 84940
rect 12577 82963 12600 83940
rect 9570 82940 12600 82963
rect 12760 82963 12783 83940
rect 15767 84940 15790 85947
rect 15950 85947 18980 85970
rect 15950 84940 15973 85947
rect 15767 83940 15973 84940
rect 15767 82963 15790 83940
rect 12760 82940 15790 82963
rect 15950 82963 15973 83940
rect 18957 84940 18980 85947
rect 19140 85947 22170 85970
rect 19140 84940 19163 85947
rect 18957 83940 19163 84940
rect 18957 82963 18980 83940
rect 15950 82940 18980 82963
rect 19140 82963 19163 83940
rect 22147 84940 22170 85947
rect 22330 85947 25360 85970
rect 22330 84940 22353 85947
rect 22147 83940 22353 84940
rect 22147 82963 22170 83940
rect 19140 82940 22170 82963
rect 22330 82963 22353 83940
rect 25337 84940 25360 85947
rect 25520 85947 28550 85970
rect 25520 84940 25543 85947
rect 25337 83940 25543 84940
rect 25337 82963 25360 83940
rect 22330 82940 25360 82963
rect 25520 82963 25543 83940
rect 28527 84940 28550 85947
rect 28710 85947 31740 85970
rect 28710 84940 28733 85947
rect 28527 83940 28733 84940
rect 28527 82963 28550 83940
rect 25520 82940 28550 82963
rect 28710 82963 28733 83940
rect 31717 84940 31740 85947
rect 31900 85947 34930 85970
rect 31900 84940 31923 85947
rect 31717 83940 31923 84940
rect 31717 82963 31740 83940
rect 28710 82940 31740 82963
rect 31900 82963 31923 83940
rect 34907 84940 34930 85947
rect 35090 85947 38120 85970
rect 35090 84940 35113 85947
rect 34907 83940 35113 84940
rect 34907 82963 34930 83940
rect 31900 82940 34930 82963
rect 35090 82963 35113 83940
rect 38097 84940 38120 85947
rect 38280 85947 41310 85970
rect 38280 84940 38303 85947
rect 38097 83940 38303 84940
rect 38097 82963 38120 83940
rect 35090 82940 38120 82963
rect 38280 82963 38303 83940
rect 41287 84940 41310 85947
rect 41470 85947 44500 85970
rect 41470 84940 41493 85947
rect 41287 83940 41493 84940
rect 41287 82963 41310 83940
rect 38280 82940 41310 82963
rect 41470 82963 41493 83940
rect 44477 84940 44500 85947
rect 44660 85947 47690 85970
rect 44660 84940 44683 85947
rect 44477 83940 44683 84940
rect 44477 82963 44500 83940
rect 41470 82940 44500 82963
rect 44660 82963 44683 83940
rect 47667 84940 47690 85947
rect 47850 85947 50880 85970
rect 47850 84940 47873 85947
rect 47667 83940 47873 84940
rect 47667 82963 47690 83940
rect 44660 82940 47690 82963
rect 47850 82963 47873 83940
rect 50857 84940 50880 85947
rect 51040 85947 54070 85970
rect 51040 84940 51063 85947
rect 50857 83940 51063 84940
rect 50857 82963 50880 83940
rect 47850 82940 50880 82963
rect 51040 82963 51063 83940
rect 54047 84940 54070 85947
rect 54230 85947 57260 85970
rect 54230 84940 54253 85947
rect 54047 83940 54253 84940
rect 54047 82963 54070 83940
rect 51040 82940 54070 82963
rect 54230 82963 54253 83940
rect 57237 84940 57260 85947
rect 57420 85947 60450 85970
rect 57420 84940 57443 85947
rect 57237 83940 57443 84940
rect 57237 82963 57260 83940
rect 54230 82940 57260 82963
rect 57420 82963 57443 83940
rect 60427 84940 60450 85947
rect 60610 85947 63640 85970
rect 60610 84940 60633 85947
rect 60427 83940 60633 84940
rect 60427 82963 60450 83940
rect 57420 82940 60450 82963
rect 60610 82963 60633 83940
rect 63617 84940 63640 85947
rect 63800 85947 66830 85970
rect 63800 84940 63823 85947
rect 63617 83940 63823 84940
rect 63617 82963 63640 83940
rect 60610 82940 63640 82963
rect 63800 82963 63823 83940
rect 66807 84940 66830 85947
rect 66990 85947 70020 85970
rect 66990 84940 67013 85947
rect 66807 83940 67013 84940
rect 66807 82963 66830 83940
rect 63800 82940 66830 82963
rect 66990 82963 67013 83940
rect 69997 84940 70020 85947
rect 70180 85947 73210 85970
rect 70180 84940 70203 85947
rect 69997 83940 70203 84940
rect 69997 82963 70020 83940
rect 66990 82940 70020 82963
rect 70180 82963 70203 83940
rect 73187 84940 73210 85947
rect 73370 85947 76400 85970
rect 73370 84940 73393 85947
rect 73187 83940 73393 84940
rect 73187 82963 73210 83940
rect 70180 82940 73210 82963
rect 73370 82963 73393 83940
rect 76377 84940 76400 85947
rect 76560 85947 79590 85970
rect 76560 84940 76583 85947
rect 76377 83940 76583 84940
rect 76377 82963 76400 83940
rect 73370 82940 76400 82963
rect 76560 82963 76583 83940
rect 79567 84940 79590 85947
rect 79750 85947 82780 85970
rect 79750 84940 79773 85947
rect 79567 83940 79773 84940
rect 79567 82963 79590 83940
rect 76560 82940 79590 82963
rect 79750 82963 79773 83940
rect 82757 84940 82780 85947
rect 82940 85947 85970 85970
rect 82940 84940 82963 85947
rect 82757 83940 82963 84940
rect 82757 82963 82780 83940
rect 79750 82940 82780 82963
rect 82940 82963 82963 83940
rect 85947 84940 85970 85947
rect 86130 85947 89160 85970
rect 86130 84940 86153 85947
rect 85947 83940 86153 84940
rect 85947 82963 85970 83940
rect 82940 82940 85970 82963
rect 86130 82963 86153 83940
rect 89137 84940 89160 85947
rect 89320 85947 92350 85970
rect 89320 84940 89343 85947
rect 89137 83940 89343 84940
rect 89137 82963 89160 83940
rect 86130 82940 89160 82963
rect 89320 82963 89343 83940
rect 92327 84940 92350 85947
rect 92510 85947 95540 85970
rect 92510 84940 92533 85947
rect 92327 83940 92533 84940
rect 92327 82963 92350 83940
rect 89320 82940 92350 82963
rect 92510 82963 92533 83940
rect 95517 84940 95540 85947
rect 95700 85947 98730 85970
rect 95700 84940 95723 85947
rect 95517 83940 95723 84940
rect 95517 82963 95540 83940
rect 92510 82940 95540 82963
rect 95700 82963 95723 83940
rect 98707 84940 98730 85947
rect 98890 85947 101920 85970
rect 98890 84940 98913 85947
rect 98707 83940 98913 84940
rect 98707 82963 98730 83940
rect 95700 82940 98730 82963
rect 98890 82963 98913 83940
rect 101897 84940 101920 85947
rect 102080 85947 105110 85970
rect 102080 84940 102103 85947
rect 101897 83940 102103 84940
rect 101897 82963 101920 83940
rect 98890 82940 101920 82963
rect 102080 82963 102103 83940
rect 105087 84940 105110 85947
rect 105270 85947 108300 85970
rect 105270 84940 105293 85947
rect 105087 83940 105293 84940
rect 105087 82963 105110 83940
rect 102080 82940 105110 82963
rect 105270 82963 105293 83940
rect 108277 84940 108300 85947
rect 108460 85947 111490 85970
rect 108460 84940 108483 85947
rect 108277 83940 108483 84940
rect 108277 82963 108300 83940
rect 105270 82940 108300 82963
rect 108460 82963 108483 83940
rect 111467 84940 111490 85947
rect 111650 85947 114680 85970
rect 111650 84940 111673 85947
rect 111467 83940 111673 84940
rect 111467 82963 111490 83940
rect 108460 82940 111490 82963
rect 111650 82963 111673 83940
rect 114657 84940 114680 85947
rect 114840 85947 117870 85970
rect 114840 84940 114863 85947
rect 114657 83940 114863 84940
rect 114657 82963 114680 83940
rect 111650 82940 114680 82963
rect 114840 82963 114863 83940
rect 117847 84940 117870 85947
rect 118030 85947 121060 85970
rect 118030 84940 118053 85947
rect 117847 83940 118053 84940
rect 117847 82963 117870 83940
rect 114840 82940 117870 82963
rect 118030 82963 118053 83940
rect 121037 84940 121060 85947
rect 121220 85947 124250 85970
rect 121220 84940 121243 85947
rect 121037 83940 121243 84940
rect 121037 82963 121060 83940
rect 118030 82940 121060 82963
rect 121220 82963 121243 83940
rect 124227 84940 124250 85947
rect 124410 85947 127440 85970
rect 124410 84940 124433 85947
rect 124227 83940 124433 84940
rect 124227 82963 124250 83940
rect 121220 82940 124250 82963
rect 124410 82963 124433 83940
rect 127417 84940 127440 85947
rect 127600 85947 130630 85970
rect 127600 84940 127623 85947
rect 127417 83940 127623 84940
rect 127417 82963 127440 83940
rect 124410 82940 127440 82963
rect 127600 82963 127623 83940
rect 130607 84940 130630 85947
rect 130790 85947 133820 85970
rect 130790 84940 130813 85947
rect 130607 83940 130813 84940
rect 130607 82963 130630 83940
rect 127600 82940 130630 82963
rect 130790 82963 130813 83940
rect 133797 84940 133820 85947
rect 133980 85947 137010 85970
rect 133980 84940 134003 85947
rect 133797 83940 134003 84940
rect 133797 82963 133820 83940
rect 130790 82940 133820 82963
rect 133980 82963 134003 83940
rect 136987 84940 137010 85947
rect 136987 83940 137170 84940
rect 136987 82963 137010 83940
rect 133980 82940 137010 82963
rect 10570 82780 11570 82940
rect 13760 82780 14760 82940
rect 16950 82780 17950 82940
rect 20140 82780 21140 82940
rect 23330 82780 24330 82940
rect 26520 82780 27520 82940
rect 29710 82780 30710 82940
rect 32900 82780 33900 82940
rect 36090 82780 37090 82940
rect 39280 82780 40280 82940
rect 42470 82780 43470 82940
rect 45660 82780 46660 82940
rect 48850 82780 49850 82940
rect 52040 82780 53040 82940
rect 55230 82780 56230 82940
rect 58420 82780 59420 82940
rect 61610 82780 62610 82940
rect 64800 82780 65800 82940
rect 67990 82780 68990 82940
rect 71180 82780 72180 82940
rect 74370 82780 75370 82940
rect 77560 82780 78560 82940
rect 80750 82780 81750 82940
rect 83940 82780 84940 82940
rect 87130 82780 88130 82940
rect 90320 82780 91320 82940
rect 93510 82780 94510 82940
rect 96700 82780 97700 82940
rect 99890 82780 100890 82940
rect 103080 82780 104080 82940
rect 106270 82780 107270 82940
rect 109460 82780 110460 82940
rect 112650 82780 113650 82940
rect 115840 82780 116840 82940
rect 119030 82780 120030 82940
rect 122220 82780 123220 82940
rect 125410 82780 126410 82940
rect 128600 82780 129600 82940
rect 131790 82780 132790 82940
rect 134980 82780 135980 82940
rect 0 79789 9370 79839
rect 9570 82757 12600 82780
rect 9570 79773 9593 82757
rect 12577 81750 12600 82757
rect 12760 82757 15790 82780
rect 12760 81750 12783 82757
rect 12577 80750 12783 81750
rect 12577 79773 12600 80750
rect 9570 79750 12600 79773
rect 12760 79773 12783 80750
rect 15767 81750 15790 82757
rect 15950 82757 18980 82780
rect 15950 81750 15973 82757
rect 15767 80750 15973 81750
rect 15767 79773 15790 80750
rect 12760 79750 15790 79773
rect 15950 79773 15973 80750
rect 18957 81750 18980 82757
rect 19140 82757 22170 82780
rect 19140 81750 19163 82757
rect 18957 80750 19163 81750
rect 18957 79773 18980 80750
rect 15950 79750 18980 79773
rect 19140 79773 19163 80750
rect 22147 81750 22170 82757
rect 22330 82757 25360 82780
rect 22330 81750 22353 82757
rect 22147 80750 22353 81750
rect 22147 79773 22170 80750
rect 19140 79750 22170 79773
rect 22330 79773 22353 80750
rect 25337 81750 25360 82757
rect 25520 82757 28550 82780
rect 25520 81750 25543 82757
rect 25337 80750 25543 81750
rect 25337 79773 25360 80750
rect 22330 79750 25360 79773
rect 25520 79773 25543 80750
rect 28527 81750 28550 82757
rect 28710 82757 31740 82780
rect 28710 81750 28733 82757
rect 28527 80750 28733 81750
rect 28527 79773 28550 80750
rect 25520 79750 28550 79773
rect 28710 79773 28733 80750
rect 31717 81750 31740 82757
rect 31900 82757 34930 82780
rect 31900 81750 31923 82757
rect 31717 80750 31923 81750
rect 31717 79773 31740 80750
rect 28710 79750 31740 79773
rect 31900 79773 31923 80750
rect 34907 81750 34930 82757
rect 35090 82757 38120 82780
rect 35090 81750 35113 82757
rect 34907 80750 35113 81750
rect 34907 79773 34930 80750
rect 31900 79750 34930 79773
rect 35090 79773 35113 80750
rect 38097 81750 38120 82757
rect 38280 82757 41310 82780
rect 38280 81750 38303 82757
rect 38097 80750 38303 81750
rect 38097 79773 38120 80750
rect 35090 79750 38120 79773
rect 38280 79773 38303 80750
rect 41287 81750 41310 82757
rect 41470 82757 44500 82780
rect 41470 81750 41493 82757
rect 41287 80750 41493 81750
rect 41287 79773 41310 80750
rect 38280 79750 41310 79773
rect 41470 79773 41493 80750
rect 44477 81750 44500 82757
rect 44660 82757 47690 82780
rect 44660 81750 44683 82757
rect 44477 80750 44683 81750
rect 44477 79773 44500 80750
rect 41470 79750 44500 79773
rect 44660 79773 44683 80750
rect 47667 81750 47690 82757
rect 47850 82757 50880 82780
rect 47850 81750 47873 82757
rect 47667 80750 47873 81750
rect 47667 79773 47690 80750
rect 44660 79750 47690 79773
rect 47850 79773 47873 80750
rect 50857 81750 50880 82757
rect 51040 82757 54070 82780
rect 51040 81750 51063 82757
rect 50857 80750 51063 81750
rect 50857 79773 50880 80750
rect 47850 79750 50880 79773
rect 51040 79773 51063 80750
rect 54047 81750 54070 82757
rect 54230 82757 57260 82780
rect 54230 81750 54253 82757
rect 54047 80750 54253 81750
rect 54047 79773 54070 80750
rect 51040 79750 54070 79773
rect 54230 79773 54253 80750
rect 57237 81750 57260 82757
rect 57420 82757 60450 82780
rect 57420 81750 57443 82757
rect 57237 80750 57443 81750
rect 57237 79773 57260 80750
rect 54230 79750 57260 79773
rect 57420 79773 57443 80750
rect 60427 81750 60450 82757
rect 60610 82757 63640 82780
rect 60610 81750 60633 82757
rect 60427 80750 60633 81750
rect 60427 79773 60450 80750
rect 57420 79750 60450 79773
rect 60610 79773 60633 80750
rect 63617 81750 63640 82757
rect 63800 82757 66830 82780
rect 63800 81750 63823 82757
rect 63617 80750 63823 81750
rect 63617 79773 63640 80750
rect 60610 79750 63640 79773
rect 63800 79773 63823 80750
rect 66807 81750 66830 82757
rect 66990 82757 70020 82780
rect 66990 81750 67013 82757
rect 66807 80750 67013 81750
rect 66807 79773 66830 80750
rect 63800 79750 66830 79773
rect 66990 79773 67013 80750
rect 69997 81750 70020 82757
rect 70180 82757 73210 82780
rect 70180 81750 70203 82757
rect 69997 80750 70203 81750
rect 69997 79773 70020 80750
rect 66990 79750 70020 79773
rect 70180 79773 70203 80750
rect 73187 81750 73210 82757
rect 73370 82757 76400 82780
rect 73370 81750 73393 82757
rect 73187 80750 73393 81750
rect 73187 79773 73210 80750
rect 70180 79750 73210 79773
rect 73370 79773 73393 80750
rect 76377 81750 76400 82757
rect 76560 82757 79590 82780
rect 76560 81750 76583 82757
rect 76377 80750 76583 81750
rect 76377 79773 76400 80750
rect 73370 79750 76400 79773
rect 76560 79773 76583 80750
rect 79567 81750 79590 82757
rect 79750 82757 82780 82780
rect 79750 81750 79773 82757
rect 79567 80750 79773 81750
rect 79567 79773 79590 80750
rect 76560 79750 79590 79773
rect 79750 79773 79773 80750
rect 82757 81750 82780 82757
rect 82940 82757 85970 82780
rect 82940 81750 82963 82757
rect 82757 80750 82963 81750
rect 82757 79773 82780 80750
rect 79750 79750 82780 79773
rect 82940 79773 82963 80750
rect 85947 81750 85970 82757
rect 86130 82757 89160 82780
rect 86130 81750 86153 82757
rect 85947 80750 86153 81750
rect 85947 79773 85970 80750
rect 82940 79750 85970 79773
rect 86130 79773 86153 80750
rect 89137 81750 89160 82757
rect 89320 82757 92350 82780
rect 89320 81750 89343 82757
rect 89137 80750 89343 81750
rect 89137 79773 89160 80750
rect 86130 79750 89160 79773
rect 89320 79773 89343 80750
rect 92327 81750 92350 82757
rect 92510 82757 95540 82780
rect 92510 81750 92533 82757
rect 92327 80750 92533 81750
rect 92327 79773 92350 80750
rect 89320 79750 92350 79773
rect 92510 79773 92533 80750
rect 95517 81750 95540 82757
rect 95700 82757 98730 82780
rect 95700 81750 95723 82757
rect 95517 80750 95723 81750
rect 95517 79773 95540 80750
rect 92510 79750 95540 79773
rect 95700 79773 95723 80750
rect 98707 81750 98730 82757
rect 98890 82757 101920 82780
rect 98890 81750 98913 82757
rect 98707 80750 98913 81750
rect 98707 79773 98730 80750
rect 95700 79750 98730 79773
rect 98890 79773 98913 80750
rect 101897 81750 101920 82757
rect 102080 82757 105110 82780
rect 102080 81750 102103 82757
rect 101897 80750 102103 81750
rect 101897 79773 101920 80750
rect 98890 79750 101920 79773
rect 102080 79773 102103 80750
rect 105087 81750 105110 82757
rect 105270 82757 108300 82780
rect 105270 81750 105293 82757
rect 105087 80750 105293 81750
rect 105087 79773 105110 80750
rect 102080 79750 105110 79773
rect 105270 79773 105293 80750
rect 108277 81750 108300 82757
rect 108460 82757 111490 82780
rect 108460 81750 108483 82757
rect 108277 80750 108483 81750
rect 108277 79773 108300 80750
rect 105270 79750 108300 79773
rect 108460 79773 108483 80750
rect 111467 81750 111490 82757
rect 111650 82757 114680 82780
rect 111650 81750 111673 82757
rect 111467 80750 111673 81750
rect 111467 79773 111490 80750
rect 108460 79750 111490 79773
rect 111650 79773 111673 80750
rect 114657 81750 114680 82757
rect 114840 82757 117870 82780
rect 114840 81750 114863 82757
rect 114657 80750 114863 81750
rect 114657 79773 114680 80750
rect 111650 79750 114680 79773
rect 114840 79773 114863 80750
rect 117847 81750 117870 82757
rect 118030 82757 121060 82780
rect 118030 81750 118053 82757
rect 117847 80750 118053 81750
rect 117847 79773 117870 80750
rect 114840 79750 117870 79773
rect 118030 79773 118053 80750
rect 121037 81750 121060 82757
rect 121220 82757 124250 82780
rect 121220 81750 121243 82757
rect 121037 80750 121243 81750
rect 121037 79773 121060 80750
rect 118030 79750 121060 79773
rect 121220 79773 121243 80750
rect 124227 81750 124250 82757
rect 124410 82757 127440 82780
rect 124410 81750 124433 82757
rect 124227 80750 124433 81750
rect 124227 79773 124250 80750
rect 121220 79750 124250 79773
rect 124410 79773 124433 80750
rect 127417 81750 127440 82757
rect 127600 82757 130630 82780
rect 127600 81750 127623 82757
rect 127417 80750 127623 81750
rect 127417 79773 127440 80750
rect 124410 79750 127440 79773
rect 127600 79773 127623 80750
rect 130607 81750 130630 82757
rect 130790 82757 133820 82780
rect 130790 81750 130813 82757
rect 130607 80750 130813 81750
rect 130607 79773 130630 80750
rect 127600 79750 130630 79773
rect 130790 79773 130813 80750
rect 133797 81750 133820 82757
rect 133980 82757 137010 82780
rect 133980 81750 134003 82757
rect 133797 80750 134003 81750
rect 133797 79773 133820 80750
rect 130790 79750 133820 79773
rect 133980 79773 134003 80750
rect 136987 81750 137010 82757
rect 136987 80750 137170 81750
rect 136987 79773 137010 80750
rect 133980 79750 137010 79773
rect 10570 79590 11570 79750
rect 13760 79590 14760 79750
rect 16950 79590 17950 79750
rect 20140 79590 21140 79750
rect 23330 79590 24330 79750
rect 26520 79590 27520 79750
rect 29710 79590 30710 79750
rect 32900 79590 33900 79750
rect 36090 79590 37090 79750
rect 39280 79590 40280 79750
rect 42470 79590 43470 79750
rect 45660 79590 46660 79750
rect 48850 79590 49850 79750
rect 52040 79590 53040 79750
rect 55230 79590 56230 79750
rect 58420 79590 59420 79750
rect 61610 79590 62610 79750
rect 64800 79590 65800 79750
rect 67990 79590 68990 79750
rect 71180 79590 72180 79750
rect 74370 79590 75370 79750
rect 77560 79590 78560 79750
rect 80750 79590 81750 79750
rect 83940 79590 84940 79750
rect 87130 79590 88130 79750
rect 90320 79590 91320 79750
rect 93510 79590 94510 79750
rect 96700 79590 97700 79750
rect 99890 79590 100890 79750
rect 103080 79590 104080 79750
rect 106270 79590 107270 79750
rect 109460 79590 110460 79750
rect 112650 79590 113650 79750
rect 115840 79590 116840 79750
rect 119030 79590 120030 79750
rect 122220 79590 123220 79750
rect 125410 79590 126410 79750
rect 128600 79590 129600 79750
rect 131790 79590 132790 79750
rect 134980 79590 135980 79750
rect 0 79567 3030 79589
rect 0 76583 23 79567
rect 3007 78560 3030 79567
rect 3190 79567 6220 79589
rect 3190 78560 3213 79567
rect 3007 77560 3213 78560
rect 3007 76583 3030 77560
rect 0 76560 3030 76583
rect 3190 76583 3213 77560
rect 6197 78560 6220 79567
rect 6380 79567 9410 79589
rect 6380 78560 6403 79567
rect 6197 77560 6403 78560
rect 6197 76583 6220 77560
rect 3190 76560 6220 76583
rect 6380 76583 6403 77560
rect 9387 78560 9410 79567
rect 9570 79567 12600 79590
rect 9570 78560 9593 79567
rect 9387 77560 9593 78560
rect 9387 76583 9410 77560
rect 6380 76560 9410 76583
rect 9570 76583 9593 77560
rect 12577 78560 12600 79567
rect 12760 79567 15790 79590
rect 12760 78560 12783 79567
rect 12577 77560 12783 78560
rect 12577 76583 12600 77560
rect 9570 76560 12600 76583
rect 12760 76583 12783 77560
rect 15767 78560 15790 79567
rect 15950 79567 18980 79590
rect 15950 78560 15973 79567
rect 15767 77560 15973 78560
rect 15767 76583 15790 77560
rect 12760 76560 15790 76583
rect 15950 76583 15973 77560
rect 18957 78560 18980 79567
rect 19140 79567 22170 79590
rect 19140 78560 19163 79567
rect 18957 77560 19163 78560
rect 18957 76583 18980 77560
rect 15950 76560 18980 76583
rect 19140 76583 19163 77560
rect 22147 78560 22170 79567
rect 22330 79567 25360 79590
rect 22330 78560 22353 79567
rect 22147 77560 22353 78560
rect 22147 76583 22170 77560
rect 19140 76560 22170 76583
rect 22330 76583 22353 77560
rect 25337 78560 25360 79567
rect 25520 79567 28550 79590
rect 25520 78560 25543 79567
rect 25337 77560 25543 78560
rect 25337 76583 25360 77560
rect 22330 76560 25360 76583
rect 25520 76583 25543 77560
rect 28527 78560 28550 79567
rect 28710 79567 31740 79590
rect 28710 78560 28733 79567
rect 28527 77560 28733 78560
rect 28527 76583 28550 77560
rect 25520 76560 28550 76583
rect 28710 76583 28733 77560
rect 31717 78560 31740 79567
rect 31900 79567 34930 79590
rect 31900 78560 31923 79567
rect 31717 77560 31923 78560
rect 31717 76583 31740 77560
rect 28710 76560 31740 76583
rect 31900 76583 31923 77560
rect 34907 78560 34930 79567
rect 35090 79567 38120 79590
rect 35090 78560 35113 79567
rect 34907 77560 35113 78560
rect 34907 76583 34930 77560
rect 31900 76560 34930 76583
rect 35090 76583 35113 77560
rect 38097 78560 38120 79567
rect 38280 79567 41310 79590
rect 38280 78560 38303 79567
rect 38097 77560 38303 78560
rect 38097 76583 38120 77560
rect 35090 76560 38120 76583
rect 38280 76583 38303 77560
rect 41287 78560 41310 79567
rect 41470 79567 44500 79590
rect 41470 78560 41493 79567
rect 41287 77560 41493 78560
rect 41287 76583 41310 77560
rect 38280 76560 41310 76583
rect 41470 76583 41493 77560
rect 44477 78560 44500 79567
rect 44660 79567 47690 79590
rect 44660 78560 44683 79567
rect 44477 77560 44683 78560
rect 44477 76583 44500 77560
rect 41470 76560 44500 76583
rect 44660 76583 44683 77560
rect 47667 78560 47690 79567
rect 47850 79567 50880 79590
rect 47850 78560 47873 79567
rect 47667 77560 47873 78560
rect 47667 76583 47690 77560
rect 44660 76560 47690 76583
rect 47850 76583 47873 77560
rect 50857 78560 50880 79567
rect 51040 79567 54070 79590
rect 51040 78560 51063 79567
rect 50857 77560 51063 78560
rect 50857 76583 50880 77560
rect 47850 76560 50880 76583
rect 51040 76583 51063 77560
rect 54047 78560 54070 79567
rect 54230 79567 57260 79590
rect 54230 78560 54253 79567
rect 54047 77560 54253 78560
rect 54047 76583 54070 77560
rect 51040 76560 54070 76583
rect 54230 76583 54253 77560
rect 57237 78560 57260 79567
rect 57420 79567 60450 79590
rect 57420 78560 57443 79567
rect 57237 77560 57443 78560
rect 57237 76583 57260 77560
rect 54230 76560 57260 76583
rect 57420 76583 57443 77560
rect 60427 78560 60450 79567
rect 60610 79567 63640 79590
rect 60610 78560 60633 79567
rect 60427 77560 60633 78560
rect 60427 76583 60450 77560
rect 57420 76560 60450 76583
rect 60610 76583 60633 77560
rect 63617 78560 63640 79567
rect 63800 79567 66830 79590
rect 63800 78560 63823 79567
rect 63617 77560 63823 78560
rect 63617 76583 63640 77560
rect 60610 76560 63640 76583
rect 63800 76583 63823 77560
rect 66807 78560 66830 79567
rect 66990 79567 70020 79590
rect 66990 78560 67013 79567
rect 66807 77560 67013 78560
rect 66807 76583 66830 77560
rect 63800 76560 66830 76583
rect 66990 76583 67013 77560
rect 69997 78560 70020 79567
rect 70180 79567 73210 79590
rect 70180 78560 70203 79567
rect 69997 77560 70203 78560
rect 69997 76583 70020 77560
rect 66990 76560 70020 76583
rect 70180 76583 70203 77560
rect 73187 78560 73210 79567
rect 73370 79567 76400 79590
rect 73370 78560 73393 79567
rect 73187 77560 73393 78560
rect 73187 76583 73210 77560
rect 70180 76560 73210 76583
rect 73370 76583 73393 77560
rect 76377 78560 76400 79567
rect 76560 79567 79590 79590
rect 76560 78560 76583 79567
rect 76377 77560 76583 78560
rect 76377 76583 76400 77560
rect 73370 76560 76400 76583
rect 76560 76583 76583 77560
rect 79567 78560 79590 79567
rect 79750 79567 82780 79590
rect 79750 78560 79773 79567
rect 79567 77560 79773 78560
rect 79567 76583 79590 77560
rect 76560 76560 79590 76583
rect 79750 76583 79773 77560
rect 82757 78560 82780 79567
rect 82940 79567 85970 79590
rect 82940 78560 82963 79567
rect 82757 77560 82963 78560
rect 82757 76583 82780 77560
rect 79750 76560 82780 76583
rect 82940 76583 82963 77560
rect 85947 78560 85970 79567
rect 86130 79567 89160 79590
rect 86130 78560 86153 79567
rect 85947 77560 86153 78560
rect 85947 76583 85970 77560
rect 82940 76560 85970 76583
rect 86130 76583 86153 77560
rect 89137 78560 89160 79567
rect 89320 79567 92350 79590
rect 89320 78560 89343 79567
rect 89137 77560 89343 78560
rect 89137 76583 89160 77560
rect 86130 76560 89160 76583
rect 89320 76583 89343 77560
rect 92327 78560 92350 79567
rect 92510 79567 95540 79590
rect 92510 78560 92533 79567
rect 92327 77560 92533 78560
rect 92327 76583 92350 77560
rect 89320 76560 92350 76583
rect 92510 76583 92533 77560
rect 95517 78560 95540 79567
rect 95700 79567 98730 79590
rect 95700 78560 95723 79567
rect 95517 77560 95723 78560
rect 95517 76583 95540 77560
rect 92510 76560 95540 76583
rect 95700 76583 95723 77560
rect 98707 78560 98730 79567
rect 98890 79567 101920 79590
rect 98890 78560 98913 79567
rect 98707 77560 98913 78560
rect 98707 76583 98730 77560
rect 95700 76560 98730 76583
rect 98890 76583 98913 77560
rect 101897 78560 101920 79567
rect 102080 79567 105110 79590
rect 102080 78560 102103 79567
rect 101897 77560 102103 78560
rect 101897 76583 101920 77560
rect 98890 76560 101920 76583
rect 102080 76583 102103 77560
rect 105087 78560 105110 79567
rect 105270 79567 108300 79590
rect 105270 78560 105293 79567
rect 105087 77560 105293 78560
rect 105087 76583 105110 77560
rect 102080 76560 105110 76583
rect 105270 76583 105293 77560
rect 108277 78560 108300 79567
rect 108460 79567 111490 79590
rect 108460 78560 108483 79567
rect 108277 77560 108483 78560
rect 108277 76583 108300 77560
rect 105270 76560 108300 76583
rect 108460 76583 108483 77560
rect 111467 78560 111490 79567
rect 111650 79567 114680 79590
rect 111650 78560 111673 79567
rect 111467 77560 111673 78560
rect 111467 76583 111490 77560
rect 108460 76560 111490 76583
rect 111650 76583 111673 77560
rect 114657 78560 114680 79567
rect 114840 79567 117870 79590
rect 114840 78560 114863 79567
rect 114657 77560 114863 78560
rect 114657 76583 114680 77560
rect 111650 76560 114680 76583
rect 114840 76583 114863 77560
rect 117847 78560 117870 79567
rect 118030 79567 121060 79590
rect 118030 78560 118053 79567
rect 117847 77560 118053 78560
rect 117847 76583 117870 77560
rect 114840 76560 117870 76583
rect 118030 76583 118053 77560
rect 121037 78560 121060 79567
rect 121220 79567 124250 79590
rect 121220 78560 121243 79567
rect 121037 77560 121243 78560
rect 121037 76583 121060 77560
rect 118030 76560 121060 76583
rect 121220 76583 121243 77560
rect 124227 78560 124250 79567
rect 124410 79567 127440 79590
rect 124410 78560 124433 79567
rect 124227 77560 124433 78560
rect 124227 76583 124250 77560
rect 121220 76560 124250 76583
rect 124410 76583 124433 77560
rect 127417 78560 127440 79567
rect 127600 79567 130630 79590
rect 127600 78560 127623 79567
rect 127417 77560 127623 78560
rect 127417 76583 127440 77560
rect 124410 76560 127440 76583
rect 127600 76583 127623 77560
rect 130607 78560 130630 79567
rect 130790 79567 133820 79590
rect 130790 78560 130813 79567
rect 130607 77560 130813 78560
rect 130607 76583 130630 77560
rect 127600 76560 130630 76583
rect 130790 76583 130813 77560
rect 133797 78560 133820 79567
rect 133980 79567 137010 79590
rect 133980 78560 134003 79567
rect 133797 77560 134003 78560
rect 133797 76583 133820 77560
rect 130790 76560 133820 76583
rect 133980 76583 134003 77560
rect 136987 78560 137010 79567
rect 136987 77560 137170 78560
rect 136987 76583 137010 77560
rect 133980 76560 137010 76583
rect 1000 76400 2000 76560
rect 4190 76400 5190 76560
rect 7380 76400 8380 76560
rect 10570 76400 11570 76560
rect 13760 76400 14760 76560
rect 16950 76400 17950 76560
rect 20140 76400 21140 76560
rect 23330 76400 24330 76560
rect 26520 76400 27520 76560
rect 29710 76400 30710 76560
rect 32900 76400 33900 76560
rect 36090 76400 37090 76560
rect 39280 76400 40280 76560
rect 42470 76400 43470 76560
rect 45660 76400 46660 76560
rect 48850 76400 49850 76560
rect 52040 76400 53040 76560
rect 55230 76400 56230 76560
rect 58420 76400 59420 76560
rect 61610 76400 62610 76560
rect 64800 76400 65800 76560
rect 67990 76400 68990 76560
rect 71180 76400 72180 76560
rect 74370 76400 75370 76560
rect 77560 76400 78560 76560
rect 80750 76400 81750 76560
rect 83940 76400 84940 76560
rect 87130 76400 88130 76560
rect 90320 76400 91320 76560
rect 93510 76400 94510 76560
rect 96700 76400 97700 76560
rect 99890 76400 100890 76560
rect 103080 76400 104080 76560
rect 106270 76400 107270 76560
rect 109460 76400 110460 76560
rect 112650 76400 113650 76560
rect 115840 76400 116840 76560
rect 119030 76400 120030 76560
rect 122220 76400 123220 76560
rect 125410 76400 126410 76560
rect 128600 76400 129600 76560
rect 131790 76400 132790 76560
rect 134980 76400 135980 76560
rect 0 76377 3030 76400
rect 0 73393 23 76377
rect 3007 75370 3030 76377
rect 3190 76377 6220 76400
rect 3190 75370 3213 76377
rect 3007 74370 3213 75370
rect 3007 73393 3030 74370
rect 0 73370 3030 73393
rect 3190 73393 3213 74370
rect 6197 75370 6220 76377
rect 6380 76377 9410 76400
rect 6380 75370 6403 76377
rect 6197 74370 6403 75370
rect 6197 73393 6220 74370
rect 3190 73370 6220 73393
rect 6380 73393 6403 74370
rect 9387 75370 9410 76377
rect 9570 76377 12600 76400
rect 9570 75370 9593 76377
rect 9387 74370 9593 75370
rect 9387 73393 9410 74370
rect 6380 73370 9410 73393
rect 9570 73393 9593 74370
rect 12577 75370 12600 76377
rect 12760 76377 15790 76400
rect 12760 75370 12783 76377
rect 12577 74370 12783 75370
rect 12577 73393 12600 74370
rect 9570 73370 12600 73393
rect 12760 73393 12783 74370
rect 15767 75370 15790 76377
rect 15950 76377 18980 76400
rect 15950 75370 15973 76377
rect 15767 74370 15973 75370
rect 15767 73393 15790 74370
rect 12760 73370 15790 73393
rect 15950 73393 15973 74370
rect 18957 75370 18980 76377
rect 19140 76377 22170 76400
rect 19140 75370 19163 76377
rect 18957 74370 19163 75370
rect 18957 73393 18980 74370
rect 15950 73370 18980 73393
rect 19140 73393 19163 74370
rect 22147 75370 22170 76377
rect 22330 76377 25360 76400
rect 22330 75370 22353 76377
rect 22147 74370 22353 75370
rect 22147 73393 22170 74370
rect 19140 73370 22170 73393
rect 22330 73393 22353 74370
rect 25337 75370 25360 76377
rect 25520 76377 28550 76400
rect 25520 75370 25543 76377
rect 25337 74370 25543 75370
rect 25337 73393 25360 74370
rect 22330 73370 25360 73393
rect 25520 73393 25543 74370
rect 28527 75370 28550 76377
rect 28710 76377 31740 76400
rect 28710 75370 28733 76377
rect 28527 74370 28733 75370
rect 28527 73393 28550 74370
rect 25520 73370 28550 73393
rect 28710 73393 28733 74370
rect 31717 75370 31740 76377
rect 31900 76377 34930 76400
rect 31900 75370 31923 76377
rect 31717 74370 31923 75370
rect 31717 73393 31740 74370
rect 28710 73370 31740 73393
rect 31900 73393 31923 74370
rect 34907 75370 34930 76377
rect 35090 76377 38120 76400
rect 35090 75370 35113 76377
rect 34907 74370 35113 75370
rect 34907 73393 34930 74370
rect 31900 73370 34930 73393
rect 35090 73393 35113 74370
rect 38097 75370 38120 76377
rect 38280 76377 41310 76400
rect 38280 75370 38303 76377
rect 38097 74370 38303 75370
rect 38097 73393 38120 74370
rect 35090 73370 38120 73393
rect 38280 73393 38303 74370
rect 41287 75370 41310 76377
rect 41470 76377 44500 76400
rect 41470 75370 41493 76377
rect 41287 74370 41493 75370
rect 41287 73393 41310 74370
rect 38280 73370 41310 73393
rect 41470 73393 41493 74370
rect 44477 75370 44500 76377
rect 44660 76377 47690 76400
rect 44660 75370 44683 76377
rect 44477 74370 44683 75370
rect 44477 73393 44500 74370
rect 41470 73370 44500 73393
rect 44660 73393 44683 74370
rect 47667 75370 47690 76377
rect 47850 76377 50880 76400
rect 47850 75370 47873 76377
rect 47667 74370 47873 75370
rect 47667 73393 47690 74370
rect 44660 73370 47690 73393
rect 47850 73393 47873 74370
rect 50857 75370 50880 76377
rect 51040 76377 54070 76400
rect 51040 75370 51063 76377
rect 50857 74370 51063 75370
rect 50857 73393 50880 74370
rect 47850 73370 50880 73393
rect 51040 73393 51063 74370
rect 54047 75370 54070 76377
rect 54230 76377 57260 76400
rect 54230 75370 54253 76377
rect 54047 74370 54253 75370
rect 54047 73393 54070 74370
rect 51040 73370 54070 73393
rect 54230 73393 54253 74370
rect 57237 75370 57260 76377
rect 57420 76377 60450 76400
rect 57420 75370 57443 76377
rect 57237 74370 57443 75370
rect 57237 73393 57260 74370
rect 54230 73370 57260 73393
rect 57420 73393 57443 74370
rect 60427 75370 60450 76377
rect 60610 76377 63640 76400
rect 60610 75370 60633 76377
rect 60427 74370 60633 75370
rect 60427 73393 60450 74370
rect 57420 73370 60450 73393
rect 60610 73393 60633 74370
rect 63617 75370 63640 76377
rect 63800 76377 66830 76400
rect 63800 75370 63823 76377
rect 63617 74370 63823 75370
rect 63617 73393 63640 74370
rect 60610 73370 63640 73393
rect 63800 73393 63823 74370
rect 66807 75370 66830 76377
rect 66990 76377 70020 76400
rect 66990 75370 67013 76377
rect 66807 74370 67013 75370
rect 66807 73393 66830 74370
rect 63800 73370 66830 73393
rect 66990 73393 67013 74370
rect 69997 75370 70020 76377
rect 70180 76377 73210 76400
rect 70180 75370 70203 76377
rect 69997 74370 70203 75370
rect 69997 73393 70020 74370
rect 66990 73370 70020 73393
rect 70180 73393 70203 74370
rect 73187 75370 73210 76377
rect 73370 76377 76400 76400
rect 73370 75370 73393 76377
rect 73187 74370 73393 75370
rect 73187 73393 73210 74370
rect 70180 73370 73210 73393
rect 73370 73393 73393 74370
rect 76377 75370 76400 76377
rect 76560 76377 79590 76400
rect 76560 75370 76583 76377
rect 76377 74370 76583 75370
rect 76377 73393 76400 74370
rect 73370 73370 76400 73393
rect 76560 73393 76583 74370
rect 79567 75370 79590 76377
rect 79750 76377 82780 76400
rect 79750 75370 79773 76377
rect 79567 74370 79773 75370
rect 79567 73393 79590 74370
rect 76560 73370 79590 73393
rect 79750 73393 79773 74370
rect 82757 75370 82780 76377
rect 82940 76377 85970 76400
rect 82940 75370 82963 76377
rect 82757 74370 82963 75370
rect 82757 73393 82780 74370
rect 79750 73370 82780 73393
rect 82940 73393 82963 74370
rect 85947 75370 85970 76377
rect 86130 76377 89160 76400
rect 86130 75370 86153 76377
rect 85947 74370 86153 75370
rect 85947 73393 85970 74370
rect 82940 73370 85970 73393
rect 86130 73393 86153 74370
rect 89137 75370 89160 76377
rect 89320 76377 92350 76400
rect 89320 75370 89343 76377
rect 89137 74370 89343 75370
rect 89137 73393 89160 74370
rect 86130 73370 89160 73393
rect 89320 73393 89343 74370
rect 92327 75370 92350 76377
rect 92510 76377 95540 76400
rect 92510 75370 92533 76377
rect 92327 74370 92533 75370
rect 92327 73393 92350 74370
rect 89320 73370 92350 73393
rect 92510 73393 92533 74370
rect 95517 75370 95540 76377
rect 95700 76377 98730 76400
rect 95700 75370 95723 76377
rect 95517 74370 95723 75370
rect 95517 73393 95540 74370
rect 92510 73370 95540 73393
rect 95700 73393 95723 74370
rect 98707 75370 98730 76377
rect 98890 76377 101920 76400
rect 98890 75370 98913 76377
rect 98707 74370 98913 75370
rect 98707 73393 98730 74370
rect 95700 73370 98730 73393
rect 98890 73393 98913 74370
rect 101897 75370 101920 76377
rect 102080 76377 105110 76400
rect 102080 75370 102103 76377
rect 101897 74370 102103 75370
rect 101897 73393 101920 74370
rect 98890 73370 101920 73393
rect 102080 73393 102103 74370
rect 105087 75370 105110 76377
rect 105270 76377 108300 76400
rect 105270 75370 105293 76377
rect 105087 74370 105293 75370
rect 105087 73393 105110 74370
rect 102080 73370 105110 73393
rect 105270 73393 105293 74370
rect 108277 75370 108300 76377
rect 108460 76377 111490 76400
rect 108460 75370 108483 76377
rect 108277 74370 108483 75370
rect 108277 73393 108300 74370
rect 105270 73370 108300 73393
rect 108460 73393 108483 74370
rect 111467 75370 111490 76377
rect 111650 76377 114680 76400
rect 111650 75370 111673 76377
rect 111467 74370 111673 75370
rect 111467 73393 111490 74370
rect 108460 73370 111490 73393
rect 111650 73393 111673 74370
rect 114657 75370 114680 76377
rect 114840 76377 117870 76400
rect 114840 75370 114863 76377
rect 114657 74370 114863 75370
rect 114657 73393 114680 74370
rect 111650 73370 114680 73393
rect 114840 73393 114863 74370
rect 117847 75370 117870 76377
rect 118030 76377 121060 76400
rect 118030 75370 118053 76377
rect 117847 74370 118053 75370
rect 117847 73393 117870 74370
rect 114840 73370 117870 73393
rect 118030 73393 118053 74370
rect 121037 75370 121060 76377
rect 121220 76377 124250 76400
rect 121220 75370 121243 76377
rect 121037 74370 121243 75370
rect 121037 73393 121060 74370
rect 118030 73370 121060 73393
rect 121220 73393 121243 74370
rect 124227 75370 124250 76377
rect 124410 76377 127440 76400
rect 124410 75370 124433 76377
rect 124227 74370 124433 75370
rect 124227 73393 124250 74370
rect 121220 73370 124250 73393
rect 124410 73393 124433 74370
rect 127417 75370 127440 76377
rect 127600 76377 130630 76400
rect 127600 75370 127623 76377
rect 127417 74370 127623 75370
rect 127417 73393 127440 74370
rect 124410 73370 127440 73393
rect 127600 73393 127623 74370
rect 130607 75370 130630 76377
rect 130790 76377 133820 76400
rect 130790 75370 130813 76377
rect 130607 74370 130813 75370
rect 130607 73393 130630 74370
rect 127600 73370 130630 73393
rect 130790 73393 130813 74370
rect 133797 75370 133820 76377
rect 133980 76377 137010 76400
rect 133980 75370 134003 76377
rect 133797 74370 134003 75370
rect 133797 73393 133820 74370
rect 130790 73370 133820 73393
rect 133980 73393 134003 74370
rect 136987 75370 137010 76377
rect 136987 74370 137170 75370
rect 136987 73393 137010 74370
rect 133980 73370 137010 73393
rect 1000 73210 2000 73370
rect 4190 73210 5190 73370
rect 7380 73210 8380 73370
rect 10570 73210 11570 73370
rect 13760 73210 14760 73370
rect 16950 73210 17950 73370
rect 20140 73210 21140 73370
rect 23330 73210 24330 73370
rect 26520 73210 27520 73370
rect 29710 73210 30710 73370
rect 32900 73210 33900 73370
rect 36090 73210 37090 73370
rect 39280 73210 40280 73370
rect 42470 73210 43470 73370
rect 45660 73210 46660 73370
rect 48850 73210 49850 73370
rect 52040 73210 53040 73370
rect 55230 73210 56230 73370
rect 58420 73210 59420 73370
rect 61610 73210 62610 73370
rect 64800 73210 65800 73370
rect 67990 73210 68990 73370
rect 71180 73210 72180 73370
rect 74370 73210 75370 73370
rect 77560 73210 78560 73370
rect 80750 73210 81750 73370
rect 83940 73210 84940 73370
rect 87130 73210 88130 73370
rect 90320 73210 91320 73370
rect 93510 73210 94510 73370
rect 96700 73210 97700 73370
rect 99890 73210 100890 73370
rect 103080 73210 104080 73370
rect 106270 73210 107270 73370
rect 109460 73210 110460 73370
rect 112650 73210 113650 73370
rect 115840 73210 116840 73370
rect 119030 73210 120030 73370
rect 122220 73210 123220 73370
rect 125410 73210 126410 73370
rect 128600 73210 129600 73370
rect 131790 73210 132790 73370
rect 134980 73210 135980 73370
rect 0 73187 3030 73210
rect 0 70203 23 73187
rect 3007 72180 3030 73187
rect 3190 73187 6220 73210
rect 3190 72180 3213 73187
rect 3007 71180 3213 72180
rect 3007 70203 3030 71180
rect 0 70180 3030 70203
rect 3190 70203 3213 71180
rect 6197 72180 6220 73187
rect 6380 73187 9410 73210
rect 6380 72180 6403 73187
rect 6197 71180 6403 72180
rect 6197 70203 6220 71180
rect 3190 70180 6220 70203
rect 6380 70203 6403 71180
rect 9387 72180 9410 73187
rect 9570 73187 12600 73210
rect 9570 72180 9593 73187
rect 9387 71180 9593 72180
rect 9387 70203 9410 71180
rect 6380 70180 9410 70203
rect 9570 70203 9593 71180
rect 12577 72180 12600 73187
rect 12760 73187 15790 73210
rect 12760 72180 12783 73187
rect 12577 71180 12783 72180
rect 12577 70203 12600 71180
rect 9570 70180 12600 70203
rect 12760 70203 12783 71180
rect 15767 72180 15790 73187
rect 15950 73187 18980 73210
rect 15950 72180 15973 73187
rect 15767 71180 15973 72180
rect 15767 70203 15790 71180
rect 12760 70180 15790 70203
rect 15950 70203 15973 71180
rect 18957 72180 18980 73187
rect 19140 73187 22170 73210
rect 19140 72180 19163 73187
rect 18957 71180 19163 72180
rect 18957 70203 18980 71180
rect 15950 70180 18980 70203
rect 19140 70203 19163 71180
rect 22147 72180 22170 73187
rect 22330 73187 25360 73210
rect 22330 72180 22353 73187
rect 22147 71180 22353 72180
rect 22147 70203 22170 71180
rect 19140 70180 22170 70203
rect 22330 70203 22353 71180
rect 25337 72180 25360 73187
rect 25520 73187 28550 73210
rect 25520 72180 25543 73187
rect 25337 71180 25543 72180
rect 25337 70203 25360 71180
rect 22330 70180 25360 70203
rect 25520 70203 25543 71180
rect 28527 72180 28550 73187
rect 28710 73187 31740 73210
rect 28710 72180 28733 73187
rect 28527 71180 28733 72180
rect 28527 70203 28550 71180
rect 25520 70180 28550 70203
rect 28710 70203 28733 71180
rect 31717 72180 31740 73187
rect 31900 73187 34930 73210
rect 31900 72180 31923 73187
rect 31717 71180 31923 72180
rect 31717 70203 31740 71180
rect 28710 70180 31740 70203
rect 31900 70203 31923 71180
rect 34907 72180 34930 73187
rect 35090 73187 38120 73210
rect 35090 72180 35113 73187
rect 34907 71180 35113 72180
rect 34907 70203 34930 71180
rect 31900 70180 34930 70203
rect 35090 70203 35113 71180
rect 38097 72180 38120 73187
rect 38280 73187 41310 73210
rect 38280 72180 38303 73187
rect 38097 71180 38303 72180
rect 38097 70203 38120 71180
rect 35090 70180 38120 70203
rect 38280 70203 38303 71180
rect 41287 72180 41310 73187
rect 41470 73187 44500 73210
rect 41470 72180 41493 73187
rect 41287 71180 41493 72180
rect 41287 70203 41310 71180
rect 38280 70180 41310 70203
rect 41470 70203 41493 71180
rect 44477 72180 44500 73187
rect 44660 73187 47690 73210
rect 44660 72180 44683 73187
rect 44477 71180 44683 72180
rect 44477 70203 44500 71180
rect 41470 70180 44500 70203
rect 44660 70203 44683 71180
rect 47667 72180 47690 73187
rect 47850 73187 50880 73210
rect 47850 72180 47873 73187
rect 47667 71180 47873 72180
rect 47667 70203 47690 71180
rect 44660 70180 47690 70203
rect 47850 70203 47873 71180
rect 50857 72180 50880 73187
rect 51040 73187 54070 73210
rect 51040 72180 51063 73187
rect 50857 71180 51063 72180
rect 50857 70203 50880 71180
rect 47850 70180 50880 70203
rect 51040 70203 51063 71180
rect 54047 72180 54070 73187
rect 54230 73187 57260 73210
rect 54230 72180 54253 73187
rect 54047 71180 54253 72180
rect 54047 70203 54070 71180
rect 51040 70180 54070 70203
rect 54230 70203 54253 71180
rect 57237 72180 57260 73187
rect 57420 73187 60450 73210
rect 57420 72180 57443 73187
rect 57237 71180 57443 72180
rect 57237 70203 57260 71180
rect 54230 70180 57260 70203
rect 57420 70203 57443 71180
rect 60427 72180 60450 73187
rect 60610 73187 63640 73210
rect 60610 72180 60633 73187
rect 60427 71180 60633 72180
rect 60427 70203 60450 71180
rect 57420 70180 60450 70203
rect 60610 70203 60633 71180
rect 63617 72180 63640 73187
rect 63800 73187 66830 73210
rect 63800 72180 63823 73187
rect 63617 71180 63823 72180
rect 63617 70203 63640 71180
rect 60610 70180 63640 70203
rect 63800 70203 63823 71180
rect 66807 72180 66830 73187
rect 66990 73187 70020 73210
rect 66990 72180 67013 73187
rect 66807 71180 67013 72180
rect 66807 70203 66830 71180
rect 63800 70180 66830 70203
rect 66990 70203 67013 71180
rect 69997 72180 70020 73187
rect 70180 73187 73210 73210
rect 70180 72180 70203 73187
rect 69997 71180 70203 72180
rect 69997 70203 70020 71180
rect 66990 70180 70020 70203
rect 70180 70203 70203 71180
rect 73187 72180 73210 73187
rect 73370 73187 76400 73210
rect 73370 72180 73393 73187
rect 73187 71180 73393 72180
rect 73187 70203 73210 71180
rect 70180 70180 73210 70203
rect 73370 70203 73393 71180
rect 76377 72180 76400 73187
rect 76560 73187 79590 73210
rect 76560 72180 76583 73187
rect 76377 71180 76583 72180
rect 76377 70203 76400 71180
rect 73370 70180 76400 70203
rect 76560 70203 76583 71180
rect 79567 72180 79590 73187
rect 79750 73187 82780 73210
rect 79750 72180 79773 73187
rect 79567 71180 79773 72180
rect 79567 70203 79590 71180
rect 76560 70180 79590 70203
rect 79750 70203 79773 71180
rect 82757 72180 82780 73187
rect 82940 73187 85970 73210
rect 82940 72180 82963 73187
rect 82757 71180 82963 72180
rect 82757 70203 82780 71180
rect 79750 70180 82780 70203
rect 82940 70203 82963 71180
rect 85947 72180 85970 73187
rect 86130 73187 89160 73210
rect 86130 72180 86153 73187
rect 85947 71180 86153 72180
rect 85947 70203 85970 71180
rect 82940 70180 85970 70203
rect 86130 70203 86153 71180
rect 89137 72180 89160 73187
rect 89320 73187 92350 73210
rect 89320 72180 89343 73187
rect 89137 71180 89343 72180
rect 89137 70203 89160 71180
rect 86130 70180 89160 70203
rect 89320 70203 89343 71180
rect 92327 72180 92350 73187
rect 92510 73187 95540 73210
rect 92510 72180 92533 73187
rect 92327 71180 92533 72180
rect 92327 70203 92350 71180
rect 89320 70180 92350 70203
rect 92510 70203 92533 71180
rect 95517 72180 95540 73187
rect 95700 73187 98730 73210
rect 95700 72180 95723 73187
rect 95517 71180 95723 72180
rect 95517 70203 95540 71180
rect 92510 70180 95540 70203
rect 95700 70203 95723 71180
rect 98707 72180 98730 73187
rect 98890 73187 101920 73210
rect 98890 72180 98913 73187
rect 98707 71180 98913 72180
rect 98707 70203 98730 71180
rect 95700 70180 98730 70203
rect 98890 70203 98913 71180
rect 101897 72180 101920 73187
rect 102080 73187 105110 73210
rect 102080 72180 102103 73187
rect 101897 71180 102103 72180
rect 101897 70203 101920 71180
rect 98890 70180 101920 70203
rect 102080 70203 102103 71180
rect 105087 72180 105110 73187
rect 105270 73187 108300 73210
rect 105270 72180 105293 73187
rect 105087 71180 105293 72180
rect 105087 70203 105110 71180
rect 102080 70180 105110 70203
rect 105270 70203 105293 71180
rect 108277 72180 108300 73187
rect 108460 73187 111490 73210
rect 108460 72180 108483 73187
rect 108277 71180 108483 72180
rect 108277 70203 108300 71180
rect 105270 70180 108300 70203
rect 108460 70203 108483 71180
rect 111467 72180 111490 73187
rect 111650 73187 114680 73210
rect 111650 72180 111673 73187
rect 111467 71180 111673 72180
rect 111467 70203 111490 71180
rect 108460 70180 111490 70203
rect 111650 70203 111673 71180
rect 114657 72180 114680 73187
rect 114840 73187 117870 73210
rect 114840 72180 114863 73187
rect 114657 71180 114863 72180
rect 114657 70203 114680 71180
rect 111650 70180 114680 70203
rect 114840 70203 114863 71180
rect 117847 72180 117870 73187
rect 118030 73187 121060 73210
rect 118030 72180 118053 73187
rect 117847 71180 118053 72180
rect 117847 70203 117870 71180
rect 114840 70180 117870 70203
rect 118030 70203 118053 71180
rect 121037 72180 121060 73187
rect 121220 73187 124250 73210
rect 121220 72180 121243 73187
rect 121037 71180 121243 72180
rect 121037 70203 121060 71180
rect 118030 70180 121060 70203
rect 121220 70203 121243 71180
rect 124227 72180 124250 73187
rect 124410 73187 127440 73210
rect 124410 72180 124433 73187
rect 124227 71180 124433 72180
rect 124227 70203 124250 71180
rect 121220 70180 124250 70203
rect 124410 70203 124433 71180
rect 127417 72180 127440 73187
rect 127600 73187 130630 73210
rect 127600 72180 127623 73187
rect 127417 71180 127623 72180
rect 127417 70203 127440 71180
rect 124410 70180 127440 70203
rect 127600 70203 127623 71180
rect 130607 72180 130630 73187
rect 130790 73187 133820 73210
rect 130790 72180 130813 73187
rect 130607 71180 130813 72180
rect 130607 70203 130630 71180
rect 127600 70180 130630 70203
rect 130790 70203 130813 71180
rect 133797 72180 133820 73187
rect 133980 73187 137010 73210
rect 133980 72180 134003 73187
rect 133797 71180 134003 72180
rect 133797 70203 133820 71180
rect 130790 70180 133820 70203
rect 133980 70203 134003 71180
rect 136987 72180 137010 73187
rect 136987 71180 137170 72180
rect 136987 70203 137010 71180
rect 133980 70180 137010 70203
rect 1000 70020 2000 70180
rect 4190 70020 5190 70180
rect 7380 70020 8380 70180
rect 10570 70020 11570 70180
rect 13760 70020 14760 70180
rect 16950 70020 17950 70180
rect 20140 70020 21140 70180
rect 23330 70020 24330 70180
rect 26520 70020 27520 70180
rect 29710 70020 30710 70180
rect 32900 70020 33900 70180
rect 36090 70020 37090 70180
rect 39280 70020 40280 70180
rect 42470 70020 43470 70180
rect 45660 70020 46660 70180
rect 48850 70020 49850 70180
rect 52040 70020 53040 70180
rect 55230 70020 56230 70180
rect 58420 70020 59420 70180
rect 61610 70020 62610 70180
rect 64800 70020 65800 70180
rect 67990 70020 68990 70180
rect 71180 70020 72180 70180
rect 74370 70020 75370 70180
rect 77560 70020 78560 70180
rect 80750 70020 81750 70180
rect 83940 70020 84940 70180
rect 87130 70020 88130 70180
rect 90320 70020 91320 70180
rect 93510 70020 94510 70180
rect 96700 70020 97700 70180
rect 99890 70020 100890 70180
rect 103080 70020 104080 70180
rect 106270 70020 107270 70180
rect 109460 70020 110460 70180
rect 112650 70020 113650 70180
rect 115840 70020 116840 70180
rect 119030 70020 120030 70180
rect 122220 70020 123220 70180
rect 125410 70020 126410 70180
rect 128600 70020 129600 70180
rect 131790 70020 132790 70180
rect 134980 70020 135980 70180
rect 0 69997 3030 70020
rect 0 67013 23 69997
rect 3007 68990 3030 69997
rect 3190 69997 6220 70020
rect 3190 68990 3213 69997
rect 3007 67990 3213 68990
rect 3007 67013 3030 67990
rect 0 66990 3030 67013
rect 3190 67013 3213 67990
rect 6197 68990 6220 69997
rect 6380 69997 9410 70020
rect 6380 68990 6403 69997
rect 6197 67990 6403 68990
rect 6197 67013 6220 67990
rect 3190 66990 6220 67013
rect 6380 67013 6403 67990
rect 9387 68990 9410 69997
rect 9570 69997 12600 70020
rect 9570 68990 9593 69997
rect 9387 67990 9593 68990
rect 9387 67013 9410 67990
rect 6380 66990 9410 67013
rect 9570 67013 9593 67990
rect 12577 68990 12600 69997
rect 12760 69997 15790 70020
rect 12760 68990 12783 69997
rect 12577 67990 12783 68990
rect 12577 67013 12600 67990
rect 9570 66990 12600 67013
rect 12760 67013 12783 67990
rect 15767 68990 15790 69997
rect 15950 69997 18980 70020
rect 15950 68990 15973 69997
rect 15767 67990 15973 68990
rect 15767 67013 15790 67990
rect 12760 66990 15790 67013
rect 15950 67013 15973 67990
rect 18957 68990 18980 69997
rect 19140 69997 22170 70020
rect 19140 68990 19163 69997
rect 18957 67990 19163 68990
rect 18957 67013 18980 67990
rect 15950 66990 18980 67013
rect 19140 67013 19163 67990
rect 22147 68990 22170 69997
rect 22330 69997 25360 70020
rect 22330 68990 22353 69997
rect 22147 67990 22353 68990
rect 22147 67013 22170 67990
rect 19140 66990 22170 67013
rect 22330 67013 22353 67990
rect 25337 68990 25360 69997
rect 25520 69997 28550 70020
rect 25520 68990 25543 69997
rect 25337 67990 25543 68990
rect 25337 67013 25360 67990
rect 22330 66990 25360 67013
rect 25520 67013 25543 67990
rect 28527 68990 28550 69997
rect 28710 69997 31740 70020
rect 28710 68990 28733 69997
rect 28527 67990 28733 68990
rect 28527 67013 28550 67990
rect 25520 66990 28550 67013
rect 28710 67013 28733 67990
rect 31717 68990 31740 69997
rect 31900 69997 34930 70020
rect 31900 68990 31923 69997
rect 31717 67990 31923 68990
rect 31717 67013 31740 67990
rect 28710 66990 31740 67013
rect 31900 67013 31923 67990
rect 34907 68990 34930 69997
rect 35090 69997 38120 70020
rect 35090 68990 35113 69997
rect 34907 67990 35113 68990
rect 34907 67013 34930 67990
rect 31900 66990 34930 67013
rect 35090 67013 35113 67990
rect 38097 68990 38120 69997
rect 38280 69997 41310 70020
rect 38280 68990 38303 69997
rect 38097 67990 38303 68990
rect 38097 67013 38120 67990
rect 35090 66990 38120 67013
rect 38280 67013 38303 67990
rect 41287 68990 41310 69997
rect 41470 69997 44500 70020
rect 41470 68990 41493 69997
rect 41287 67990 41493 68990
rect 41287 67013 41310 67990
rect 38280 66990 41310 67013
rect 41470 67013 41493 67990
rect 44477 68990 44500 69997
rect 44660 69997 47690 70020
rect 44660 68990 44683 69997
rect 44477 67990 44683 68990
rect 44477 67013 44500 67990
rect 41470 66990 44500 67013
rect 44660 67013 44683 67990
rect 47667 68990 47690 69997
rect 47850 69997 50880 70020
rect 47850 68990 47873 69997
rect 47667 67990 47873 68990
rect 47667 67013 47690 67990
rect 44660 66990 47690 67013
rect 47850 67013 47873 67990
rect 50857 68990 50880 69997
rect 51040 69997 54070 70020
rect 51040 68990 51063 69997
rect 50857 67990 51063 68990
rect 50857 67013 50880 67990
rect 47850 66990 50880 67013
rect 51040 67013 51063 67990
rect 54047 68990 54070 69997
rect 54230 69997 57260 70020
rect 54230 68990 54253 69997
rect 54047 67990 54253 68990
rect 54047 67013 54070 67990
rect 51040 66990 54070 67013
rect 54230 67013 54253 67990
rect 57237 68990 57260 69997
rect 57420 69997 60450 70020
rect 57420 68990 57443 69997
rect 57237 67990 57443 68990
rect 57237 67013 57260 67990
rect 54230 66990 57260 67013
rect 57420 67013 57443 67990
rect 60427 68990 60450 69997
rect 60610 69997 63640 70020
rect 60610 68990 60633 69997
rect 60427 67990 60633 68990
rect 60427 67013 60450 67990
rect 57420 66990 60450 67013
rect 60610 67013 60633 67990
rect 63617 68990 63640 69997
rect 63800 69997 66830 70020
rect 63800 68990 63823 69997
rect 63617 67990 63823 68990
rect 63617 67013 63640 67990
rect 60610 66990 63640 67013
rect 63800 67013 63823 67990
rect 66807 68990 66830 69997
rect 66990 69997 70020 70020
rect 66990 68990 67013 69997
rect 66807 67990 67013 68990
rect 66807 67013 66830 67990
rect 63800 66990 66830 67013
rect 66990 67013 67013 67990
rect 69997 68990 70020 69997
rect 70180 69997 73210 70020
rect 70180 68990 70203 69997
rect 69997 67990 70203 68990
rect 69997 67013 70020 67990
rect 66990 66990 70020 67013
rect 70180 67013 70203 67990
rect 73187 68990 73210 69997
rect 73370 69997 76400 70020
rect 73370 68990 73393 69997
rect 73187 67990 73393 68990
rect 73187 67013 73210 67990
rect 70180 66990 73210 67013
rect 73370 67013 73393 67990
rect 76377 68990 76400 69997
rect 76560 69997 79590 70020
rect 76560 68990 76583 69997
rect 76377 67990 76583 68990
rect 76377 67013 76400 67990
rect 73370 66990 76400 67013
rect 76560 67013 76583 67990
rect 79567 68990 79590 69997
rect 79750 69997 82780 70020
rect 79750 68990 79773 69997
rect 79567 67990 79773 68990
rect 79567 67013 79590 67990
rect 76560 66990 79590 67013
rect 79750 67013 79773 67990
rect 82757 68990 82780 69997
rect 82940 69997 85970 70020
rect 82940 68990 82963 69997
rect 82757 67990 82963 68990
rect 82757 67013 82780 67990
rect 79750 66990 82780 67013
rect 82940 67013 82963 67990
rect 85947 68990 85970 69997
rect 86130 69997 89160 70020
rect 86130 68990 86153 69997
rect 85947 67990 86153 68990
rect 85947 67013 85970 67990
rect 82940 66990 85970 67013
rect 86130 67013 86153 67990
rect 89137 68990 89160 69997
rect 89320 69997 92350 70020
rect 89320 68990 89343 69997
rect 89137 67990 89343 68990
rect 89137 67013 89160 67990
rect 86130 66990 89160 67013
rect 89320 67013 89343 67990
rect 92327 68990 92350 69997
rect 92510 69997 95540 70020
rect 92510 68990 92533 69997
rect 92327 67990 92533 68990
rect 92327 67013 92350 67990
rect 89320 66990 92350 67013
rect 92510 67013 92533 67990
rect 95517 68990 95540 69997
rect 95700 69997 98730 70020
rect 95700 68990 95723 69997
rect 95517 67990 95723 68990
rect 95517 67013 95540 67990
rect 92510 66990 95540 67013
rect 95700 67013 95723 67990
rect 98707 68990 98730 69997
rect 98890 69997 101920 70020
rect 98890 68990 98913 69997
rect 98707 67990 98913 68990
rect 98707 67013 98730 67990
rect 95700 66990 98730 67013
rect 98890 67013 98913 67990
rect 101897 68990 101920 69997
rect 102080 69997 105110 70020
rect 102080 68990 102103 69997
rect 101897 67990 102103 68990
rect 101897 67013 101920 67990
rect 98890 66990 101920 67013
rect 102080 67013 102103 67990
rect 105087 68990 105110 69997
rect 105270 69997 108300 70020
rect 105270 68990 105293 69997
rect 105087 67990 105293 68990
rect 105087 67013 105110 67990
rect 102080 66990 105110 67013
rect 105270 67013 105293 67990
rect 108277 68990 108300 69997
rect 108460 69997 111490 70020
rect 108460 68990 108483 69997
rect 108277 67990 108483 68990
rect 108277 67013 108300 67990
rect 105270 66990 108300 67013
rect 108460 67013 108483 67990
rect 111467 68990 111490 69997
rect 111650 69997 114680 70020
rect 111650 68990 111673 69997
rect 111467 67990 111673 68990
rect 111467 67013 111490 67990
rect 108460 66990 111490 67013
rect 111650 67013 111673 67990
rect 114657 68990 114680 69997
rect 114840 69997 117870 70020
rect 114840 68990 114863 69997
rect 114657 67990 114863 68990
rect 114657 67013 114680 67990
rect 111650 66990 114680 67013
rect 114840 67013 114863 67990
rect 117847 68990 117870 69997
rect 118030 69997 121060 70020
rect 118030 68990 118053 69997
rect 117847 67990 118053 68990
rect 117847 67013 117870 67990
rect 114840 66990 117870 67013
rect 118030 67013 118053 67990
rect 121037 68990 121060 69997
rect 121220 69997 124250 70020
rect 121220 68990 121243 69997
rect 121037 67990 121243 68990
rect 121037 67013 121060 67990
rect 118030 66990 121060 67013
rect 121220 67013 121243 67990
rect 124227 68990 124250 69997
rect 124410 69997 127440 70020
rect 124410 68990 124433 69997
rect 124227 67990 124433 68990
rect 124227 67013 124250 67990
rect 121220 66990 124250 67013
rect 124410 67013 124433 67990
rect 127417 68990 127440 69997
rect 127600 69997 130630 70020
rect 127600 68990 127623 69997
rect 127417 67990 127623 68990
rect 127417 67013 127440 67990
rect 124410 66990 127440 67013
rect 127600 67013 127623 67990
rect 130607 68990 130630 69997
rect 130790 69997 133820 70020
rect 130790 68990 130813 69997
rect 130607 67990 130813 68990
rect 130607 67013 130630 67990
rect 127600 66990 130630 67013
rect 130790 67013 130813 67990
rect 133797 68990 133820 69997
rect 133980 69997 137010 70020
rect 133980 68990 134003 69997
rect 133797 67990 134003 68990
rect 133797 67013 133820 67990
rect 130790 66990 133820 67013
rect 133980 67013 134003 67990
rect 136987 68990 137010 69997
rect 136987 67990 137170 68990
rect 136987 67013 137010 67990
rect 133980 66990 137010 67013
rect 1000 66830 2000 66990
rect 4190 66830 5190 66990
rect 7380 66830 8380 66990
rect 10570 66830 11570 66990
rect 13760 66830 14760 66990
rect 16950 66830 17950 66990
rect 20140 66830 21140 66990
rect 23330 66830 24330 66990
rect 26520 66830 27520 66990
rect 29710 66830 30710 66990
rect 32900 66830 33900 66990
rect 36090 66830 37090 66990
rect 39280 66830 40280 66990
rect 42470 66830 43470 66990
rect 45660 66830 46660 66990
rect 48850 66830 49850 66990
rect 52040 66830 53040 66990
rect 55230 66830 56230 66990
rect 58420 66830 59420 66990
rect 61610 66830 62610 66990
rect 64800 66830 65800 66990
rect 67990 66830 68990 66990
rect 71180 66830 72180 66990
rect 74370 66830 75370 66990
rect 77560 66830 78560 66990
rect 80750 66830 81750 66990
rect 83940 66830 84940 66990
rect 87130 66830 88130 66990
rect 90320 66830 91320 66990
rect 93510 66830 94510 66990
rect 96700 66830 97700 66990
rect 99890 66830 100890 66990
rect 103080 66830 104080 66990
rect 106270 66830 107270 66990
rect 109460 66830 110460 66990
rect 112650 66830 113650 66990
rect 115840 66830 116840 66990
rect 119030 66830 120030 66990
rect 122220 66830 123220 66990
rect 125410 66830 126410 66990
rect 128600 66830 129600 66990
rect 131790 66830 132790 66990
rect 134980 66830 135980 66990
rect 0 66807 3030 66830
rect 0 63823 23 66807
rect 3007 65800 3030 66807
rect 3190 66807 6220 66830
rect 3190 65800 3213 66807
rect 3007 64800 3213 65800
rect 3007 63823 3030 64800
rect 0 63800 3030 63823
rect 3190 63823 3213 64800
rect 6197 65800 6220 66807
rect 6380 66807 9410 66830
rect 6380 65800 6403 66807
rect 6197 64800 6403 65800
rect 6197 63823 6220 64800
rect 3190 63800 6220 63823
rect 6380 63823 6403 64800
rect 9387 65800 9410 66807
rect 9570 66807 12600 66830
rect 9570 65800 9593 66807
rect 9387 64800 9593 65800
rect 9387 63823 9410 64800
rect 6380 63800 9410 63823
rect 9570 63823 9593 64800
rect 12577 65800 12600 66807
rect 12760 66807 15790 66830
rect 12760 65800 12783 66807
rect 12577 64800 12783 65800
rect 12577 63823 12600 64800
rect 9570 63800 12600 63823
rect 12760 63823 12783 64800
rect 15767 65800 15790 66807
rect 15950 66807 18980 66830
rect 15950 65800 15973 66807
rect 15767 64800 15973 65800
rect 15767 63823 15790 64800
rect 12760 63800 15790 63823
rect 15950 63823 15973 64800
rect 18957 65800 18980 66807
rect 19140 66807 22170 66830
rect 19140 65800 19163 66807
rect 18957 64800 19163 65800
rect 18957 63823 18980 64800
rect 15950 63800 18980 63823
rect 19140 63823 19163 64800
rect 22147 65800 22170 66807
rect 22330 66807 25360 66830
rect 22330 65800 22353 66807
rect 22147 64800 22353 65800
rect 22147 63823 22170 64800
rect 19140 63800 22170 63823
rect 22330 63823 22353 64800
rect 25337 65800 25360 66807
rect 25520 66807 28550 66830
rect 25520 65800 25543 66807
rect 25337 64800 25543 65800
rect 25337 63823 25360 64800
rect 22330 63800 25360 63823
rect 25520 63823 25543 64800
rect 28527 65800 28550 66807
rect 28710 66807 31740 66830
rect 28710 65800 28733 66807
rect 28527 64800 28733 65800
rect 28527 63823 28550 64800
rect 25520 63800 28550 63823
rect 28710 63823 28733 64800
rect 31717 65800 31740 66807
rect 31900 66807 34930 66830
rect 31900 65800 31923 66807
rect 31717 64800 31923 65800
rect 31717 63823 31740 64800
rect 28710 63800 31740 63823
rect 31900 63823 31923 64800
rect 34907 65800 34930 66807
rect 35090 66807 38120 66830
rect 35090 65800 35113 66807
rect 34907 64800 35113 65800
rect 34907 63823 34930 64800
rect 31900 63800 34930 63823
rect 35090 63823 35113 64800
rect 38097 65800 38120 66807
rect 38280 66807 41310 66830
rect 38280 65800 38303 66807
rect 38097 64800 38303 65800
rect 38097 63823 38120 64800
rect 35090 63800 38120 63823
rect 38280 63823 38303 64800
rect 41287 65800 41310 66807
rect 41470 66807 44500 66830
rect 41470 65800 41493 66807
rect 41287 64800 41493 65800
rect 41287 63823 41310 64800
rect 38280 63800 41310 63823
rect 41470 63823 41493 64800
rect 44477 65800 44500 66807
rect 44660 66807 47690 66830
rect 44660 65800 44683 66807
rect 44477 64800 44683 65800
rect 44477 63823 44500 64800
rect 41470 63800 44500 63823
rect 44660 63823 44683 64800
rect 47667 65800 47690 66807
rect 47850 66807 50880 66830
rect 47850 65800 47873 66807
rect 47667 64800 47873 65800
rect 47667 63823 47690 64800
rect 44660 63800 47690 63823
rect 47850 63823 47873 64800
rect 50857 65800 50880 66807
rect 51040 66807 54070 66830
rect 51040 65800 51063 66807
rect 50857 64800 51063 65800
rect 50857 63823 50880 64800
rect 47850 63800 50880 63823
rect 51040 63823 51063 64800
rect 54047 65800 54070 66807
rect 54230 66807 57260 66830
rect 54230 65800 54253 66807
rect 54047 64800 54253 65800
rect 54047 63823 54070 64800
rect 51040 63800 54070 63823
rect 54230 63823 54253 64800
rect 57237 65800 57260 66807
rect 57420 66807 60450 66830
rect 57420 65800 57443 66807
rect 57237 64800 57443 65800
rect 57237 63823 57260 64800
rect 54230 63800 57260 63823
rect 57420 63823 57443 64800
rect 60427 65800 60450 66807
rect 60610 66807 63640 66830
rect 60610 65800 60633 66807
rect 60427 64800 60633 65800
rect 60427 63823 60450 64800
rect 57420 63800 60450 63823
rect 60610 63823 60633 64800
rect 63617 65800 63640 66807
rect 63800 66807 66830 66830
rect 63800 65800 63823 66807
rect 63617 64800 63823 65800
rect 63617 63823 63640 64800
rect 60610 63800 63640 63823
rect 63800 63823 63823 64800
rect 66807 65800 66830 66807
rect 66990 66807 70020 66830
rect 66990 65800 67013 66807
rect 66807 64800 67013 65800
rect 66807 63823 66830 64800
rect 63800 63800 66830 63823
rect 66990 63823 67013 64800
rect 69997 65800 70020 66807
rect 70180 66807 73210 66830
rect 70180 65800 70203 66807
rect 69997 64800 70203 65800
rect 69997 63823 70020 64800
rect 66990 63800 70020 63823
rect 70180 63823 70203 64800
rect 73187 65800 73210 66807
rect 73370 66807 76400 66830
rect 73370 65800 73393 66807
rect 73187 64800 73393 65800
rect 73187 63823 73210 64800
rect 70180 63800 73210 63823
rect 73370 63823 73393 64800
rect 76377 65800 76400 66807
rect 76560 66807 79590 66830
rect 76560 65800 76583 66807
rect 76377 64800 76583 65800
rect 76377 63823 76400 64800
rect 73370 63800 76400 63823
rect 76560 63823 76583 64800
rect 79567 65800 79590 66807
rect 79750 66807 82780 66830
rect 79750 65800 79773 66807
rect 79567 64800 79773 65800
rect 79567 63823 79590 64800
rect 76560 63800 79590 63823
rect 79750 63823 79773 64800
rect 82757 65800 82780 66807
rect 82940 66807 85970 66830
rect 82940 65800 82963 66807
rect 82757 64800 82963 65800
rect 82757 63823 82780 64800
rect 79750 63800 82780 63823
rect 82940 63823 82963 64800
rect 85947 65800 85970 66807
rect 86130 66807 89160 66830
rect 86130 65800 86153 66807
rect 85947 64800 86153 65800
rect 85947 63823 85970 64800
rect 82940 63800 85970 63823
rect 86130 63823 86153 64800
rect 89137 65800 89160 66807
rect 89320 66807 92350 66830
rect 89320 65800 89343 66807
rect 89137 64800 89343 65800
rect 89137 63823 89160 64800
rect 86130 63800 89160 63823
rect 89320 63823 89343 64800
rect 92327 65800 92350 66807
rect 92510 66807 95540 66830
rect 92510 65800 92533 66807
rect 92327 64800 92533 65800
rect 92327 63823 92350 64800
rect 89320 63800 92350 63823
rect 92510 63823 92533 64800
rect 95517 65800 95540 66807
rect 95700 66807 98730 66830
rect 95700 65800 95723 66807
rect 95517 64800 95723 65800
rect 95517 63823 95540 64800
rect 92510 63800 95540 63823
rect 95700 63823 95723 64800
rect 98707 65800 98730 66807
rect 98890 66807 101920 66830
rect 98890 65800 98913 66807
rect 98707 64800 98913 65800
rect 98707 63823 98730 64800
rect 95700 63800 98730 63823
rect 98890 63823 98913 64800
rect 101897 65800 101920 66807
rect 102080 66807 105110 66830
rect 102080 65800 102103 66807
rect 101897 64800 102103 65800
rect 101897 63823 101920 64800
rect 98890 63800 101920 63823
rect 102080 63823 102103 64800
rect 105087 65800 105110 66807
rect 105270 66807 108300 66830
rect 105270 65800 105293 66807
rect 105087 64800 105293 65800
rect 105087 63823 105110 64800
rect 102080 63800 105110 63823
rect 105270 63823 105293 64800
rect 108277 65800 108300 66807
rect 108460 66807 111490 66830
rect 108460 65800 108483 66807
rect 108277 64800 108483 65800
rect 108277 63823 108300 64800
rect 105270 63800 108300 63823
rect 108460 63823 108483 64800
rect 111467 65800 111490 66807
rect 111650 66807 114680 66830
rect 111650 65800 111673 66807
rect 111467 64800 111673 65800
rect 111467 63823 111490 64800
rect 108460 63800 111490 63823
rect 111650 63823 111673 64800
rect 114657 65800 114680 66807
rect 114840 66807 117870 66830
rect 114840 65800 114863 66807
rect 114657 64800 114863 65800
rect 114657 63823 114680 64800
rect 111650 63800 114680 63823
rect 114840 63823 114863 64800
rect 117847 65800 117870 66807
rect 118030 66807 121060 66830
rect 118030 65800 118053 66807
rect 117847 64800 118053 65800
rect 117847 63823 117870 64800
rect 114840 63800 117870 63823
rect 118030 63823 118053 64800
rect 121037 65800 121060 66807
rect 121220 66807 124250 66830
rect 121220 65800 121243 66807
rect 121037 64800 121243 65800
rect 121037 63823 121060 64800
rect 118030 63800 121060 63823
rect 121220 63823 121243 64800
rect 124227 65800 124250 66807
rect 124410 66807 127440 66830
rect 124410 65800 124433 66807
rect 124227 64800 124433 65800
rect 124227 63823 124250 64800
rect 121220 63800 124250 63823
rect 124410 63823 124433 64800
rect 127417 65800 127440 66807
rect 127600 66807 130630 66830
rect 127600 65800 127623 66807
rect 127417 64800 127623 65800
rect 127417 63823 127440 64800
rect 124410 63800 127440 63823
rect 127600 63823 127623 64800
rect 130607 65800 130630 66807
rect 130790 66807 133820 66830
rect 130790 65800 130813 66807
rect 130607 64800 130813 65800
rect 130607 63823 130630 64800
rect 127600 63800 130630 63823
rect 130790 63823 130813 64800
rect 133797 65800 133820 66807
rect 133980 66807 137010 66830
rect 133980 65800 134003 66807
rect 133797 64800 134003 65800
rect 133797 63823 133820 64800
rect 130790 63800 133820 63823
rect 133980 63823 134003 64800
rect 136987 65800 137010 66807
rect 136987 64800 137170 65800
rect 136987 63823 137010 64800
rect 133980 63800 137010 63823
rect 1000 63640 2000 63800
rect 4190 63640 5190 63800
rect 7380 63640 8380 63800
rect 10570 63640 11570 63800
rect 13760 63640 14760 63800
rect 16950 63640 17950 63800
rect 20140 63640 21140 63800
rect 23330 63640 24330 63800
rect 26520 63640 27520 63800
rect 29710 63640 30710 63800
rect 32900 63640 33900 63800
rect 36090 63640 37090 63800
rect 39280 63640 40280 63800
rect 42470 63640 43470 63800
rect 45660 63640 46660 63800
rect 48850 63640 49850 63800
rect 52040 63640 53040 63800
rect 55230 63640 56230 63800
rect 58420 63640 59420 63800
rect 61610 63640 62610 63800
rect 64800 63640 65800 63800
rect 67990 63640 68990 63800
rect 71180 63640 72180 63800
rect 74370 63640 75370 63800
rect 77560 63640 78560 63800
rect 80750 63640 81750 63800
rect 83940 63640 84940 63800
rect 87130 63640 88130 63800
rect 90320 63640 91320 63800
rect 93510 63640 94510 63800
rect 96700 63640 97700 63800
rect 99890 63640 100890 63800
rect 103080 63640 104080 63800
rect 106270 63640 107270 63800
rect 109460 63640 110460 63800
rect 112650 63640 113650 63800
rect 115840 63640 116840 63800
rect 119030 63640 120030 63800
rect 122220 63640 123220 63800
rect 125410 63640 126410 63800
rect 128600 63640 129600 63800
rect 131790 63640 132790 63800
rect 134980 63640 135980 63800
rect 0 63617 3030 63640
rect 0 60633 23 63617
rect 3007 62610 3030 63617
rect 3190 63617 6220 63640
rect 3190 62610 3213 63617
rect 3007 61610 3213 62610
rect 3007 60633 3030 61610
rect 0 60610 3030 60633
rect 3190 60633 3213 61610
rect 6197 62610 6220 63617
rect 6380 63617 9410 63640
rect 6380 62610 6403 63617
rect 6197 61610 6403 62610
rect 6197 60633 6220 61610
rect 3190 60610 6220 60633
rect 6380 60633 6403 61610
rect 9387 62610 9410 63617
rect 9570 63617 12600 63640
rect 9570 62610 9593 63617
rect 9387 61610 9593 62610
rect 9387 60633 9410 61610
rect 6380 60610 9410 60633
rect 9570 60633 9593 61610
rect 12577 62610 12600 63617
rect 12760 63617 15790 63640
rect 12760 62610 12783 63617
rect 12577 61610 12783 62610
rect 12577 60633 12600 61610
rect 9570 60610 12600 60633
rect 12760 60633 12783 61610
rect 15767 62610 15790 63617
rect 15950 63617 18980 63640
rect 15950 62610 15973 63617
rect 15767 61610 15973 62610
rect 15767 60633 15790 61610
rect 12760 60610 15790 60633
rect 15950 60633 15973 61610
rect 18957 62610 18980 63617
rect 19140 63617 22170 63640
rect 19140 62610 19163 63617
rect 18957 61610 19163 62610
rect 18957 60633 18980 61610
rect 15950 60610 18980 60633
rect 19140 60633 19163 61610
rect 22147 62610 22170 63617
rect 22330 63617 25360 63640
rect 22330 62610 22353 63617
rect 22147 61610 22353 62610
rect 22147 60633 22170 61610
rect 19140 60610 22170 60633
rect 22330 60633 22353 61610
rect 25337 62610 25360 63617
rect 25520 63617 28550 63640
rect 25520 62610 25543 63617
rect 25337 61610 25543 62610
rect 25337 60633 25360 61610
rect 22330 60610 25360 60633
rect 25520 60633 25543 61610
rect 28527 62610 28550 63617
rect 28710 63617 31740 63640
rect 28710 62610 28733 63617
rect 28527 61610 28733 62610
rect 28527 60633 28550 61610
rect 25520 60610 28550 60633
rect 28710 60633 28733 61610
rect 31717 62610 31740 63617
rect 31900 63617 34930 63640
rect 31900 62610 31923 63617
rect 31717 61610 31923 62610
rect 31717 60633 31740 61610
rect 28710 60610 31740 60633
rect 31900 60633 31923 61610
rect 34907 62610 34930 63617
rect 35090 63617 38120 63640
rect 35090 62610 35113 63617
rect 34907 61610 35113 62610
rect 34907 60633 34930 61610
rect 31900 60610 34930 60633
rect 35090 60633 35113 61610
rect 38097 62610 38120 63617
rect 38280 63617 41310 63640
rect 38280 62610 38303 63617
rect 38097 61610 38303 62610
rect 38097 60633 38120 61610
rect 35090 60610 38120 60633
rect 38280 60633 38303 61610
rect 41287 62610 41310 63617
rect 41470 63617 44500 63640
rect 41470 62610 41493 63617
rect 41287 61610 41493 62610
rect 41287 60633 41310 61610
rect 38280 60610 41310 60633
rect 41470 60633 41493 61610
rect 44477 62610 44500 63617
rect 44660 63617 47690 63640
rect 44660 62610 44683 63617
rect 44477 61610 44683 62610
rect 44477 60633 44500 61610
rect 41470 60610 44500 60633
rect 44660 60633 44683 61610
rect 47667 62610 47690 63617
rect 47850 63617 50880 63640
rect 47850 62610 47873 63617
rect 47667 61610 47873 62610
rect 47667 60633 47690 61610
rect 44660 60610 47690 60633
rect 47850 60633 47873 61610
rect 50857 62610 50880 63617
rect 51040 63617 54070 63640
rect 51040 62610 51063 63617
rect 50857 61610 51063 62610
rect 50857 60633 50880 61610
rect 47850 60610 50880 60633
rect 51040 60633 51063 61610
rect 54047 62610 54070 63617
rect 54230 63617 57260 63640
rect 54230 62610 54253 63617
rect 54047 61610 54253 62610
rect 54047 60633 54070 61610
rect 51040 60610 54070 60633
rect 54230 60633 54253 61610
rect 57237 62610 57260 63617
rect 57420 63617 60450 63640
rect 57420 62610 57443 63617
rect 57237 61610 57443 62610
rect 57237 60633 57260 61610
rect 54230 60610 57260 60633
rect 57420 60633 57443 61610
rect 60427 62610 60450 63617
rect 60610 63617 63640 63640
rect 60610 62610 60633 63617
rect 60427 61610 60633 62610
rect 60427 60633 60450 61610
rect 57420 60610 60450 60633
rect 60610 60633 60633 61610
rect 63617 62610 63640 63617
rect 63800 63617 66830 63640
rect 63800 62610 63823 63617
rect 63617 61610 63823 62610
rect 63617 60633 63640 61610
rect 60610 60610 63640 60633
rect 63800 60633 63823 61610
rect 66807 62610 66830 63617
rect 66990 63617 70020 63640
rect 66990 62610 67013 63617
rect 66807 61610 67013 62610
rect 66807 60633 66830 61610
rect 63800 60610 66830 60633
rect 66990 60633 67013 61610
rect 69997 62610 70020 63617
rect 70180 63617 73210 63640
rect 70180 62610 70203 63617
rect 69997 61610 70203 62610
rect 69997 60633 70020 61610
rect 66990 60610 70020 60633
rect 70180 60633 70203 61610
rect 73187 62610 73210 63617
rect 73370 63617 76400 63640
rect 73370 62610 73393 63617
rect 73187 61610 73393 62610
rect 73187 60633 73210 61610
rect 70180 60610 73210 60633
rect 73370 60633 73393 61610
rect 76377 62610 76400 63617
rect 76560 63617 79590 63640
rect 76560 62610 76583 63617
rect 76377 61610 76583 62610
rect 76377 60633 76400 61610
rect 73370 60610 76400 60633
rect 76560 60633 76583 61610
rect 79567 62610 79590 63617
rect 79750 63617 82780 63640
rect 79750 62610 79773 63617
rect 79567 61610 79773 62610
rect 79567 60633 79590 61610
rect 76560 60610 79590 60633
rect 79750 60633 79773 61610
rect 82757 62610 82780 63617
rect 82940 63617 85970 63640
rect 82940 62610 82963 63617
rect 82757 61610 82963 62610
rect 82757 60633 82780 61610
rect 79750 60610 82780 60633
rect 82940 60633 82963 61610
rect 85947 62610 85970 63617
rect 86130 63617 89160 63640
rect 86130 62610 86153 63617
rect 85947 61610 86153 62610
rect 85947 60633 85970 61610
rect 82940 60610 85970 60633
rect 86130 60633 86153 61610
rect 89137 62610 89160 63617
rect 89320 63617 92350 63640
rect 89320 62610 89343 63617
rect 89137 61610 89343 62610
rect 89137 60633 89160 61610
rect 86130 60610 89160 60633
rect 89320 60633 89343 61610
rect 92327 62610 92350 63617
rect 92510 63617 95540 63640
rect 92510 62610 92533 63617
rect 92327 61610 92533 62610
rect 92327 60633 92350 61610
rect 89320 60610 92350 60633
rect 92510 60633 92533 61610
rect 95517 62610 95540 63617
rect 95700 63617 98730 63640
rect 95700 62610 95723 63617
rect 95517 61610 95723 62610
rect 95517 60633 95540 61610
rect 92510 60610 95540 60633
rect 95700 60633 95723 61610
rect 98707 62610 98730 63617
rect 98890 63617 101920 63640
rect 98890 62610 98913 63617
rect 98707 61610 98913 62610
rect 98707 60633 98730 61610
rect 95700 60610 98730 60633
rect 98890 60633 98913 61610
rect 101897 62610 101920 63617
rect 102080 63617 105110 63640
rect 102080 62610 102103 63617
rect 101897 61610 102103 62610
rect 101897 60633 101920 61610
rect 98890 60610 101920 60633
rect 102080 60633 102103 61610
rect 105087 62610 105110 63617
rect 105270 63617 108300 63640
rect 105270 62610 105293 63617
rect 105087 61610 105293 62610
rect 105087 60633 105110 61610
rect 102080 60610 105110 60633
rect 105270 60633 105293 61610
rect 108277 62610 108300 63617
rect 108460 63617 111490 63640
rect 108460 62610 108483 63617
rect 108277 61610 108483 62610
rect 108277 60633 108300 61610
rect 105270 60610 108300 60633
rect 108460 60633 108483 61610
rect 111467 62610 111490 63617
rect 111650 63617 114680 63640
rect 111650 62610 111673 63617
rect 111467 61610 111673 62610
rect 111467 60633 111490 61610
rect 108460 60610 111490 60633
rect 111650 60633 111673 61610
rect 114657 62610 114680 63617
rect 114840 63617 117870 63640
rect 114840 62610 114863 63617
rect 114657 61610 114863 62610
rect 114657 60633 114680 61610
rect 111650 60610 114680 60633
rect 114840 60633 114863 61610
rect 117847 62610 117870 63617
rect 118030 63617 121060 63640
rect 118030 62610 118053 63617
rect 117847 61610 118053 62610
rect 117847 60633 117870 61610
rect 114840 60610 117870 60633
rect 118030 60633 118053 61610
rect 121037 62610 121060 63617
rect 121220 63617 124250 63640
rect 121220 62610 121243 63617
rect 121037 61610 121243 62610
rect 121037 60633 121060 61610
rect 118030 60610 121060 60633
rect 121220 60633 121243 61610
rect 124227 62610 124250 63617
rect 124410 63617 127440 63640
rect 124410 62610 124433 63617
rect 124227 61610 124433 62610
rect 124227 60633 124250 61610
rect 121220 60610 124250 60633
rect 124410 60633 124433 61610
rect 127417 62610 127440 63617
rect 127600 63617 130630 63640
rect 127600 62610 127623 63617
rect 127417 61610 127623 62610
rect 127417 60633 127440 61610
rect 124410 60610 127440 60633
rect 127600 60633 127623 61610
rect 130607 62610 130630 63617
rect 130790 63617 133820 63640
rect 130790 62610 130813 63617
rect 130607 61610 130813 62610
rect 130607 60633 130630 61610
rect 127600 60610 130630 60633
rect 130790 60633 130813 61610
rect 133797 62610 133820 63617
rect 133980 63617 137010 63640
rect 133980 62610 134003 63617
rect 133797 61610 134003 62610
rect 133797 60633 133820 61610
rect 130790 60610 133820 60633
rect 133980 60633 134003 61610
rect 136987 62610 137010 63617
rect 136987 61610 137170 62610
rect 136987 60633 137010 61610
rect 133980 60610 137010 60633
rect 1000 60450 2000 60610
rect 4190 60450 5190 60610
rect 7380 60450 8380 60610
rect 10570 60450 11570 60610
rect 13760 60450 14760 60610
rect 16950 60450 17950 60610
rect 20140 60450 21140 60610
rect 23330 60450 24330 60610
rect 26520 60450 27520 60610
rect 29710 60450 30710 60610
rect 32900 60450 33900 60610
rect 36090 60450 37090 60610
rect 39280 60450 40280 60610
rect 42470 60450 43470 60610
rect 45660 60450 46660 60610
rect 48850 60450 49850 60610
rect 52040 60450 53040 60610
rect 55230 60450 56230 60610
rect 58420 60450 59420 60610
rect 61610 60450 62610 60610
rect 64800 60450 65800 60610
rect 67990 60450 68990 60610
rect 71180 60450 72180 60610
rect 74370 60450 75370 60610
rect 77560 60450 78560 60610
rect 80750 60450 81750 60610
rect 83940 60450 84940 60610
rect 87130 60450 88130 60610
rect 90320 60450 91320 60610
rect 93510 60450 94510 60610
rect 96700 60450 97700 60610
rect 99890 60450 100890 60610
rect 103080 60450 104080 60610
rect 106270 60450 107270 60610
rect 109460 60450 110460 60610
rect 112650 60450 113650 60610
rect 115840 60450 116840 60610
rect 119030 60450 120030 60610
rect 122220 60450 123220 60610
rect 125410 60450 126410 60610
rect 128600 60450 129600 60610
rect 131790 60450 132790 60610
rect 134980 60450 135980 60610
rect 0 60427 3030 60450
rect 0 57443 23 60427
rect 3007 59420 3030 60427
rect 3190 60427 6220 60450
rect 3190 59420 3213 60427
rect 3007 58420 3213 59420
rect 3007 57443 3030 58420
rect 0 57420 3030 57443
rect 3190 57443 3213 58420
rect 6197 59420 6220 60427
rect 6380 60427 9410 60450
rect 6380 59420 6403 60427
rect 6197 58420 6403 59420
rect 6197 57443 6220 58420
rect 3190 57420 6220 57443
rect 6380 57443 6403 58420
rect 9387 59420 9410 60427
rect 9570 60427 12600 60450
rect 9570 59420 9593 60427
rect 9387 58420 9593 59420
rect 9387 57443 9410 58420
rect 6380 57420 9410 57443
rect 9570 57443 9593 58420
rect 12577 59420 12600 60427
rect 12760 60427 15790 60450
rect 12760 59420 12783 60427
rect 12577 58420 12783 59420
rect 12577 57443 12600 58420
rect 9570 57420 12600 57443
rect 12760 57443 12783 58420
rect 15767 59420 15790 60427
rect 15950 60427 18980 60450
rect 15950 59420 15973 60427
rect 15767 58420 15973 59420
rect 15767 57443 15790 58420
rect 12760 57420 15790 57443
rect 15950 57443 15973 58420
rect 18957 59420 18980 60427
rect 19140 60427 22170 60450
rect 19140 59420 19163 60427
rect 18957 58420 19163 59420
rect 18957 57443 18980 58420
rect 15950 57420 18980 57443
rect 19140 57443 19163 58420
rect 22147 59420 22170 60427
rect 22330 60427 25360 60450
rect 22330 59420 22353 60427
rect 22147 58420 22353 59420
rect 22147 57443 22170 58420
rect 19140 57420 22170 57443
rect 22330 57443 22353 58420
rect 25337 59420 25360 60427
rect 25520 60427 28550 60450
rect 25520 59420 25543 60427
rect 25337 58420 25543 59420
rect 25337 57443 25360 58420
rect 22330 57420 25360 57443
rect 25520 57443 25543 58420
rect 28527 59420 28550 60427
rect 28710 60427 31740 60450
rect 28710 59420 28733 60427
rect 28527 58420 28733 59420
rect 28527 57443 28550 58420
rect 25520 57420 28550 57443
rect 28710 57443 28733 58420
rect 31717 59420 31740 60427
rect 31900 60427 34930 60450
rect 31900 59420 31923 60427
rect 31717 58420 31923 59420
rect 31717 57443 31740 58420
rect 28710 57420 31740 57443
rect 31900 57443 31923 58420
rect 34907 59420 34930 60427
rect 35090 60427 38120 60450
rect 35090 59420 35113 60427
rect 34907 58420 35113 59420
rect 34907 57443 34930 58420
rect 31900 57420 34930 57443
rect 35090 57443 35113 58420
rect 38097 59420 38120 60427
rect 38280 60427 41310 60450
rect 38280 59420 38303 60427
rect 38097 58420 38303 59420
rect 38097 57443 38120 58420
rect 35090 57420 38120 57443
rect 38280 57443 38303 58420
rect 41287 59420 41310 60427
rect 41470 60427 44500 60450
rect 41470 59420 41493 60427
rect 41287 58420 41493 59420
rect 41287 57443 41310 58420
rect 38280 57420 41310 57443
rect 41470 57443 41493 58420
rect 44477 59420 44500 60427
rect 44660 60427 47690 60450
rect 44660 59420 44683 60427
rect 44477 58420 44683 59420
rect 44477 57443 44500 58420
rect 41470 57420 44500 57443
rect 44660 57443 44683 58420
rect 47667 59420 47690 60427
rect 47850 60427 50880 60450
rect 47850 59420 47873 60427
rect 47667 58420 47873 59420
rect 47667 57443 47690 58420
rect 44660 57420 47690 57443
rect 47850 57443 47873 58420
rect 50857 59420 50880 60427
rect 51040 60427 54070 60450
rect 51040 59420 51063 60427
rect 50857 58420 51063 59420
rect 50857 57443 50880 58420
rect 47850 57420 50880 57443
rect 51040 57443 51063 58420
rect 54047 59420 54070 60427
rect 54230 60427 57260 60450
rect 54230 59420 54253 60427
rect 54047 58420 54253 59420
rect 54047 57443 54070 58420
rect 51040 57420 54070 57443
rect 54230 57443 54253 58420
rect 57237 59420 57260 60427
rect 57420 60427 60450 60450
rect 57420 59420 57443 60427
rect 57237 58420 57443 59420
rect 57237 57443 57260 58420
rect 54230 57420 57260 57443
rect 57420 57443 57443 58420
rect 60427 59420 60450 60427
rect 60610 60427 63640 60450
rect 60610 59420 60633 60427
rect 60427 58420 60633 59420
rect 60427 57443 60450 58420
rect 57420 57420 60450 57443
rect 60610 57443 60633 58420
rect 63617 59420 63640 60427
rect 63800 60427 66830 60450
rect 63800 59420 63823 60427
rect 63617 58420 63823 59420
rect 63617 57443 63640 58420
rect 60610 57420 63640 57443
rect 63800 57443 63823 58420
rect 66807 59420 66830 60427
rect 66990 60427 70020 60450
rect 66990 59420 67013 60427
rect 66807 58420 67013 59420
rect 66807 57443 66830 58420
rect 63800 57420 66830 57443
rect 66990 57443 67013 58420
rect 69997 59420 70020 60427
rect 70180 60427 73210 60450
rect 70180 59420 70203 60427
rect 69997 58420 70203 59420
rect 69997 57443 70020 58420
rect 66990 57420 70020 57443
rect 70180 57443 70203 58420
rect 73187 59420 73210 60427
rect 73370 60427 76400 60450
rect 73370 59420 73393 60427
rect 73187 58420 73393 59420
rect 73187 57443 73210 58420
rect 70180 57420 73210 57443
rect 73370 57443 73393 58420
rect 76377 59420 76400 60427
rect 76560 60427 79590 60450
rect 76560 59420 76583 60427
rect 76377 58420 76583 59420
rect 76377 57443 76400 58420
rect 73370 57420 76400 57443
rect 76560 57443 76583 58420
rect 79567 59420 79590 60427
rect 79750 60427 82780 60450
rect 79750 59420 79773 60427
rect 79567 58420 79773 59420
rect 79567 57443 79590 58420
rect 76560 57420 79590 57443
rect 79750 57443 79773 58420
rect 82757 59420 82780 60427
rect 82940 60427 85970 60450
rect 82940 59420 82963 60427
rect 82757 58420 82963 59420
rect 82757 57443 82780 58420
rect 79750 57420 82780 57443
rect 82940 57443 82963 58420
rect 85947 59420 85970 60427
rect 86130 60427 89160 60450
rect 86130 59420 86153 60427
rect 85947 58420 86153 59420
rect 85947 57443 85970 58420
rect 82940 57420 85970 57443
rect 86130 57443 86153 58420
rect 89137 59420 89160 60427
rect 89320 60427 92350 60450
rect 89320 59420 89343 60427
rect 89137 58420 89343 59420
rect 89137 57443 89160 58420
rect 86130 57420 89160 57443
rect 89320 57443 89343 58420
rect 92327 59420 92350 60427
rect 92510 60427 95540 60450
rect 92510 59420 92533 60427
rect 92327 58420 92533 59420
rect 92327 57443 92350 58420
rect 89320 57420 92350 57443
rect 92510 57443 92533 58420
rect 95517 59420 95540 60427
rect 95700 60427 98730 60450
rect 95700 59420 95723 60427
rect 95517 58420 95723 59420
rect 95517 57443 95540 58420
rect 92510 57420 95540 57443
rect 95700 57443 95723 58420
rect 98707 59420 98730 60427
rect 98890 60427 101920 60450
rect 98890 59420 98913 60427
rect 98707 58420 98913 59420
rect 98707 57443 98730 58420
rect 95700 57420 98730 57443
rect 98890 57443 98913 58420
rect 101897 59420 101920 60427
rect 102080 60427 105110 60450
rect 102080 59420 102103 60427
rect 101897 58420 102103 59420
rect 101897 57443 101920 58420
rect 98890 57420 101920 57443
rect 102080 57443 102103 58420
rect 105087 59420 105110 60427
rect 105270 60427 108300 60450
rect 105270 59420 105293 60427
rect 105087 58420 105293 59420
rect 105087 57443 105110 58420
rect 102080 57420 105110 57443
rect 105270 57443 105293 58420
rect 108277 59420 108300 60427
rect 108460 60427 111490 60450
rect 108460 59420 108483 60427
rect 108277 58420 108483 59420
rect 108277 57443 108300 58420
rect 105270 57420 108300 57443
rect 108460 57443 108483 58420
rect 111467 59420 111490 60427
rect 111650 60427 114680 60450
rect 111650 59420 111673 60427
rect 111467 58420 111673 59420
rect 111467 57443 111490 58420
rect 108460 57420 111490 57443
rect 111650 57443 111673 58420
rect 114657 59420 114680 60427
rect 114840 60427 117870 60450
rect 114840 59420 114863 60427
rect 114657 58420 114863 59420
rect 114657 57443 114680 58420
rect 111650 57420 114680 57443
rect 114840 57443 114863 58420
rect 117847 59420 117870 60427
rect 118030 60427 121060 60450
rect 118030 59420 118053 60427
rect 117847 58420 118053 59420
rect 117847 57443 117870 58420
rect 114840 57420 117870 57443
rect 118030 57443 118053 58420
rect 121037 59420 121060 60427
rect 121220 60427 124250 60450
rect 121220 59420 121243 60427
rect 121037 58420 121243 59420
rect 121037 57443 121060 58420
rect 118030 57420 121060 57443
rect 121220 57443 121243 58420
rect 124227 59420 124250 60427
rect 124410 60427 127440 60450
rect 124410 59420 124433 60427
rect 124227 58420 124433 59420
rect 124227 57443 124250 58420
rect 121220 57420 124250 57443
rect 124410 57443 124433 58420
rect 127417 59420 127440 60427
rect 127600 60427 130630 60450
rect 127600 59420 127623 60427
rect 127417 58420 127623 59420
rect 127417 57443 127440 58420
rect 124410 57420 127440 57443
rect 127600 57443 127623 58420
rect 130607 59420 130630 60427
rect 130790 60427 133820 60450
rect 130790 59420 130813 60427
rect 130607 58420 130813 59420
rect 130607 57443 130630 58420
rect 127600 57420 130630 57443
rect 130790 57443 130813 58420
rect 133797 59420 133820 60427
rect 133980 60427 137010 60450
rect 133980 59420 134003 60427
rect 133797 58420 134003 59420
rect 133797 57443 133820 58420
rect 130790 57420 133820 57443
rect 133980 57443 134003 58420
rect 136987 59420 137010 60427
rect 136987 58420 137170 59420
rect 136987 57443 137010 58420
rect 133980 57420 137010 57443
rect 1000 57260 2000 57420
rect 4190 57260 5190 57420
rect 7380 57260 8380 57420
rect 10570 57260 11570 57420
rect 13760 57260 14760 57420
rect 16950 57260 17950 57420
rect 20140 57260 21140 57420
rect 23330 57260 24330 57420
rect 26520 57260 27520 57420
rect 29710 57260 30710 57420
rect 32900 57260 33900 57420
rect 36090 57260 37090 57420
rect 39280 57260 40280 57420
rect 42470 57260 43470 57420
rect 45660 57260 46660 57420
rect 48850 57260 49850 57420
rect 52040 57260 53040 57420
rect 55230 57260 56230 57420
rect 58420 57260 59420 57420
rect 61610 57260 62610 57420
rect 64800 57260 65800 57420
rect 67990 57260 68990 57420
rect 71180 57260 72180 57420
rect 74370 57260 75370 57420
rect 77560 57260 78560 57420
rect 80750 57260 81750 57420
rect 83940 57260 84940 57420
rect 87130 57260 88130 57420
rect 90320 57260 91320 57420
rect 93510 57260 94510 57420
rect 96700 57260 97700 57420
rect 99890 57260 100890 57420
rect 103080 57260 104080 57420
rect 106270 57260 107270 57420
rect 109460 57260 110460 57420
rect 112650 57260 113650 57420
rect 115840 57260 116840 57420
rect 119030 57260 120030 57420
rect 122220 57260 123220 57420
rect 125410 57260 126410 57420
rect 128600 57260 129600 57420
rect 131790 57260 132790 57420
rect 134980 57260 135980 57420
rect 0 57237 3030 57260
rect 0 54253 23 57237
rect 3007 56230 3030 57237
rect 3190 57237 6220 57260
rect 3190 56230 3213 57237
rect 3007 55230 3213 56230
rect 3007 54253 3030 55230
rect 0 54230 3030 54253
rect 3190 54253 3213 55230
rect 6197 56230 6220 57237
rect 6380 57237 9410 57260
rect 6380 56230 6403 57237
rect 6197 55230 6403 56230
rect 6197 54253 6220 55230
rect 3190 54230 6220 54253
rect 6380 54253 6403 55230
rect 9387 56230 9410 57237
rect 9570 57237 12600 57260
rect 9570 56230 9593 57237
rect 9387 55230 9593 56230
rect 9387 54253 9410 55230
rect 6380 54230 9410 54253
rect 9570 54253 9593 55230
rect 12577 56230 12600 57237
rect 12760 57237 15790 57260
rect 12760 56230 12783 57237
rect 12577 55230 12783 56230
rect 12577 54253 12600 55230
rect 9570 54230 12600 54253
rect 12760 54253 12783 55230
rect 15767 56230 15790 57237
rect 15950 57237 18980 57260
rect 15950 56230 15973 57237
rect 15767 55230 15973 56230
rect 15767 54253 15790 55230
rect 12760 54230 15790 54253
rect 15950 54253 15973 55230
rect 18957 56230 18980 57237
rect 19140 57237 22170 57260
rect 19140 56230 19163 57237
rect 18957 55230 19163 56230
rect 18957 54253 18980 55230
rect 15950 54230 18980 54253
rect 19140 54253 19163 55230
rect 22147 56230 22170 57237
rect 22330 57237 25360 57260
rect 22330 56230 22353 57237
rect 22147 55230 22353 56230
rect 22147 54253 22170 55230
rect 19140 54230 22170 54253
rect 22330 54253 22353 55230
rect 25337 56230 25360 57237
rect 25520 57237 28550 57260
rect 25520 56230 25543 57237
rect 25337 55230 25543 56230
rect 25337 54253 25360 55230
rect 22330 54230 25360 54253
rect 25520 54253 25543 55230
rect 28527 56230 28550 57237
rect 28710 57237 31740 57260
rect 28710 56230 28733 57237
rect 28527 55230 28733 56230
rect 28527 54253 28550 55230
rect 25520 54230 28550 54253
rect 28710 54253 28733 55230
rect 31717 56230 31740 57237
rect 31900 57237 34930 57260
rect 31900 56230 31923 57237
rect 31717 55230 31923 56230
rect 31717 54253 31740 55230
rect 28710 54230 31740 54253
rect 31900 54253 31923 55230
rect 34907 56230 34930 57237
rect 35090 57237 38120 57260
rect 35090 56230 35113 57237
rect 34907 55230 35113 56230
rect 34907 54253 34930 55230
rect 31900 54230 34930 54253
rect 35090 54253 35113 55230
rect 38097 56230 38120 57237
rect 38280 57237 41310 57260
rect 38280 56230 38303 57237
rect 38097 55230 38303 56230
rect 38097 54253 38120 55230
rect 35090 54230 38120 54253
rect 38280 54253 38303 55230
rect 41287 56230 41310 57237
rect 41470 57237 44500 57260
rect 41470 56230 41493 57237
rect 41287 55230 41493 56230
rect 41287 54253 41310 55230
rect 38280 54230 41310 54253
rect 41470 54253 41493 55230
rect 44477 56230 44500 57237
rect 44660 57237 47690 57260
rect 44660 56230 44683 57237
rect 44477 55230 44683 56230
rect 44477 54253 44500 55230
rect 41470 54230 44500 54253
rect 44660 54253 44683 55230
rect 47667 56230 47690 57237
rect 47850 57237 50880 57260
rect 47850 56230 47873 57237
rect 47667 55230 47873 56230
rect 47667 54253 47690 55230
rect 44660 54230 47690 54253
rect 47850 54253 47873 55230
rect 50857 56230 50880 57237
rect 51040 57237 54070 57260
rect 51040 56230 51063 57237
rect 50857 55230 51063 56230
rect 50857 54253 50880 55230
rect 47850 54230 50880 54253
rect 51040 54253 51063 55230
rect 54047 56230 54070 57237
rect 54230 57237 57260 57260
rect 54230 56230 54253 57237
rect 54047 55230 54253 56230
rect 54047 54253 54070 55230
rect 51040 54230 54070 54253
rect 54230 54253 54253 55230
rect 57237 56230 57260 57237
rect 57420 57237 60450 57260
rect 57420 56230 57443 57237
rect 57237 55230 57443 56230
rect 57237 54253 57260 55230
rect 54230 54230 57260 54253
rect 57420 54253 57443 55230
rect 60427 56230 60450 57237
rect 60610 57237 63640 57260
rect 60610 56230 60633 57237
rect 60427 55230 60633 56230
rect 60427 54253 60450 55230
rect 57420 54230 60450 54253
rect 60610 54253 60633 55230
rect 63617 56230 63640 57237
rect 63800 57237 66830 57260
rect 63800 56230 63823 57237
rect 63617 55230 63823 56230
rect 63617 54253 63640 55230
rect 60610 54230 63640 54253
rect 63800 54253 63823 55230
rect 66807 56230 66830 57237
rect 66990 57237 70020 57260
rect 66990 56230 67013 57237
rect 66807 55230 67013 56230
rect 66807 54253 66830 55230
rect 63800 54230 66830 54253
rect 66990 54253 67013 55230
rect 69997 56230 70020 57237
rect 70180 57237 73210 57260
rect 70180 56230 70203 57237
rect 69997 55230 70203 56230
rect 69997 54253 70020 55230
rect 66990 54230 70020 54253
rect 70180 54253 70203 55230
rect 73187 56230 73210 57237
rect 73370 57237 76400 57260
rect 73370 56230 73393 57237
rect 73187 55230 73393 56230
rect 73187 54253 73210 55230
rect 70180 54230 73210 54253
rect 73370 54253 73393 55230
rect 76377 56230 76400 57237
rect 76560 57237 79590 57260
rect 76560 56230 76583 57237
rect 76377 55230 76583 56230
rect 76377 54253 76400 55230
rect 73370 54230 76400 54253
rect 76560 54253 76583 55230
rect 79567 56230 79590 57237
rect 79750 57237 82780 57260
rect 79750 56230 79773 57237
rect 79567 55230 79773 56230
rect 79567 54253 79590 55230
rect 76560 54230 79590 54253
rect 79750 54253 79773 55230
rect 82757 56230 82780 57237
rect 82940 57237 85970 57260
rect 82940 56230 82963 57237
rect 82757 55230 82963 56230
rect 82757 54253 82780 55230
rect 79750 54230 82780 54253
rect 82940 54253 82963 55230
rect 85947 56230 85970 57237
rect 86130 57237 89160 57260
rect 86130 56230 86153 57237
rect 85947 55230 86153 56230
rect 85947 54253 85970 55230
rect 82940 54230 85970 54253
rect 86130 54253 86153 55230
rect 89137 56230 89160 57237
rect 89320 57237 92350 57260
rect 89320 56230 89343 57237
rect 89137 55230 89343 56230
rect 89137 54253 89160 55230
rect 86130 54230 89160 54253
rect 89320 54253 89343 55230
rect 92327 56230 92350 57237
rect 92510 57237 95540 57260
rect 92510 56230 92533 57237
rect 92327 55230 92533 56230
rect 92327 54253 92350 55230
rect 89320 54230 92350 54253
rect 92510 54253 92533 55230
rect 95517 56230 95540 57237
rect 95700 57237 98730 57260
rect 95700 56230 95723 57237
rect 95517 55230 95723 56230
rect 95517 54253 95540 55230
rect 92510 54230 95540 54253
rect 95700 54253 95723 55230
rect 98707 56230 98730 57237
rect 98890 57237 101920 57260
rect 98890 56230 98913 57237
rect 98707 55230 98913 56230
rect 98707 54253 98730 55230
rect 95700 54230 98730 54253
rect 98890 54253 98913 55230
rect 101897 56230 101920 57237
rect 102080 57237 105110 57260
rect 102080 56230 102103 57237
rect 101897 55230 102103 56230
rect 101897 54253 101920 55230
rect 98890 54230 101920 54253
rect 102080 54253 102103 55230
rect 105087 56230 105110 57237
rect 105270 57237 108300 57260
rect 105270 56230 105293 57237
rect 105087 55230 105293 56230
rect 105087 54253 105110 55230
rect 102080 54230 105110 54253
rect 105270 54253 105293 55230
rect 108277 56230 108300 57237
rect 108460 57237 111490 57260
rect 108460 56230 108483 57237
rect 108277 55230 108483 56230
rect 108277 54253 108300 55230
rect 105270 54230 108300 54253
rect 108460 54253 108483 55230
rect 111467 56230 111490 57237
rect 111650 57237 114680 57260
rect 111650 56230 111673 57237
rect 111467 55230 111673 56230
rect 111467 54253 111490 55230
rect 108460 54230 111490 54253
rect 111650 54253 111673 55230
rect 114657 56230 114680 57237
rect 114840 57237 117870 57260
rect 114840 56230 114863 57237
rect 114657 55230 114863 56230
rect 114657 54253 114680 55230
rect 111650 54230 114680 54253
rect 114840 54253 114863 55230
rect 117847 56230 117870 57237
rect 118030 57237 121060 57260
rect 118030 56230 118053 57237
rect 117847 55230 118053 56230
rect 117847 54253 117870 55230
rect 114840 54230 117870 54253
rect 118030 54253 118053 55230
rect 121037 56230 121060 57237
rect 121220 57237 124250 57260
rect 121220 56230 121243 57237
rect 121037 55230 121243 56230
rect 121037 54253 121060 55230
rect 118030 54230 121060 54253
rect 121220 54253 121243 55230
rect 124227 56230 124250 57237
rect 124410 57237 127440 57260
rect 124410 56230 124433 57237
rect 124227 55230 124433 56230
rect 124227 54253 124250 55230
rect 121220 54230 124250 54253
rect 124410 54253 124433 55230
rect 127417 56230 127440 57237
rect 127600 57237 130630 57260
rect 127600 56230 127623 57237
rect 127417 55230 127623 56230
rect 127417 54253 127440 55230
rect 124410 54230 127440 54253
rect 127600 54253 127623 55230
rect 130607 56230 130630 57237
rect 130790 57237 133820 57260
rect 130790 56230 130813 57237
rect 130607 55230 130813 56230
rect 130607 54253 130630 55230
rect 127600 54230 130630 54253
rect 130790 54253 130813 55230
rect 133797 56230 133820 57237
rect 133980 57237 137010 57260
rect 133980 56230 134003 57237
rect 133797 55230 134003 56230
rect 133797 54253 133820 55230
rect 130790 54230 133820 54253
rect 133980 54253 134003 55230
rect 136987 56230 137010 57237
rect 136987 55230 137170 56230
rect 136987 54253 137010 55230
rect 133980 54230 137010 54253
rect 1000 54070 2000 54230
rect 4190 54070 5190 54230
rect 7380 54070 8380 54230
rect 10570 54070 11570 54230
rect 13760 54070 14760 54230
rect 16950 54070 17950 54230
rect 20140 54070 21140 54230
rect 23330 54070 24330 54230
rect 26520 54070 27520 54230
rect 29710 54070 30710 54230
rect 32900 54070 33900 54230
rect 36090 54070 37090 54230
rect 39280 54070 40280 54230
rect 42470 54070 43470 54230
rect 45660 54070 46660 54230
rect 48850 54070 49850 54230
rect 52040 54070 53040 54230
rect 55230 54070 56230 54230
rect 58420 54070 59420 54230
rect 61610 54070 62610 54230
rect 64800 54070 65800 54230
rect 67990 54070 68990 54230
rect 71180 54070 72180 54230
rect 74370 54070 75370 54230
rect 77560 54070 78560 54230
rect 80750 54070 81750 54230
rect 83940 54070 84940 54230
rect 87130 54070 88130 54230
rect 90320 54070 91320 54230
rect 93510 54070 94510 54230
rect 96700 54070 97700 54230
rect 99890 54070 100890 54230
rect 103080 54070 104080 54230
rect 106270 54070 107270 54230
rect 109460 54070 110460 54230
rect 112650 54070 113650 54230
rect 115840 54070 116840 54230
rect 119030 54070 120030 54230
rect 122220 54070 123220 54230
rect 125410 54070 126410 54230
rect 128600 54070 129600 54230
rect 131790 54070 132790 54230
rect 134980 54070 135980 54230
rect 0 54047 3030 54070
rect 0 51063 23 54047
rect 3007 53040 3030 54047
rect 3190 54047 6220 54070
rect 3190 53040 3213 54047
rect 3007 52040 3213 53040
rect 3007 51063 3030 52040
rect 0 51040 3030 51063
rect 3190 51063 3213 52040
rect 6197 53040 6220 54047
rect 6380 54047 9410 54070
rect 6380 53040 6403 54047
rect 6197 52040 6403 53040
rect 6197 51063 6220 52040
rect 3190 51040 6220 51063
rect 6380 51063 6403 52040
rect 9387 53040 9410 54047
rect 9570 54047 12600 54070
rect 9570 53040 9593 54047
rect 9387 52040 9593 53040
rect 9387 51063 9410 52040
rect 6380 51040 9410 51063
rect 9570 51063 9593 52040
rect 12577 53040 12600 54047
rect 12760 54047 15790 54070
rect 12760 53040 12783 54047
rect 12577 52040 12783 53040
rect 12577 51063 12600 52040
rect 9570 51040 12600 51063
rect 12760 51063 12783 52040
rect 15767 53040 15790 54047
rect 15950 54047 18980 54070
rect 15950 53040 15973 54047
rect 15767 52040 15973 53040
rect 15767 51063 15790 52040
rect 12760 51040 15790 51063
rect 15950 51063 15973 52040
rect 18957 53040 18980 54047
rect 19140 54047 22170 54070
rect 19140 53040 19163 54047
rect 18957 52040 19163 53040
rect 18957 51063 18980 52040
rect 15950 51040 18980 51063
rect 19140 51063 19163 52040
rect 22147 53040 22170 54047
rect 22330 54047 25360 54070
rect 22330 53040 22353 54047
rect 22147 52040 22353 53040
rect 22147 51063 22170 52040
rect 19140 51040 22170 51063
rect 22330 51063 22353 52040
rect 25337 53040 25360 54047
rect 25520 54047 28550 54070
rect 25520 53040 25543 54047
rect 25337 52040 25543 53040
rect 25337 51063 25360 52040
rect 22330 51040 25360 51063
rect 25520 51063 25543 52040
rect 28527 53040 28550 54047
rect 28710 54047 31740 54070
rect 28710 53040 28733 54047
rect 28527 52040 28733 53040
rect 28527 51063 28550 52040
rect 25520 51040 28550 51063
rect 28710 51063 28733 52040
rect 31717 53040 31740 54047
rect 31900 54047 34930 54070
rect 31900 53040 31923 54047
rect 31717 52040 31923 53040
rect 31717 51063 31740 52040
rect 28710 51040 31740 51063
rect 31900 51063 31923 52040
rect 34907 53040 34930 54047
rect 35090 54047 38120 54070
rect 35090 53040 35113 54047
rect 34907 52040 35113 53040
rect 34907 51063 34930 52040
rect 31900 51040 34930 51063
rect 35090 51063 35113 52040
rect 38097 53040 38120 54047
rect 38280 54047 41310 54070
rect 38280 53040 38303 54047
rect 38097 52040 38303 53040
rect 38097 51063 38120 52040
rect 35090 51040 38120 51063
rect 38280 51063 38303 52040
rect 41287 53040 41310 54047
rect 41470 54047 44500 54070
rect 41470 53040 41493 54047
rect 41287 52040 41493 53040
rect 41287 51063 41310 52040
rect 38280 51040 41310 51063
rect 41470 51063 41493 52040
rect 44477 53040 44500 54047
rect 44660 54047 47690 54070
rect 44660 53040 44683 54047
rect 44477 52040 44683 53040
rect 44477 51063 44500 52040
rect 41470 51040 44500 51063
rect 44660 51063 44683 52040
rect 47667 53040 47690 54047
rect 47850 54047 50880 54070
rect 47850 53040 47873 54047
rect 47667 52040 47873 53040
rect 47667 51063 47690 52040
rect 44660 51040 47690 51063
rect 47850 51063 47873 52040
rect 50857 53040 50880 54047
rect 51040 54047 54070 54070
rect 51040 53040 51063 54047
rect 50857 52040 51063 53040
rect 50857 51063 50880 52040
rect 47850 51040 50880 51063
rect 51040 51063 51063 52040
rect 54047 53040 54070 54047
rect 54230 54047 57260 54070
rect 54230 53040 54253 54047
rect 54047 52040 54253 53040
rect 54047 51063 54070 52040
rect 51040 51040 54070 51063
rect 54230 51063 54253 52040
rect 57237 53040 57260 54047
rect 57420 54047 60450 54070
rect 57420 53040 57443 54047
rect 57237 52040 57443 53040
rect 57237 51063 57260 52040
rect 54230 51040 57260 51063
rect 57420 51063 57443 52040
rect 60427 53040 60450 54047
rect 60610 54047 63640 54070
rect 60610 53040 60633 54047
rect 60427 52040 60633 53040
rect 60427 51063 60450 52040
rect 57420 51040 60450 51063
rect 60610 51063 60633 52040
rect 63617 53040 63640 54047
rect 63800 54047 66830 54070
rect 63800 53040 63823 54047
rect 63617 52040 63823 53040
rect 63617 51063 63640 52040
rect 60610 51040 63640 51063
rect 63800 51063 63823 52040
rect 66807 53040 66830 54047
rect 66990 54047 70020 54070
rect 66990 53040 67013 54047
rect 66807 52040 67013 53040
rect 66807 51063 66830 52040
rect 63800 51040 66830 51063
rect 66990 51063 67013 52040
rect 69997 53040 70020 54047
rect 70180 54047 73210 54070
rect 70180 53040 70203 54047
rect 69997 52040 70203 53040
rect 69997 51063 70020 52040
rect 66990 51040 70020 51063
rect 70180 51063 70203 52040
rect 73187 53040 73210 54047
rect 73370 54047 76400 54070
rect 73370 53040 73393 54047
rect 73187 52040 73393 53040
rect 73187 51063 73210 52040
rect 70180 51040 73210 51063
rect 73370 51063 73393 52040
rect 76377 53040 76400 54047
rect 76560 54047 79590 54070
rect 76560 53040 76583 54047
rect 76377 52040 76583 53040
rect 76377 51063 76400 52040
rect 73370 51040 76400 51063
rect 76560 51063 76583 52040
rect 79567 53040 79590 54047
rect 79750 54047 82780 54070
rect 79750 53040 79773 54047
rect 79567 52040 79773 53040
rect 79567 51063 79590 52040
rect 76560 51040 79590 51063
rect 79750 51063 79773 52040
rect 82757 53040 82780 54047
rect 82940 54047 85970 54070
rect 82940 53040 82963 54047
rect 82757 52040 82963 53040
rect 82757 51063 82780 52040
rect 79750 51040 82780 51063
rect 82940 51063 82963 52040
rect 85947 53040 85970 54047
rect 86130 54047 89160 54070
rect 86130 53040 86153 54047
rect 85947 52040 86153 53040
rect 85947 51063 85970 52040
rect 82940 51040 85970 51063
rect 86130 51063 86153 52040
rect 89137 53040 89160 54047
rect 89320 54047 92350 54070
rect 89320 53040 89343 54047
rect 89137 52040 89343 53040
rect 89137 51063 89160 52040
rect 86130 51040 89160 51063
rect 89320 51063 89343 52040
rect 92327 53040 92350 54047
rect 92510 54047 95540 54070
rect 92510 53040 92533 54047
rect 92327 52040 92533 53040
rect 92327 51063 92350 52040
rect 89320 51040 92350 51063
rect 92510 51063 92533 52040
rect 95517 53040 95540 54047
rect 95700 54047 98730 54070
rect 95700 53040 95723 54047
rect 95517 52040 95723 53040
rect 95517 51063 95540 52040
rect 92510 51040 95540 51063
rect 95700 51063 95723 52040
rect 98707 53040 98730 54047
rect 98890 54047 101920 54070
rect 98890 53040 98913 54047
rect 98707 52040 98913 53040
rect 98707 51063 98730 52040
rect 95700 51040 98730 51063
rect 98890 51063 98913 52040
rect 101897 53040 101920 54047
rect 102080 54047 105110 54070
rect 102080 53040 102103 54047
rect 101897 52040 102103 53040
rect 101897 51063 101920 52040
rect 98890 51040 101920 51063
rect 102080 51063 102103 52040
rect 105087 53040 105110 54047
rect 105270 54047 108300 54070
rect 105270 53040 105293 54047
rect 105087 52040 105293 53040
rect 105087 51063 105110 52040
rect 102080 51040 105110 51063
rect 105270 51063 105293 52040
rect 108277 53040 108300 54047
rect 108460 54047 111490 54070
rect 108460 53040 108483 54047
rect 108277 52040 108483 53040
rect 108277 51063 108300 52040
rect 105270 51040 108300 51063
rect 108460 51063 108483 52040
rect 111467 53040 111490 54047
rect 111650 54047 114680 54070
rect 111650 53040 111673 54047
rect 111467 52040 111673 53040
rect 111467 51063 111490 52040
rect 108460 51040 111490 51063
rect 111650 51063 111673 52040
rect 114657 53040 114680 54047
rect 114840 54047 117870 54070
rect 114840 53040 114863 54047
rect 114657 52040 114863 53040
rect 114657 51063 114680 52040
rect 111650 51040 114680 51063
rect 114840 51063 114863 52040
rect 117847 53040 117870 54047
rect 118030 54047 121060 54070
rect 118030 53040 118053 54047
rect 117847 52040 118053 53040
rect 117847 51063 117870 52040
rect 114840 51040 117870 51063
rect 118030 51063 118053 52040
rect 121037 53040 121060 54047
rect 121220 54047 124250 54070
rect 121220 53040 121243 54047
rect 121037 52040 121243 53040
rect 121037 51063 121060 52040
rect 118030 51040 121060 51063
rect 121220 51063 121243 52040
rect 124227 53040 124250 54047
rect 124410 54047 127440 54070
rect 124410 53040 124433 54047
rect 124227 52040 124433 53040
rect 124227 51063 124250 52040
rect 121220 51040 124250 51063
rect 124410 51063 124433 52040
rect 127417 53040 127440 54047
rect 127600 54047 130630 54070
rect 127600 53040 127623 54047
rect 127417 52040 127623 53040
rect 127417 51063 127440 52040
rect 124410 51040 127440 51063
rect 127600 51063 127623 52040
rect 130607 53040 130630 54047
rect 130790 54047 133820 54070
rect 130790 53040 130813 54047
rect 130607 52040 130813 53040
rect 130607 51063 130630 52040
rect 127600 51040 130630 51063
rect 130790 51063 130813 52040
rect 133797 53040 133820 54047
rect 133980 54047 137010 54070
rect 133980 53040 134003 54047
rect 133797 52040 134003 53040
rect 133797 51063 133820 52040
rect 130790 51040 133820 51063
rect 133980 51063 134003 52040
rect 136987 53040 137010 54047
rect 136987 52040 137170 53040
rect 136987 51063 137010 52040
rect 133980 51040 137010 51063
rect 1000 50880 2000 51040
rect 4190 50880 5190 51040
rect 7380 50880 8380 51040
rect 10570 50880 11570 51040
rect 13760 50880 14760 51040
rect 16950 50880 17950 51040
rect 20140 50880 21140 51040
rect 23330 50880 24330 51040
rect 26520 50880 27520 51040
rect 29710 50880 30710 51040
rect 32900 50880 33900 51040
rect 36090 50880 37090 51040
rect 39280 50880 40280 51040
rect 42470 50880 43470 51040
rect 45660 50880 46660 51040
rect 48850 50880 49850 51040
rect 52040 50880 53040 51040
rect 55230 50880 56230 51040
rect 58420 50880 59420 51040
rect 61610 50880 62610 51040
rect 64800 50880 65800 51040
rect 67990 50880 68990 51040
rect 71180 50880 72180 51040
rect 74370 50880 75370 51040
rect 77560 50880 78560 51040
rect 80750 50880 81750 51040
rect 83940 50880 84940 51040
rect 87130 50880 88130 51040
rect 90320 50880 91320 51040
rect 93510 50880 94510 51040
rect 96700 50880 97700 51040
rect 99890 50880 100890 51040
rect 103080 50880 104080 51040
rect 106270 50880 107270 51040
rect 109460 50880 110460 51040
rect 112650 50880 113650 51040
rect 115840 50880 116840 51040
rect 119030 50880 120030 51040
rect 122220 50880 123220 51040
rect 125410 50880 126410 51040
rect 128600 50880 129600 51040
rect 131790 50880 132790 51040
rect 134980 50880 135980 51040
rect 0 50857 3030 50880
rect 0 47873 23 50857
rect 3007 49850 3030 50857
rect 3190 50857 6220 50880
rect 3190 49850 3213 50857
rect 3007 48850 3213 49850
rect 3007 47873 3030 48850
rect 0 47850 3030 47873
rect 3190 47873 3213 48850
rect 6197 49850 6220 50857
rect 6380 50857 9410 50880
rect 6380 49850 6403 50857
rect 6197 48850 6403 49850
rect 6197 47873 6220 48850
rect 3190 47850 6220 47873
rect 6380 47873 6403 48850
rect 9387 49850 9410 50857
rect 9570 50857 12600 50880
rect 9570 49850 9593 50857
rect 9387 48850 9593 49850
rect 9387 47873 9410 48850
rect 6380 47850 9410 47873
rect 9570 47873 9593 48850
rect 12577 49850 12600 50857
rect 12760 50857 15790 50880
rect 12760 49850 12783 50857
rect 12577 48850 12783 49850
rect 12577 47873 12600 48850
rect 9570 47850 12600 47873
rect 12760 47873 12783 48850
rect 15767 49850 15790 50857
rect 15950 50857 18980 50880
rect 15950 49850 15973 50857
rect 15767 48850 15973 49850
rect 15767 47873 15790 48850
rect 12760 47850 15790 47873
rect 15950 47873 15973 48850
rect 18957 49850 18980 50857
rect 19140 50857 22170 50880
rect 19140 49850 19163 50857
rect 18957 48850 19163 49850
rect 18957 47873 18980 48850
rect 15950 47850 18980 47873
rect 19140 47873 19163 48850
rect 22147 49850 22170 50857
rect 22330 50857 25360 50880
rect 22330 49850 22353 50857
rect 22147 48850 22353 49850
rect 22147 47873 22170 48850
rect 19140 47850 22170 47873
rect 22330 47873 22353 48850
rect 25337 49850 25360 50857
rect 25520 50857 28550 50880
rect 25520 49850 25543 50857
rect 25337 48850 25543 49850
rect 25337 47873 25360 48850
rect 22330 47850 25360 47873
rect 25520 47873 25543 48850
rect 28527 49850 28550 50857
rect 28710 50857 31740 50880
rect 28710 49850 28733 50857
rect 28527 48850 28733 49850
rect 28527 47873 28550 48850
rect 25520 47850 28550 47873
rect 28710 47873 28733 48850
rect 31717 49850 31740 50857
rect 31900 50857 34930 50880
rect 31900 49850 31923 50857
rect 31717 48850 31923 49850
rect 31717 47873 31740 48850
rect 28710 47850 31740 47873
rect 31900 47873 31923 48850
rect 34907 49850 34930 50857
rect 35090 50857 38120 50880
rect 35090 49850 35113 50857
rect 34907 48850 35113 49850
rect 34907 47873 34930 48850
rect 31900 47850 34930 47873
rect 35090 47873 35113 48850
rect 38097 49850 38120 50857
rect 38280 50857 41310 50880
rect 38280 49850 38303 50857
rect 38097 48850 38303 49850
rect 38097 47873 38120 48850
rect 35090 47850 38120 47873
rect 38280 47873 38303 48850
rect 41287 49850 41310 50857
rect 41470 50857 44500 50880
rect 41470 49850 41493 50857
rect 41287 48850 41493 49850
rect 41287 47873 41310 48850
rect 38280 47850 41310 47873
rect 41470 47873 41493 48850
rect 44477 49850 44500 50857
rect 44660 50857 47690 50880
rect 44660 49850 44683 50857
rect 44477 48850 44683 49850
rect 44477 47873 44500 48850
rect 41470 47850 44500 47873
rect 44660 47873 44683 48850
rect 47667 49850 47690 50857
rect 47850 50857 50880 50880
rect 47850 49850 47873 50857
rect 47667 48850 47873 49850
rect 47667 47873 47690 48850
rect 44660 47850 47690 47873
rect 47850 47873 47873 48850
rect 50857 49850 50880 50857
rect 51040 50857 54070 50880
rect 51040 49850 51063 50857
rect 50857 48850 51063 49850
rect 50857 47873 50880 48850
rect 47850 47850 50880 47873
rect 51040 47873 51063 48850
rect 54047 49850 54070 50857
rect 54230 50857 57260 50880
rect 54230 49850 54253 50857
rect 54047 48850 54253 49850
rect 54047 47873 54070 48850
rect 51040 47850 54070 47873
rect 54230 47873 54253 48850
rect 57237 49850 57260 50857
rect 57420 50857 60450 50880
rect 57420 49850 57443 50857
rect 57237 48850 57443 49850
rect 57237 47873 57260 48850
rect 54230 47850 57260 47873
rect 57420 47873 57443 48850
rect 60427 49850 60450 50857
rect 60610 50857 63640 50880
rect 60610 49850 60633 50857
rect 60427 48850 60633 49850
rect 60427 47873 60450 48850
rect 57420 47850 60450 47873
rect 60610 47873 60633 48850
rect 63617 49850 63640 50857
rect 63800 50857 66830 50880
rect 63800 49850 63823 50857
rect 63617 48850 63823 49850
rect 63617 47873 63640 48850
rect 60610 47850 63640 47873
rect 63800 47873 63823 48850
rect 66807 49850 66830 50857
rect 66990 50857 70020 50880
rect 66990 49850 67013 50857
rect 66807 48850 67013 49850
rect 66807 47873 66830 48850
rect 63800 47850 66830 47873
rect 66990 47873 67013 48850
rect 69997 49850 70020 50857
rect 70180 50857 73210 50880
rect 70180 49850 70203 50857
rect 69997 48850 70203 49850
rect 69997 47873 70020 48850
rect 66990 47850 70020 47873
rect 70180 47873 70203 48850
rect 73187 49850 73210 50857
rect 73370 50857 76400 50880
rect 73370 49850 73393 50857
rect 73187 48850 73393 49850
rect 73187 47873 73210 48850
rect 70180 47850 73210 47873
rect 73370 47873 73393 48850
rect 76377 49850 76400 50857
rect 76560 50857 79590 50880
rect 76560 49850 76583 50857
rect 76377 48850 76583 49850
rect 76377 47873 76400 48850
rect 73370 47850 76400 47873
rect 76560 47873 76583 48850
rect 79567 49850 79590 50857
rect 79750 50857 82780 50880
rect 79750 49850 79773 50857
rect 79567 48850 79773 49850
rect 79567 47873 79590 48850
rect 76560 47850 79590 47873
rect 79750 47873 79773 48850
rect 82757 49850 82780 50857
rect 82940 50857 85970 50880
rect 82940 49850 82963 50857
rect 82757 48850 82963 49850
rect 82757 47873 82780 48850
rect 79750 47850 82780 47873
rect 82940 47873 82963 48850
rect 85947 49850 85970 50857
rect 86130 50857 89160 50880
rect 86130 49850 86153 50857
rect 85947 48850 86153 49850
rect 85947 47873 85970 48850
rect 82940 47850 85970 47873
rect 86130 47873 86153 48850
rect 89137 49850 89160 50857
rect 89320 50857 92350 50880
rect 89320 49850 89343 50857
rect 89137 48850 89343 49850
rect 89137 47873 89160 48850
rect 86130 47850 89160 47873
rect 89320 47873 89343 48850
rect 92327 49850 92350 50857
rect 92510 50857 95540 50880
rect 92510 49850 92533 50857
rect 92327 48850 92533 49850
rect 92327 47873 92350 48850
rect 89320 47850 92350 47873
rect 92510 47873 92533 48850
rect 95517 49850 95540 50857
rect 95700 50857 98730 50880
rect 95700 49850 95723 50857
rect 95517 48850 95723 49850
rect 95517 47873 95540 48850
rect 92510 47850 95540 47873
rect 95700 47873 95723 48850
rect 98707 49850 98730 50857
rect 98890 50857 101920 50880
rect 98890 49850 98913 50857
rect 98707 48850 98913 49850
rect 98707 47873 98730 48850
rect 95700 47850 98730 47873
rect 98890 47873 98913 48850
rect 101897 49850 101920 50857
rect 102080 50857 105110 50880
rect 102080 49850 102103 50857
rect 101897 48850 102103 49850
rect 101897 47873 101920 48850
rect 98890 47850 101920 47873
rect 102080 47873 102103 48850
rect 105087 49850 105110 50857
rect 105270 50857 108300 50880
rect 105270 49850 105293 50857
rect 105087 48850 105293 49850
rect 105087 47873 105110 48850
rect 102080 47850 105110 47873
rect 105270 47873 105293 48850
rect 108277 49850 108300 50857
rect 108460 50857 111490 50880
rect 108460 49850 108483 50857
rect 108277 48850 108483 49850
rect 108277 47873 108300 48850
rect 105270 47850 108300 47873
rect 108460 47873 108483 48850
rect 111467 49850 111490 50857
rect 111650 50857 114680 50880
rect 111650 49850 111673 50857
rect 111467 48850 111673 49850
rect 111467 47873 111490 48850
rect 108460 47850 111490 47873
rect 111650 47873 111673 48850
rect 114657 49850 114680 50857
rect 114840 50857 117870 50880
rect 114840 49850 114863 50857
rect 114657 48850 114863 49850
rect 114657 47873 114680 48850
rect 111650 47850 114680 47873
rect 114840 47873 114863 48850
rect 117847 49850 117870 50857
rect 118030 50857 121060 50880
rect 118030 49850 118053 50857
rect 117847 48850 118053 49850
rect 117847 47873 117870 48850
rect 114840 47850 117870 47873
rect 118030 47873 118053 48850
rect 121037 49850 121060 50857
rect 121220 50857 124250 50880
rect 121220 49850 121243 50857
rect 121037 48850 121243 49850
rect 121037 47873 121060 48850
rect 118030 47850 121060 47873
rect 121220 47873 121243 48850
rect 124227 49850 124250 50857
rect 124410 50857 127440 50880
rect 124410 49850 124433 50857
rect 124227 48850 124433 49850
rect 124227 47873 124250 48850
rect 121220 47850 124250 47873
rect 124410 47873 124433 48850
rect 127417 49850 127440 50857
rect 127600 50857 130630 50880
rect 127600 49850 127623 50857
rect 127417 48850 127623 49850
rect 127417 47873 127440 48850
rect 124410 47850 127440 47873
rect 127600 47873 127623 48850
rect 130607 49850 130630 50857
rect 130790 50857 133820 50880
rect 130790 49850 130813 50857
rect 130607 48850 130813 49850
rect 130607 47873 130630 48850
rect 127600 47850 130630 47873
rect 130790 47873 130813 48850
rect 133797 49850 133820 50857
rect 133980 50857 137010 50880
rect 133980 49850 134003 50857
rect 133797 48850 134003 49850
rect 133797 47873 133820 48850
rect 130790 47850 133820 47873
rect 133980 47873 134003 48850
rect 136987 49850 137010 50857
rect 136987 48850 137170 49850
rect 136987 47873 137010 48850
rect 133980 47850 137010 47873
rect 1000 47690 2000 47850
rect 4190 47690 5190 47850
rect 7380 47690 8380 47850
rect 10570 47690 11570 47850
rect 13760 47690 14760 47850
rect 16950 47690 17950 47850
rect 20140 47690 21140 47850
rect 23330 47690 24330 47850
rect 26520 47690 27520 47850
rect 29710 47690 30710 47850
rect 32900 47690 33900 47850
rect 36090 47690 37090 47850
rect 39280 47690 40280 47850
rect 42470 47690 43470 47850
rect 45660 47690 46660 47850
rect 48850 47690 49850 47850
rect 52040 47690 53040 47850
rect 55230 47690 56230 47850
rect 58420 47690 59420 47850
rect 61610 47690 62610 47850
rect 64800 47690 65800 47850
rect 67990 47690 68990 47850
rect 71180 47690 72180 47850
rect 74370 47690 75370 47850
rect 77560 47690 78560 47850
rect 80750 47690 81750 47850
rect 83940 47690 84940 47850
rect 87130 47690 88130 47850
rect 90320 47690 91320 47850
rect 93510 47690 94510 47850
rect 96700 47690 97700 47850
rect 99890 47690 100890 47850
rect 103080 47690 104080 47850
rect 106270 47690 107270 47850
rect 109460 47690 110460 47850
rect 112650 47690 113650 47850
rect 115840 47690 116840 47850
rect 119030 47690 120030 47850
rect 122220 47690 123220 47850
rect 125410 47690 126410 47850
rect 128600 47690 129600 47850
rect 131790 47690 132790 47850
rect 134980 47690 135980 47850
rect 0 47667 3030 47690
rect 0 44683 23 47667
rect 3007 46660 3030 47667
rect 3190 47667 6220 47690
rect 3190 46660 3213 47667
rect 3007 45660 3213 46660
rect 3007 44683 3030 45660
rect 0 44660 3030 44683
rect 3190 44683 3213 45660
rect 6197 46660 6220 47667
rect 6380 47667 9410 47690
rect 6380 46660 6403 47667
rect 6197 45660 6403 46660
rect 6197 44683 6220 45660
rect 3190 44660 6220 44683
rect 6380 44683 6403 45660
rect 9387 46660 9410 47667
rect 9570 47667 12600 47690
rect 9570 46660 9593 47667
rect 9387 45660 9593 46660
rect 9387 44683 9410 45660
rect 6380 44660 9410 44683
rect 9570 44683 9593 45660
rect 12577 46660 12600 47667
rect 12760 47667 15790 47690
rect 12760 46660 12783 47667
rect 12577 45660 12783 46660
rect 12577 44683 12600 45660
rect 9570 44660 12600 44683
rect 12760 44683 12783 45660
rect 15767 46660 15790 47667
rect 15950 47667 18980 47690
rect 15950 46660 15973 47667
rect 15767 45660 15973 46660
rect 15767 44683 15790 45660
rect 12760 44660 15790 44683
rect 15950 44683 15973 45660
rect 18957 46660 18980 47667
rect 19140 47667 22170 47690
rect 19140 46660 19163 47667
rect 18957 45660 19163 46660
rect 18957 44683 18980 45660
rect 15950 44660 18980 44683
rect 19140 44683 19163 45660
rect 22147 46660 22170 47667
rect 22330 47667 25360 47690
rect 22330 46660 22353 47667
rect 22147 45660 22353 46660
rect 22147 44683 22170 45660
rect 19140 44660 22170 44683
rect 22330 44683 22353 45660
rect 25337 46660 25360 47667
rect 25520 47667 28550 47690
rect 25520 46660 25543 47667
rect 25337 45660 25543 46660
rect 25337 44683 25360 45660
rect 22330 44660 25360 44683
rect 25520 44683 25543 45660
rect 28527 46660 28550 47667
rect 28710 47667 31740 47690
rect 28710 46660 28733 47667
rect 28527 45660 28733 46660
rect 28527 44683 28550 45660
rect 25520 44660 28550 44683
rect 28710 44683 28733 45660
rect 31717 46660 31740 47667
rect 31900 47667 34930 47690
rect 31900 46660 31923 47667
rect 31717 45660 31923 46660
rect 31717 44683 31740 45660
rect 28710 44660 31740 44683
rect 31900 44683 31923 45660
rect 34907 46660 34930 47667
rect 35090 47667 38120 47690
rect 35090 46660 35113 47667
rect 34907 45660 35113 46660
rect 34907 44683 34930 45660
rect 31900 44660 34930 44683
rect 35090 44683 35113 45660
rect 38097 46660 38120 47667
rect 38280 47667 41310 47690
rect 38280 46660 38303 47667
rect 38097 45660 38303 46660
rect 38097 44683 38120 45660
rect 35090 44660 38120 44683
rect 38280 44683 38303 45660
rect 41287 46660 41310 47667
rect 41470 47667 44500 47690
rect 41470 46660 41493 47667
rect 41287 45660 41493 46660
rect 41287 44683 41310 45660
rect 38280 44660 41310 44683
rect 41470 44683 41493 45660
rect 44477 46660 44500 47667
rect 44660 47667 47690 47690
rect 44660 46660 44683 47667
rect 44477 45660 44683 46660
rect 44477 44683 44500 45660
rect 41470 44660 44500 44683
rect 44660 44683 44683 45660
rect 47667 46660 47690 47667
rect 47850 47667 50880 47690
rect 47850 46660 47873 47667
rect 47667 45660 47873 46660
rect 47667 44683 47690 45660
rect 44660 44660 47690 44683
rect 47850 44683 47873 45660
rect 50857 46660 50880 47667
rect 51040 47667 54070 47690
rect 51040 46660 51063 47667
rect 50857 45660 51063 46660
rect 50857 44683 50880 45660
rect 47850 44660 50880 44683
rect 51040 44683 51063 45660
rect 54047 46660 54070 47667
rect 54230 47667 57260 47690
rect 54230 46660 54253 47667
rect 54047 45660 54253 46660
rect 54047 44683 54070 45660
rect 51040 44660 54070 44683
rect 54230 44683 54253 45660
rect 57237 46660 57260 47667
rect 57420 47667 60450 47690
rect 57420 46660 57443 47667
rect 57237 45660 57443 46660
rect 57237 44683 57260 45660
rect 54230 44660 57260 44683
rect 57420 44683 57443 45660
rect 60427 46660 60450 47667
rect 60610 47667 63640 47690
rect 60610 46660 60633 47667
rect 60427 45660 60633 46660
rect 60427 44683 60450 45660
rect 57420 44660 60450 44683
rect 60610 44683 60633 45660
rect 63617 46660 63640 47667
rect 63800 47667 66830 47690
rect 63800 46660 63823 47667
rect 63617 45660 63823 46660
rect 63617 44683 63640 45660
rect 60610 44660 63640 44683
rect 63800 44683 63823 45660
rect 66807 46660 66830 47667
rect 66990 47667 70020 47690
rect 66990 46660 67013 47667
rect 66807 45660 67013 46660
rect 66807 44683 66830 45660
rect 63800 44660 66830 44683
rect 66990 44683 67013 45660
rect 69997 46660 70020 47667
rect 70180 47667 73210 47690
rect 70180 46660 70203 47667
rect 69997 45660 70203 46660
rect 69997 44683 70020 45660
rect 66990 44660 70020 44683
rect 70180 44683 70203 45660
rect 73187 46660 73210 47667
rect 73370 47667 76400 47690
rect 73370 46660 73393 47667
rect 73187 45660 73393 46660
rect 73187 44683 73210 45660
rect 70180 44660 73210 44683
rect 73370 44683 73393 45660
rect 76377 46660 76400 47667
rect 76560 47667 79590 47690
rect 76560 46660 76583 47667
rect 76377 45660 76583 46660
rect 76377 44683 76400 45660
rect 73370 44660 76400 44683
rect 76560 44683 76583 45660
rect 79567 46660 79590 47667
rect 79750 47667 82780 47690
rect 79750 46660 79773 47667
rect 79567 45660 79773 46660
rect 79567 44683 79590 45660
rect 76560 44660 79590 44683
rect 79750 44683 79773 45660
rect 82757 46660 82780 47667
rect 82940 47667 85970 47690
rect 82940 46660 82963 47667
rect 82757 45660 82963 46660
rect 82757 44683 82780 45660
rect 79750 44660 82780 44683
rect 82940 44683 82963 45660
rect 85947 46660 85970 47667
rect 86130 47667 89160 47690
rect 86130 46660 86153 47667
rect 85947 45660 86153 46660
rect 85947 44683 85970 45660
rect 82940 44660 85970 44683
rect 86130 44683 86153 45660
rect 89137 46660 89160 47667
rect 89320 47667 92350 47690
rect 89320 46660 89343 47667
rect 89137 45660 89343 46660
rect 89137 44683 89160 45660
rect 86130 44660 89160 44683
rect 89320 44683 89343 45660
rect 92327 46660 92350 47667
rect 92510 47667 95540 47690
rect 92510 46660 92533 47667
rect 92327 45660 92533 46660
rect 92327 44683 92350 45660
rect 89320 44660 92350 44683
rect 92510 44683 92533 45660
rect 95517 46660 95540 47667
rect 95700 47667 98730 47690
rect 95700 46660 95723 47667
rect 95517 45660 95723 46660
rect 95517 44683 95540 45660
rect 92510 44660 95540 44683
rect 95700 44683 95723 45660
rect 98707 46660 98730 47667
rect 98890 47667 101920 47690
rect 98890 46660 98913 47667
rect 98707 45660 98913 46660
rect 98707 44683 98730 45660
rect 95700 44660 98730 44683
rect 98890 44683 98913 45660
rect 101897 46660 101920 47667
rect 102080 47667 105110 47690
rect 102080 46660 102103 47667
rect 101897 45660 102103 46660
rect 101897 44683 101920 45660
rect 98890 44660 101920 44683
rect 102080 44683 102103 45660
rect 105087 46660 105110 47667
rect 105270 47667 108300 47690
rect 105270 46660 105293 47667
rect 105087 45660 105293 46660
rect 105087 44683 105110 45660
rect 102080 44660 105110 44683
rect 105270 44683 105293 45660
rect 108277 46660 108300 47667
rect 108460 47667 111490 47690
rect 108460 46660 108483 47667
rect 108277 45660 108483 46660
rect 108277 44683 108300 45660
rect 105270 44660 108300 44683
rect 108460 44683 108483 45660
rect 111467 46660 111490 47667
rect 111650 47667 114680 47690
rect 111650 46660 111673 47667
rect 111467 45660 111673 46660
rect 111467 44683 111490 45660
rect 108460 44660 111490 44683
rect 111650 44683 111673 45660
rect 114657 46660 114680 47667
rect 114840 47667 117870 47690
rect 114840 46660 114863 47667
rect 114657 45660 114863 46660
rect 114657 44683 114680 45660
rect 111650 44660 114680 44683
rect 114840 44683 114863 45660
rect 117847 46660 117870 47667
rect 118030 47667 121060 47690
rect 118030 46660 118053 47667
rect 117847 45660 118053 46660
rect 117847 44683 117870 45660
rect 114840 44660 117870 44683
rect 118030 44683 118053 45660
rect 121037 46660 121060 47667
rect 121220 47667 124250 47690
rect 121220 46660 121243 47667
rect 121037 45660 121243 46660
rect 121037 44683 121060 45660
rect 118030 44660 121060 44683
rect 121220 44683 121243 45660
rect 124227 46660 124250 47667
rect 124410 47667 127440 47690
rect 124410 46660 124433 47667
rect 124227 45660 124433 46660
rect 124227 44683 124250 45660
rect 121220 44660 124250 44683
rect 124410 44683 124433 45660
rect 127417 46660 127440 47667
rect 127600 47667 130630 47690
rect 127600 46660 127623 47667
rect 127417 45660 127623 46660
rect 127417 44683 127440 45660
rect 124410 44660 127440 44683
rect 127600 44683 127623 45660
rect 130607 46660 130630 47667
rect 130790 47667 133820 47690
rect 130790 46660 130813 47667
rect 130607 45660 130813 46660
rect 130607 44683 130630 45660
rect 127600 44660 130630 44683
rect 130790 44683 130813 45660
rect 133797 46660 133820 47667
rect 133980 47667 137010 47690
rect 133980 46660 134003 47667
rect 133797 45660 134003 46660
rect 133797 44683 133820 45660
rect 130790 44660 133820 44683
rect 133980 44683 134003 45660
rect 136987 46660 137010 47667
rect 136987 45660 137170 46660
rect 136987 44683 137010 45660
rect 133980 44660 137010 44683
rect 1000 44500 2000 44660
rect 4190 44500 5190 44660
rect 7380 44500 8380 44660
rect 10570 44500 11570 44660
rect 13760 44500 14760 44660
rect 16950 44500 17950 44660
rect 20140 44500 21140 44660
rect 23330 44500 24330 44660
rect 26520 44500 27520 44660
rect 29710 44500 30710 44660
rect 32900 44500 33900 44660
rect 36090 44500 37090 44660
rect 39280 44500 40280 44660
rect 42470 44500 43470 44660
rect 45660 44500 46660 44660
rect 48850 44500 49850 44660
rect 52040 44500 53040 44660
rect 55230 44500 56230 44660
rect 58420 44500 59420 44660
rect 61610 44500 62610 44660
rect 64800 44500 65800 44660
rect 67990 44500 68990 44660
rect 71180 44500 72180 44660
rect 74370 44500 75370 44660
rect 77560 44500 78560 44660
rect 80750 44500 81750 44660
rect 83940 44500 84940 44660
rect 87130 44500 88130 44660
rect 90320 44500 91320 44660
rect 93510 44500 94510 44660
rect 96700 44500 97700 44660
rect 99890 44500 100890 44660
rect 103080 44500 104080 44660
rect 106270 44500 107270 44660
rect 109460 44500 110460 44660
rect 112650 44500 113650 44660
rect 115840 44500 116840 44660
rect 119030 44500 120030 44660
rect 122220 44500 123220 44660
rect 125410 44500 126410 44660
rect 128600 44500 129600 44660
rect 131790 44500 132790 44660
rect 134980 44500 135980 44660
rect 0 44477 3030 44500
rect 0 41493 23 44477
rect 3007 43470 3030 44477
rect 3190 44477 6220 44500
rect 3190 43470 3213 44477
rect 3007 42470 3213 43470
rect 3007 41493 3030 42470
rect 0 41470 3030 41493
rect 3190 41493 3213 42470
rect 6197 43470 6220 44477
rect 6380 44477 9410 44500
rect 6380 43470 6403 44477
rect 6197 42470 6403 43470
rect 6197 41493 6220 42470
rect 3190 41470 6220 41493
rect 6380 41493 6403 42470
rect 9387 43470 9410 44477
rect 9570 44477 12600 44500
rect 9570 43470 9593 44477
rect 9387 42470 9593 43470
rect 9387 41493 9410 42470
rect 6380 41470 9410 41493
rect 9570 41493 9593 42470
rect 12577 43470 12600 44477
rect 12760 44477 15790 44500
rect 12760 43470 12783 44477
rect 12577 42470 12783 43470
rect 12577 41493 12600 42470
rect 9570 41470 12600 41493
rect 12760 41493 12783 42470
rect 15767 43470 15790 44477
rect 15950 44477 18980 44500
rect 15950 43470 15973 44477
rect 15767 42470 15973 43470
rect 15767 41493 15790 42470
rect 12760 41470 15790 41493
rect 15950 41493 15973 42470
rect 18957 43470 18980 44477
rect 19140 44477 22170 44500
rect 19140 43470 19163 44477
rect 18957 42470 19163 43470
rect 18957 41493 18980 42470
rect 15950 41470 18980 41493
rect 19140 41493 19163 42470
rect 22147 43470 22170 44477
rect 22330 44477 25360 44500
rect 22330 43470 22353 44477
rect 22147 42470 22353 43470
rect 22147 41493 22170 42470
rect 19140 41470 22170 41493
rect 22330 41493 22353 42470
rect 25337 43470 25360 44477
rect 25520 44477 28550 44500
rect 25520 43470 25543 44477
rect 25337 42470 25543 43470
rect 25337 41493 25360 42470
rect 22330 41470 25360 41493
rect 25520 41493 25543 42470
rect 28527 43470 28550 44477
rect 28710 44477 31740 44500
rect 28710 43470 28733 44477
rect 28527 42470 28733 43470
rect 28527 41493 28550 42470
rect 25520 41470 28550 41493
rect 28710 41493 28733 42470
rect 31717 43470 31740 44477
rect 31900 44477 34930 44500
rect 31900 43470 31923 44477
rect 31717 42470 31923 43470
rect 31717 41493 31740 42470
rect 28710 41470 31740 41493
rect 31900 41493 31923 42470
rect 34907 43470 34930 44477
rect 35090 44477 38120 44500
rect 35090 43470 35113 44477
rect 34907 42470 35113 43470
rect 34907 41493 34930 42470
rect 31900 41470 34930 41493
rect 35090 41493 35113 42470
rect 38097 43470 38120 44477
rect 38280 44477 41310 44500
rect 38280 43470 38303 44477
rect 38097 42470 38303 43470
rect 38097 41493 38120 42470
rect 35090 41470 38120 41493
rect 38280 41493 38303 42470
rect 41287 43470 41310 44477
rect 41470 44477 44500 44500
rect 41470 43470 41493 44477
rect 41287 42470 41493 43470
rect 41287 41493 41310 42470
rect 38280 41470 41310 41493
rect 41470 41493 41493 42470
rect 44477 43470 44500 44477
rect 44660 44477 47690 44500
rect 44660 43470 44683 44477
rect 44477 42470 44683 43470
rect 44477 41493 44500 42470
rect 41470 41470 44500 41493
rect 44660 41493 44683 42470
rect 47667 43470 47690 44477
rect 47850 44477 50880 44500
rect 47850 43470 47873 44477
rect 47667 42470 47873 43470
rect 47667 41493 47690 42470
rect 44660 41470 47690 41493
rect 47850 41493 47873 42470
rect 50857 43470 50880 44477
rect 51040 44477 54070 44500
rect 51040 43470 51063 44477
rect 50857 42470 51063 43470
rect 50857 41493 50880 42470
rect 47850 41470 50880 41493
rect 51040 41493 51063 42470
rect 54047 43470 54070 44477
rect 54230 44477 57260 44500
rect 54230 43470 54253 44477
rect 54047 42470 54253 43470
rect 54047 41493 54070 42470
rect 51040 41470 54070 41493
rect 54230 41493 54253 42470
rect 57237 43470 57260 44477
rect 57420 44477 60450 44500
rect 57420 43470 57443 44477
rect 57237 42470 57443 43470
rect 57237 41493 57260 42470
rect 54230 41470 57260 41493
rect 57420 41493 57443 42470
rect 60427 43470 60450 44477
rect 60610 44477 63640 44500
rect 60610 43470 60633 44477
rect 60427 42470 60633 43470
rect 60427 41493 60450 42470
rect 57420 41470 60450 41493
rect 60610 41493 60633 42470
rect 63617 43470 63640 44477
rect 63800 44477 66830 44500
rect 63800 43470 63823 44477
rect 63617 42470 63823 43470
rect 63617 41493 63640 42470
rect 60610 41470 63640 41493
rect 63800 41493 63823 42470
rect 66807 43470 66830 44477
rect 66990 44477 70020 44500
rect 66990 43470 67013 44477
rect 66807 42470 67013 43470
rect 66807 41493 66830 42470
rect 63800 41470 66830 41493
rect 66990 41493 67013 42470
rect 69997 43470 70020 44477
rect 70180 44477 73210 44500
rect 70180 43470 70203 44477
rect 69997 42470 70203 43470
rect 69997 41493 70020 42470
rect 66990 41470 70020 41493
rect 70180 41493 70203 42470
rect 73187 43470 73210 44477
rect 73370 44477 76400 44500
rect 73370 43470 73393 44477
rect 73187 42470 73393 43470
rect 73187 41493 73210 42470
rect 70180 41470 73210 41493
rect 73370 41493 73393 42470
rect 76377 43470 76400 44477
rect 76560 44477 79590 44500
rect 76560 43470 76583 44477
rect 76377 42470 76583 43470
rect 76377 41493 76400 42470
rect 73370 41470 76400 41493
rect 76560 41493 76583 42470
rect 79567 43470 79590 44477
rect 79750 44477 82780 44500
rect 79750 43470 79773 44477
rect 79567 42470 79773 43470
rect 79567 41493 79590 42470
rect 76560 41470 79590 41493
rect 79750 41493 79773 42470
rect 82757 43470 82780 44477
rect 82940 44477 85970 44500
rect 82940 43470 82963 44477
rect 82757 42470 82963 43470
rect 82757 41493 82780 42470
rect 79750 41470 82780 41493
rect 82940 41493 82963 42470
rect 85947 43470 85970 44477
rect 86130 44477 89160 44500
rect 86130 43470 86153 44477
rect 85947 42470 86153 43470
rect 85947 41493 85970 42470
rect 82940 41470 85970 41493
rect 86130 41493 86153 42470
rect 89137 43470 89160 44477
rect 89320 44477 92350 44500
rect 89320 43470 89343 44477
rect 89137 42470 89343 43470
rect 89137 41493 89160 42470
rect 86130 41470 89160 41493
rect 89320 41493 89343 42470
rect 92327 43470 92350 44477
rect 92510 44477 95540 44500
rect 92510 43470 92533 44477
rect 92327 42470 92533 43470
rect 92327 41493 92350 42470
rect 89320 41470 92350 41493
rect 92510 41493 92533 42470
rect 95517 43470 95540 44477
rect 95700 44477 98730 44500
rect 95700 43470 95723 44477
rect 95517 42470 95723 43470
rect 95517 41493 95540 42470
rect 92510 41470 95540 41493
rect 95700 41493 95723 42470
rect 98707 43470 98730 44477
rect 98890 44477 101920 44500
rect 98890 43470 98913 44477
rect 98707 42470 98913 43470
rect 98707 41493 98730 42470
rect 95700 41470 98730 41493
rect 98890 41493 98913 42470
rect 101897 43470 101920 44477
rect 102080 44477 105110 44500
rect 102080 43470 102103 44477
rect 101897 42470 102103 43470
rect 101897 41493 101920 42470
rect 98890 41470 101920 41493
rect 102080 41493 102103 42470
rect 105087 43470 105110 44477
rect 105270 44477 108300 44500
rect 105270 43470 105293 44477
rect 105087 42470 105293 43470
rect 105087 41493 105110 42470
rect 102080 41470 105110 41493
rect 105270 41493 105293 42470
rect 108277 43470 108300 44477
rect 108460 44477 111490 44500
rect 108460 43470 108483 44477
rect 108277 42470 108483 43470
rect 108277 41493 108300 42470
rect 105270 41470 108300 41493
rect 108460 41493 108483 42470
rect 111467 43470 111490 44477
rect 111650 44477 114680 44500
rect 111650 43470 111673 44477
rect 111467 42470 111673 43470
rect 111467 41493 111490 42470
rect 108460 41470 111490 41493
rect 111650 41493 111673 42470
rect 114657 43470 114680 44477
rect 114840 44477 117870 44500
rect 114840 43470 114863 44477
rect 114657 42470 114863 43470
rect 114657 41493 114680 42470
rect 111650 41470 114680 41493
rect 114840 41493 114863 42470
rect 117847 43470 117870 44477
rect 118030 44477 121060 44500
rect 118030 43470 118053 44477
rect 117847 42470 118053 43470
rect 117847 41493 117870 42470
rect 114840 41470 117870 41493
rect 118030 41493 118053 42470
rect 121037 43470 121060 44477
rect 121220 44477 124250 44500
rect 121220 43470 121243 44477
rect 121037 42470 121243 43470
rect 121037 41493 121060 42470
rect 118030 41470 121060 41493
rect 121220 41493 121243 42470
rect 124227 43470 124250 44477
rect 124410 44477 127440 44500
rect 124410 43470 124433 44477
rect 124227 42470 124433 43470
rect 124227 41493 124250 42470
rect 121220 41470 124250 41493
rect 124410 41493 124433 42470
rect 127417 43470 127440 44477
rect 127600 44477 130630 44500
rect 127600 43470 127623 44477
rect 127417 42470 127623 43470
rect 127417 41493 127440 42470
rect 124410 41470 127440 41493
rect 127600 41493 127623 42470
rect 130607 43470 130630 44477
rect 130790 44477 133820 44500
rect 130790 43470 130813 44477
rect 130607 42470 130813 43470
rect 130607 41493 130630 42470
rect 127600 41470 130630 41493
rect 130790 41493 130813 42470
rect 133797 43470 133820 44477
rect 133980 44477 137010 44500
rect 133980 43470 134003 44477
rect 133797 42470 134003 43470
rect 133797 41493 133820 42470
rect 130790 41470 133820 41493
rect 133980 41493 134003 42470
rect 136987 43470 137010 44477
rect 136987 42470 137170 43470
rect 136987 41493 137010 42470
rect 133980 41470 137010 41493
rect 1000 41310 2000 41470
rect 4190 41310 5190 41470
rect 7380 41310 8380 41470
rect 10570 41310 11570 41470
rect 13760 41310 14760 41470
rect 16950 41310 17950 41470
rect 20140 41310 21140 41470
rect 23330 41310 24330 41470
rect 26520 41310 27520 41470
rect 29710 41310 30710 41470
rect 32900 41310 33900 41470
rect 36090 41310 37090 41470
rect 39280 41310 40280 41470
rect 42470 41310 43470 41470
rect 45660 41310 46660 41470
rect 48850 41310 49850 41470
rect 52040 41310 53040 41470
rect 55230 41310 56230 41470
rect 58420 41310 59420 41470
rect 61610 41310 62610 41470
rect 64800 41310 65800 41470
rect 67990 41310 68990 41470
rect 71180 41310 72180 41470
rect 74370 41310 75370 41470
rect 77560 41310 78560 41470
rect 80750 41310 81750 41470
rect 83940 41310 84940 41470
rect 87130 41310 88130 41470
rect 90320 41310 91320 41470
rect 93510 41310 94510 41470
rect 96700 41310 97700 41470
rect 99890 41310 100890 41470
rect 103080 41310 104080 41470
rect 106270 41310 107270 41470
rect 109460 41310 110460 41470
rect 112650 41310 113650 41470
rect 115840 41310 116840 41470
rect 119030 41310 120030 41470
rect 122220 41310 123220 41470
rect 125410 41310 126410 41470
rect 128600 41310 129600 41470
rect 131790 41310 132790 41470
rect 134980 41310 135980 41470
rect 0 41287 3030 41310
rect 0 38303 23 41287
rect 3007 40280 3030 41287
rect 3190 41287 6220 41310
rect 3190 40280 3213 41287
rect 3007 39280 3213 40280
rect 3007 38303 3030 39280
rect 0 38280 3030 38303
rect 3190 38303 3213 39280
rect 6197 40280 6220 41287
rect 6380 41287 9410 41310
rect 6380 40280 6403 41287
rect 6197 39280 6403 40280
rect 6197 38303 6220 39280
rect 3190 38280 6220 38303
rect 6380 38303 6403 39280
rect 9387 40280 9410 41287
rect 9570 41287 12600 41310
rect 9570 40280 9593 41287
rect 9387 39280 9593 40280
rect 9387 38303 9410 39280
rect 6380 38280 9410 38303
rect 9570 38303 9593 39280
rect 12577 40280 12600 41287
rect 12760 41287 15790 41310
rect 12760 40280 12783 41287
rect 12577 39280 12783 40280
rect 12577 38303 12600 39280
rect 9570 38280 12600 38303
rect 12760 38303 12783 39280
rect 15767 40280 15790 41287
rect 15950 41287 18980 41310
rect 15950 40280 15973 41287
rect 15767 39280 15973 40280
rect 15767 38303 15790 39280
rect 12760 38280 15790 38303
rect 15950 38303 15973 39280
rect 18957 40280 18980 41287
rect 19140 41287 22170 41310
rect 19140 40280 19163 41287
rect 18957 39280 19163 40280
rect 18957 38303 18980 39280
rect 15950 38280 18980 38303
rect 19140 38303 19163 39280
rect 22147 40280 22170 41287
rect 22330 41287 25360 41310
rect 22330 40280 22353 41287
rect 22147 39280 22353 40280
rect 22147 38303 22170 39280
rect 19140 38280 22170 38303
rect 22330 38303 22353 39280
rect 25337 40280 25360 41287
rect 25520 41287 28550 41310
rect 25520 40280 25543 41287
rect 25337 39280 25543 40280
rect 25337 38303 25360 39280
rect 22330 38280 25360 38303
rect 25520 38303 25543 39280
rect 28527 40280 28550 41287
rect 28710 41287 31740 41310
rect 28710 40280 28733 41287
rect 28527 39280 28733 40280
rect 28527 38303 28550 39280
rect 25520 38280 28550 38303
rect 28710 38303 28733 39280
rect 31717 40280 31740 41287
rect 31900 41287 34930 41310
rect 31900 40280 31923 41287
rect 31717 39280 31923 40280
rect 31717 38303 31740 39280
rect 28710 38280 31740 38303
rect 31900 38303 31923 39280
rect 34907 40280 34930 41287
rect 35090 41287 38120 41310
rect 35090 40280 35113 41287
rect 34907 39280 35113 40280
rect 34907 38303 34930 39280
rect 31900 38280 34930 38303
rect 35090 38303 35113 39280
rect 38097 40280 38120 41287
rect 38280 41287 41310 41310
rect 38280 40280 38303 41287
rect 38097 39280 38303 40280
rect 38097 38303 38120 39280
rect 35090 38280 38120 38303
rect 38280 38303 38303 39280
rect 41287 40280 41310 41287
rect 41470 41287 44500 41310
rect 41470 40280 41493 41287
rect 41287 39280 41493 40280
rect 41287 38303 41310 39280
rect 38280 38280 41310 38303
rect 41470 38303 41493 39280
rect 44477 40280 44500 41287
rect 44660 41287 47690 41310
rect 44660 40280 44683 41287
rect 44477 39280 44683 40280
rect 44477 38303 44500 39280
rect 41470 38280 44500 38303
rect 44660 38303 44683 39280
rect 47667 40280 47690 41287
rect 47850 41287 50880 41310
rect 47850 40280 47873 41287
rect 47667 39280 47873 40280
rect 47667 38303 47690 39280
rect 44660 38280 47690 38303
rect 47850 38303 47873 39280
rect 50857 40280 50880 41287
rect 51040 41287 54070 41310
rect 51040 40280 51063 41287
rect 50857 39280 51063 40280
rect 50857 38303 50880 39280
rect 47850 38280 50880 38303
rect 51040 38303 51063 39280
rect 54047 40280 54070 41287
rect 54230 41287 57260 41310
rect 54230 40280 54253 41287
rect 54047 39280 54253 40280
rect 54047 38303 54070 39280
rect 51040 38280 54070 38303
rect 54230 38303 54253 39280
rect 57237 40280 57260 41287
rect 57420 41287 60450 41310
rect 57420 40280 57443 41287
rect 57237 39280 57443 40280
rect 57237 38303 57260 39280
rect 54230 38280 57260 38303
rect 57420 38303 57443 39280
rect 60427 40280 60450 41287
rect 60610 41287 63640 41310
rect 60610 40280 60633 41287
rect 60427 39280 60633 40280
rect 60427 38303 60450 39280
rect 57420 38280 60450 38303
rect 60610 38303 60633 39280
rect 63617 40280 63640 41287
rect 63800 41287 66830 41310
rect 63800 40280 63823 41287
rect 63617 39280 63823 40280
rect 63617 38303 63640 39280
rect 60610 38280 63640 38303
rect 63800 38303 63823 39280
rect 66807 40280 66830 41287
rect 66990 41287 70020 41310
rect 66990 40280 67013 41287
rect 66807 39280 67013 40280
rect 66807 38303 66830 39280
rect 63800 38280 66830 38303
rect 66990 38303 67013 39280
rect 69997 40280 70020 41287
rect 70180 41287 73210 41310
rect 70180 40280 70203 41287
rect 69997 39280 70203 40280
rect 69997 38303 70020 39280
rect 66990 38280 70020 38303
rect 70180 38303 70203 39280
rect 73187 40280 73210 41287
rect 73370 41287 76400 41310
rect 73370 40280 73393 41287
rect 73187 39280 73393 40280
rect 73187 38303 73210 39280
rect 70180 38280 73210 38303
rect 73370 38303 73393 39280
rect 76377 40280 76400 41287
rect 76560 41287 79590 41310
rect 76560 40280 76583 41287
rect 76377 39280 76583 40280
rect 76377 38303 76400 39280
rect 73370 38280 76400 38303
rect 76560 38303 76583 39280
rect 79567 40280 79590 41287
rect 79750 41287 82780 41310
rect 79750 40280 79773 41287
rect 79567 39280 79773 40280
rect 79567 38303 79590 39280
rect 76560 38280 79590 38303
rect 79750 38303 79773 39280
rect 82757 40280 82780 41287
rect 82940 41287 85970 41310
rect 82940 40280 82963 41287
rect 82757 39280 82963 40280
rect 82757 38303 82780 39280
rect 79750 38280 82780 38303
rect 82940 38303 82963 39280
rect 85947 40280 85970 41287
rect 86130 41287 89160 41310
rect 86130 40280 86153 41287
rect 85947 39280 86153 40280
rect 85947 38303 85970 39280
rect 82940 38280 85970 38303
rect 86130 38303 86153 39280
rect 89137 40280 89160 41287
rect 89320 41287 92350 41310
rect 89320 40280 89343 41287
rect 89137 39280 89343 40280
rect 89137 38303 89160 39280
rect 86130 38280 89160 38303
rect 89320 38303 89343 39280
rect 92327 40280 92350 41287
rect 92510 41287 95540 41310
rect 92510 40280 92533 41287
rect 92327 39280 92533 40280
rect 92327 38303 92350 39280
rect 89320 38280 92350 38303
rect 92510 38303 92533 39280
rect 95517 40280 95540 41287
rect 95700 41287 98730 41310
rect 95700 40280 95723 41287
rect 95517 39280 95723 40280
rect 95517 38303 95540 39280
rect 92510 38280 95540 38303
rect 95700 38303 95723 39280
rect 98707 40280 98730 41287
rect 98890 41287 101920 41310
rect 98890 40280 98913 41287
rect 98707 39280 98913 40280
rect 98707 38303 98730 39280
rect 95700 38280 98730 38303
rect 98890 38303 98913 39280
rect 101897 40280 101920 41287
rect 102080 41287 105110 41310
rect 102080 40280 102103 41287
rect 101897 39280 102103 40280
rect 101897 38303 101920 39280
rect 98890 38280 101920 38303
rect 102080 38303 102103 39280
rect 105087 40280 105110 41287
rect 105270 41287 108300 41310
rect 105270 40280 105293 41287
rect 105087 39280 105293 40280
rect 105087 38303 105110 39280
rect 102080 38280 105110 38303
rect 105270 38303 105293 39280
rect 108277 40280 108300 41287
rect 108460 41287 111490 41310
rect 108460 40280 108483 41287
rect 108277 39280 108483 40280
rect 108277 38303 108300 39280
rect 105270 38280 108300 38303
rect 108460 38303 108483 39280
rect 111467 40280 111490 41287
rect 111650 41287 114680 41310
rect 111650 40280 111673 41287
rect 111467 39280 111673 40280
rect 111467 38303 111490 39280
rect 108460 38280 111490 38303
rect 111650 38303 111673 39280
rect 114657 40280 114680 41287
rect 114840 41287 117870 41310
rect 114840 40280 114863 41287
rect 114657 39280 114863 40280
rect 114657 38303 114680 39280
rect 111650 38280 114680 38303
rect 114840 38303 114863 39280
rect 117847 40280 117870 41287
rect 118030 41287 121060 41310
rect 118030 40280 118053 41287
rect 117847 39280 118053 40280
rect 117847 38303 117870 39280
rect 114840 38280 117870 38303
rect 118030 38303 118053 39280
rect 121037 40280 121060 41287
rect 121220 41287 124250 41310
rect 121220 40280 121243 41287
rect 121037 39280 121243 40280
rect 121037 38303 121060 39280
rect 118030 38280 121060 38303
rect 121220 38303 121243 39280
rect 124227 40280 124250 41287
rect 124410 41287 127440 41310
rect 124410 40280 124433 41287
rect 124227 39280 124433 40280
rect 124227 38303 124250 39280
rect 121220 38280 124250 38303
rect 124410 38303 124433 39280
rect 127417 40280 127440 41287
rect 127600 41287 130630 41310
rect 127600 40280 127623 41287
rect 127417 39280 127623 40280
rect 127417 38303 127440 39280
rect 124410 38280 127440 38303
rect 127600 38303 127623 39280
rect 130607 40280 130630 41287
rect 130790 41287 133820 41310
rect 130790 40280 130813 41287
rect 130607 39280 130813 40280
rect 130607 38303 130630 39280
rect 127600 38280 130630 38303
rect 130790 38303 130813 39280
rect 133797 40280 133820 41287
rect 133980 41287 137010 41310
rect 133980 40280 134003 41287
rect 133797 39280 134003 40280
rect 133797 38303 133820 39280
rect 130790 38280 133820 38303
rect 133980 38303 134003 39280
rect 136987 40280 137010 41287
rect 136987 39280 137170 40280
rect 136987 38303 137010 39280
rect 133980 38280 137010 38303
rect 1000 38120 2000 38280
rect 4190 38120 5190 38280
rect 7380 38120 8380 38280
rect 10570 38120 11570 38280
rect 13760 38120 14760 38280
rect 16950 38120 17950 38280
rect 20140 38120 21140 38280
rect 23330 38120 24330 38280
rect 26520 38120 27520 38280
rect 29710 38120 30710 38280
rect 32900 38120 33900 38280
rect 36090 38120 37090 38280
rect 39280 38120 40280 38280
rect 42470 38120 43470 38280
rect 45660 38120 46660 38280
rect 48850 38120 49850 38280
rect 52040 38120 53040 38280
rect 55230 38120 56230 38280
rect 58420 38120 59420 38280
rect 61610 38120 62610 38280
rect 64800 38120 65800 38280
rect 67990 38120 68990 38280
rect 71180 38120 72180 38280
rect 74370 38120 75370 38280
rect 77560 38120 78560 38280
rect 80750 38120 81750 38280
rect 83940 38120 84940 38280
rect 87130 38120 88130 38280
rect 90320 38120 91320 38280
rect 93510 38120 94510 38280
rect 96700 38120 97700 38280
rect 99890 38120 100890 38280
rect 103080 38120 104080 38280
rect 106270 38120 107270 38280
rect 109460 38120 110460 38280
rect 112650 38120 113650 38280
rect 115840 38120 116840 38280
rect 119030 38120 120030 38280
rect 122220 38120 123220 38280
rect 125410 38120 126410 38280
rect 128600 38120 129600 38280
rect 131790 38120 132790 38280
rect 134980 38120 135980 38280
rect 0 38097 3030 38120
rect 0 35113 23 38097
rect 3007 37090 3030 38097
rect 3190 38097 6220 38120
rect 3190 37090 3213 38097
rect 3007 36090 3213 37090
rect 3007 35113 3030 36090
rect 0 35090 3030 35113
rect 3190 35113 3213 36090
rect 6197 37090 6220 38097
rect 6380 38097 9410 38120
rect 6380 37090 6403 38097
rect 6197 36090 6403 37090
rect 6197 35113 6220 36090
rect 3190 35090 6220 35113
rect 6380 35113 6403 36090
rect 9387 37090 9410 38097
rect 9570 38097 12600 38120
rect 9570 37090 9593 38097
rect 9387 36090 9593 37090
rect 9387 35113 9410 36090
rect 6380 35090 9410 35113
rect 9570 35113 9593 36090
rect 12577 37090 12600 38097
rect 12760 38097 15790 38120
rect 12760 37090 12783 38097
rect 12577 36090 12783 37090
rect 12577 35113 12600 36090
rect 9570 35090 12600 35113
rect 12760 35113 12783 36090
rect 15767 37090 15790 38097
rect 15950 38097 18980 38120
rect 15950 37090 15973 38097
rect 15767 36090 15973 37090
rect 15767 35113 15790 36090
rect 12760 35090 15790 35113
rect 15950 35113 15973 36090
rect 18957 37090 18980 38097
rect 19140 38097 22170 38120
rect 19140 37090 19163 38097
rect 18957 36090 19163 37090
rect 18957 35113 18980 36090
rect 15950 35090 18980 35113
rect 19140 35113 19163 36090
rect 22147 37090 22170 38097
rect 22330 38097 25360 38120
rect 22330 37090 22353 38097
rect 22147 36090 22353 37090
rect 22147 35113 22170 36090
rect 19140 35090 22170 35113
rect 22330 35113 22353 36090
rect 25337 37090 25360 38097
rect 25520 38097 28550 38120
rect 25520 37090 25543 38097
rect 25337 36090 25543 37090
rect 25337 35113 25360 36090
rect 22330 35090 25360 35113
rect 25520 35113 25543 36090
rect 28527 37090 28550 38097
rect 28710 38097 31740 38120
rect 28710 37090 28733 38097
rect 28527 36090 28733 37090
rect 28527 35113 28550 36090
rect 25520 35090 28550 35113
rect 28710 35113 28733 36090
rect 31717 37090 31740 38097
rect 31900 38097 34930 38120
rect 31900 37090 31923 38097
rect 31717 36090 31923 37090
rect 31717 35113 31740 36090
rect 28710 35090 31740 35113
rect 31900 35113 31923 36090
rect 34907 37090 34930 38097
rect 35090 38097 38120 38120
rect 35090 37090 35113 38097
rect 34907 36090 35113 37090
rect 34907 35113 34930 36090
rect 31900 35090 34930 35113
rect 35090 35113 35113 36090
rect 38097 37090 38120 38097
rect 38280 38097 41310 38120
rect 38280 37090 38303 38097
rect 38097 36090 38303 37090
rect 38097 35113 38120 36090
rect 35090 35090 38120 35113
rect 38280 35113 38303 36090
rect 41287 37090 41310 38097
rect 41470 38097 44500 38120
rect 41470 37090 41493 38097
rect 41287 36090 41493 37090
rect 41287 35113 41310 36090
rect 38280 35090 41310 35113
rect 41470 35113 41493 36090
rect 44477 37090 44500 38097
rect 44660 38097 47690 38120
rect 44660 37090 44683 38097
rect 44477 36090 44683 37090
rect 44477 35113 44500 36090
rect 41470 35090 44500 35113
rect 44660 35113 44683 36090
rect 47667 37090 47690 38097
rect 47850 38097 50880 38120
rect 47850 37090 47873 38097
rect 47667 36090 47873 37090
rect 47667 35113 47690 36090
rect 44660 35090 47690 35113
rect 47850 35113 47873 36090
rect 50857 37090 50880 38097
rect 51040 38097 54070 38120
rect 51040 37090 51063 38097
rect 50857 36090 51063 37090
rect 50857 35113 50880 36090
rect 47850 35090 50880 35113
rect 51040 35113 51063 36090
rect 54047 37090 54070 38097
rect 54230 38097 57260 38120
rect 54230 37090 54253 38097
rect 54047 36090 54253 37090
rect 54047 35113 54070 36090
rect 51040 35090 54070 35113
rect 54230 35113 54253 36090
rect 57237 37090 57260 38097
rect 57420 38097 60450 38120
rect 57420 37090 57443 38097
rect 57237 36090 57443 37090
rect 57237 35113 57260 36090
rect 54230 35090 57260 35113
rect 57420 35113 57443 36090
rect 60427 37090 60450 38097
rect 60610 38097 63640 38120
rect 60610 37090 60633 38097
rect 60427 36090 60633 37090
rect 60427 35113 60450 36090
rect 57420 35090 60450 35113
rect 60610 35113 60633 36090
rect 63617 37090 63640 38097
rect 63800 38097 66830 38120
rect 63800 37090 63823 38097
rect 63617 36090 63823 37090
rect 63617 35113 63640 36090
rect 60610 35090 63640 35113
rect 63800 35113 63823 36090
rect 66807 37090 66830 38097
rect 66990 38097 70020 38120
rect 66990 37090 67013 38097
rect 66807 36090 67013 37090
rect 66807 35113 66830 36090
rect 63800 35090 66830 35113
rect 66990 35113 67013 36090
rect 69997 37090 70020 38097
rect 70180 38097 73210 38120
rect 70180 37090 70203 38097
rect 69997 36090 70203 37090
rect 69997 35113 70020 36090
rect 66990 35090 70020 35113
rect 70180 35113 70203 36090
rect 73187 37090 73210 38097
rect 73370 38097 76400 38120
rect 73370 37090 73393 38097
rect 73187 36090 73393 37090
rect 73187 35113 73210 36090
rect 70180 35090 73210 35113
rect 73370 35113 73393 36090
rect 76377 37090 76400 38097
rect 76560 38097 79590 38120
rect 76560 37090 76583 38097
rect 76377 36090 76583 37090
rect 76377 35113 76400 36090
rect 73370 35090 76400 35113
rect 76560 35113 76583 36090
rect 79567 37090 79590 38097
rect 79750 38097 82780 38120
rect 79750 37090 79773 38097
rect 79567 36090 79773 37090
rect 79567 35113 79590 36090
rect 76560 35090 79590 35113
rect 79750 35113 79773 36090
rect 82757 37090 82780 38097
rect 82940 38097 85970 38120
rect 82940 37090 82963 38097
rect 82757 36090 82963 37090
rect 82757 35113 82780 36090
rect 79750 35090 82780 35113
rect 82940 35113 82963 36090
rect 85947 37090 85970 38097
rect 86130 38097 89160 38120
rect 86130 37090 86153 38097
rect 85947 36090 86153 37090
rect 85947 35113 85970 36090
rect 82940 35090 85970 35113
rect 86130 35113 86153 36090
rect 89137 37090 89160 38097
rect 89320 38097 92350 38120
rect 89320 37090 89343 38097
rect 89137 36090 89343 37090
rect 89137 35113 89160 36090
rect 86130 35090 89160 35113
rect 89320 35113 89343 36090
rect 92327 37090 92350 38097
rect 92510 38097 95540 38120
rect 92510 37090 92533 38097
rect 92327 36090 92533 37090
rect 92327 35113 92350 36090
rect 89320 35090 92350 35113
rect 92510 35113 92533 36090
rect 95517 37090 95540 38097
rect 95700 38097 98730 38120
rect 95700 37090 95723 38097
rect 95517 36090 95723 37090
rect 95517 35113 95540 36090
rect 92510 35090 95540 35113
rect 95700 35113 95723 36090
rect 98707 37090 98730 38097
rect 98890 38097 101920 38120
rect 98890 37090 98913 38097
rect 98707 36090 98913 37090
rect 98707 35113 98730 36090
rect 95700 35090 98730 35113
rect 98890 35113 98913 36090
rect 101897 37090 101920 38097
rect 102080 38097 105110 38120
rect 102080 37090 102103 38097
rect 101897 36090 102103 37090
rect 101897 35113 101920 36090
rect 98890 35090 101920 35113
rect 102080 35113 102103 36090
rect 105087 37090 105110 38097
rect 105270 38097 108300 38120
rect 105270 37090 105293 38097
rect 105087 36090 105293 37090
rect 105087 35113 105110 36090
rect 102080 35090 105110 35113
rect 105270 35113 105293 36090
rect 108277 37090 108300 38097
rect 108460 38097 111490 38120
rect 108460 37090 108483 38097
rect 108277 36090 108483 37090
rect 108277 35113 108300 36090
rect 105270 35090 108300 35113
rect 108460 35113 108483 36090
rect 111467 37090 111490 38097
rect 111650 38097 114680 38120
rect 111650 37090 111673 38097
rect 111467 36090 111673 37090
rect 111467 35113 111490 36090
rect 108460 35090 111490 35113
rect 111650 35113 111673 36090
rect 114657 37090 114680 38097
rect 114840 38097 117870 38120
rect 114840 37090 114863 38097
rect 114657 36090 114863 37090
rect 114657 35113 114680 36090
rect 111650 35090 114680 35113
rect 114840 35113 114863 36090
rect 117847 37090 117870 38097
rect 118030 38097 121060 38120
rect 118030 37090 118053 38097
rect 117847 36090 118053 37090
rect 117847 35113 117870 36090
rect 114840 35090 117870 35113
rect 118030 35113 118053 36090
rect 121037 37090 121060 38097
rect 121220 38097 124250 38120
rect 121220 37090 121243 38097
rect 121037 36090 121243 37090
rect 121037 35113 121060 36090
rect 118030 35090 121060 35113
rect 121220 35113 121243 36090
rect 124227 37090 124250 38097
rect 124410 38097 127440 38120
rect 124410 37090 124433 38097
rect 124227 36090 124433 37090
rect 124227 35113 124250 36090
rect 121220 35090 124250 35113
rect 124410 35113 124433 36090
rect 127417 37090 127440 38097
rect 127600 38097 130630 38120
rect 127600 37090 127623 38097
rect 127417 36090 127623 37090
rect 127417 35113 127440 36090
rect 124410 35090 127440 35113
rect 127600 35113 127623 36090
rect 130607 37090 130630 38097
rect 130790 38097 133820 38120
rect 130790 37090 130813 38097
rect 130607 36090 130813 37090
rect 130607 35113 130630 36090
rect 127600 35090 130630 35113
rect 130790 35113 130813 36090
rect 133797 37090 133820 38097
rect 133980 38097 137010 38120
rect 133980 37090 134003 38097
rect 133797 36090 134003 37090
rect 133797 35113 133820 36090
rect 130790 35090 133820 35113
rect 133980 35113 134003 36090
rect 136987 37090 137010 38097
rect 136987 36090 137170 37090
rect 136987 35113 137010 36090
rect 133980 35090 137010 35113
rect 1000 34930 2000 35090
rect 4190 34930 5190 35090
rect 7380 34930 8380 35090
rect 10570 34930 11570 35090
rect 13760 34930 14760 35090
rect 16950 34930 17950 35090
rect 20140 34930 21140 35090
rect 23330 34930 24330 35090
rect 26520 34930 27520 35090
rect 29710 34930 30710 35090
rect 32900 34930 33900 35090
rect 36090 34930 37090 35090
rect 39280 34930 40280 35090
rect 42470 34930 43470 35090
rect 45660 34930 46660 35090
rect 48850 34930 49850 35090
rect 52040 34930 53040 35090
rect 55230 34930 56230 35090
rect 58420 34930 59420 35090
rect 61610 34930 62610 35090
rect 64800 34930 65800 35090
rect 67990 34930 68990 35090
rect 71180 34930 72180 35090
rect 74370 34930 75370 35090
rect 77560 34930 78560 35090
rect 80750 34930 81750 35090
rect 83940 34930 84940 35090
rect 87130 34930 88130 35090
rect 90320 34930 91320 35090
rect 93510 34930 94510 35090
rect 96700 34930 97700 35090
rect 99890 34930 100890 35090
rect 103080 34930 104080 35090
rect 106270 34930 107270 35090
rect 109460 34930 110460 35090
rect 112650 34930 113650 35090
rect 115840 34930 116840 35090
rect 119030 34930 120030 35090
rect 122220 34930 123220 35090
rect 125410 34930 126410 35090
rect 128600 34930 129600 35090
rect 131790 34930 132790 35090
rect 134980 34930 135980 35090
rect 0 34907 3030 34930
rect 0 31923 23 34907
rect 3007 33900 3030 34907
rect 3190 34907 6220 34930
rect 3190 33900 3213 34907
rect 3007 32900 3213 33900
rect 3007 31923 3030 32900
rect 0 31900 3030 31923
rect 3190 31923 3213 32900
rect 6197 33900 6220 34907
rect 6380 34907 9410 34930
rect 6380 33900 6403 34907
rect 6197 32900 6403 33900
rect 6197 31923 6220 32900
rect 3190 31900 6220 31923
rect 6380 31923 6403 32900
rect 9387 33900 9410 34907
rect 9570 34907 12600 34930
rect 9570 33900 9593 34907
rect 9387 32900 9593 33900
rect 9387 31923 9410 32900
rect 6380 31900 9410 31923
rect 9570 31923 9593 32900
rect 12577 33900 12600 34907
rect 12760 34907 15790 34930
rect 12760 33900 12783 34907
rect 12577 32900 12783 33900
rect 12577 31923 12600 32900
rect 9570 31900 12600 31923
rect 12760 31923 12783 32900
rect 15767 33900 15790 34907
rect 15950 34907 18980 34930
rect 15950 33900 15973 34907
rect 15767 32900 15973 33900
rect 15767 31923 15790 32900
rect 12760 31900 15790 31923
rect 15950 31923 15973 32900
rect 18957 33900 18980 34907
rect 19140 34907 22170 34930
rect 19140 33900 19163 34907
rect 18957 32900 19163 33900
rect 18957 31923 18980 32900
rect 15950 31900 18980 31923
rect 19140 31923 19163 32900
rect 22147 33900 22170 34907
rect 22330 34907 25360 34930
rect 22330 33900 22353 34907
rect 22147 32900 22353 33900
rect 22147 31923 22170 32900
rect 19140 31900 22170 31923
rect 22330 31923 22353 32900
rect 25337 33900 25360 34907
rect 25520 34907 28550 34930
rect 25520 33900 25543 34907
rect 25337 32900 25543 33900
rect 25337 31923 25360 32900
rect 22330 31900 25360 31923
rect 25520 31923 25543 32900
rect 28527 33900 28550 34907
rect 28710 34907 31740 34930
rect 28710 33900 28733 34907
rect 28527 32900 28733 33900
rect 28527 31923 28550 32900
rect 25520 31900 28550 31923
rect 28710 31923 28733 32900
rect 31717 33900 31740 34907
rect 31900 34907 34930 34930
rect 31900 33900 31923 34907
rect 31717 32900 31923 33900
rect 31717 31923 31740 32900
rect 28710 31900 31740 31923
rect 31900 31923 31923 32900
rect 34907 33900 34930 34907
rect 35090 34907 38120 34930
rect 35090 33900 35113 34907
rect 34907 32900 35113 33900
rect 34907 31923 34930 32900
rect 31900 31900 34930 31923
rect 35090 31923 35113 32900
rect 38097 33900 38120 34907
rect 38280 34907 41310 34930
rect 38280 33900 38303 34907
rect 38097 32900 38303 33900
rect 38097 31923 38120 32900
rect 35090 31900 38120 31923
rect 38280 31923 38303 32900
rect 41287 33900 41310 34907
rect 41470 34907 44500 34930
rect 41470 33900 41493 34907
rect 41287 32900 41493 33900
rect 41287 31923 41310 32900
rect 38280 31900 41310 31923
rect 41470 31923 41493 32900
rect 44477 33900 44500 34907
rect 44660 34907 47690 34930
rect 44660 33900 44683 34907
rect 44477 32900 44683 33900
rect 44477 31923 44500 32900
rect 41470 31900 44500 31923
rect 44660 31923 44683 32900
rect 47667 33900 47690 34907
rect 47850 34907 50880 34930
rect 47850 33900 47873 34907
rect 47667 32900 47873 33900
rect 47667 31923 47690 32900
rect 44660 31900 47690 31923
rect 47850 31923 47873 32900
rect 50857 33900 50880 34907
rect 51040 34907 54070 34930
rect 51040 33900 51063 34907
rect 50857 32900 51063 33900
rect 50857 31923 50880 32900
rect 47850 31900 50880 31923
rect 51040 31923 51063 32900
rect 54047 33900 54070 34907
rect 54230 34907 57260 34930
rect 54230 33900 54253 34907
rect 54047 32900 54253 33900
rect 54047 31923 54070 32900
rect 51040 31900 54070 31923
rect 54230 31923 54253 32900
rect 57237 33900 57260 34907
rect 57420 34907 60450 34930
rect 57420 33900 57443 34907
rect 57237 32900 57443 33900
rect 57237 31923 57260 32900
rect 54230 31900 57260 31923
rect 57420 31923 57443 32900
rect 60427 33900 60450 34907
rect 60610 34907 63640 34930
rect 60610 33900 60633 34907
rect 60427 32900 60633 33900
rect 60427 31923 60450 32900
rect 57420 31900 60450 31923
rect 60610 31923 60633 32900
rect 63617 33900 63640 34907
rect 63800 34907 66830 34930
rect 63800 33900 63823 34907
rect 63617 32900 63823 33900
rect 63617 31923 63640 32900
rect 60610 31900 63640 31923
rect 63800 31923 63823 32900
rect 66807 33900 66830 34907
rect 66990 34907 70020 34930
rect 66990 33900 67013 34907
rect 66807 32900 67013 33900
rect 66807 31923 66830 32900
rect 63800 31900 66830 31923
rect 66990 31923 67013 32900
rect 69997 33900 70020 34907
rect 70180 34907 73210 34930
rect 70180 33900 70203 34907
rect 69997 32900 70203 33900
rect 69997 31923 70020 32900
rect 66990 31900 70020 31923
rect 70180 31923 70203 32900
rect 73187 33900 73210 34907
rect 73370 34907 76400 34930
rect 73370 33900 73393 34907
rect 73187 32900 73393 33900
rect 73187 31923 73210 32900
rect 70180 31900 73210 31923
rect 73370 31923 73393 32900
rect 76377 33900 76400 34907
rect 76560 34907 79590 34930
rect 76560 33900 76583 34907
rect 76377 32900 76583 33900
rect 76377 31923 76400 32900
rect 73370 31900 76400 31923
rect 76560 31923 76583 32900
rect 79567 33900 79590 34907
rect 79750 34907 82780 34930
rect 79750 33900 79773 34907
rect 79567 32900 79773 33900
rect 79567 31923 79590 32900
rect 76560 31900 79590 31923
rect 79750 31923 79773 32900
rect 82757 33900 82780 34907
rect 82940 34907 85970 34930
rect 82940 33900 82963 34907
rect 82757 32900 82963 33900
rect 82757 31923 82780 32900
rect 79750 31900 82780 31923
rect 82940 31923 82963 32900
rect 85947 33900 85970 34907
rect 86130 34907 89160 34930
rect 86130 33900 86153 34907
rect 85947 32900 86153 33900
rect 85947 31923 85970 32900
rect 82940 31900 85970 31923
rect 86130 31923 86153 32900
rect 89137 33900 89160 34907
rect 89320 34907 92350 34930
rect 89320 33900 89343 34907
rect 89137 32900 89343 33900
rect 89137 31923 89160 32900
rect 86130 31900 89160 31923
rect 89320 31923 89343 32900
rect 92327 33900 92350 34907
rect 92510 34907 95540 34930
rect 92510 33900 92533 34907
rect 92327 32900 92533 33900
rect 92327 31923 92350 32900
rect 89320 31900 92350 31923
rect 92510 31923 92533 32900
rect 95517 33900 95540 34907
rect 95700 34907 98730 34930
rect 95700 33900 95723 34907
rect 95517 32900 95723 33900
rect 95517 31923 95540 32900
rect 92510 31900 95540 31923
rect 95700 31923 95723 32900
rect 98707 33900 98730 34907
rect 98890 34907 101920 34930
rect 98890 33900 98913 34907
rect 98707 32900 98913 33900
rect 98707 31923 98730 32900
rect 95700 31900 98730 31923
rect 98890 31923 98913 32900
rect 101897 33900 101920 34907
rect 102080 34907 105110 34930
rect 102080 33900 102103 34907
rect 101897 32900 102103 33900
rect 101897 31923 101920 32900
rect 98890 31900 101920 31923
rect 102080 31923 102103 32900
rect 105087 33900 105110 34907
rect 105270 34907 108300 34930
rect 105270 33900 105293 34907
rect 105087 32900 105293 33900
rect 105087 31923 105110 32900
rect 102080 31900 105110 31923
rect 105270 31923 105293 32900
rect 108277 33900 108300 34907
rect 108460 34907 111490 34930
rect 108460 33900 108483 34907
rect 108277 32900 108483 33900
rect 108277 31923 108300 32900
rect 105270 31900 108300 31923
rect 108460 31923 108483 32900
rect 111467 33900 111490 34907
rect 111650 34907 114680 34930
rect 111650 33900 111673 34907
rect 111467 32900 111673 33900
rect 111467 31923 111490 32900
rect 108460 31900 111490 31923
rect 111650 31923 111673 32900
rect 114657 33900 114680 34907
rect 114840 34907 117870 34930
rect 114840 33900 114863 34907
rect 114657 32900 114863 33900
rect 114657 31923 114680 32900
rect 111650 31900 114680 31923
rect 114840 31923 114863 32900
rect 117847 33900 117870 34907
rect 118030 34907 121060 34930
rect 118030 33900 118053 34907
rect 117847 32900 118053 33900
rect 117847 31923 117870 32900
rect 114840 31900 117870 31923
rect 118030 31923 118053 32900
rect 121037 33900 121060 34907
rect 121220 34907 124250 34930
rect 121220 33900 121243 34907
rect 121037 32900 121243 33900
rect 121037 31923 121060 32900
rect 118030 31900 121060 31923
rect 121220 31923 121243 32900
rect 124227 33900 124250 34907
rect 124410 34907 127440 34930
rect 124410 33900 124433 34907
rect 124227 32900 124433 33900
rect 124227 31923 124250 32900
rect 121220 31900 124250 31923
rect 124410 31923 124433 32900
rect 127417 33900 127440 34907
rect 127600 34907 130630 34930
rect 127600 33900 127623 34907
rect 127417 32900 127623 33900
rect 127417 31923 127440 32900
rect 124410 31900 127440 31923
rect 127600 31923 127623 32900
rect 130607 33900 130630 34907
rect 130790 34907 133820 34930
rect 130790 33900 130813 34907
rect 130607 32900 130813 33900
rect 130607 31923 130630 32900
rect 127600 31900 130630 31923
rect 130790 31923 130813 32900
rect 133797 33900 133820 34907
rect 133980 34907 137010 34930
rect 133980 33900 134003 34907
rect 133797 32900 134003 33900
rect 133797 31923 133820 32900
rect 130790 31900 133820 31923
rect 133980 31923 134003 32900
rect 136987 33900 137010 34907
rect 136987 32900 137170 33900
rect 136987 31923 137010 32900
rect 133980 31900 137010 31923
rect 1000 31740 2000 31900
rect 4190 31740 5190 31900
rect 7380 31740 8380 31900
rect 10570 31740 11570 31900
rect 13760 31740 14760 31900
rect 16950 31740 17950 31900
rect 20140 31740 21140 31900
rect 23330 31740 24330 31900
rect 26520 31740 27520 31900
rect 29710 31740 30710 31900
rect 32900 31740 33900 31900
rect 36090 31740 37090 31900
rect 39280 31740 40280 31900
rect 42470 31740 43470 31900
rect 45660 31740 46660 31900
rect 48850 31740 49850 31900
rect 52040 31740 53040 31900
rect 55230 31740 56230 31900
rect 58420 31740 59420 31900
rect 61610 31740 62610 31900
rect 64800 31740 65800 31900
rect 67990 31740 68990 31900
rect 71180 31740 72180 31900
rect 74370 31740 75370 31900
rect 77560 31740 78560 31900
rect 80750 31740 81750 31900
rect 83940 31740 84940 31900
rect 87130 31740 88130 31900
rect 90320 31740 91320 31900
rect 93510 31740 94510 31900
rect 96700 31740 97700 31900
rect 99890 31740 100890 31900
rect 103080 31740 104080 31900
rect 106270 31740 107270 31900
rect 109460 31740 110460 31900
rect 112650 31740 113650 31900
rect 115840 31740 116840 31900
rect 119030 31740 120030 31900
rect 122220 31740 123220 31900
rect 125410 31740 126410 31900
rect 128600 31740 129600 31900
rect 131790 31740 132790 31900
rect 134980 31740 135980 31900
rect 0 31717 3030 31740
rect 0 28733 23 31717
rect 3007 30710 3030 31717
rect 3190 31717 6220 31740
rect 3190 30710 3213 31717
rect 3007 29710 3213 30710
rect 3007 28733 3030 29710
rect 0 28710 3030 28733
rect 3190 28733 3213 29710
rect 6197 30710 6220 31717
rect 6380 31717 9410 31740
rect 6380 30710 6403 31717
rect 6197 29710 6403 30710
rect 6197 28733 6220 29710
rect 3190 28710 6220 28733
rect 6380 28733 6403 29710
rect 9387 30710 9410 31717
rect 9570 31717 12600 31740
rect 9570 30710 9593 31717
rect 9387 29710 9593 30710
rect 9387 28733 9410 29710
rect 6380 28710 9410 28733
rect 9570 28733 9593 29710
rect 12577 30710 12600 31717
rect 12760 31717 15790 31740
rect 12760 30710 12783 31717
rect 12577 29710 12783 30710
rect 12577 28733 12600 29710
rect 9570 28710 12600 28733
rect 12760 28733 12783 29710
rect 15767 30710 15790 31717
rect 15950 31717 18980 31740
rect 15950 30710 15973 31717
rect 15767 29710 15973 30710
rect 15767 28733 15790 29710
rect 12760 28710 15790 28733
rect 15950 28733 15973 29710
rect 18957 30710 18980 31717
rect 19140 31717 22170 31740
rect 19140 30710 19163 31717
rect 18957 29710 19163 30710
rect 18957 28733 18980 29710
rect 15950 28710 18980 28733
rect 19140 28733 19163 29710
rect 22147 30710 22170 31717
rect 22330 31717 25360 31740
rect 22330 30710 22353 31717
rect 22147 29710 22353 30710
rect 22147 28733 22170 29710
rect 19140 28710 22170 28733
rect 22330 28733 22353 29710
rect 25337 30710 25360 31717
rect 25520 31717 28550 31740
rect 25520 30710 25543 31717
rect 25337 29710 25543 30710
rect 25337 28733 25360 29710
rect 22330 28710 25360 28733
rect 25520 28733 25543 29710
rect 28527 30710 28550 31717
rect 28710 31717 31740 31740
rect 28710 30710 28733 31717
rect 28527 29710 28733 30710
rect 28527 28733 28550 29710
rect 25520 28710 28550 28733
rect 28710 28733 28733 29710
rect 31717 30710 31740 31717
rect 31900 31717 34930 31740
rect 31900 30710 31923 31717
rect 31717 29710 31923 30710
rect 31717 28733 31740 29710
rect 28710 28710 31740 28733
rect 31900 28733 31923 29710
rect 34907 30710 34930 31717
rect 35090 31717 38120 31740
rect 35090 30710 35113 31717
rect 34907 29710 35113 30710
rect 34907 28733 34930 29710
rect 31900 28710 34930 28733
rect 35090 28733 35113 29710
rect 38097 30710 38120 31717
rect 38280 31717 41310 31740
rect 38280 30710 38303 31717
rect 38097 29710 38303 30710
rect 38097 28733 38120 29710
rect 35090 28710 38120 28733
rect 38280 28733 38303 29710
rect 41287 30710 41310 31717
rect 41470 31717 44500 31740
rect 41470 30710 41493 31717
rect 41287 29710 41493 30710
rect 41287 28733 41310 29710
rect 38280 28710 41310 28733
rect 41470 28733 41493 29710
rect 44477 30710 44500 31717
rect 44660 31717 47690 31740
rect 44660 30710 44683 31717
rect 44477 29710 44683 30710
rect 44477 28733 44500 29710
rect 41470 28710 44500 28733
rect 44660 28733 44683 29710
rect 47667 30710 47690 31717
rect 47850 31717 50880 31740
rect 47850 30710 47873 31717
rect 47667 29710 47873 30710
rect 47667 28733 47690 29710
rect 44660 28710 47690 28733
rect 47850 28733 47873 29710
rect 50857 30710 50880 31717
rect 51040 31717 54070 31740
rect 51040 30710 51063 31717
rect 50857 29710 51063 30710
rect 50857 28733 50880 29710
rect 47850 28710 50880 28733
rect 51040 28733 51063 29710
rect 54047 30710 54070 31717
rect 54230 31717 57260 31740
rect 54230 30710 54253 31717
rect 54047 29710 54253 30710
rect 54047 28733 54070 29710
rect 51040 28710 54070 28733
rect 54230 28733 54253 29710
rect 57237 30710 57260 31717
rect 57420 31717 60450 31740
rect 57420 30710 57443 31717
rect 57237 29710 57443 30710
rect 57237 28733 57260 29710
rect 54230 28710 57260 28733
rect 57420 28733 57443 29710
rect 60427 30710 60450 31717
rect 60610 31717 63640 31740
rect 60610 30710 60633 31717
rect 60427 29710 60633 30710
rect 60427 28733 60450 29710
rect 57420 28710 60450 28733
rect 60610 28733 60633 29710
rect 63617 30710 63640 31717
rect 63800 31717 66830 31740
rect 63800 30710 63823 31717
rect 63617 29710 63823 30710
rect 63617 28733 63640 29710
rect 60610 28710 63640 28733
rect 63800 28733 63823 29710
rect 66807 30710 66830 31717
rect 66990 31717 70020 31740
rect 66990 30710 67013 31717
rect 66807 29710 67013 30710
rect 66807 28733 66830 29710
rect 63800 28710 66830 28733
rect 66990 28733 67013 29710
rect 69997 30710 70020 31717
rect 70180 31717 73210 31740
rect 70180 30710 70203 31717
rect 69997 29710 70203 30710
rect 69997 28733 70020 29710
rect 66990 28710 70020 28733
rect 70180 28733 70203 29710
rect 73187 30710 73210 31717
rect 73370 31717 76400 31740
rect 73370 30710 73393 31717
rect 73187 29710 73393 30710
rect 73187 28733 73210 29710
rect 70180 28710 73210 28733
rect 73370 28733 73393 29710
rect 76377 30710 76400 31717
rect 76560 31717 79590 31740
rect 76560 30710 76583 31717
rect 76377 29710 76583 30710
rect 76377 28733 76400 29710
rect 73370 28710 76400 28733
rect 76560 28733 76583 29710
rect 79567 30710 79590 31717
rect 79750 31717 82780 31740
rect 79750 30710 79773 31717
rect 79567 29710 79773 30710
rect 79567 28733 79590 29710
rect 76560 28710 79590 28733
rect 79750 28733 79773 29710
rect 82757 30710 82780 31717
rect 82940 31717 85970 31740
rect 82940 30710 82963 31717
rect 82757 29710 82963 30710
rect 82757 28733 82780 29710
rect 79750 28710 82780 28733
rect 82940 28733 82963 29710
rect 85947 30710 85970 31717
rect 86130 31717 89160 31740
rect 86130 30710 86153 31717
rect 85947 29710 86153 30710
rect 85947 28733 85970 29710
rect 82940 28710 85970 28733
rect 86130 28733 86153 29710
rect 89137 30710 89160 31717
rect 89320 31717 92350 31740
rect 89320 30710 89343 31717
rect 89137 29710 89343 30710
rect 89137 28733 89160 29710
rect 86130 28710 89160 28733
rect 89320 28733 89343 29710
rect 92327 30710 92350 31717
rect 92510 31717 95540 31740
rect 92510 30710 92533 31717
rect 92327 29710 92533 30710
rect 92327 28733 92350 29710
rect 89320 28710 92350 28733
rect 92510 28733 92533 29710
rect 95517 30710 95540 31717
rect 95700 31717 98730 31740
rect 95700 30710 95723 31717
rect 95517 29710 95723 30710
rect 95517 28733 95540 29710
rect 92510 28710 95540 28733
rect 95700 28733 95723 29710
rect 98707 30710 98730 31717
rect 98890 31717 101920 31740
rect 98890 30710 98913 31717
rect 98707 29710 98913 30710
rect 98707 28733 98730 29710
rect 95700 28710 98730 28733
rect 98890 28733 98913 29710
rect 101897 30710 101920 31717
rect 102080 31717 105110 31740
rect 102080 30710 102103 31717
rect 101897 29710 102103 30710
rect 101897 28733 101920 29710
rect 98890 28710 101920 28733
rect 102080 28733 102103 29710
rect 105087 30710 105110 31717
rect 105270 31717 108300 31740
rect 105270 30710 105293 31717
rect 105087 29710 105293 30710
rect 105087 28733 105110 29710
rect 102080 28710 105110 28733
rect 105270 28733 105293 29710
rect 108277 30710 108300 31717
rect 108460 31717 111490 31740
rect 108460 30710 108483 31717
rect 108277 29710 108483 30710
rect 108277 28733 108300 29710
rect 105270 28710 108300 28733
rect 108460 28733 108483 29710
rect 111467 30710 111490 31717
rect 111650 31717 114680 31740
rect 111650 30710 111673 31717
rect 111467 29710 111673 30710
rect 111467 28733 111490 29710
rect 108460 28710 111490 28733
rect 111650 28733 111673 29710
rect 114657 30710 114680 31717
rect 114840 31717 117870 31740
rect 114840 30710 114863 31717
rect 114657 29710 114863 30710
rect 114657 28733 114680 29710
rect 111650 28710 114680 28733
rect 114840 28733 114863 29710
rect 117847 30710 117870 31717
rect 118030 31717 121060 31740
rect 118030 30710 118053 31717
rect 117847 29710 118053 30710
rect 117847 28733 117870 29710
rect 114840 28710 117870 28733
rect 118030 28733 118053 29710
rect 121037 30710 121060 31717
rect 121220 31717 124250 31740
rect 121220 30710 121243 31717
rect 121037 29710 121243 30710
rect 121037 28733 121060 29710
rect 118030 28710 121060 28733
rect 121220 28733 121243 29710
rect 124227 30710 124250 31717
rect 124410 31717 127440 31740
rect 124410 30710 124433 31717
rect 124227 29710 124433 30710
rect 124227 28733 124250 29710
rect 121220 28710 124250 28733
rect 124410 28733 124433 29710
rect 127417 30710 127440 31717
rect 127600 31717 130630 31740
rect 127600 30710 127623 31717
rect 127417 29710 127623 30710
rect 127417 28733 127440 29710
rect 124410 28710 127440 28733
rect 127600 28733 127623 29710
rect 130607 30710 130630 31717
rect 130790 31717 133820 31740
rect 130790 30710 130813 31717
rect 130607 29710 130813 30710
rect 130607 28733 130630 29710
rect 127600 28710 130630 28733
rect 130790 28733 130813 29710
rect 133797 30710 133820 31717
rect 133980 31717 137010 31740
rect 133980 30710 134003 31717
rect 133797 29710 134003 30710
rect 133797 28733 133820 29710
rect 130790 28710 133820 28733
rect 133980 28733 134003 29710
rect 136987 30710 137010 31717
rect 136987 29710 137170 30710
rect 136987 28733 137010 29710
rect 133980 28710 137010 28733
rect 1000 28550 2000 28710
rect 4190 28550 5190 28710
rect 7380 28550 8380 28710
rect 10570 28550 11570 28710
rect 13760 28550 14760 28710
rect 16950 28550 17950 28710
rect 20140 28550 21140 28710
rect 23330 28550 24330 28710
rect 26520 28550 27520 28710
rect 29710 28550 30710 28710
rect 32900 28550 33900 28710
rect 36090 28550 37090 28710
rect 39280 28550 40280 28710
rect 42470 28550 43470 28710
rect 45660 28550 46660 28710
rect 48850 28550 49850 28710
rect 52040 28550 53040 28710
rect 55230 28550 56230 28710
rect 58420 28550 59420 28710
rect 61610 28550 62610 28710
rect 64800 28550 65800 28710
rect 67990 28550 68990 28710
rect 71180 28550 72180 28710
rect 74370 28550 75370 28710
rect 77560 28550 78560 28710
rect 80750 28550 81750 28710
rect 83940 28550 84940 28710
rect 87130 28550 88130 28710
rect 90320 28550 91320 28710
rect 93510 28550 94510 28710
rect 96700 28550 97700 28710
rect 99890 28550 100890 28710
rect 103080 28550 104080 28710
rect 106270 28550 107270 28710
rect 109460 28550 110460 28710
rect 112650 28550 113650 28710
rect 115840 28550 116840 28710
rect 119030 28550 120030 28710
rect 122220 28550 123220 28710
rect 125410 28550 126410 28710
rect 128600 28550 129600 28710
rect 131790 28550 132790 28710
rect 134980 28550 135980 28710
rect 0 28527 3030 28550
rect 0 25543 23 28527
rect 3007 27520 3030 28527
rect 3190 28527 6220 28550
rect 3190 27520 3213 28527
rect 3007 26520 3213 27520
rect 3007 25543 3030 26520
rect 0 25520 3030 25543
rect 3190 25543 3213 26520
rect 6197 27520 6220 28527
rect 6380 28527 9410 28550
rect 6380 27520 6403 28527
rect 6197 26520 6403 27520
rect 6197 25543 6220 26520
rect 3190 25520 6220 25543
rect 6380 25543 6403 26520
rect 9387 27520 9410 28527
rect 9570 28527 12600 28550
rect 9570 27520 9593 28527
rect 9387 26520 9593 27520
rect 9387 25543 9410 26520
rect 6380 25520 9410 25543
rect 9570 25543 9593 26520
rect 12577 27520 12600 28527
rect 12760 28527 15790 28550
rect 12760 27520 12783 28527
rect 12577 26520 12783 27520
rect 12577 25543 12600 26520
rect 9570 25520 12600 25543
rect 12760 25543 12783 26520
rect 15767 27520 15790 28527
rect 15950 28527 18980 28550
rect 15950 27520 15973 28527
rect 15767 26520 15973 27520
rect 15767 25543 15790 26520
rect 12760 25520 15790 25543
rect 15950 25543 15973 26520
rect 18957 27520 18980 28527
rect 19140 28527 22170 28550
rect 19140 27520 19163 28527
rect 18957 26520 19163 27520
rect 18957 25543 18980 26520
rect 15950 25520 18980 25543
rect 19140 25543 19163 26520
rect 22147 27520 22170 28527
rect 22330 28527 25360 28550
rect 22330 27520 22353 28527
rect 22147 26520 22353 27520
rect 22147 25543 22170 26520
rect 19140 25520 22170 25543
rect 22330 25543 22353 26520
rect 25337 27520 25360 28527
rect 25520 28527 28550 28550
rect 25520 27520 25543 28527
rect 25337 26520 25543 27520
rect 25337 25543 25360 26520
rect 22330 25520 25360 25543
rect 25520 25543 25543 26520
rect 28527 27520 28550 28527
rect 28710 28527 31740 28550
rect 28710 27520 28733 28527
rect 28527 26520 28733 27520
rect 28527 25543 28550 26520
rect 25520 25520 28550 25543
rect 28710 25543 28733 26520
rect 31717 27520 31740 28527
rect 31900 28527 34930 28550
rect 31900 27520 31923 28527
rect 31717 26520 31923 27520
rect 31717 25543 31740 26520
rect 28710 25520 31740 25543
rect 31900 25543 31923 26520
rect 34907 27520 34930 28527
rect 35090 28527 38120 28550
rect 35090 27520 35113 28527
rect 34907 26520 35113 27520
rect 34907 25543 34930 26520
rect 31900 25520 34930 25543
rect 35090 25543 35113 26520
rect 38097 27520 38120 28527
rect 38280 28527 41310 28550
rect 38280 27520 38303 28527
rect 38097 26520 38303 27520
rect 38097 25543 38120 26520
rect 35090 25520 38120 25543
rect 38280 25543 38303 26520
rect 41287 27520 41310 28527
rect 41470 28527 44500 28550
rect 41470 27520 41493 28527
rect 41287 26520 41493 27520
rect 41287 25543 41310 26520
rect 38280 25520 41310 25543
rect 41470 25543 41493 26520
rect 44477 27520 44500 28527
rect 44660 28527 47690 28550
rect 44660 27520 44683 28527
rect 44477 26520 44683 27520
rect 44477 25543 44500 26520
rect 41470 25520 44500 25543
rect 44660 25543 44683 26520
rect 47667 27520 47690 28527
rect 47850 28527 50880 28550
rect 47850 27520 47873 28527
rect 47667 26520 47873 27520
rect 47667 25543 47690 26520
rect 44660 25520 47690 25543
rect 47850 25543 47873 26520
rect 50857 27520 50880 28527
rect 51040 28527 54070 28550
rect 51040 27520 51063 28527
rect 50857 26520 51063 27520
rect 50857 25543 50880 26520
rect 47850 25520 50880 25543
rect 51040 25543 51063 26520
rect 54047 27520 54070 28527
rect 54230 28527 57260 28550
rect 54230 27520 54253 28527
rect 54047 26520 54253 27520
rect 54047 25543 54070 26520
rect 51040 25520 54070 25543
rect 54230 25543 54253 26520
rect 57237 27520 57260 28527
rect 57420 28527 60450 28550
rect 57420 27520 57443 28527
rect 57237 26520 57443 27520
rect 57237 25543 57260 26520
rect 54230 25520 57260 25543
rect 57420 25543 57443 26520
rect 60427 27520 60450 28527
rect 60610 28527 63640 28550
rect 60610 27520 60633 28527
rect 60427 26520 60633 27520
rect 60427 25543 60450 26520
rect 57420 25520 60450 25543
rect 60610 25543 60633 26520
rect 63617 27520 63640 28527
rect 63800 28527 66830 28550
rect 63800 27520 63823 28527
rect 63617 26520 63823 27520
rect 63617 25543 63640 26520
rect 60610 25520 63640 25543
rect 63800 25543 63823 26520
rect 66807 27520 66830 28527
rect 66990 28527 70020 28550
rect 66990 27520 67013 28527
rect 66807 26520 67013 27520
rect 66807 25543 66830 26520
rect 63800 25520 66830 25543
rect 66990 25543 67013 26520
rect 69997 27520 70020 28527
rect 70180 28527 73210 28550
rect 70180 27520 70203 28527
rect 69997 26520 70203 27520
rect 69997 25543 70020 26520
rect 66990 25520 70020 25543
rect 70180 25543 70203 26520
rect 73187 27520 73210 28527
rect 73370 28527 76400 28550
rect 73370 27520 73393 28527
rect 73187 26520 73393 27520
rect 73187 25543 73210 26520
rect 70180 25520 73210 25543
rect 73370 25543 73393 26520
rect 76377 27520 76400 28527
rect 76560 28527 79590 28550
rect 76560 27520 76583 28527
rect 76377 26520 76583 27520
rect 76377 25543 76400 26520
rect 73370 25520 76400 25543
rect 76560 25543 76583 26520
rect 79567 27520 79590 28527
rect 79750 28527 82780 28550
rect 79750 27520 79773 28527
rect 79567 26520 79773 27520
rect 79567 25543 79590 26520
rect 76560 25520 79590 25543
rect 79750 25543 79773 26520
rect 82757 27520 82780 28527
rect 82940 28527 85970 28550
rect 82940 27520 82963 28527
rect 82757 26520 82963 27520
rect 82757 25543 82780 26520
rect 79750 25520 82780 25543
rect 82940 25543 82963 26520
rect 85947 27520 85970 28527
rect 86130 28527 89160 28550
rect 86130 27520 86153 28527
rect 85947 26520 86153 27520
rect 85947 25543 85970 26520
rect 82940 25520 85970 25543
rect 86130 25543 86153 26520
rect 89137 27520 89160 28527
rect 89320 28527 92350 28550
rect 89320 27520 89343 28527
rect 89137 26520 89343 27520
rect 89137 25543 89160 26520
rect 86130 25520 89160 25543
rect 89320 25543 89343 26520
rect 92327 27520 92350 28527
rect 92510 28527 95540 28550
rect 92510 27520 92533 28527
rect 92327 26520 92533 27520
rect 92327 25543 92350 26520
rect 89320 25520 92350 25543
rect 92510 25543 92533 26520
rect 95517 27520 95540 28527
rect 95700 28527 98730 28550
rect 95700 27520 95723 28527
rect 95517 26520 95723 27520
rect 95517 25543 95540 26520
rect 92510 25520 95540 25543
rect 95700 25543 95723 26520
rect 98707 27520 98730 28527
rect 98890 28527 101920 28550
rect 98890 27520 98913 28527
rect 98707 26520 98913 27520
rect 98707 25543 98730 26520
rect 95700 25520 98730 25543
rect 98890 25543 98913 26520
rect 101897 27520 101920 28527
rect 102080 28527 105110 28550
rect 102080 27520 102103 28527
rect 101897 26520 102103 27520
rect 101897 25543 101920 26520
rect 98890 25520 101920 25543
rect 102080 25543 102103 26520
rect 105087 27520 105110 28527
rect 105270 28527 108300 28550
rect 105270 27520 105293 28527
rect 105087 26520 105293 27520
rect 105087 25543 105110 26520
rect 102080 25520 105110 25543
rect 105270 25543 105293 26520
rect 108277 27520 108300 28527
rect 108460 28527 111490 28550
rect 108460 27520 108483 28527
rect 108277 26520 108483 27520
rect 108277 25543 108300 26520
rect 105270 25520 108300 25543
rect 108460 25543 108483 26520
rect 111467 27520 111490 28527
rect 111650 28527 114680 28550
rect 111650 27520 111673 28527
rect 111467 26520 111673 27520
rect 111467 25543 111490 26520
rect 108460 25520 111490 25543
rect 111650 25543 111673 26520
rect 114657 27520 114680 28527
rect 114840 28527 117870 28550
rect 114840 27520 114863 28527
rect 114657 26520 114863 27520
rect 114657 25543 114680 26520
rect 111650 25520 114680 25543
rect 114840 25543 114863 26520
rect 117847 27520 117870 28527
rect 118030 28527 121060 28550
rect 118030 27520 118053 28527
rect 117847 26520 118053 27520
rect 117847 25543 117870 26520
rect 114840 25520 117870 25543
rect 118030 25543 118053 26520
rect 121037 27520 121060 28527
rect 121220 28527 124250 28550
rect 121220 27520 121243 28527
rect 121037 26520 121243 27520
rect 121037 25543 121060 26520
rect 118030 25520 121060 25543
rect 121220 25543 121243 26520
rect 124227 27520 124250 28527
rect 124410 28527 127440 28550
rect 124410 27520 124433 28527
rect 124227 26520 124433 27520
rect 124227 25543 124250 26520
rect 121220 25520 124250 25543
rect 124410 25543 124433 26520
rect 127417 27520 127440 28527
rect 127600 28527 130630 28550
rect 127600 27520 127623 28527
rect 127417 26520 127623 27520
rect 127417 25543 127440 26520
rect 124410 25520 127440 25543
rect 127600 25543 127623 26520
rect 130607 27520 130630 28527
rect 130790 28527 133820 28550
rect 130790 27520 130813 28527
rect 130607 26520 130813 27520
rect 130607 25543 130630 26520
rect 127600 25520 130630 25543
rect 130790 25543 130813 26520
rect 133797 27520 133820 28527
rect 133980 28527 137010 28550
rect 133980 27520 134003 28527
rect 133797 26520 134003 27520
rect 133797 25543 133820 26520
rect 130790 25520 133820 25543
rect 133980 25543 134003 26520
rect 136987 27520 137010 28527
rect 136987 26520 137170 27520
rect 136987 25543 137010 26520
rect 133980 25520 137010 25543
rect 1000 25360 2000 25520
rect 4190 25360 5190 25520
rect 7380 25360 8380 25520
rect 10570 25360 11570 25520
rect 13760 25360 14760 25520
rect 16950 25360 17950 25520
rect 20140 25360 21140 25520
rect 23330 25360 24330 25520
rect 26520 25360 27520 25520
rect 29710 25360 30710 25520
rect 32900 25360 33900 25520
rect 36090 25360 37090 25520
rect 39280 25360 40280 25520
rect 42470 25360 43470 25520
rect 45660 25360 46660 25520
rect 48850 25360 49850 25520
rect 52040 25360 53040 25520
rect 55230 25360 56230 25520
rect 58420 25360 59420 25520
rect 61610 25360 62610 25520
rect 64800 25360 65800 25520
rect 67990 25360 68990 25520
rect 71180 25360 72180 25520
rect 74370 25360 75370 25520
rect 77560 25360 78560 25520
rect 80750 25360 81750 25520
rect 83940 25360 84940 25520
rect 87130 25360 88130 25520
rect 90320 25360 91320 25520
rect 93510 25360 94510 25520
rect 96700 25360 97700 25520
rect 99890 25360 100890 25520
rect 103080 25360 104080 25520
rect 106270 25360 107270 25520
rect 109460 25360 110460 25520
rect 112650 25360 113650 25520
rect 115840 25360 116840 25520
rect 119030 25360 120030 25520
rect 122220 25360 123220 25520
rect 125410 25360 126410 25520
rect 128600 25360 129600 25520
rect 131790 25360 132790 25520
rect 134980 25360 135980 25520
rect 0 25337 3030 25360
rect 0 22353 23 25337
rect 3007 24330 3030 25337
rect 3190 25337 6220 25360
rect 3190 24330 3213 25337
rect 3007 23330 3213 24330
rect 3007 22353 3030 23330
rect 0 22330 3030 22353
rect 3190 22353 3213 23330
rect 6197 24330 6220 25337
rect 6380 25337 9410 25360
rect 6380 24330 6403 25337
rect 6197 23330 6403 24330
rect 6197 22353 6220 23330
rect 3190 22330 6220 22353
rect 6380 22353 6403 23330
rect 9387 24330 9410 25337
rect 9570 25337 12600 25360
rect 9570 24330 9593 25337
rect 9387 23330 9593 24330
rect 9387 22353 9410 23330
rect 6380 22330 9410 22353
rect 9570 22353 9593 23330
rect 12577 24330 12600 25337
rect 12760 25337 15790 25360
rect 12760 24330 12783 25337
rect 12577 23330 12783 24330
rect 12577 22353 12600 23330
rect 9570 22330 12600 22353
rect 12760 22353 12783 23330
rect 15767 24330 15790 25337
rect 15950 25337 18980 25360
rect 15950 24330 15973 25337
rect 15767 23330 15973 24330
rect 15767 22353 15790 23330
rect 12760 22330 15790 22353
rect 15950 22353 15973 23330
rect 18957 24330 18980 25337
rect 19140 25337 22170 25360
rect 19140 24330 19163 25337
rect 18957 23330 19163 24330
rect 18957 22353 18980 23330
rect 15950 22330 18980 22353
rect 19140 22353 19163 23330
rect 22147 24330 22170 25337
rect 22330 25337 25360 25360
rect 22330 24330 22353 25337
rect 22147 23330 22353 24330
rect 22147 22353 22170 23330
rect 19140 22330 22170 22353
rect 22330 22353 22353 23330
rect 25337 24330 25360 25337
rect 25520 25337 28550 25360
rect 25520 24330 25543 25337
rect 25337 23330 25543 24330
rect 25337 22353 25360 23330
rect 22330 22330 25360 22353
rect 25520 22353 25543 23330
rect 28527 24330 28550 25337
rect 28710 25337 31740 25360
rect 28710 24330 28733 25337
rect 28527 23330 28733 24330
rect 28527 22353 28550 23330
rect 25520 22330 28550 22353
rect 28710 22353 28733 23330
rect 31717 24330 31740 25337
rect 31900 25337 34930 25360
rect 31900 24330 31923 25337
rect 31717 23330 31923 24330
rect 31717 22353 31740 23330
rect 28710 22330 31740 22353
rect 31900 22353 31923 23330
rect 34907 24330 34930 25337
rect 35090 25337 38120 25360
rect 35090 24330 35113 25337
rect 34907 23330 35113 24330
rect 34907 22353 34930 23330
rect 31900 22330 34930 22353
rect 35090 22353 35113 23330
rect 38097 24330 38120 25337
rect 38280 25337 41310 25360
rect 38280 24330 38303 25337
rect 38097 23330 38303 24330
rect 38097 22353 38120 23330
rect 35090 22330 38120 22353
rect 38280 22353 38303 23330
rect 41287 24330 41310 25337
rect 41470 25337 44500 25360
rect 41470 24330 41493 25337
rect 41287 23330 41493 24330
rect 41287 22353 41310 23330
rect 38280 22330 41310 22353
rect 41470 22353 41493 23330
rect 44477 24330 44500 25337
rect 44660 25337 47690 25360
rect 44660 24330 44683 25337
rect 44477 23330 44683 24330
rect 44477 22353 44500 23330
rect 41470 22330 44500 22353
rect 44660 22353 44683 23330
rect 47667 24330 47690 25337
rect 47850 25337 50880 25360
rect 47850 24330 47873 25337
rect 47667 23330 47873 24330
rect 47667 22353 47690 23330
rect 44660 22330 47690 22353
rect 47850 22353 47873 23330
rect 50857 24330 50880 25337
rect 51040 25337 54070 25360
rect 51040 24330 51063 25337
rect 50857 23330 51063 24330
rect 50857 22353 50880 23330
rect 47850 22330 50880 22353
rect 51040 22353 51063 23330
rect 54047 24330 54070 25337
rect 54230 25337 57260 25360
rect 54230 24330 54253 25337
rect 54047 23330 54253 24330
rect 54047 22353 54070 23330
rect 51040 22330 54070 22353
rect 54230 22353 54253 23330
rect 57237 24330 57260 25337
rect 57420 25337 60450 25360
rect 57420 24330 57443 25337
rect 57237 23330 57443 24330
rect 57237 22353 57260 23330
rect 54230 22330 57260 22353
rect 57420 22353 57443 23330
rect 60427 24330 60450 25337
rect 60610 25337 63640 25360
rect 60610 24330 60633 25337
rect 60427 23330 60633 24330
rect 60427 22353 60450 23330
rect 57420 22330 60450 22353
rect 60610 22353 60633 23330
rect 63617 24330 63640 25337
rect 63800 25337 66830 25360
rect 63800 24330 63823 25337
rect 63617 23330 63823 24330
rect 63617 22353 63640 23330
rect 60610 22330 63640 22353
rect 63800 22353 63823 23330
rect 66807 24330 66830 25337
rect 66990 25337 70020 25360
rect 66990 24330 67013 25337
rect 66807 23330 67013 24330
rect 66807 22353 66830 23330
rect 63800 22330 66830 22353
rect 66990 22353 67013 23330
rect 69997 24330 70020 25337
rect 70180 25337 73210 25360
rect 70180 24330 70203 25337
rect 69997 23330 70203 24330
rect 69997 22353 70020 23330
rect 66990 22330 70020 22353
rect 70180 22353 70203 23330
rect 73187 24330 73210 25337
rect 73370 25337 76400 25360
rect 73370 24330 73393 25337
rect 73187 23330 73393 24330
rect 73187 22353 73210 23330
rect 70180 22330 73210 22353
rect 73370 22353 73393 23330
rect 76377 24330 76400 25337
rect 76560 25337 79590 25360
rect 76560 24330 76583 25337
rect 76377 23330 76583 24330
rect 76377 22353 76400 23330
rect 73370 22330 76400 22353
rect 76560 22353 76583 23330
rect 79567 24330 79590 25337
rect 79750 25337 82780 25360
rect 79750 24330 79773 25337
rect 79567 23330 79773 24330
rect 79567 22353 79590 23330
rect 76560 22330 79590 22353
rect 79750 22353 79773 23330
rect 82757 24330 82780 25337
rect 82940 25337 85970 25360
rect 82940 24330 82963 25337
rect 82757 23330 82963 24330
rect 82757 22353 82780 23330
rect 79750 22330 82780 22353
rect 82940 22353 82963 23330
rect 85947 24330 85970 25337
rect 86130 25337 89160 25360
rect 86130 24330 86153 25337
rect 85947 23330 86153 24330
rect 85947 22353 85970 23330
rect 82940 22330 85970 22353
rect 86130 22353 86153 23330
rect 89137 24330 89160 25337
rect 89320 25337 92350 25360
rect 89320 24330 89343 25337
rect 89137 23330 89343 24330
rect 89137 22353 89160 23330
rect 86130 22330 89160 22353
rect 89320 22353 89343 23330
rect 92327 24330 92350 25337
rect 92510 25337 95540 25360
rect 92510 24330 92533 25337
rect 92327 23330 92533 24330
rect 92327 22353 92350 23330
rect 89320 22330 92350 22353
rect 92510 22353 92533 23330
rect 95517 24330 95540 25337
rect 95700 25337 98730 25360
rect 95700 24330 95723 25337
rect 95517 23330 95723 24330
rect 95517 22353 95540 23330
rect 92510 22330 95540 22353
rect 95700 22353 95723 23330
rect 98707 24330 98730 25337
rect 98890 25337 101920 25360
rect 98890 24330 98913 25337
rect 98707 23330 98913 24330
rect 98707 22353 98730 23330
rect 95700 22330 98730 22353
rect 98890 22353 98913 23330
rect 101897 24330 101920 25337
rect 102080 25337 105110 25360
rect 102080 24330 102103 25337
rect 101897 23330 102103 24330
rect 101897 22353 101920 23330
rect 98890 22330 101920 22353
rect 102080 22353 102103 23330
rect 105087 24330 105110 25337
rect 105270 25337 108300 25360
rect 105270 24330 105293 25337
rect 105087 23330 105293 24330
rect 105087 22353 105110 23330
rect 102080 22330 105110 22353
rect 105270 22353 105293 23330
rect 108277 24330 108300 25337
rect 108460 25337 111490 25360
rect 108460 24330 108483 25337
rect 108277 23330 108483 24330
rect 108277 22353 108300 23330
rect 105270 22330 108300 22353
rect 108460 22353 108483 23330
rect 111467 24330 111490 25337
rect 111650 25337 114680 25360
rect 111650 24330 111673 25337
rect 111467 23330 111673 24330
rect 111467 22353 111490 23330
rect 108460 22330 111490 22353
rect 111650 22353 111673 23330
rect 114657 24330 114680 25337
rect 114840 25337 117870 25360
rect 114840 24330 114863 25337
rect 114657 23330 114863 24330
rect 114657 22353 114680 23330
rect 111650 22330 114680 22353
rect 114840 22353 114863 23330
rect 117847 24330 117870 25337
rect 118030 25337 121060 25360
rect 118030 24330 118053 25337
rect 117847 23330 118053 24330
rect 117847 22353 117870 23330
rect 114840 22330 117870 22353
rect 118030 22353 118053 23330
rect 121037 24330 121060 25337
rect 121220 25337 124250 25360
rect 121220 24330 121243 25337
rect 121037 23330 121243 24330
rect 121037 22353 121060 23330
rect 118030 22330 121060 22353
rect 121220 22353 121243 23330
rect 124227 24330 124250 25337
rect 124410 25337 127440 25360
rect 124410 24330 124433 25337
rect 124227 23330 124433 24330
rect 124227 22353 124250 23330
rect 121220 22330 124250 22353
rect 124410 22353 124433 23330
rect 127417 24330 127440 25337
rect 127600 25337 130630 25360
rect 127600 24330 127623 25337
rect 127417 23330 127623 24330
rect 127417 22353 127440 23330
rect 124410 22330 127440 22353
rect 127600 22353 127623 23330
rect 130607 24330 130630 25337
rect 130790 25337 133820 25360
rect 130790 24330 130813 25337
rect 130607 23330 130813 24330
rect 130607 22353 130630 23330
rect 127600 22330 130630 22353
rect 130790 22353 130813 23330
rect 133797 24330 133820 25337
rect 133980 25337 137010 25360
rect 133980 24330 134003 25337
rect 133797 23330 134003 24330
rect 133797 22353 133820 23330
rect 130790 22330 133820 22353
rect 133980 22353 134003 23330
rect 136987 24330 137010 25337
rect 136987 23330 137170 24330
rect 136987 22353 137010 23330
rect 133980 22330 137010 22353
rect 1000 22170 2000 22330
rect 4190 22170 5190 22330
rect 7380 22170 8380 22330
rect 10570 22170 11570 22330
rect 13760 22170 14760 22330
rect 16950 22170 17950 22330
rect 20140 22170 21140 22330
rect 23330 22170 24330 22330
rect 26520 22170 27520 22330
rect 29710 22170 30710 22330
rect 32900 22170 33900 22330
rect 36090 22170 37090 22330
rect 39280 22170 40280 22330
rect 42470 22170 43470 22330
rect 45660 22170 46660 22330
rect 48850 22170 49850 22330
rect 52040 22170 53040 22330
rect 55230 22170 56230 22330
rect 58420 22170 59420 22330
rect 61610 22170 62610 22330
rect 64800 22170 65800 22330
rect 67990 22170 68990 22330
rect 71180 22170 72180 22330
rect 74370 22170 75370 22330
rect 77560 22170 78560 22330
rect 80750 22170 81750 22330
rect 83940 22170 84940 22330
rect 87130 22170 88130 22330
rect 90320 22170 91320 22330
rect 93510 22170 94510 22330
rect 96700 22170 97700 22330
rect 99890 22170 100890 22330
rect 103080 22170 104080 22330
rect 106270 22170 107270 22330
rect 109460 22170 110460 22330
rect 112650 22170 113650 22330
rect 115840 22170 116840 22330
rect 119030 22170 120030 22330
rect 122220 22170 123220 22330
rect 125410 22170 126410 22330
rect 128600 22170 129600 22330
rect 131790 22170 132790 22330
rect 134980 22170 135980 22330
rect 0 22147 3030 22170
rect 0 19163 23 22147
rect 3007 21140 3030 22147
rect 3190 22147 6220 22170
rect 3190 21140 3213 22147
rect 3007 20140 3213 21140
rect 3007 19163 3030 20140
rect 0 19140 3030 19163
rect 3190 19163 3213 20140
rect 6197 21140 6220 22147
rect 6380 22147 9410 22170
rect 6380 21140 6403 22147
rect 6197 20140 6403 21140
rect 6197 19163 6220 20140
rect 3190 19140 6220 19163
rect 6380 19163 6403 20140
rect 9387 21140 9410 22147
rect 9570 22147 12600 22170
rect 9570 21140 9593 22147
rect 9387 20140 9593 21140
rect 9387 19163 9410 20140
rect 6380 19140 9410 19163
rect 9570 19163 9593 20140
rect 12577 21140 12600 22147
rect 12760 22147 15790 22170
rect 12760 21140 12783 22147
rect 12577 20140 12783 21140
rect 12577 19163 12600 20140
rect 9570 19140 12600 19163
rect 12760 19163 12783 20140
rect 15767 21140 15790 22147
rect 15950 22147 18980 22170
rect 15950 21140 15973 22147
rect 15767 20140 15973 21140
rect 15767 19163 15790 20140
rect 12760 19140 15790 19163
rect 15950 19163 15973 20140
rect 18957 21140 18980 22147
rect 19140 22147 22170 22170
rect 19140 21140 19163 22147
rect 18957 20140 19163 21140
rect 18957 19163 18980 20140
rect 15950 19140 18980 19163
rect 19140 19163 19163 20140
rect 22147 21140 22170 22147
rect 22330 22147 25360 22170
rect 22330 21140 22353 22147
rect 22147 20140 22353 21140
rect 22147 19163 22170 20140
rect 19140 19140 22170 19163
rect 22330 19163 22353 20140
rect 25337 21140 25360 22147
rect 25520 22147 28550 22170
rect 25520 21140 25543 22147
rect 25337 20140 25543 21140
rect 25337 19163 25360 20140
rect 22330 19140 25360 19163
rect 25520 19163 25543 20140
rect 28527 21140 28550 22147
rect 28710 22147 31740 22170
rect 28710 21140 28733 22147
rect 28527 20140 28733 21140
rect 28527 19163 28550 20140
rect 25520 19140 28550 19163
rect 28710 19163 28733 20140
rect 31717 21140 31740 22147
rect 31900 22147 34930 22170
rect 31900 21140 31923 22147
rect 31717 20140 31923 21140
rect 31717 19163 31740 20140
rect 28710 19140 31740 19163
rect 31900 19163 31923 20140
rect 34907 21140 34930 22147
rect 35090 22147 38120 22170
rect 35090 21140 35113 22147
rect 34907 20140 35113 21140
rect 34907 19163 34930 20140
rect 31900 19140 34930 19163
rect 35090 19163 35113 20140
rect 38097 21140 38120 22147
rect 38280 22147 41310 22170
rect 38280 21140 38303 22147
rect 38097 20140 38303 21140
rect 38097 19163 38120 20140
rect 35090 19140 38120 19163
rect 38280 19163 38303 20140
rect 41287 21140 41310 22147
rect 41470 22147 44500 22170
rect 41470 21140 41493 22147
rect 41287 20140 41493 21140
rect 41287 19163 41310 20140
rect 38280 19140 41310 19163
rect 41470 19163 41493 20140
rect 44477 21140 44500 22147
rect 44660 22147 47690 22170
rect 44660 21140 44683 22147
rect 44477 20140 44683 21140
rect 44477 19163 44500 20140
rect 41470 19140 44500 19163
rect 44660 19163 44683 20140
rect 47667 21140 47690 22147
rect 47850 22147 50880 22170
rect 47850 21140 47873 22147
rect 47667 20140 47873 21140
rect 47667 19163 47690 20140
rect 44660 19140 47690 19163
rect 47850 19163 47873 20140
rect 50857 21140 50880 22147
rect 51040 22147 54070 22170
rect 51040 21140 51063 22147
rect 50857 20140 51063 21140
rect 50857 19163 50880 20140
rect 47850 19140 50880 19163
rect 51040 19163 51063 20140
rect 54047 21140 54070 22147
rect 54230 22147 57260 22170
rect 54230 21140 54253 22147
rect 54047 20140 54253 21140
rect 54047 19163 54070 20140
rect 51040 19140 54070 19163
rect 54230 19163 54253 20140
rect 57237 21140 57260 22147
rect 57420 22147 60450 22170
rect 57420 21140 57443 22147
rect 57237 20140 57443 21140
rect 57237 19163 57260 20140
rect 54230 19140 57260 19163
rect 57420 19163 57443 20140
rect 60427 21140 60450 22147
rect 60610 22147 63640 22170
rect 60610 21140 60633 22147
rect 60427 20140 60633 21140
rect 60427 19163 60450 20140
rect 57420 19140 60450 19163
rect 60610 19163 60633 20140
rect 63617 21140 63640 22147
rect 63800 22147 66830 22170
rect 63800 21140 63823 22147
rect 63617 20140 63823 21140
rect 63617 19163 63640 20140
rect 60610 19140 63640 19163
rect 63800 19163 63823 20140
rect 66807 21140 66830 22147
rect 66990 22147 70020 22170
rect 66990 21140 67013 22147
rect 66807 20140 67013 21140
rect 66807 19163 66830 20140
rect 63800 19140 66830 19163
rect 66990 19163 67013 20140
rect 69997 21140 70020 22147
rect 70180 22147 73210 22170
rect 70180 21140 70203 22147
rect 69997 20140 70203 21140
rect 69997 19163 70020 20140
rect 66990 19140 70020 19163
rect 70180 19163 70203 20140
rect 73187 21140 73210 22147
rect 73370 22147 76400 22170
rect 73370 21140 73393 22147
rect 73187 20140 73393 21140
rect 73187 19163 73210 20140
rect 70180 19140 73210 19163
rect 73370 19163 73393 20140
rect 76377 21140 76400 22147
rect 76560 22147 79590 22170
rect 76560 21140 76583 22147
rect 76377 20140 76583 21140
rect 76377 19163 76400 20140
rect 73370 19140 76400 19163
rect 76560 19163 76583 20140
rect 79567 21140 79590 22147
rect 79750 22147 82780 22170
rect 79750 21140 79773 22147
rect 79567 20140 79773 21140
rect 79567 19163 79590 20140
rect 76560 19140 79590 19163
rect 79750 19163 79773 20140
rect 82757 21140 82780 22147
rect 82940 22147 85970 22170
rect 82940 21140 82963 22147
rect 82757 20140 82963 21140
rect 82757 19163 82780 20140
rect 79750 19140 82780 19163
rect 82940 19163 82963 20140
rect 85947 21140 85970 22147
rect 86130 22147 89160 22170
rect 86130 21140 86153 22147
rect 85947 20140 86153 21140
rect 85947 19163 85970 20140
rect 82940 19140 85970 19163
rect 86130 19163 86153 20140
rect 89137 21140 89160 22147
rect 89320 22147 92350 22170
rect 89320 21140 89343 22147
rect 89137 20140 89343 21140
rect 89137 19163 89160 20140
rect 86130 19140 89160 19163
rect 89320 19163 89343 20140
rect 92327 21140 92350 22147
rect 92510 22147 95540 22170
rect 92510 21140 92533 22147
rect 92327 20140 92533 21140
rect 92327 19163 92350 20140
rect 89320 19140 92350 19163
rect 92510 19163 92533 20140
rect 95517 21140 95540 22147
rect 95700 22147 98730 22170
rect 95700 21140 95723 22147
rect 95517 20140 95723 21140
rect 95517 19163 95540 20140
rect 92510 19140 95540 19163
rect 95700 19163 95723 20140
rect 98707 21140 98730 22147
rect 98890 22147 101920 22170
rect 98890 21140 98913 22147
rect 98707 20140 98913 21140
rect 98707 19163 98730 20140
rect 95700 19140 98730 19163
rect 98890 19163 98913 20140
rect 101897 21140 101920 22147
rect 102080 22147 105110 22170
rect 102080 21140 102103 22147
rect 101897 20140 102103 21140
rect 101897 19163 101920 20140
rect 98890 19140 101920 19163
rect 102080 19163 102103 20140
rect 105087 21140 105110 22147
rect 105270 22147 108300 22170
rect 105270 21140 105293 22147
rect 105087 20140 105293 21140
rect 105087 19163 105110 20140
rect 102080 19140 105110 19163
rect 105270 19163 105293 20140
rect 108277 21140 108300 22147
rect 108460 22147 111490 22170
rect 108460 21140 108483 22147
rect 108277 20140 108483 21140
rect 108277 19163 108300 20140
rect 105270 19140 108300 19163
rect 108460 19163 108483 20140
rect 111467 21140 111490 22147
rect 111650 22147 114680 22170
rect 111650 21140 111673 22147
rect 111467 20140 111673 21140
rect 111467 19163 111490 20140
rect 108460 19140 111490 19163
rect 111650 19163 111673 20140
rect 114657 21140 114680 22147
rect 114840 22147 117870 22170
rect 114840 21140 114863 22147
rect 114657 20140 114863 21140
rect 114657 19163 114680 20140
rect 111650 19140 114680 19163
rect 114840 19163 114863 20140
rect 117847 21140 117870 22147
rect 118030 22147 121060 22170
rect 118030 21140 118053 22147
rect 117847 20140 118053 21140
rect 117847 19163 117870 20140
rect 114840 19140 117870 19163
rect 118030 19163 118053 20140
rect 121037 21140 121060 22147
rect 121220 22147 124250 22170
rect 121220 21140 121243 22147
rect 121037 20140 121243 21140
rect 121037 19163 121060 20140
rect 118030 19140 121060 19163
rect 121220 19163 121243 20140
rect 124227 21140 124250 22147
rect 124410 22147 127440 22170
rect 124410 21140 124433 22147
rect 124227 20140 124433 21140
rect 124227 19163 124250 20140
rect 121220 19140 124250 19163
rect 124410 19163 124433 20140
rect 127417 21140 127440 22147
rect 127600 22147 130630 22170
rect 127600 21140 127623 22147
rect 127417 20140 127623 21140
rect 127417 19163 127440 20140
rect 124410 19140 127440 19163
rect 127600 19163 127623 20140
rect 130607 21140 130630 22147
rect 130790 22147 133820 22170
rect 130790 21140 130813 22147
rect 130607 20140 130813 21140
rect 130607 19163 130630 20140
rect 127600 19140 130630 19163
rect 130790 19163 130813 20140
rect 133797 21140 133820 22147
rect 133980 22147 137010 22170
rect 133980 21140 134003 22147
rect 133797 20140 134003 21140
rect 133797 19163 133820 20140
rect 130790 19140 133820 19163
rect 133980 19163 134003 20140
rect 136987 21140 137010 22147
rect 136987 20140 137170 21140
rect 136987 19163 137010 20140
rect 133980 19140 137010 19163
rect 1000 18980 2000 19140
rect 4190 18980 5190 19140
rect 7380 18980 8380 19140
rect 10570 18980 11570 19140
rect 13760 18980 14760 19140
rect 16950 18980 17950 19140
rect 20140 18980 21140 19140
rect 23330 18980 24330 19140
rect 26520 18980 27520 19140
rect 29710 18980 30710 19140
rect 32900 18980 33900 19140
rect 36090 18980 37090 19140
rect 39280 18980 40280 19140
rect 42470 18980 43470 19140
rect 45660 18980 46660 19140
rect 48850 18980 49850 19140
rect 52040 18980 53040 19140
rect 55230 18980 56230 19140
rect 58420 18980 59420 19140
rect 61610 18980 62610 19140
rect 64800 18980 65800 19140
rect 67990 18980 68990 19140
rect 71180 18980 72180 19140
rect 74370 18980 75370 19140
rect 77560 18980 78560 19140
rect 80750 18980 81750 19140
rect 83940 18980 84940 19140
rect 87130 18980 88130 19140
rect 90320 18980 91320 19140
rect 93510 18980 94510 19140
rect 96700 18980 97700 19140
rect 99890 18980 100890 19140
rect 103080 18980 104080 19140
rect 106270 18980 107270 19140
rect 109460 18980 110460 19140
rect 112650 18980 113650 19140
rect 115840 18980 116840 19140
rect 119030 18980 120030 19140
rect 122220 18980 123220 19140
rect 125410 18980 126410 19140
rect 128600 18980 129600 19140
rect 131790 18980 132790 19140
rect 134980 18980 135980 19140
rect 0 18957 3030 18980
rect 0 15973 23 18957
rect 3007 17950 3030 18957
rect 3190 18957 6220 18980
rect 3190 17950 3213 18957
rect 3007 16950 3213 17950
rect 3007 15973 3030 16950
rect 0 15950 3030 15973
rect 3190 15973 3213 16950
rect 6197 17950 6220 18957
rect 6380 18957 9410 18980
rect 6380 17950 6403 18957
rect 6197 16950 6403 17950
rect 6197 15973 6220 16950
rect 3190 15950 6220 15973
rect 6380 15973 6403 16950
rect 9387 17950 9410 18957
rect 9570 18957 12600 18980
rect 9570 17950 9593 18957
rect 9387 16950 9593 17950
rect 9387 15973 9410 16950
rect 6380 15950 9410 15973
rect 9570 15973 9593 16950
rect 12577 17950 12600 18957
rect 12760 18957 15790 18980
rect 12760 17950 12783 18957
rect 12577 16950 12783 17950
rect 12577 15973 12600 16950
rect 9570 15950 12600 15973
rect 12760 15973 12783 16950
rect 15767 17950 15790 18957
rect 15950 18957 18980 18980
rect 15950 17950 15973 18957
rect 15767 16950 15973 17950
rect 15767 15973 15790 16950
rect 12760 15950 15790 15973
rect 15950 15973 15973 16950
rect 18957 17950 18980 18957
rect 19140 18957 22170 18980
rect 19140 17950 19163 18957
rect 18957 16950 19163 17950
rect 18957 15973 18980 16950
rect 15950 15950 18980 15973
rect 19140 15973 19163 16950
rect 22147 17950 22170 18957
rect 22330 18957 25360 18980
rect 22330 17950 22353 18957
rect 22147 16950 22353 17950
rect 22147 15973 22170 16950
rect 19140 15950 22170 15973
rect 22330 15973 22353 16950
rect 25337 17950 25360 18957
rect 25520 18957 28550 18980
rect 25520 17950 25543 18957
rect 25337 16950 25543 17950
rect 25337 15973 25360 16950
rect 22330 15950 25360 15973
rect 25520 15973 25543 16950
rect 28527 17950 28550 18957
rect 28710 18957 31740 18980
rect 28710 17950 28733 18957
rect 28527 16950 28733 17950
rect 28527 15973 28550 16950
rect 25520 15950 28550 15973
rect 28710 15973 28733 16950
rect 31717 17950 31740 18957
rect 31900 18957 34930 18980
rect 31900 17950 31923 18957
rect 31717 16950 31923 17950
rect 31717 15973 31740 16950
rect 28710 15950 31740 15973
rect 31900 15973 31923 16950
rect 34907 17950 34930 18957
rect 35090 18957 38120 18980
rect 35090 17950 35113 18957
rect 34907 16950 35113 17950
rect 34907 15973 34930 16950
rect 31900 15950 34930 15973
rect 35090 15973 35113 16950
rect 38097 17950 38120 18957
rect 38280 18957 41310 18980
rect 38280 17950 38303 18957
rect 38097 16950 38303 17950
rect 38097 15973 38120 16950
rect 35090 15950 38120 15973
rect 38280 15973 38303 16950
rect 41287 17950 41310 18957
rect 41470 18957 44500 18980
rect 41470 17950 41493 18957
rect 41287 16950 41493 17950
rect 41287 15973 41310 16950
rect 38280 15950 41310 15973
rect 41470 15973 41493 16950
rect 44477 17950 44500 18957
rect 44660 18957 47690 18980
rect 44660 17950 44683 18957
rect 44477 16950 44683 17950
rect 44477 15973 44500 16950
rect 41470 15950 44500 15973
rect 44660 15973 44683 16950
rect 47667 17950 47690 18957
rect 47850 18957 50880 18980
rect 47850 17950 47873 18957
rect 47667 16950 47873 17950
rect 47667 15973 47690 16950
rect 44660 15950 47690 15973
rect 47850 15973 47873 16950
rect 50857 17950 50880 18957
rect 51040 18957 54070 18980
rect 51040 17950 51063 18957
rect 50857 16950 51063 17950
rect 50857 15973 50880 16950
rect 47850 15950 50880 15973
rect 51040 15973 51063 16950
rect 54047 17950 54070 18957
rect 54230 18957 57260 18980
rect 54230 17950 54253 18957
rect 54047 16950 54253 17950
rect 54047 15973 54070 16950
rect 51040 15950 54070 15973
rect 54230 15973 54253 16950
rect 57237 17950 57260 18957
rect 57420 18957 60450 18980
rect 57420 17950 57443 18957
rect 57237 16950 57443 17950
rect 57237 15973 57260 16950
rect 54230 15950 57260 15973
rect 57420 15973 57443 16950
rect 60427 17950 60450 18957
rect 60610 18957 63640 18980
rect 60610 17950 60633 18957
rect 60427 16950 60633 17950
rect 60427 15973 60450 16950
rect 57420 15950 60450 15973
rect 60610 15973 60633 16950
rect 63617 17950 63640 18957
rect 63800 18957 66830 18980
rect 63800 17950 63823 18957
rect 63617 16950 63823 17950
rect 63617 15973 63640 16950
rect 60610 15950 63640 15973
rect 63800 15973 63823 16950
rect 66807 17950 66830 18957
rect 66990 18957 70020 18980
rect 66990 17950 67013 18957
rect 66807 16950 67013 17950
rect 66807 15973 66830 16950
rect 63800 15950 66830 15973
rect 66990 15973 67013 16950
rect 69997 17950 70020 18957
rect 70180 18957 73210 18980
rect 70180 17950 70203 18957
rect 69997 16950 70203 17950
rect 69997 15973 70020 16950
rect 66990 15950 70020 15973
rect 70180 15973 70203 16950
rect 73187 17950 73210 18957
rect 73370 18957 76400 18980
rect 73370 17950 73393 18957
rect 73187 16950 73393 17950
rect 73187 15973 73210 16950
rect 70180 15950 73210 15973
rect 73370 15973 73393 16950
rect 76377 17950 76400 18957
rect 76560 18957 79590 18980
rect 76560 17950 76583 18957
rect 76377 16950 76583 17950
rect 76377 15973 76400 16950
rect 73370 15950 76400 15973
rect 76560 15973 76583 16950
rect 79567 17950 79590 18957
rect 79750 18957 82780 18980
rect 79750 17950 79773 18957
rect 79567 16950 79773 17950
rect 79567 15973 79590 16950
rect 76560 15950 79590 15973
rect 79750 15973 79773 16950
rect 82757 17950 82780 18957
rect 82940 18957 85970 18980
rect 82940 17950 82963 18957
rect 82757 16950 82963 17950
rect 82757 15973 82780 16950
rect 79750 15950 82780 15973
rect 82940 15973 82963 16950
rect 85947 17950 85970 18957
rect 86130 18957 89160 18980
rect 86130 17950 86153 18957
rect 85947 16950 86153 17950
rect 85947 15973 85970 16950
rect 82940 15950 85970 15973
rect 86130 15973 86153 16950
rect 89137 17950 89160 18957
rect 89320 18957 92350 18980
rect 89320 17950 89343 18957
rect 89137 16950 89343 17950
rect 89137 15973 89160 16950
rect 86130 15950 89160 15973
rect 89320 15973 89343 16950
rect 92327 17950 92350 18957
rect 92510 18957 95540 18980
rect 92510 17950 92533 18957
rect 92327 16950 92533 17950
rect 92327 15973 92350 16950
rect 89320 15950 92350 15973
rect 92510 15973 92533 16950
rect 95517 17950 95540 18957
rect 95700 18957 98730 18980
rect 95700 17950 95723 18957
rect 95517 16950 95723 17950
rect 95517 15973 95540 16950
rect 92510 15950 95540 15973
rect 95700 15973 95723 16950
rect 98707 17950 98730 18957
rect 98890 18957 101920 18980
rect 98890 17950 98913 18957
rect 98707 16950 98913 17950
rect 98707 15973 98730 16950
rect 95700 15950 98730 15973
rect 98890 15973 98913 16950
rect 101897 17950 101920 18957
rect 102080 18957 105110 18980
rect 102080 17950 102103 18957
rect 101897 16950 102103 17950
rect 101897 15973 101920 16950
rect 98890 15950 101920 15973
rect 102080 15973 102103 16950
rect 105087 17950 105110 18957
rect 105270 18957 108300 18980
rect 105270 17950 105293 18957
rect 105087 16950 105293 17950
rect 105087 15973 105110 16950
rect 102080 15950 105110 15973
rect 105270 15973 105293 16950
rect 108277 17950 108300 18957
rect 108460 18957 111490 18980
rect 108460 17950 108483 18957
rect 108277 16950 108483 17950
rect 108277 15973 108300 16950
rect 105270 15950 108300 15973
rect 108460 15973 108483 16950
rect 111467 17950 111490 18957
rect 111650 18957 114680 18980
rect 111650 17950 111673 18957
rect 111467 16950 111673 17950
rect 111467 15973 111490 16950
rect 108460 15950 111490 15973
rect 111650 15973 111673 16950
rect 114657 17950 114680 18957
rect 114840 18957 117870 18980
rect 114840 17950 114863 18957
rect 114657 16950 114863 17950
rect 114657 15973 114680 16950
rect 111650 15950 114680 15973
rect 114840 15973 114863 16950
rect 117847 17950 117870 18957
rect 118030 18957 121060 18980
rect 118030 17950 118053 18957
rect 117847 16950 118053 17950
rect 117847 15973 117870 16950
rect 114840 15950 117870 15973
rect 118030 15973 118053 16950
rect 121037 17950 121060 18957
rect 121220 18957 124250 18980
rect 121220 17950 121243 18957
rect 121037 16950 121243 17950
rect 121037 15973 121060 16950
rect 118030 15950 121060 15973
rect 121220 15973 121243 16950
rect 124227 17950 124250 18957
rect 124410 18957 127440 18980
rect 124410 17950 124433 18957
rect 124227 16950 124433 17950
rect 124227 15973 124250 16950
rect 121220 15950 124250 15973
rect 124410 15973 124433 16950
rect 127417 17950 127440 18957
rect 127600 18957 130630 18980
rect 127600 17950 127623 18957
rect 127417 16950 127623 17950
rect 127417 15973 127440 16950
rect 124410 15950 127440 15973
rect 127600 15973 127623 16950
rect 130607 17950 130630 18957
rect 130790 18957 133820 18980
rect 130790 17950 130813 18957
rect 130607 16950 130813 17950
rect 130607 15973 130630 16950
rect 127600 15950 130630 15973
rect 130790 15973 130813 16950
rect 133797 17950 133820 18957
rect 133980 18957 137010 18980
rect 133980 17950 134003 18957
rect 133797 16950 134003 17950
rect 133797 15973 133820 16950
rect 130790 15950 133820 15973
rect 133980 15973 134003 16950
rect 136987 17950 137010 18957
rect 136987 16950 137170 17950
rect 136987 15973 137010 16950
rect 133980 15950 137010 15973
rect 1000 15790 2000 15950
rect 4190 15790 5190 15950
rect 7380 15790 8380 15950
rect 10570 15790 11570 15950
rect 13760 15790 14760 15950
rect 16950 15790 17950 15950
rect 20140 15790 21140 15950
rect 23330 15790 24330 15950
rect 26520 15790 27520 15950
rect 29710 15790 30710 15950
rect 32900 15790 33900 15950
rect 36090 15790 37090 15950
rect 39280 15790 40280 15950
rect 42470 15790 43470 15950
rect 45660 15790 46660 15950
rect 48850 15790 49850 15950
rect 52040 15790 53040 15950
rect 55230 15790 56230 15950
rect 58420 15790 59420 15950
rect 61610 15790 62610 15950
rect 64800 15790 65800 15950
rect 67990 15790 68990 15950
rect 71180 15790 72180 15950
rect 74370 15790 75370 15950
rect 77560 15790 78560 15950
rect 80750 15790 81750 15950
rect 83940 15790 84940 15950
rect 87130 15790 88130 15950
rect 90320 15790 91320 15950
rect 93510 15790 94510 15950
rect 96700 15790 97700 15950
rect 99890 15790 100890 15950
rect 103080 15790 104080 15950
rect 106270 15790 107270 15950
rect 109460 15790 110460 15950
rect 112650 15790 113650 15950
rect 115840 15790 116840 15950
rect 119030 15790 120030 15950
rect 122220 15790 123220 15950
rect 125410 15790 126410 15950
rect 128600 15790 129600 15950
rect 131790 15790 132790 15950
rect 134980 15790 135980 15950
rect 0 15767 3030 15790
rect 0 12783 23 15767
rect 3007 14760 3030 15767
rect 3190 15767 6220 15790
rect 3190 14760 3213 15767
rect 3007 13760 3213 14760
rect 3007 12783 3030 13760
rect 0 12760 3030 12783
rect 3190 12783 3213 13760
rect 6197 14760 6220 15767
rect 6380 15767 9410 15790
rect 6380 14760 6403 15767
rect 6197 13760 6403 14760
rect 6197 12783 6220 13760
rect 3190 12760 6220 12783
rect 6380 12783 6403 13760
rect 9387 14760 9410 15767
rect 9570 15767 12600 15790
rect 9570 14760 9593 15767
rect 9387 13760 9593 14760
rect 9387 12783 9410 13760
rect 6380 12760 9410 12783
rect 9570 12783 9593 13760
rect 12577 14760 12600 15767
rect 12760 15767 15790 15790
rect 12760 14760 12783 15767
rect 12577 13760 12783 14760
rect 12577 12783 12600 13760
rect 9570 12760 12600 12783
rect 12760 12783 12783 13760
rect 15767 14760 15790 15767
rect 15950 15767 18980 15790
rect 15950 14760 15973 15767
rect 15767 13760 15973 14760
rect 15767 12783 15790 13760
rect 12760 12760 15790 12783
rect 15950 12783 15973 13760
rect 18957 14760 18980 15767
rect 19140 15767 22170 15790
rect 19140 14760 19163 15767
rect 18957 13760 19163 14760
rect 18957 12783 18980 13760
rect 15950 12760 18980 12783
rect 19140 12783 19163 13760
rect 22147 14760 22170 15767
rect 22330 15767 25360 15790
rect 22330 14760 22353 15767
rect 22147 13760 22353 14760
rect 22147 12783 22170 13760
rect 19140 12760 22170 12783
rect 22330 12783 22353 13760
rect 25337 14760 25360 15767
rect 25520 15767 28550 15790
rect 25520 14760 25543 15767
rect 25337 13760 25543 14760
rect 25337 12783 25360 13760
rect 22330 12760 25360 12783
rect 25520 12783 25543 13760
rect 28527 14760 28550 15767
rect 28710 15767 31740 15790
rect 28710 14760 28733 15767
rect 28527 13760 28733 14760
rect 28527 12783 28550 13760
rect 25520 12760 28550 12783
rect 28710 12783 28733 13760
rect 31717 14760 31740 15767
rect 31900 15767 34930 15790
rect 31900 14760 31923 15767
rect 31717 13760 31923 14760
rect 31717 12783 31740 13760
rect 28710 12760 31740 12783
rect 31900 12783 31923 13760
rect 34907 14760 34930 15767
rect 35090 15767 38120 15790
rect 35090 14760 35113 15767
rect 34907 13760 35113 14760
rect 34907 12783 34930 13760
rect 31900 12760 34930 12783
rect 35090 12783 35113 13760
rect 38097 14760 38120 15767
rect 38280 15767 41310 15790
rect 38280 14760 38303 15767
rect 38097 13760 38303 14760
rect 38097 12783 38120 13760
rect 35090 12760 38120 12783
rect 38280 12783 38303 13760
rect 41287 14760 41310 15767
rect 41470 15767 44500 15790
rect 41470 14760 41493 15767
rect 41287 13760 41493 14760
rect 41287 12783 41310 13760
rect 38280 12760 41310 12783
rect 41470 12783 41493 13760
rect 44477 14760 44500 15767
rect 44660 15767 47690 15790
rect 44660 14760 44683 15767
rect 44477 13760 44683 14760
rect 44477 12783 44500 13760
rect 41470 12760 44500 12783
rect 44660 12783 44683 13760
rect 47667 14760 47690 15767
rect 47850 15767 50880 15790
rect 47850 14760 47873 15767
rect 47667 13760 47873 14760
rect 47667 12783 47690 13760
rect 44660 12760 47690 12783
rect 47850 12783 47873 13760
rect 50857 14760 50880 15767
rect 51040 15767 54070 15790
rect 51040 14760 51063 15767
rect 50857 13760 51063 14760
rect 50857 12783 50880 13760
rect 47850 12760 50880 12783
rect 51040 12783 51063 13760
rect 54047 14760 54070 15767
rect 54230 15767 57260 15790
rect 54230 14760 54253 15767
rect 54047 13760 54253 14760
rect 54047 12783 54070 13760
rect 51040 12760 54070 12783
rect 54230 12783 54253 13760
rect 57237 14760 57260 15767
rect 57420 15767 60450 15790
rect 57420 14760 57443 15767
rect 57237 13760 57443 14760
rect 57237 12783 57260 13760
rect 54230 12760 57260 12783
rect 57420 12783 57443 13760
rect 60427 14760 60450 15767
rect 60610 15767 63640 15790
rect 60610 14760 60633 15767
rect 60427 13760 60633 14760
rect 60427 12783 60450 13760
rect 57420 12760 60450 12783
rect 60610 12783 60633 13760
rect 63617 14760 63640 15767
rect 63800 15767 66830 15790
rect 63800 14760 63823 15767
rect 63617 13760 63823 14760
rect 63617 12783 63640 13760
rect 60610 12760 63640 12783
rect 63800 12783 63823 13760
rect 66807 14760 66830 15767
rect 66990 15767 70020 15790
rect 66990 14760 67013 15767
rect 66807 13760 67013 14760
rect 66807 12783 66830 13760
rect 63800 12760 66830 12783
rect 66990 12783 67013 13760
rect 69997 14760 70020 15767
rect 70180 15767 73210 15790
rect 70180 14760 70203 15767
rect 69997 13760 70203 14760
rect 69997 12783 70020 13760
rect 66990 12760 70020 12783
rect 70180 12783 70203 13760
rect 73187 14760 73210 15767
rect 73370 15767 76400 15790
rect 73370 14760 73393 15767
rect 73187 13760 73393 14760
rect 73187 12783 73210 13760
rect 70180 12760 73210 12783
rect 73370 12783 73393 13760
rect 76377 14760 76400 15767
rect 76560 15767 79590 15790
rect 76560 14760 76583 15767
rect 76377 13760 76583 14760
rect 76377 12783 76400 13760
rect 73370 12760 76400 12783
rect 76560 12783 76583 13760
rect 79567 14760 79590 15767
rect 79750 15767 82780 15790
rect 79750 14760 79773 15767
rect 79567 13760 79773 14760
rect 79567 12783 79590 13760
rect 76560 12760 79590 12783
rect 79750 12783 79773 13760
rect 82757 14760 82780 15767
rect 82940 15767 85970 15790
rect 82940 14760 82963 15767
rect 82757 13760 82963 14760
rect 82757 12783 82780 13760
rect 79750 12760 82780 12783
rect 82940 12783 82963 13760
rect 85947 14760 85970 15767
rect 86130 15767 89160 15790
rect 86130 14760 86153 15767
rect 85947 13760 86153 14760
rect 85947 12783 85970 13760
rect 82940 12760 85970 12783
rect 86130 12783 86153 13760
rect 89137 14760 89160 15767
rect 89320 15767 92350 15790
rect 89320 14760 89343 15767
rect 89137 13760 89343 14760
rect 89137 12783 89160 13760
rect 86130 12760 89160 12783
rect 89320 12783 89343 13760
rect 92327 14760 92350 15767
rect 92510 15767 95540 15790
rect 92510 14760 92533 15767
rect 92327 13760 92533 14760
rect 92327 12783 92350 13760
rect 89320 12760 92350 12783
rect 92510 12783 92533 13760
rect 95517 14760 95540 15767
rect 95700 15767 98730 15790
rect 95700 14760 95723 15767
rect 95517 13760 95723 14760
rect 95517 12783 95540 13760
rect 92510 12760 95540 12783
rect 95700 12783 95723 13760
rect 98707 14760 98730 15767
rect 98890 15767 101920 15790
rect 98890 14760 98913 15767
rect 98707 13760 98913 14760
rect 98707 12783 98730 13760
rect 95700 12760 98730 12783
rect 98890 12783 98913 13760
rect 101897 14760 101920 15767
rect 102080 15767 105110 15790
rect 102080 14760 102103 15767
rect 101897 13760 102103 14760
rect 101897 12783 101920 13760
rect 98890 12760 101920 12783
rect 102080 12783 102103 13760
rect 105087 14760 105110 15767
rect 105270 15767 108300 15790
rect 105270 14760 105293 15767
rect 105087 13760 105293 14760
rect 105087 12783 105110 13760
rect 102080 12760 105110 12783
rect 105270 12783 105293 13760
rect 108277 14760 108300 15767
rect 108460 15767 111490 15790
rect 108460 14760 108483 15767
rect 108277 13760 108483 14760
rect 108277 12783 108300 13760
rect 105270 12760 108300 12783
rect 108460 12783 108483 13760
rect 111467 14760 111490 15767
rect 111650 15767 114680 15790
rect 111650 14760 111673 15767
rect 111467 13760 111673 14760
rect 111467 12783 111490 13760
rect 108460 12760 111490 12783
rect 111650 12783 111673 13760
rect 114657 14760 114680 15767
rect 114840 15767 117870 15790
rect 114840 14760 114863 15767
rect 114657 13760 114863 14760
rect 114657 12783 114680 13760
rect 111650 12760 114680 12783
rect 114840 12783 114863 13760
rect 117847 14760 117870 15767
rect 118030 15767 121060 15790
rect 118030 14760 118053 15767
rect 117847 13760 118053 14760
rect 117847 12783 117870 13760
rect 114840 12760 117870 12783
rect 118030 12783 118053 13760
rect 121037 14760 121060 15767
rect 121220 15767 124250 15790
rect 121220 14760 121243 15767
rect 121037 13760 121243 14760
rect 121037 12783 121060 13760
rect 118030 12760 121060 12783
rect 121220 12783 121243 13760
rect 124227 14760 124250 15767
rect 124410 15767 127440 15790
rect 124410 14760 124433 15767
rect 124227 13760 124433 14760
rect 124227 12783 124250 13760
rect 121220 12760 124250 12783
rect 124410 12783 124433 13760
rect 127417 14760 127440 15767
rect 127600 15767 130630 15790
rect 127600 14760 127623 15767
rect 127417 13760 127623 14760
rect 127417 12783 127440 13760
rect 124410 12760 127440 12783
rect 127600 12783 127623 13760
rect 130607 14760 130630 15767
rect 130790 15767 133820 15790
rect 130790 14760 130813 15767
rect 130607 13760 130813 14760
rect 130607 12783 130630 13760
rect 127600 12760 130630 12783
rect 130790 12783 130813 13760
rect 133797 14760 133820 15767
rect 133980 15767 137010 15790
rect 133980 14760 134003 15767
rect 133797 13760 134003 14760
rect 133797 12783 133820 13760
rect 130790 12760 133820 12783
rect 133980 12783 134003 13760
rect 136987 14760 137010 15767
rect 136987 13760 137170 14760
rect 136987 12783 137010 13760
rect 133980 12760 137010 12783
rect 1000 12600 2000 12760
rect 4190 12600 5190 12760
rect 7380 12600 8380 12760
rect 10570 12600 11570 12760
rect 13760 12600 14760 12760
rect 16950 12600 17950 12760
rect 20140 12600 21140 12760
rect 23330 12600 24330 12760
rect 26520 12600 27520 12760
rect 29710 12600 30710 12760
rect 32900 12600 33900 12760
rect 36090 12600 37090 12760
rect 39280 12600 40280 12760
rect 42470 12600 43470 12760
rect 45660 12600 46660 12760
rect 48850 12600 49850 12760
rect 52040 12600 53040 12760
rect 55230 12600 56230 12760
rect 58420 12600 59420 12760
rect 61610 12600 62610 12760
rect 64800 12600 65800 12760
rect 67990 12600 68990 12760
rect 71180 12600 72180 12760
rect 74370 12600 75370 12760
rect 77560 12600 78560 12760
rect 80750 12600 81750 12760
rect 83940 12600 84940 12760
rect 87130 12600 88130 12760
rect 90320 12600 91320 12760
rect 93510 12600 94510 12760
rect 96700 12600 97700 12760
rect 99890 12600 100890 12760
rect 103080 12600 104080 12760
rect 106270 12600 107270 12760
rect 109460 12600 110460 12760
rect 112650 12600 113650 12760
rect 115840 12600 116840 12760
rect 119030 12600 120030 12760
rect 122220 12600 123220 12760
rect 125410 12600 126410 12760
rect 128600 12600 129600 12760
rect 131790 12600 132790 12760
rect 134980 12600 135980 12760
rect 0 12577 3030 12600
rect 0 9593 23 12577
rect 3007 11570 3030 12577
rect 3190 12577 6220 12600
rect 3190 11570 3213 12577
rect 3007 10570 3213 11570
rect 3007 9593 3030 10570
rect 0 9570 3030 9593
rect 3190 9593 3213 10570
rect 6197 11570 6220 12577
rect 6380 12577 9410 12600
rect 6380 11570 6403 12577
rect 6197 10570 6403 11570
rect 6197 9593 6220 10570
rect 3190 9570 6220 9593
rect 6380 9593 6403 10570
rect 9387 11570 9410 12577
rect 9570 12577 12600 12600
rect 9570 11570 9593 12577
rect 9387 10570 9593 11570
rect 9387 9593 9410 10570
rect 6380 9570 9410 9593
rect 9570 9593 9593 10570
rect 12577 11570 12600 12577
rect 12760 12577 15790 12600
rect 12760 11570 12783 12577
rect 12577 10570 12783 11570
rect 12577 9593 12600 10570
rect 9570 9570 12600 9593
rect 12760 9593 12783 10570
rect 15767 11570 15790 12577
rect 15950 12577 18980 12600
rect 15950 11570 15973 12577
rect 15767 10570 15973 11570
rect 15767 9593 15790 10570
rect 12760 9570 15790 9593
rect 15950 9593 15973 10570
rect 18957 11570 18980 12577
rect 19140 12577 22170 12600
rect 19140 11570 19163 12577
rect 18957 10570 19163 11570
rect 18957 9593 18980 10570
rect 15950 9570 18980 9593
rect 19140 9593 19163 10570
rect 22147 11570 22170 12577
rect 22330 12577 25360 12600
rect 22330 11570 22353 12577
rect 22147 10570 22353 11570
rect 22147 9593 22170 10570
rect 19140 9570 22170 9593
rect 22330 9593 22353 10570
rect 25337 11570 25360 12577
rect 25520 12577 28550 12600
rect 25520 11570 25543 12577
rect 25337 10570 25543 11570
rect 25337 9593 25360 10570
rect 22330 9570 25360 9593
rect 25520 9593 25543 10570
rect 28527 11570 28550 12577
rect 28710 12577 31740 12600
rect 28710 11570 28733 12577
rect 28527 10570 28733 11570
rect 28527 9593 28550 10570
rect 25520 9570 28550 9593
rect 28710 9593 28733 10570
rect 31717 11570 31740 12577
rect 31900 12577 34930 12600
rect 31900 11570 31923 12577
rect 31717 10570 31923 11570
rect 31717 9593 31740 10570
rect 28710 9570 31740 9593
rect 31900 9593 31923 10570
rect 34907 11570 34930 12577
rect 35090 12577 38120 12600
rect 35090 11570 35113 12577
rect 34907 10570 35113 11570
rect 34907 9593 34930 10570
rect 31900 9570 34930 9593
rect 35090 9593 35113 10570
rect 38097 11570 38120 12577
rect 38280 12577 41310 12600
rect 38280 11570 38303 12577
rect 38097 10570 38303 11570
rect 38097 9593 38120 10570
rect 35090 9570 38120 9593
rect 38280 9593 38303 10570
rect 41287 11570 41310 12577
rect 41470 12577 44500 12600
rect 41470 11570 41493 12577
rect 41287 10570 41493 11570
rect 41287 9593 41310 10570
rect 38280 9570 41310 9593
rect 41470 9593 41493 10570
rect 44477 11570 44500 12577
rect 44660 12577 47690 12600
rect 44660 11570 44683 12577
rect 44477 10570 44683 11570
rect 44477 9593 44500 10570
rect 41470 9570 44500 9593
rect 44660 9593 44683 10570
rect 47667 11570 47690 12577
rect 47850 12577 50880 12600
rect 47850 11570 47873 12577
rect 47667 10570 47873 11570
rect 47667 9593 47690 10570
rect 44660 9570 47690 9593
rect 47850 9593 47873 10570
rect 50857 11570 50880 12577
rect 51040 12577 54070 12600
rect 51040 11570 51063 12577
rect 50857 10570 51063 11570
rect 50857 9593 50880 10570
rect 47850 9570 50880 9593
rect 51040 9593 51063 10570
rect 54047 11570 54070 12577
rect 54230 12577 57260 12600
rect 54230 11570 54253 12577
rect 54047 10570 54253 11570
rect 54047 9593 54070 10570
rect 51040 9570 54070 9593
rect 54230 9593 54253 10570
rect 57237 11570 57260 12577
rect 57420 12577 60450 12600
rect 57420 11570 57443 12577
rect 57237 10570 57443 11570
rect 57237 9593 57260 10570
rect 54230 9570 57260 9593
rect 57420 9593 57443 10570
rect 60427 11570 60450 12577
rect 60610 12577 63640 12600
rect 60610 11570 60633 12577
rect 60427 10570 60633 11570
rect 60427 9593 60450 10570
rect 57420 9570 60450 9593
rect 60610 9593 60633 10570
rect 63617 11570 63640 12577
rect 63800 12577 66830 12600
rect 63800 11570 63823 12577
rect 63617 10570 63823 11570
rect 63617 9593 63640 10570
rect 60610 9570 63640 9593
rect 63800 9593 63823 10570
rect 66807 11570 66830 12577
rect 66990 12577 70020 12600
rect 66990 11570 67013 12577
rect 66807 10570 67013 11570
rect 66807 9593 66830 10570
rect 63800 9570 66830 9593
rect 66990 9593 67013 10570
rect 69997 11570 70020 12577
rect 70180 12577 73210 12600
rect 70180 11570 70203 12577
rect 69997 10570 70203 11570
rect 69997 9593 70020 10570
rect 66990 9570 70020 9593
rect 70180 9593 70203 10570
rect 73187 11570 73210 12577
rect 73370 12577 76400 12600
rect 73370 11570 73393 12577
rect 73187 10570 73393 11570
rect 73187 9593 73210 10570
rect 70180 9570 73210 9593
rect 73370 9593 73393 10570
rect 76377 11570 76400 12577
rect 76560 12577 79590 12600
rect 76560 11570 76583 12577
rect 76377 10570 76583 11570
rect 76377 9593 76400 10570
rect 73370 9570 76400 9593
rect 76560 9593 76583 10570
rect 79567 11570 79590 12577
rect 79750 12577 82780 12600
rect 79750 11570 79773 12577
rect 79567 10570 79773 11570
rect 79567 9593 79590 10570
rect 76560 9570 79590 9593
rect 79750 9593 79773 10570
rect 82757 11570 82780 12577
rect 82940 12577 85970 12600
rect 82940 11570 82963 12577
rect 82757 10570 82963 11570
rect 82757 9593 82780 10570
rect 79750 9570 82780 9593
rect 82940 9593 82963 10570
rect 85947 11570 85970 12577
rect 86130 12577 89160 12600
rect 86130 11570 86153 12577
rect 85947 10570 86153 11570
rect 85947 9593 85970 10570
rect 82940 9570 85970 9593
rect 86130 9593 86153 10570
rect 89137 11570 89160 12577
rect 89320 12577 92350 12600
rect 89320 11570 89343 12577
rect 89137 10570 89343 11570
rect 89137 9593 89160 10570
rect 86130 9570 89160 9593
rect 89320 9593 89343 10570
rect 92327 11570 92350 12577
rect 92510 12577 95540 12600
rect 92510 11570 92533 12577
rect 92327 10570 92533 11570
rect 92327 9593 92350 10570
rect 89320 9570 92350 9593
rect 92510 9593 92533 10570
rect 95517 11570 95540 12577
rect 95700 12577 98730 12600
rect 95700 11570 95723 12577
rect 95517 10570 95723 11570
rect 95517 9593 95540 10570
rect 92510 9570 95540 9593
rect 95700 9593 95723 10570
rect 98707 11570 98730 12577
rect 98890 12577 101920 12600
rect 98890 11570 98913 12577
rect 98707 10570 98913 11570
rect 98707 9593 98730 10570
rect 95700 9570 98730 9593
rect 98890 9593 98913 10570
rect 101897 11570 101920 12577
rect 102080 12577 105110 12600
rect 102080 11570 102103 12577
rect 101897 10570 102103 11570
rect 101897 9593 101920 10570
rect 98890 9570 101920 9593
rect 102080 9593 102103 10570
rect 105087 11570 105110 12577
rect 105270 12577 108300 12600
rect 105270 11570 105293 12577
rect 105087 10570 105293 11570
rect 105087 9593 105110 10570
rect 102080 9570 105110 9593
rect 105270 9593 105293 10570
rect 108277 11570 108300 12577
rect 108460 12577 111490 12600
rect 108460 11570 108483 12577
rect 108277 10570 108483 11570
rect 108277 9593 108300 10570
rect 105270 9570 108300 9593
rect 108460 9593 108483 10570
rect 111467 11570 111490 12577
rect 111650 12577 114680 12600
rect 111650 11570 111673 12577
rect 111467 10570 111673 11570
rect 111467 9593 111490 10570
rect 108460 9570 111490 9593
rect 111650 9593 111673 10570
rect 114657 11570 114680 12577
rect 114840 12577 117870 12600
rect 114840 11570 114863 12577
rect 114657 10570 114863 11570
rect 114657 9593 114680 10570
rect 111650 9570 114680 9593
rect 114840 9593 114863 10570
rect 117847 11570 117870 12577
rect 118030 12577 121060 12600
rect 118030 11570 118053 12577
rect 117847 10570 118053 11570
rect 117847 9593 117870 10570
rect 114840 9570 117870 9593
rect 118030 9593 118053 10570
rect 121037 11570 121060 12577
rect 121220 12577 124250 12600
rect 121220 11570 121243 12577
rect 121037 10570 121243 11570
rect 121037 9593 121060 10570
rect 118030 9570 121060 9593
rect 121220 9593 121243 10570
rect 124227 11570 124250 12577
rect 124410 12577 127440 12600
rect 124410 11570 124433 12577
rect 124227 10570 124433 11570
rect 124227 9593 124250 10570
rect 121220 9570 124250 9593
rect 124410 9593 124433 10570
rect 127417 11570 127440 12577
rect 127600 12577 130630 12600
rect 127600 11570 127623 12577
rect 127417 10570 127623 11570
rect 127417 9593 127440 10570
rect 124410 9570 127440 9593
rect 127600 9593 127623 10570
rect 130607 11570 130630 12577
rect 130790 12577 133820 12600
rect 130790 11570 130813 12577
rect 130607 10570 130813 11570
rect 130607 9593 130630 10570
rect 127600 9570 130630 9593
rect 130790 9593 130813 10570
rect 133797 11570 133820 12577
rect 133980 12577 137010 12600
rect 133980 11570 134003 12577
rect 133797 10570 134003 11570
rect 133797 9593 133820 10570
rect 130790 9570 133820 9593
rect 133980 9593 134003 10570
rect 136987 11570 137010 12577
rect 136987 10570 137170 11570
rect 136987 9593 137010 10570
rect 133980 9570 137010 9593
rect 1000 9410 2000 9570
rect 4190 9410 5190 9570
rect 7380 9410 8380 9570
rect 10570 9410 11570 9570
rect 13760 9410 14760 9570
rect 16950 9410 17950 9570
rect 20140 9410 21140 9570
rect 23330 9410 24330 9570
rect 26520 9410 27520 9570
rect 29710 9410 30710 9570
rect 32900 9410 33900 9570
rect 36090 9410 37090 9570
rect 39280 9410 40280 9570
rect 42470 9410 43470 9570
rect 45660 9410 46660 9570
rect 48850 9410 49850 9570
rect 52040 9410 53040 9570
rect 55230 9410 56230 9570
rect 58420 9410 59420 9570
rect 61610 9410 62610 9570
rect 64800 9410 65800 9570
rect 67990 9410 68990 9570
rect 71180 9410 72180 9570
rect 74370 9410 75370 9570
rect 77560 9410 78560 9570
rect 80750 9410 81750 9570
rect 83940 9410 84940 9570
rect 87130 9410 88130 9570
rect 90320 9410 91320 9570
rect 93510 9410 94510 9570
rect 96700 9410 97700 9570
rect 99890 9410 100890 9570
rect 103080 9410 104080 9570
rect 106270 9410 107270 9570
rect 109460 9410 110460 9570
rect 112650 9410 113650 9570
rect 115840 9410 116840 9570
rect 119030 9410 120030 9570
rect 122220 9410 123220 9570
rect 125410 9410 126410 9570
rect 128600 9410 129600 9570
rect 131790 9410 132790 9570
rect 134980 9410 135980 9570
rect 0 9387 3030 9410
rect 0 6403 23 9387
rect 3007 8380 3030 9387
rect 3190 9387 6220 9410
rect 3190 8380 3213 9387
rect 3007 7380 3213 8380
rect 3007 6403 3030 7380
rect 0 6380 3030 6403
rect 3190 6403 3213 7380
rect 6197 8380 6220 9387
rect 6380 9387 9410 9410
rect 6380 8380 6403 9387
rect 6197 7380 6403 8380
rect 6197 6403 6220 7380
rect 3190 6380 6220 6403
rect 6380 6403 6403 7380
rect 9387 8380 9410 9387
rect 9570 9387 12600 9410
rect 9570 8380 9593 9387
rect 9387 7380 9593 8380
rect 9387 6403 9410 7380
rect 6380 6380 9410 6403
rect 9570 6403 9593 7380
rect 12577 8380 12600 9387
rect 12760 9387 15790 9410
rect 12760 8380 12783 9387
rect 12577 7380 12783 8380
rect 12577 6403 12600 7380
rect 9570 6380 12600 6403
rect 12760 6403 12783 7380
rect 15767 8380 15790 9387
rect 15950 9387 18980 9410
rect 15950 8380 15973 9387
rect 15767 7380 15973 8380
rect 15767 6403 15790 7380
rect 12760 6380 15790 6403
rect 15950 6403 15973 7380
rect 18957 8380 18980 9387
rect 19140 9387 22170 9410
rect 19140 8380 19163 9387
rect 18957 7380 19163 8380
rect 18957 6403 18980 7380
rect 15950 6380 18980 6403
rect 19140 6403 19163 7380
rect 22147 8380 22170 9387
rect 22330 9387 25360 9410
rect 22330 8380 22353 9387
rect 22147 7380 22353 8380
rect 22147 6403 22170 7380
rect 19140 6380 22170 6403
rect 22330 6403 22353 7380
rect 25337 8380 25360 9387
rect 25520 9387 28550 9410
rect 25520 8380 25543 9387
rect 25337 7380 25543 8380
rect 25337 6403 25360 7380
rect 22330 6380 25360 6403
rect 25520 6403 25543 7380
rect 28527 8380 28550 9387
rect 28710 9387 31740 9410
rect 28710 8380 28733 9387
rect 28527 7380 28733 8380
rect 28527 6403 28550 7380
rect 25520 6380 28550 6403
rect 28710 6403 28733 7380
rect 31717 8380 31740 9387
rect 31900 9387 34930 9410
rect 31900 8380 31923 9387
rect 31717 7380 31923 8380
rect 31717 6403 31740 7380
rect 28710 6380 31740 6403
rect 31900 6403 31923 7380
rect 34907 8380 34930 9387
rect 35090 9387 38120 9410
rect 35090 8380 35113 9387
rect 34907 7380 35113 8380
rect 34907 6403 34930 7380
rect 31900 6380 34930 6403
rect 35090 6403 35113 7380
rect 38097 8380 38120 9387
rect 38280 9387 41310 9410
rect 38280 8380 38303 9387
rect 38097 7380 38303 8380
rect 38097 6403 38120 7380
rect 35090 6380 38120 6403
rect 38280 6403 38303 7380
rect 41287 8380 41310 9387
rect 41470 9387 44500 9410
rect 41470 8380 41493 9387
rect 41287 7380 41493 8380
rect 41287 6403 41310 7380
rect 38280 6380 41310 6403
rect 41470 6403 41493 7380
rect 44477 8380 44500 9387
rect 44660 9387 47690 9410
rect 44660 8380 44683 9387
rect 44477 7380 44683 8380
rect 44477 6403 44500 7380
rect 41470 6380 44500 6403
rect 44660 6403 44683 7380
rect 47667 8380 47690 9387
rect 47850 9387 50880 9410
rect 47850 8380 47873 9387
rect 47667 7380 47873 8380
rect 47667 6403 47690 7380
rect 44660 6380 47690 6403
rect 47850 6403 47873 7380
rect 50857 8380 50880 9387
rect 51040 9387 54070 9410
rect 51040 8380 51063 9387
rect 50857 7380 51063 8380
rect 50857 6403 50880 7380
rect 47850 6380 50880 6403
rect 51040 6403 51063 7380
rect 54047 8380 54070 9387
rect 54230 9387 57260 9410
rect 54230 8380 54253 9387
rect 54047 7380 54253 8380
rect 54047 6403 54070 7380
rect 51040 6380 54070 6403
rect 54230 6403 54253 7380
rect 57237 8380 57260 9387
rect 57420 9387 60450 9410
rect 57420 8380 57443 9387
rect 57237 7380 57443 8380
rect 57237 6403 57260 7380
rect 54230 6380 57260 6403
rect 57420 6403 57443 7380
rect 60427 8380 60450 9387
rect 60610 9387 63640 9410
rect 60610 8380 60633 9387
rect 60427 7380 60633 8380
rect 60427 6403 60450 7380
rect 57420 6380 60450 6403
rect 60610 6403 60633 7380
rect 63617 8380 63640 9387
rect 63800 9387 66830 9410
rect 63800 8380 63823 9387
rect 63617 7380 63823 8380
rect 63617 6403 63640 7380
rect 60610 6380 63640 6403
rect 63800 6403 63823 7380
rect 66807 8380 66830 9387
rect 66990 9387 70020 9410
rect 66990 8380 67013 9387
rect 66807 7380 67013 8380
rect 66807 6403 66830 7380
rect 63800 6380 66830 6403
rect 66990 6403 67013 7380
rect 69997 8380 70020 9387
rect 70180 9387 73210 9410
rect 70180 8380 70203 9387
rect 69997 7380 70203 8380
rect 69997 6403 70020 7380
rect 66990 6380 70020 6403
rect 70180 6403 70203 7380
rect 73187 8380 73210 9387
rect 73370 9387 76400 9410
rect 73370 8380 73393 9387
rect 73187 7380 73393 8380
rect 73187 6403 73210 7380
rect 70180 6380 73210 6403
rect 73370 6403 73393 7380
rect 76377 8380 76400 9387
rect 76560 9387 79590 9410
rect 76560 8380 76583 9387
rect 76377 7380 76583 8380
rect 76377 6403 76400 7380
rect 73370 6380 76400 6403
rect 76560 6403 76583 7380
rect 79567 8380 79590 9387
rect 79750 9387 82780 9410
rect 79750 8380 79773 9387
rect 79567 7380 79773 8380
rect 79567 6403 79590 7380
rect 76560 6380 79590 6403
rect 79750 6403 79773 7380
rect 82757 8380 82780 9387
rect 82940 9387 85970 9410
rect 82940 8380 82963 9387
rect 82757 7380 82963 8380
rect 82757 6403 82780 7380
rect 79750 6380 82780 6403
rect 82940 6403 82963 7380
rect 85947 8380 85970 9387
rect 86130 9387 89160 9410
rect 86130 8380 86153 9387
rect 85947 7380 86153 8380
rect 85947 6403 85970 7380
rect 82940 6380 85970 6403
rect 86130 6403 86153 7380
rect 89137 8380 89160 9387
rect 89320 9387 92350 9410
rect 89320 8380 89343 9387
rect 89137 7380 89343 8380
rect 89137 6403 89160 7380
rect 86130 6380 89160 6403
rect 89320 6403 89343 7380
rect 92327 8380 92350 9387
rect 92510 9387 95540 9410
rect 92510 8380 92533 9387
rect 92327 7380 92533 8380
rect 92327 6403 92350 7380
rect 89320 6380 92350 6403
rect 92510 6403 92533 7380
rect 95517 8380 95540 9387
rect 95700 9387 98730 9410
rect 95700 8380 95723 9387
rect 95517 7380 95723 8380
rect 95517 6403 95540 7380
rect 92510 6380 95540 6403
rect 95700 6403 95723 7380
rect 98707 8380 98730 9387
rect 98890 9387 101920 9410
rect 98890 8380 98913 9387
rect 98707 7380 98913 8380
rect 98707 6403 98730 7380
rect 95700 6380 98730 6403
rect 98890 6403 98913 7380
rect 101897 8380 101920 9387
rect 102080 9387 105110 9410
rect 102080 8380 102103 9387
rect 101897 7380 102103 8380
rect 101897 6403 101920 7380
rect 98890 6380 101920 6403
rect 102080 6403 102103 7380
rect 105087 8380 105110 9387
rect 105270 9387 108300 9410
rect 105270 8380 105293 9387
rect 105087 7380 105293 8380
rect 105087 6403 105110 7380
rect 102080 6380 105110 6403
rect 105270 6403 105293 7380
rect 108277 8380 108300 9387
rect 108460 9387 111490 9410
rect 108460 8380 108483 9387
rect 108277 7380 108483 8380
rect 108277 6403 108300 7380
rect 105270 6380 108300 6403
rect 108460 6403 108483 7380
rect 111467 8380 111490 9387
rect 111650 9387 114680 9410
rect 111650 8380 111673 9387
rect 111467 7380 111673 8380
rect 111467 6403 111490 7380
rect 108460 6380 111490 6403
rect 111650 6403 111673 7380
rect 114657 8380 114680 9387
rect 114840 9387 117870 9410
rect 114840 8380 114863 9387
rect 114657 7380 114863 8380
rect 114657 6403 114680 7380
rect 111650 6380 114680 6403
rect 114840 6403 114863 7380
rect 117847 8380 117870 9387
rect 118030 9387 121060 9410
rect 118030 8380 118053 9387
rect 117847 7380 118053 8380
rect 117847 6403 117870 7380
rect 114840 6380 117870 6403
rect 118030 6403 118053 7380
rect 121037 8380 121060 9387
rect 121220 9387 124250 9410
rect 121220 8380 121243 9387
rect 121037 7380 121243 8380
rect 121037 6403 121060 7380
rect 118030 6380 121060 6403
rect 121220 6403 121243 7380
rect 124227 8380 124250 9387
rect 124410 9387 127440 9410
rect 124410 8380 124433 9387
rect 124227 7380 124433 8380
rect 124227 6403 124250 7380
rect 121220 6380 124250 6403
rect 124410 6403 124433 7380
rect 127417 8380 127440 9387
rect 127600 9387 130630 9410
rect 127600 8380 127623 9387
rect 127417 7380 127623 8380
rect 127417 6403 127440 7380
rect 124410 6380 127440 6403
rect 127600 6403 127623 7380
rect 130607 8380 130630 9387
rect 130790 9387 133820 9410
rect 130790 8380 130813 9387
rect 130607 7380 130813 8380
rect 130607 6403 130630 7380
rect 127600 6380 130630 6403
rect 130790 6403 130813 7380
rect 133797 8380 133820 9387
rect 133980 9387 137010 9410
rect 133980 8380 134003 9387
rect 133797 7380 134003 8380
rect 133797 6403 133820 7380
rect 130790 6380 133820 6403
rect 133980 6403 134003 7380
rect 136987 8380 137010 9387
rect 136987 7380 137170 8380
rect 136987 6403 137010 7380
rect 133980 6380 137010 6403
rect 1000 6220 2000 6380
rect 4190 6220 5190 6380
rect 7380 6220 8380 6380
rect 10570 6220 11570 6380
rect 13760 6220 14760 6380
rect 16950 6220 17950 6380
rect 20140 6220 21140 6380
rect 23330 6220 24330 6380
rect 26520 6220 27520 6380
rect 29710 6220 30710 6380
rect 32900 6220 33900 6380
rect 36090 6220 37090 6380
rect 39280 6220 40280 6380
rect 42470 6220 43470 6380
rect 45660 6220 46660 6380
rect 48850 6220 49850 6380
rect 52040 6220 53040 6380
rect 55230 6220 56230 6380
rect 58420 6220 59420 6380
rect 61610 6220 62610 6380
rect 64800 6220 65800 6380
rect 67990 6220 68990 6380
rect 71180 6220 72180 6380
rect 74370 6220 75370 6380
rect 77560 6220 78560 6380
rect 80750 6220 81750 6380
rect 83940 6220 84940 6380
rect 87130 6220 88130 6380
rect 90320 6220 91320 6380
rect 93510 6220 94510 6380
rect 96700 6220 97700 6380
rect 99890 6220 100890 6380
rect 103080 6220 104080 6380
rect 106270 6220 107270 6380
rect 109460 6220 110460 6380
rect 112650 6220 113650 6380
rect 115840 6220 116840 6380
rect 119030 6220 120030 6380
rect 122220 6220 123220 6380
rect 125410 6220 126410 6380
rect 128600 6220 129600 6380
rect 131790 6220 132790 6380
rect 134980 6220 135980 6380
rect 0 6197 3030 6220
rect 0 3213 23 6197
rect 3007 5190 3030 6197
rect 3190 6197 6220 6220
rect 3190 5190 3213 6197
rect 3007 4190 3213 5190
rect 3007 3213 3030 4190
rect 0 3190 3030 3213
rect 3190 3213 3213 4190
rect 6197 5190 6220 6197
rect 6380 6197 9410 6220
rect 6380 5190 6403 6197
rect 6197 4190 6403 5190
rect 6197 3213 6220 4190
rect 3190 3190 6220 3213
rect 6380 3213 6403 4190
rect 9387 5190 9410 6197
rect 9570 6197 12600 6220
rect 9570 5190 9593 6197
rect 9387 4190 9593 5190
rect 9387 3213 9410 4190
rect 6380 3190 9410 3213
rect 9570 3213 9593 4190
rect 12577 5190 12600 6197
rect 12760 6197 15790 6220
rect 12760 5190 12783 6197
rect 12577 4190 12783 5190
rect 12577 3213 12600 4190
rect 9570 3190 12600 3213
rect 12760 3213 12783 4190
rect 15767 5190 15790 6197
rect 15950 6197 18980 6220
rect 15950 5190 15973 6197
rect 15767 4190 15973 5190
rect 15767 3213 15790 4190
rect 12760 3190 15790 3213
rect 15950 3213 15973 4190
rect 18957 5190 18980 6197
rect 19140 6197 22170 6220
rect 19140 5190 19163 6197
rect 18957 4190 19163 5190
rect 18957 3213 18980 4190
rect 15950 3190 18980 3213
rect 19140 3213 19163 4190
rect 22147 5190 22170 6197
rect 22330 6197 25360 6220
rect 22330 5190 22353 6197
rect 22147 4190 22353 5190
rect 22147 3213 22170 4190
rect 19140 3190 22170 3213
rect 22330 3213 22353 4190
rect 25337 5190 25360 6197
rect 25520 6197 28550 6220
rect 25520 5190 25543 6197
rect 25337 4190 25543 5190
rect 25337 3213 25360 4190
rect 22330 3190 25360 3213
rect 25520 3213 25543 4190
rect 28527 5190 28550 6197
rect 28710 6197 31740 6220
rect 28710 5190 28733 6197
rect 28527 4190 28733 5190
rect 28527 3213 28550 4190
rect 25520 3190 28550 3213
rect 28710 3213 28733 4190
rect 31717 5190 31740 6197
rect 31900 6197 34930 6220
rect 31900 5190 31923 6197
rect 31717 4190 31923 5190
rect 31717 3213 31740 4190
rect 28710 3190 31740 3213
rect 31900 3213 31923 4190
rect 34907 5190 34930 6197
rect 35090 6197 38120 6220
rect 35090 5190 35113 6197
rect 34907 4190 35113 5190
rect 34907 3213 34930 4190
rect 31900 3190 34930 3213
rect 35090 3213 35113 4190
rect 38097 5190 38120 6197
rect 38280 6197 41310 6220
rect 38280 5190 38303 6197
rect 38097 4190 38303 5190
rect 38097 3213 38120 4190
rect 35090 3190 38120 3213
rect 38280 3213 38303 4190
rect 41287 5190 41310 6197
rect 41470 6197 44500 6220
rect 41470 5190 41493 6197
rect 41287 4190 41493 5190
rect 41287 3213 41310 4190
rect 38280 3190 41310 3213
rect 41470 3213 41493 4190
rect 44477 5190 44500 6197
rect 44660 6197 47690 6220
rect 44660 5190 44683 6197
rect 44477 4190 44683 5190
rect 44477 3213 44500 4190
rect 41470 3190 44500 3213
rect 44660 3213 44683 4190
rect 47667 5190 47690 6197
rect 47850 6197 50880 6220
rect 47850 5190 47873 6197
rect 47667 4190 47873 5190
rect 47667 3213 47690 4190
rect 44660 3190 47690 3213
rect 47850 3213 47873 4190
rect 50857 5190 50880 6197
rect 51040 6197 54070 6220
rect 51040 5190 51063 6197
rect 50857 4190 51063 5190
rect 50857 3213 50880 4190
rect 47850 3190 50880 3213
rect 51040 3213 51063 4190
rect 54047 5190 54070 6197
rect 54230 6197 57260 6220
rect 54230 5190 54253 6197
rect 54047 4190 54253 5190
rect 54047 3213 54070 4190
rect 51040 3190 54070 3213
rect 54230 3213 54253 4190
rect 57237 5190 57260 6197
rect 57420 6197 60450 6220
rect 57420 5190 57443 6197
rect 57237 4190 57443 5190
rect 57237 3213 57260 4190
rect 54230 3190 57260 3213
rect 57420 3213 57443 4190
rect 60427 5190 60450 6197
rect 60610 6197 63640 6220
rect 60610 5190 60633 6197
rect 60427 4190 60633 5190
rect 60427 3213 60450 4190
rect 57420 3190 60450 3213
rect 60610 3213 60633 4190
rect 63617 5190 63640 6197
rect 63800 6197 66830 6220
rect 63800 5190 63823 6197
rect 63617 4190 63823 5190
rect 63617 3213 63640 4190
rect 60610 3190 63640 3213
rect 63800 3213 63823 4190
rect 66807 5190 66830 6197
rect 66990 6197 70020 6220
rect 66990 5190 67013 6197
rect 66807 4190 67013 5190
rect 66807 3213 66830 4190
rect 63800 3190 66830 3213
rect 66990 3213 67013 4190
rect 69997 5190 70020 6197
rect 70180 6197 73210 6220
rect 70180 5190 70203 6197
rect 69997 4190 70203 5190
rect 69997 3213 70020 4190
rect 66990 3190 70020 3213
rect 70180 3213 70203 4190
rect 73187 5190 73210 6197
rect 73370 6197 76400 6220
rect 73370 5190 73393 6197
rect 73187 4190 73393 5190
rect 73187 3213 73210 4190
rect 70180 3190 73210 3213
rect 73370 3213 73393 4190
rect 76377 5190 76400 6197
rect 76560 6197 79590 6220
rect 76560 5190 76583 6197
rect 76377 4190 76583 5190
rect 76377 3213 76400 4190
rect 73370 3190 76400 3213
rect 76560 3213 76583 4190
rect 79567 5190 79590 6197
rect 79750 6197 82780 6220
rect 79750 5190 79773 6197
rect 79567 4190 79773 5190
rect 79567 3213 79590 4190
rect 76560 3190 79590 3213
rect 79750 3213 79773 4190
rect 82757 5190 82780 6197
rect 82940 6197 85970 6220
rect 82940 5190 82963 6197
rect 82757 4190 82963 5190
rect 82757 3213 82780 4190
rect 79750 3190 82780 3213
rect 82940 3213 82963 4190
rect 85947 5190 85970 6197
rect 86130 6197 89160 6220
rect 86130 5190 86153 6197
rect 85947 4190 86153 5190
rect 85947 3213 85970 4190
rect 82940 3190 85970 3213
rect 86130 3213 86153 4190
rect 89137 5190 89160 6197
rect 89320 6197 92350 6220
rect 89320 5190 89343 6197
rect 89137 4190 89343 5190
rect 89137 3213 89160 4190
rect 86130 3190 89160 3213
rect 89320 3213 89343 4190
rect 92327 5190 92350 6197
rect 92510 6197 95540 6220
rect 92510 5190 92533 6197
rect 92327 4190 92533 5190
rect 92327 3213 92350 4190
rect 89320 3190 92350 3213
rect 92510 3213 92533 4190
rect 95517 5190 95540 6197
rect 95700 6197 98730 6220
rect 95700 5190 95723 6197
rect 95517 4190 95723 5190
rect 95517 3213 95540 4190
rect 92510 3190 95540 3213
rect 95700 3213 95723 4190
rect 98707 5190 98730 6197
rect 98890 6197 101920 6220
rect 98890 5190 98913 6197
rect 98707 4190 98913 5190
rect 98707 3213 98730 4190
rect 95700 3190 98730 3213
rect 98890 3213 98913 4190
rect 101897 5190 101920 6197
rect 102080 6197 105110 6220
rect 102080 5190 102103 6197
rect 101897 4190 102103 5190
rect 101897 3213 101920 4190
rect 98890 3190 101920 3213
rect 102080 3213 102103 4190
rect 105087 5190 105110 6197
rect 105270 6197 108300 6220
rect 105270 5190 105293 6197
rect 105087 4190 105293 5190
rect 105087 3213 105110 4190
rect 102080 3190 105110 3213
rect 105270 3213 105293 4190
rect 108277 5190 108300 6197
rect 108460 6197 111490 6220
rect 108460 5190 108483 6197
rect 108277 4190 108483 5190
rect 108277 3213 108300 4190
rect 105270 3190 108300 3213
rect 108460 3213 108483 4190
rect 111467 5190 111490 6197
rect 111650 6197 114680 6220
rect 111650 5190 111673 6197
rect 111467 4190 111673 5190
rect 111467 3213 111490 4190
rect 108460 3190 111490 3213
rect 111650 3213 111673 4190
rect 114657 5190 114680 6197
rect 114840 6197 117870 6220
rect 114840 5190 114863 6197
rect 114657 4190 114863 5190
rect 114657 3213 114680 4190
rect 111650 3190 114680 3213
rect 114840 3213 114863 4190
rect 117847 5190 117870 6197
rect 118030 6197 121060 6220
rect 118030 5190 118053 6197
rect 117847 4190 118053 5190
rect 117847 3213 117870 4190
rect 114840 3190 117870 3213
rect 118030 3213 118053 4190
rect 121037 5190 121060 6197
rect 121220 6197 124250 6220
rect 121220 5190 121243 6197
rect 121037 4190 121243 5190
rect 121037 3213 121060 4190
rect 118030 3190 121060 3213
rect 121220 3213 121243 4190
rect 124227 5190 124250 6197
rect 124410 6197 127440 6220
rect 124410 5190 124433 6197
rect 124227 4190 124433 5190
rect 124227 3213 124250 4190
rect 121220 3190 124250 3213
rect 124410 3213 124433 4190
rect 127417 5190 127440 6197
rect 127600 6197 130630 6220
rect 127600 5190 127623 6197
rect 127417 4190 127623 5190
rect 127417 3213 127440 4190
rect 124410 3190 127440 3213
rect 127600 3213 127623 4190
rect 130607 5190 130630 6197
rect 130790 6197 133820 6220
rect 130790 5190 130813 6197
rect 130607 4190 130813 5190
rect 130607 3213 130630 4190
rect 127600 3190 130630 3213
rect 130790 3213 130813 4190
rect 133797 5190 133820 6197
rect 133980 6197 137010 6220
rect 133980 5190 134003 6197
rect 133797 4190 134003 5190
rect 133797 3213 133820 4190
rect 130790 3190 133820 3213
rect 133980 3213 134003 4190
rect 136987 5190 137010 6197
rect 136987 4190 137170 5190
rect 136987 3213 137010 4190
rect 133980 3190 137010 3213
rect 1000 3030 2000 3190
rect 4190 3030 5190 3190
rect 7380 3030 8380 3190
rect 10570 3030 11570 3190
rect 13760 3030 14760 3190
rect 16950 3030 17950 3190
rect 20140 3030 21140 3190
rect 23330 3030 24330 3190
rect 26520 3030 27520 3190
rect 29710 3030 30710 3190
rect 32900 3030 33900 3190
rect 36090 3030 37090 3190
rect 39280 3030 40280 3190
rect 42470 3030 43470 3190
rect 45660 3030 46660 3190
rect 48850 3030 49850 3190
rect 52040 3030 53040 3190
rect 55230 3030 56230 3190
rect 58420 3030 59420 3190
rect 61610 3030 62610 3190
rect 64800 3030 65800 3190
rect 67990 3030 68990 3190
rect 71180 3030 72180 3190
rect 74370 3030 75370 3190
rect 77560 3030 78560 3190
rect 80750 3030 81750 3190
rect 83940 3030 84940 3190
rect 87130 3030 88130 3190
rect 90320 3030 91320 3190
rect 93510 3030 94510 3190
rect 96700 3030 97700 3190
rect 99890 3030 100890 3190
rect 103080 3030 104080 3190
rect 106270 3030 107270 3190
rect 109460 3030 110460 3190
rect 112650 3030 113650 3190
rect 115840 3030 116840 3190
rect 119030 3030 120030 3190
rect 122220 3030 123220 3190
rect 125410 3030 126410 3190
rect 128600 3030 129600 3190
rect 131790 3030 132790 3190
rect 134980 3030 135980 3190
rect 0 3007 3030 3030
rect 0 23 23 3007
rect 3007 2000 3030 3007
rect 3190 3007 6220 3030
rect 3190 2000 3213 3007
rect 3007 1000 3213 2000
rect 3007 23 3030 1000
rect 0 0 3030 23
rect 3190 23 3213 1000
rect 6197 2000 6220 3007
rect 6380 3007 9410 3030
rect 6380 2000 6403 3007
rect 6197 1000 6403 2000
rect 6197 23 6220 1000
rect 3190 0 6220 23
rect 6380 23 6403 1000
rect 9387 2000 9410 3007
rect 9570 3007 12600 3030
rect 9570 2000 9593 3007
rect 9387 1000 9593 2000
rect 9387 23 9410 1000
rect 6380 0 9410 23
rect 9570 23 9593 1000
rect 12577 2000 12600 3007
rect 12760 3007 15790 3030
rect 12760 2000 12783 3007
rect 12577 1000 12783 2000
rect 12577 23 12600 1000
rect 9570 0 12600 23
rect 12760 23 12783 1000
rect 15767 2000 15790 3007
rect 15950 3007 18980 3030
rect 15950 2000 15973 3007
rect 15767 1000 15973 2000
rect 15767 23 15790 1000
rect 12760 0 15790 23
rect 15950 23 15973 1000
rect 18957 2000 18980 3007
rect 19140 3007 22170 3030
rect 19140 2000 19163 3007
rect 18957 1000 19163 2000
rect 18957 23 18980 1000
rect 15950 0 18980 23
rect 19140 23 19163 1000
rect 22147 2000 22170 3007
rect 22330 3007 25360 3030
rect 22330 2000 22353 3007
rect 22147 1000 22353 2000
rect 22147 23 22170 1000
rect 19140 0 22170 23
rect 22330 23 22353 1000
rect 25337 2000 25360 3007
rect 25520 3007 28550 3030
rect 25520 2000 25543 3007
rect 25337 1000 25543 2000
rect 25337 23 25360 1000
rect 22330 0 25360 23
rect 25520 23 25543 1000
rect 28527 2000 28550 3007
rect 28710 3007 31740 3030
rect 28710 2000 28733 3007
rect 28527 1000 28733 2000
rect 28527 23 28550 1000
rect 25520 0 28550 23
rect 28710 23 28733 1000
rect 31717 2000 31740 3007
rect 31900 3007 34930 3030
rect 31900 2000 31923 3007
rect 31717 1000 31923 2000
rect 31717 23 31740 1000
rect 28710 0 31740 23
rect 31900 23 31923 1000
rect 34907 2000 34930 3007
rect 35090 3007 38120 3030
rect 35090 2000 35113 3007
rect 34907 1000 35113 2000
rect 34907 23 34930 1000
rect 31900 0 34930 23
rect 35090 23 35113 1000
rect 38097 2000 38120 3007
rect 38280 3007 41310 3030
rect 38280 2000 38303 3007
rect 38097 1000 38303 2000
rect 38097 23 38120 1000
rect 35090 0 38120 23
rect 38280 23 38303 1000
rect 41287 2000 41310 3007
rect 41470 3007 44500 3030
rect 41470 2000 41493 3007
rect 41287 1000 41493 2000
rect 41287 23 41310 1000
rect 38280 0 41310 23
rect 41470 23 41493 1000
rect 44477 2000 44500 3007
rect 44660 3007 47690 3030
rect 44660 2000 44683 3007
rect 44477 1000 44683 2000
rect 44477 23 44500 1000
rect 41470 0 44500 23
rect 44660 23 44683 1000
rect 47667 2000 47690 3007
rect 47850 3007 50880 3030
rect 47850 2000 47873 3007
rect 47667 1000 47873 2000
rect 47667 23 47690 1000
rect 44660 0 47690 23
rect 47850 23 47873 1000
rect 50857 2000 50880 3007
rect 51040 3007 54070 3030
rect 51040 2000 51063 3007
rect 50857 1000 51063 2000
rect 50857 23 50880 1000
rect 47850 0 50880 23
rect 51040 23 51063 1000
rect 54047 2000 54070 3007
rect 54230 3007 57260 3030
rect 54230 2000 54253 3007
rect 54047 1000 54253 2000
rect 54047 23 54070 1000
rect 51040 0 54070 23
rect 54230 23 54253 1000
rect 57237 2000 57260 3007
rect 57420 3007 60450 3030
rect 57420 2000 57443 3007
rect 57237 1000 57443 2000
rect 57237 23 57260 1000
rect 54230 0 57260 23
rect 57420 23 57443 1000
rect 60427 2000 60450 3007
rect 60610 3007 63640 3030
rect 60610 2000 60633 3007
rect 60427 1000 60633 2000
rect 60427 23 60450 1000
rect 57420 0 60450 23
rect 60610 23 60633 1000
rect 63617 2000 63640 3007
rect 63800 3007 66830 3030
rect 63800 2000 63823 3007
rect 63617 1000 63823 2000
rect 63617 23 63640 1000
rect 60610 0 63640 23
rect 63800 23 63823 1000
rect 66807 2000 66830 3007
rect 66990 3007 70020 3030
rect 66990 2000 67013 3007
rect 66807 1000 67013 2000
rect 66807 23 66830 1000
rect 63800 0 66830 23
rect 66990 23 67013 1000
rect 69997 2000 70020 3007
rect 70180 3007 73210 3030
rect 70180 2000 70203 3007
rect 69997 1000 70203 2000
rect 69997 23 70020 1000
rect 66990 0 70020 23
rect 70180 23 70203 1000
rect 73187 2000 73210 3007
rect 73370 3007 76400 3030
rect 73370 2000 73393 3007
rect 73187 1000 73393 2000
rect 73187 23 73210 1000
rect 70180 0 73210 23
rect 73370 23 73393 1000
rect 76377 2000 76400 3007
rect 76560 3007 79590 3030
rect 76560 2000 76583 3007
rect 76377 1000 76583 2000
rect 76377 23 76400 1000
rect 73370 0 76400 23
rect 76560 23 76583 1000
rect 79567 2000 79590 3007
rect 79750 3007 82780 3030
rect 79750 2000 79773 3007
rect 79567 1000 79773 2000
rect 79567 23 79590 1000
rect 76560 0 79590 23
rect 79750 23 79773 1000
rect 82757 2000 82780 3007
rect 82940 3007 85970 3030
rect 82940 2000 82963 3007
rect 82757 1000 82963 2000
rect 82757 23 82780 1000
rect 79750 0 82780 23
rect 82940 23 82963 1000
rect 85947 2000 85970 3007
rect 86130 3007 89160 3030
rect 86130 2000 86153 3007
rect 85947 1000 86153 2000
rect 85947 23 85970 1000
rect 82940 0 85970 23
rect 86130 23 86153 1000
rect 89137 2000 89160 3007
rect 89320 3007 92350 3030
rect 89320 2000 89343 3007
rect 89137 1000 89343 2000
rect 89137 23 89160 1000
rect 86130 0 89160 23
rect 89320 23 89343 1000
rect 92327 2000 92350 3007
rect 92510 3007 95540 3030
rect 92510 2000 92533 3007
rect 92327 1000 92533 2000
rect 92327 23 92350 1000
rect 89320 0 92350 23
rect 92510 23 92533 1000
rect 95517 2000 95540 3007
rect 95700 3007 98730 3030
rect 95700 2000 95723 3007
rect 95517 1000 95723 2000
rect 95517 23 95540 1000
rect 92510 0 95540 23
rect 95700 23 95723 1000
rect 98707 2000 98730 3007
rect 98890 3007 101920 3030
rect 98890 2000 98913 3007
rect 98707 1000 98913 2000
rect 98707 23 98730 1000
rect 95700 0 98730 23
rect 98890 23 98913 1000
rect 101897 2000 101920 3007
rect 102080 3007 105110 3030
rect 102080 2000 102103 3007
rect 101897 1000 102103 2000
rect 101897 23 101920 1000
rect 98890 0 101920 23
rect 102080 23 102103 1000
rect 105087 2000 105110 3007
rect 105270 3007 108300 3030
rect 105270 2000 105293 3007
rect 105087 1000 105293 2000
rect 105087 23 105110 1000
rect 102080 0 105110 23
rect 105270 23 105293 1000
rect 108277 2000 108300 3007
rect 108460 3007 111490 3030
rect 108460 2000 108483 3007
rect 108277 1000 108483 2000
rect 108277 23 108300 1000
rect 105270 0 108300 23
rect 108460 23 108483 1000
rect 111467 2000 111490 3007
rect 111650 3007 114680 3030
rect 111650 2000 111673 3007
rect 111467 1000 111673 2000
rect 111467 23 111490 1000
rect 108460 0 111490 23
rect 111650 23 111673 1000
rect 114657 2000 114680 3007
rect 114840 3007 117870 3030
rect 114840 2000 114863 3007
rect 114657 1000 114863 2000
rect 114657 23 114680 1000
rect 111650 0 114680 23
rect 114840 23 114863 1000
rect 117847 2000 117870 3007
rect 118030 3007 121060 3030
rect 118030 2000 118053 3007
rect 117847 1000 118053 2000
rect 117847 23 117870 1000
rect 114840 0 117870 23
rect 118030 23 118053 1000
rect 121037 2000 121060 3007
rect 121220 3007 124250 3030
rect 121220 2000 121243 3007
rect 121037 1000 121243 2000
rect 121037 23 121060 1000
rect 118030 0 121060 23
rect 121220 23 121243 1000
rect 124227 2000 124250 3007
rect 124410 3007 127440 3030
rect 124410 2000 124433 3007
rect 124227 1000 124433 2000
rect 124227 23 124250 1000
rect 121220 0 124250 23
rect 124410 23 124433 1000
rect 127417 2000 127440 3007
rect 127600 3007 130630 3030
rect 127600 2000 127623 3007
rect 127417 1000 127623 2000
rect 127417 23 127440 1000
rect 124410 0 127440 23
rect 127600 23 127623 1000
rect 130607 2000 130630 3007
rect 130790 3007 133820 3030
rect 130790 2000 130813 3007
rect 130607 1000 130813 2000
rect 130607 23 130630 1000
rect 127600 0 130630 23
rect 130790 23 130813 1000
rect 133797 2000 133820 3007
rect 133980 3007 137010 3030
rect 133980 2000 134003 3007
rect 133797 1000 134003 2000
rect 133797 23 133820 1000
rect 130790 0 133820 23
rect 133980 23 134003 1000
rect 136987 2000 137010 3007
rect 136987 1000 137170 2000
rect 136987 23 137010 1000
rect 133980 0 137010 23
<< end >>
