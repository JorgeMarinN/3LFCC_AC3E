magic
tech sky130A
timestamp 1666620395
<< checkpaint >>
rect -134766 223166 -49634 226366
rect -137966 216966 -49634 223166
rect -27666 220166 27666 226366
rect -27666 216966 137966 220166
rect -137966 216234 137966 216966
rect -137966 213034 -124634 216234
rect -137966 209966 -127834 213034
rect -59766 210566 137966 216234
rect -94966 210034 137966 210566
rect -94966 209966 94966 210034
rect 127834 209966 137966 210034
rect -139966 -1966 139966 209966
<< metal1 >>
rect -25700 224385 -300 224400
rect -25700 221415 -25685 224385
rect -315 221415 -300 224385
rect -25700 221400 -300 221415
rect -25700 221200 -22700 221400
rect -22500 221200 -19500 221400
rect -19300 221200 -16300 221400
rect -16100 221200 -13100 221400
rect -12900 221200 -9900 221400
rect -9700 221200 -6700 221400
rect -6500 221200 -3500 221400
rect -3300 221200 -300 221400
rect -25700 221185 -300 221200
rect -25700 218215 -25685 221185
rect -315 218215 -300 221185
rect -25700 218200 -300 218215
rect -25700 202200 -22700 218200
rect -22500 202200 -19500 218200
rect -19300 202200 -16300 218200
rect -16100 202200 -13100 218200
rect -12900 202200 -9900 218200
rect -9700 202200 -6700 218200
rect -6500 202200 -3500 218200
rect -3300 202200 -300 218200
rect 300 224385 25700 224400
rect 300 221415 315 224385
rect 25685 221415 25700 224385
rect 300 221400 25700 221415
rect 300 221200 3300 221400
rect 3500 221200 6500 221400
rect 6700 221200 9700 221400
rect 9900 221200 12900 221400
rect 13100 221200 16100 221400
rect 16300 221200 19300 221400
rect 19500 221200 22500 221400
rect 22700 221200 25700 221400
rect 300 221185 25700 221200
rect 300 218215 315 221185
rect 25685 218215 25700 221185
rect 300 218200 25700 218215
rect 300 208600 3300 218200
rect 3500 208600 6500 218200
rect 6700 208600 9700 218200
rect 9900 208600 12900 218200
rect 13100 208600 16100 218200
rect 16300 208600 19300 218200
rect 19500 208600 22500 218200
rect 22700 208600 25700 218200
rect 300 208585 25700 208600
rect 300 205615 315 208585
rect 25685 205615 25700 208585
rect 300 205600 25700 205615
rect 300 205400 3300 205600
rect 3500 205400 6500 205600
rect 6700 205400 9700 205600
rect 9900 205400 12900 205600
rect 13100 205400 16100 205600
rect 16300 205400 19300 205600
rect 19500 205400 22500 205600
rect 22700 205400 25700 205600
rect 300 205385 25700 205400
rect 300 202415 315 205385
rect 25685 202415 25700 205385
rect 300 202400 25700 202415
rect -26000 202185 0 202200
rect -26000 201215 -25985 202185
rect -15 201215 0 202185
rect -26000 201200 0 201215
rect -129000 168995 -70000 169000
rect -129000 168005 -128995 168995
rect -70005 168005 -70000 168995
rect -129000 168000 -70000 168005
rect -55000 168995 -9000 169000
rect -55000 168015 -54995 168995
rect -9015 168015 -9000 168995
rect -55000 168000 -9000 168015
rect 9000 168995 55000 169000
rect 9000 168005 9005 168995
rect 54995 168005 55000 168995
rect 9000 168000 55000 168005
rect 70000 168995 129000 169000
rect 70000 168005 70005 168995
rect 128995 168005 129000 168995
rect 70000 168000 129000 168005
rect -2000 166950 2000 167150
rect -138000 166295 138000 166300
rect -138000 165305 -137995 166295
rect 137995 165305 138000 166295
rect -138000 165300 138000 165305
<< via1 >>
rect -25685 221415 -315 224385
rect -25685 218215 -315 221185
rect 315 221415 25685 224385
rect 315 218215 25685 221185
rect 315 205615 25685 208585
rect 315 202415 25685 205385
rect -25985 201215 -15 202185
rect -128995 168005 -70005 168995
rect -54995 168015 -9015 168995
rect 9005 168005 54995 168995
rect 70005 168005 128995 168995
rect -137995 165305 137995 166295
<< metal2 >>
rect -25700 224385 -300 224400
rect -25700 221415 -25685 224385
rect -315 221415 -300 224385
rect -25700 221400 -300 221415
rect -25700 221200 -22700 221400
rect -22500 221200 -19500 221400
rect -19300 221200 -16300 221400
rect -16100 221200 -13100 221400
rect -12900 221200 -9900 221400
rect -9700 221200 -6700 221400
rect -6500 221200 -3500 221400
rect -3300 221200 -300 221400
rect -25700 221185 -300 221200
rect -25700 218215 -25685 221185
rect -315 218215 -300 221185
rect -25700 218200 -300 218215
rect -32500 214985 -30500 215000
rect -32500 212015 -32485 214985
rect -30505 212015 -30500 214985
rect -32500 211785 -30500 212015
rect -32500 208815 -32485 211785
rect -30505 208815 -30500 211785
rect -32500 197000 -30500 208815
rect -25700 202200 -22700 218200
rect -22500 202200 -19500 218200
rect -19300 202200 -16300 218200
rect -16100 202200 -13100 218200
rect -12900 202200 -9900 218200
rect -9700 202200 -6700 218200
rect -6500 202200 -3500 218200
rect -3300 202200 -300 218200
rect 300 224385 25700 224400
rect 300 221415 315 224385
rect 25685 221415 25700 224385
rect 300 221400 25700 221415
rect 300 221200 3300 221400
rect 3500 221200 6500 221400
rect 6700 221200 9700 221400
rect 9900 221200 12900 221400
rect 13100 221200 16100 221400
rect 16300 221200 19300 221400
rect 19500 221200 22500 221400
rect 22700 221200 25700 221400
rect 300 221185 25700 221200
rect 300 218215 315 221185
rect 25685 218215 25700 221185
rect 300 218200 25700 218215
rect 300 208600 3300 218200
rect 3500 208600 6500 218200
rect 6700 208600 9700 218200
rect 9900 208600 12900 218200
rect 13100 208600 16100 218200
rect 16300 208600 19300 218200
rect 19500 208600 22500 218200
rect 22700 208600 25700 218200
rect 300 208585 25700 208600
rect 300 205615 315 208585
rect 25685 205615 25700 208585
rect 300 205600 25700 205615
rect 300 205400 3300 205600
rect 3500 205400 6500 205600
rect 6700 205400 9700 205600
rect 9900 205400 12900 205600
rect 13100 205400 16100 205600
rect 16300 205400 19300 205600
rect 19500 205400 22500 205600
rect 22700 205400 25700 205600
rect 300 205385 25700 205400
rect 300 202415 315 205385
rect 25685 202415 25700 205385
rect 300 202400 25700 202415
rect 30200 214985 32200 215000
rect 30200 212015 30215 214985
rect 32185 212015 32200 214985
rect 30200 211785 32200 212015
rect 30200 208815 30215 211785
rect 32185 208815 32200 211785
rect -26000 202185 0 202200
rect -26000 201215 -25985 202185
rect -15 201215 0 202185
rect -26000 201200 0 201215
rect 30200 197000 32200 208815
rect -129000 168995 -70000 173000
rect -2000 171995 2000 172000
rect -2000 171005 -1995 171995
rect 1995 171005 2000 171995
rect -129000 168005 -128995 168995
rect -70005 168005 -70000 168995
rect -129000 166300 -70000 168005
rect -55000 168995 -9000 170000
rect -55000 168015 -54995 168995
rect -9015 168015 -9000 168995
rect -55000 166300 -9000 168015
rect -2000 166300 2000 171005
rect 9000 168995 55000 170000
rect 9000 168005 9005 168995
rect 54995 168005 55000 168995
rect 9000 166300 55000 168005
rect 70000 168995 129000 173000
rect 70000 168005 70005 168995
rect 128995 168005 129000 168995
rect 70000 166300 129000 168005
rect -138000 166295 138000 166300
rect -138000 165305 -137995 166295
rect 137995 165305 138000 166295
rect -138000 165300 138000 165305
<< via2 >>
rect -25685 221415 -315 224385
rect -25685 218215 -315 221185
rect -32485 212015 -30505 214985
rect -32485 208815 -30505 211785
rect 315 221415 25685 224385
rect 315 218215 25685 221185
rect 315 205615 25685 208585
rect 315 202415 25685 205385
rect 30215 212015 32185 214985
rect 30215 208815 32185 211785
rect -25985 201215 -15 202185
rect -1995 171005 1995 171995
<< metal3 >>
rect -132800 221400 -51600 224400
rect -25700 224385 -300 224400
rect -25700 221415 -25685 224385
rect -315 221415 -300 224385
rect -25700 221400 -300 221415
rect 300 224385 25700 224400
rect 300 221415 315 224385
rect 25685 221415 25700 224385
rect 300 221400 25700 221415
rect -132800 221200 -129800 221400
rect -129600 221200 -126600 221400
rect -57800 221200 -54800 221400
rect -54600 221200 -51600 221400
rect -136000 218200 -51600 221200
rect -25700 221185 -300 221200
rect -25700 218215 -25685 221185
rect -315 218215 -300 221185
rect -25700 218200 -300 218215
rect 300 221185 25700 221200
rect 300 218215 315 221185
rect 25685 218215 25700 221185
rect 300 218200 25700 218215
rect -136000 218000 -133000 218200
rect -132800 218000 -129800 218200
rect -129600 218000 -126600 218200
rect -136000 215000 -126600 218000
rect -57800 215000 -54800 218200
rect -54600 215000 -51600 218200
rect 26000 215200 136000 218200
rect 26000 215000 29000 215200
rect 29200 215000 32200 215200
rect 129800 215000 132800 215200
rect 133000 215000 136000 215200
rect -136000 206000 -133000 215000
rect -132800 206000 -129800 215000
rect -57800 214985 136000 215000
rect -57800 212015 -32485 214985
rect -30505 212015 30215 214985
rect 32185 212015 136000 214985
rect -57800 212000 136000 212015
rect -57800 211800 -54800 212000
rect -54600 211800 -51600 212000
rect 26000 211800 29000 212000
rect 29200 211800 32200 212000
rect -57800 211785 32200 211800
rect -57800 208815 -32485 211785
rect -30505 208815 30215 211785
rect 32185 208815 32200 211785
rect -57800 208800 32200 208815
rect -93000 208585 93000 208600
rect -93000 205615 315 208585
rect 25685 205615 93000 208585
rect 129800 206000 132800 212000
rect 133000 206000 136000 212000
rect -93000 205600 93000 205615
rect -61000 205400 -58000 205600
rect -57800 205400 -54800 205600
rect 54800 205400 57800 205600
rect 58000 205400 61000 205600
rect -65000 205385 65000 205400
rect -65000 202415 315 205385
rect 25685 202415 65000 205385
rect -65000 202400 65000 202415
rect -61000 200000 -58000 202400
rect -57800 200000 -54800 202400
rect -26000 202185 3000 202200
rect -26000 201215 -25985 202185
rect -15 201215 3000 202185
rect -26000 200000 3000 201215
rect 54800 200000 57800 202400
rect 58000 200000 61000 202400
rect -4000 177000 4000 200000
rect -2000 171995 2000 177000
rect -2000 171005 -1995 171995
rect 1995 171005 2000 171995
rect -2000 171000 2000 171005
<< via3 >>
rect -25685 221415 -315 224385
rect 315 221415 25685 224385
rect -25685 218215 -315 221185
rect 315 218215 25685 221185
rect -32485 212015 -30505 214985
rect 30215 212015 32185 214985
rect -32485 208815 -30505 211785
rect 30215 208815 32185 211785
rect 315 205615 25685 208585
rect 315 202415 25685 205385
rect -25985 201215 -15 202185
<< metal4 >>
rect -132800 221400 -51600 224400
rect -25700 224385 -300 224400
rect -25700 221415 -25685 224385
rect -315 221415 -300 224385
rect -25700 221400 -300 221415
rect 300 224385 25700 224400
rect 300 221415 315 224385
rect 25685 221415 25700 224385
rect 300 221400 25700 221415
rect -132800 221200 -129800 221400
rect -129600 221200 -126600 221400
rect -57800 221200 -54800 221400
rect -54600 221200 -51600 221400
rect -136000 218200 -51600 221200
rect -25700 221185 -300 221200
rect -25700 218215 -25685 221185
rect -315 218215 -300 221185
rect -25700 218200 -300 218215
rect 300 221185 25700 221200
rect 300 218215 315 221185
rect 25685 218215 25700 221185
rect 300 218200 25700 218215
rect -136000 218000 -133000 218200
rect -132800 218000 -129800 218200
rect -129600 218000 -126600 218200
rect -136000 215000 -126600 218000
rect -57800 215000 -54800 218200
rect -54600 215000 -51600 218200
rect 26000 215200 136000 218200
rect 26000 215000 29000 215200
rect 29200 215000 32200 215200
rect 129800 215000 132800 215200
rect 133000 215000 136000 215200
rect -136000 206000 -133000 215000
rect -132800 206000 -129800 215000
rect -57800 214985 136000 215000
rect -57800 212015 -32485 214985
rect -30505 212015 30215 214985
rect 32185 212015 136000 214985
rect -57800 212000 136000 212015
rect -57800 211800 -54800 212000
rect -54600 211800 -51600 212000
rect 26000 211800 29000 212000
rect 29200 211800 32200 212000
rect -57800 211785 32200 211800
rect -57800 208815 -32485 211785
rect -30505 208815 30215 211785
rect 32185 208815 32200 211785
rect -57800 208800 32200 208815
rect -93000 208585 93000 208600
rect -93000 205615 315 208585
rect 25685 205615 93000 208585
rect 129800 206000 132800 212000
rect 133000 206000 136000 212000
rect -93000 205600 93000 205615
rect -61000 205400 -58000 205600
rect -57800 205400 -54800 205600
rect 54800 205400 57800 205600
rect 58000 205400 61000 205600
rect -65000 205385 65000 205400
rect -65000 202415 315 205385
rect 25685 202415 65000 205385
rect -65000 202400 65000 202415
rect -61000 200000 -58000 202400
rect -57800 200000 -54800 202400
rect -26000 202185 3000 202200
rect -26000 201215 -25985 202185
rect -15 201215 3000 202185
rect -26000 200000 3000 201215
rect 54800 200000 57800 202400
rect 58000 200000 61000 202400
rect -4000 177000 4000 200000
<< via4 >>
rect -25685 221415 -315 224385
rect 315 221415 25685 224385
rect -25685 218215 -315 221185
rect 315 218215 25685 221185
rect -32485 212015 -30505 214985
rect 30215 212015 32185 214985
rect -32485 208815 -30505 211785
rect 30215 208815 32185 211785
rect 315 205615 25685 208585
rect 315 202415 25685 205385
rect -25985 201215 -15 202185
<< metal5 >>
rect -132800 221400 -51600 224400
rect -25700 224385 -300 224400
rect -25700 221415 -25685 224385
rect -315 221415 -300 224385
rect -25700 221400 -300 221415
rect 300 224385 25700 224400
rect 300 221415 315 224385
rect 25685 221415 25700 224385
rect 300 221400 25700 221415
rect -132800 221200 -129800 221400
rect -129600 221200 -126600 221400
rect -57800 221200 -54800 221400
rect -54600 221200 -51600 221400
rect -136000 218200 -51600 221200
rect -25700 221185 -300 221200
rect -25700 218215 -25685 221185
rect -315 218215 -300 221185
rect -25700 218200 -300 218215
rect 300 221185 25700 221200
rect 300 218215 315 221185
rect 25685 218215 25700 221185
rect 300 218200 25700 218215
rect -136000 218000 -133000 218200
rect -132800 218000 -129800 218200
rect -129600 218000 -126600 218200
rect -136000 215000 -126600 218000
rect -57800 215000 -54800 218200
rect -54600 215000 -51600 218200
rect 26000 215200 136000 218200
rect 26000 215000 29000 215200
rect 29200 215000 32200 215200
rect 129800 215000 132800 215200
rect 133000 215000 136000 215200
rect -136000 206000 -133000 215000
rect -132800 206000 -129800 215000
rect -57800 214985 136000 215000
rect -57800 212015 -32485 214985
rect -30505 212015 30215 214985
rect 32185 212015 136000 214985
rect -57800 212000 136000 212015
rect -57800 211800 -54800 212000
rect -54600 211800 -51600 212000
rect 26000 211800 29000 212000
rect 29200 211800 32200 212000
rect -57800 211785 32200 211800
rect -57800 208815 -32485 211785
rect -30505 208815 30215 211785
rect 32185 208815 32200 211785
rect -57800 208800 32200 208815
rect -93000 208585 93000 208600
rect -93000 205615 315 208585
rect 25685 205615 93000 208585
rect 129800 206000 132800 212000
rect 133000 206000 136000 212000
rect -93000 205600 93000 205615
rect -61000 205400 -58000 205600
rect -57800 205400 -54800 205600
rect 54800 205400 57800 205600
rect 58000 205400 61000 205600
rect -65000 205385 65000 205400
rect -65000 202415 315 205385
rect 25685 202415 65000 205385
rect -65000 202400 65000 202415
rect -61000 200000 -58000 202400
rect -57800 200000 -54800 202400
rect -26000 202185 3000 202200
rect -26000 201215 -25985 202185
rect -15 201215 3000 202185
rect -26000 200000 3000 201215
rect 54800 200000 57800 202400
rect 58000 200000 61000 202400
rect -4000 177000 4000 200000
use core  core_0
timestamp 1666566871
transform -1 0 -800 0 -1 208000
box 0 0 137200 208000
use core  core_1
timestamp 1666566871
transform 1 0 800 0 -1 208000
box 0 0 137200 208000
<< labels >>
rlabel metal5 -25700 221400 -22700 224400 7 GND
rlabel metal5 -54600 221400 -51600 224400 3 VH
rlabel metal5 22700 221400 25700 224400 3 Vout
<< end >>
