magic
tech sky130A
timestamp 1669125526
<< dnwell >>
rect 2450 9050 28150 34750
rect 33450 9050 59150 34750
<< obsactive >>
rect 0 41215 145000 47000
rect 0 37215 2006 41215
rect 9006 37215 54006 41215
rect 61006 37215 63006 41215
rect 70006 37215 128006 41215
rect 135006 37215 145000 41215
rect 0 36800 145000 37215
rect 0 7000 400 36800
rect 30200 7000 31400 36800
rect 61200 7000 62400 36800
rect 0 400 62400 7000
rect 98800 400 100400 36800
rect 136800 400 145000 36800
rect 0 -3000 145000 400
rect 52000 -10000 145000 -3000
<< metal3 >>
rect 7000 35996 56000 42000
rect 7000 33004 7104 35996
rect 55896 33004 56000 35996
rect 7000 33000 56000 33004
rect 69100 35996 129900 36000
rect 69100 33004 69104 35996
rect 129896 33004 129900 35996
rect 69100 33000 129900 33004
<< via3 >>
rect 7104 33004 55896 35996
rect 69104 33004 129896 35996
<< metal4 >>
rect 7100 35999 55900 36000
rect 7100 35996 7121 35999
rect 55879 35996 55900 35999
rect 7100 33004 7104 35996
rect 55896 33004 55900 35996
rect 7100 33001 7121 33004
rect 55879 33001 55900 33004
rect 7100 33000 55900 33001
rect 69000 35999 130000 42000
rect 69000 35996 69121 35999
rect 129879 35996 130000 35999
rect 69000 33004 69104 35996
rect 129896 33004 130000 35996
rect 69000 33001 69121 33004
rect 129879 33001 130000 33004
rect 69000 33000 130000 33001
<< via4 >>
rect 7121 35996 55879 35999
rect 7121 33004 55879 35996
rect 7121 33001 55879 33004
rect 69121 35996 129879 35999
rect 69121 33004 129879 35996
rect 69121 33001 129879 33004
<< metal5 >>
rect 7000 35999 56000 42000
rect 7000 33001 7121 35999
rect 55879 33001 56000 35999
rect 7000 33000 56000 33001
rect 69100 35999 129900 36000
rect 69100 33001 69121 35999
rect 129879 33001 129900 35999
rect 69100 33000 129900 33001
use flying_cap  flying_cap_0
timestamp 1668351020
transform -1 0 137170 0 -1 209000
box -590 0 137170 168000
use power_stage  power_stage_0
timestamp 1663434482
transform 0 1 0 -1 0 37200
box 0 0 36813 136813
<< end >>
