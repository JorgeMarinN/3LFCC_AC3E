magic
tech sky130A
timestamp 1662147188
<< metal3 >>
rect 1030 147980 69020 148000
rect 1030 147020 1050 147980
rect 69000 147020 69020 147980
rect 1030 146740 69020 147020
rect 71210 147980 136010 148000
rect 71210 147020 71230 147980
rect 135990 147020 136010 147980
rect 71210 147000 136010 147020
<< via3 >>
rect 1050 147020 69000 147980
rect 71230 147020 135990 147980
<< metal4 >>
rect 1030 147980 69020 148000
rect 1030 147020 1050 147980
rect 69000 147020 69020 147980
rect 1030 147000 69020 147020
rect 71210 147980 136010 148000
rect 71210 147020 71230 147980
rect 135990 147020 136010 147980
rect 71210 146740 136010 147020
<< via4 >>
rect 1050 147020 69000 147980
rect 71230 147020 135990 147980
<< metal5 >>
rect 1030 147980 69020 148000
rect 1030 147020 1050 147980
rect 69000 147020 69020 147980
rect 1030 146740 69020 147020
rect 71210 147980 136010 148000
rect 71210 147020 71230 147980
rect 135990 147020 136010 147980
rect 71210 147000 136010 147020
use flying_cap  flying_cap_0
timestamp 1662145806
transform 1 0 30 0 1 0
box 0 0 137170 146740
use power_stage  power_stage_0
timestamp 1662147188
transform 0 -1 137200 1 0 150000
box 0 0 37200 137200
<< end >>
