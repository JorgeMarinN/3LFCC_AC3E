* NGSPICE file created from converter.ext - technology: sky130A

.subckt nmos_waffle_36x36 w_n1200_n1200# a_n50_n50# a_112_3350# a_112_1150#
X0 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=8.80377e+15p pd=2.14718e+10u as=3.49194e+15p ps=2.36764e+10u w=4.38e+06u l=500000u
X1 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X5 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X6 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X7 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X8 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X9 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X10 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X11 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X12 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X13 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X14 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X15 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X16 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X17 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X18 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X19 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X20 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X21 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X22 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X23 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X24 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X25 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X26 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X27 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X28 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X29 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X30 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X31 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X32 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X33 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X34 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X35 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X36 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X37 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X38 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X39 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X40 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X41 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X42 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X43 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X44 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X45 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X46 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X47 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X48 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X49 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X50 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X51 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X52 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X53 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X54 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X55 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X56 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X57 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X58 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X59 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X60 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X61 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X62 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X63 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X64 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X65 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X66 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X67 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X68 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X69 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X70 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X71 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X72 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X73 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X74 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X75 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X76 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X77 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X78 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X79 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X80 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X81 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X82 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X83 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X84 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X85 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X86 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X87 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X88 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X89 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X90 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X91 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X92 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X93 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X94 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X95 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X96 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X97 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X98 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X99 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X100 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X101 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X102 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X103 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X104 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X105 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X106 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X107 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X108 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X109 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X110 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X111 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X112 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X113 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X114 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X115 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X116 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X117 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X118 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X119 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X120 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X121 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X122 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X123 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X124 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X125 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X126 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X127 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X128 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X129 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X130 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X131 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X132 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X133 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X134 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X135 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X136 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X137 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X138 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X139 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X140 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X141 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X142 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X143 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X144 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X145 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X146 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X147 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X148 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X149 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X150 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X151 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X152 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X153 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X154 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X155 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X156 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X157 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X158 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X159 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X160 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X161 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X162 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X163 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X164 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X165 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X166 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X167 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X168 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X169 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X170 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X171 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X172 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X173 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X174 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X175 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X176 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X177 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X178 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X179 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X180 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X181 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X182 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X183 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X184 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X185 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X186 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X187 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X188 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X189 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X190 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X191 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X192 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X193 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X194 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X195 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X196 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X197 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X198 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X199 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X200 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X201 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X202 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X203 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X204 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X205 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X206 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X207 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X208 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X209 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X210 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X211 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X212 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X213 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X214 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X215 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X216 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X217 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X218 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X219 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X220 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X221 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X222 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X223 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X224 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X225 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X226 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X227 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X228 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X229 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X230 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X231 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X232 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X233 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X234 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X235 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X236 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X237 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X238 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X239 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X240 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X241 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X242 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X243 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X244 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X245 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X246 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X247 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X248 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X249 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X250 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X251 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X252 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X253 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X254 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X255 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X256 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X257 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X258 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X259 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X260 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X261 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X262 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X263 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X264 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X265 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X266 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X267 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X268 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X269 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X270 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X271 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X272 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X273 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X274 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X275 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X276 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X277 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X278 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X279 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X280 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X281 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X282 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X283 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X284 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X285 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X286 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X287 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X288 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X289 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X290 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X291 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X292 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X293 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X294 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X295 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X296 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X297 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X298 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X299 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X300 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X301 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X302 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X303 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X304 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X305 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X306 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X307 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X308 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X309 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X310 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X311 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X312 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X313 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X314 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X315 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X316 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X317 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X318 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X319 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X320 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X321 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X322 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X323 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X324 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X325 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X326 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X327 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X328 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X329 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X330 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X331 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X332 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X333 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X334 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X335 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X336 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X337 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X338 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X339 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X340 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X341 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X342 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X343 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X344 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X345 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X346 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X347 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X348 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X349 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X350 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X351 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X352 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X353 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X354 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X355 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X356 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X357 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X358 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X359 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X360 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X361 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X362 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X363 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X364 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X365 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X366 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X367 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X368 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X369 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X370 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X371 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X372 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X373 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X374 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X375 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X376 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X377 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X378 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X379 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X380 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X381 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X382 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X383 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X384 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X385 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X386 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X387 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X388 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X389 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X390 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X391 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X392 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X393 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X394 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X395 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X396 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X397 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X398 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X399 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X400 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X401 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X402 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X403 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X404 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X405 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X406 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X407 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X408 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X409 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X410 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X411 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X412 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X413 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X414 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X415 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X416 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X417 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X418 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X419 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X420 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X421 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X422 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X423 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X424 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X425 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X426 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X427 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X428 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X429 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X430 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X431 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X432 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X433 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X434 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X435 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X436 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X437 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X438 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X439 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X440 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X441 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X442 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X443 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X444 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X445 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X446 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X447 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X448 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X449 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X450 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X451 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X452 w_n1200_n1200# a_n50_n50# a_112_1150# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=8.1096e+12p ps=5.636e+07u w=4.38e+06u l=500000u
X453 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X454 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X455 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X456 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X457 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X458 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X459 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X460 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X461 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X462 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X463 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X464 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X465 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X466 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X467 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X468 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X469 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X470 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X471 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X472 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X473 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X474 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X475 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X476 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X477 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X478 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X479 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X480 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X481 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X482 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X483 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X484 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X485 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X486 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X487 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X488 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X489 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X490 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X491 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X492 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X493 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X494 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X495 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X496 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X497 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X498 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X499 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X500 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X501 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X502 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X503 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X504 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X505 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X506 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X507 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X508 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X509 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X510 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X511 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X512 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X513 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X514 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X515 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X516 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X517 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X518 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X519 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X520 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X521 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X522 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X523 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X524 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X525 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X526 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X527 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X528 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X529 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X530 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X531 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X532 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X533 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X534 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X535 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X536 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X537 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X538 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X539 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X540 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X541 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X542 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X543 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X544 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X545 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X546 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X547 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X548 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X549 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X550 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X551 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X552 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X553 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X554 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X555 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X556 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X557 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X558 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X559 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X560 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X561 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X562 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X563 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X564 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X565 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X566 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X567 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X568 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X569 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X570 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X571 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X572 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X573 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X574 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X575 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X576 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X577 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X578 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X579 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X580 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X581 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X582 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X583 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X584 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X585 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X586 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X587 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X588 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X589 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X590 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X591 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X592 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X593 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X594 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X595 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X596 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X597 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X598 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X599 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X600 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X601 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X602 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X603 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X604 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X605 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X606 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X607 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X608 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X609 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X610 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X611 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X612 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X613 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X614 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X615 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X616 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X617 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X618 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X619 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X620 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X621 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X622 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X623 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X624 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X625 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X626 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X627 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X628 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X629 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X630 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X631 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X632 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X633 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X634 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X635 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X636 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X637 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X638 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X639 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X640 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X641 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X642 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X643 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X644 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X645 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X646 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X647 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X648 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X649 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X650 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X651 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X652 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X653 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X654 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X655 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X656 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X657 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X658 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X659 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X660 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X661 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X662 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X663 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X664 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X665 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X666 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X667 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X668 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X669 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X670 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X671 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X672 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X673 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X674 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X675 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X676 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X677 w_n1200_n1200# a_n50_n50# a_112_1150# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X678 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X679 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X680 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X681 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X682 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X683 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X684 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X685 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X686 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X687 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X688 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X689 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X690 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X691 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X692 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X693 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X694 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X695 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X696 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X697 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X698 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X699 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X700 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X701 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X702 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X703 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X704 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X705 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X706 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X707 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X708 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X709 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X710 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X711 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X712 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X713 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X714 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X715 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X716 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X717 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X718 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X719 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X720 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X721 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X722 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X723 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X724 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X725 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X726 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X727 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X728 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X729 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X730 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X731 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X732 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X733 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X734 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X735 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X736 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X737 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X738 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X739 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X740 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X741 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X742 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X743 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X744 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X745 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X746 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X747 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X748 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X749 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X750 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X751 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X752 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X753 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X754 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X755 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X756 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X757 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X758 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X759 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X760 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X761 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X762 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X763 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X764 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X765 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X766 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X767 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X768 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X769 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X770 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X771 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X772 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X773 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X774 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X775 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X776 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X777 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X778 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X779 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X780 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X781 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X782 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X783 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X784 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X785 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X786 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X787 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X788 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X789 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X790 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X791 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X792 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X793 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X794 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X795 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X796 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X797 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X798 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X799 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X800 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X801 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X802 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X803 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X804 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X805 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X806 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X807 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X808 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X809 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X810 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X811 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X812 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X813 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X814 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X815 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X816 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X817 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X818 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X819 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X820 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X821 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X822 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X823 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X824 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X825 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X826 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X827 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X828 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X829 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X830 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X831 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X832 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X833 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X834 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X835 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X836 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X837 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X838 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X839 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X840 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X841 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X842 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X843 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X844 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X845 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X846 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X847 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X848 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X849 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X850 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X851 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X852 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X853 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X854 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X855 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X856 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X857 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X858 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X859 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X860 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X861 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X862 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X863 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X864 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X865 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X866 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X867 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X868 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X869 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X870 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X871 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X872 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X873 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X874 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X875 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X876 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X877 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X878 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X879 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X880 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X881 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X882 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X883 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X884 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X885 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X886 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X887 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X888 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X889 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X890 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X891 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X892 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X893 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X894 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X895 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X896 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X897 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X898 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X899 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X900 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X901 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X902 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X903 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X904 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X905 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X906 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X907 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X908 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X909 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X910 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X911 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X912 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X913 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X914 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X915 w_n1200_n1200# a_n50_n50# a_112_1150# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X916 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X917 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X918 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X919 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X920 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X921 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X922 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X923 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X924 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X925 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X926 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X927 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X928 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X929 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X930 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X931 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X932 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X933 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X934 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X935 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X936 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X937 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X938 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X939 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X940 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X941 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X942 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X943 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X944 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X945 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X946 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X947 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X948 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X949 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X950 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X951 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X952 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X953 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X954 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X955 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X956 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X957 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X958 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X959 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X960 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X961 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X962 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X963 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X964 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X965 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X966 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X967 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X968 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X969 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X970 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X971 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X972 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X973 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X974 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X975 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X976 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X977 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X978 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X979 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X980 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X981 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X982 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X983 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X984 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X985 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X986 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X987 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X988 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X989 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X990 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X991 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X992 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X993 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X994 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X995 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X996 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X997 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X998 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X999 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1000 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1001 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1002 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1003 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1004 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1005 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1006 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1007 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1008 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1009 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1010 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1011 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1012 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1013 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1014 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1015 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1016 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1017 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1018 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1019 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1020 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1021 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1022 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1023 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1024 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1025 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1026 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1027 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1028 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1029 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1030 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1031 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1032 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1033 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1034 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1035 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1036 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1037 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1038 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1039 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1040 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1041 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1042 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1043 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1044 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1045 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1046 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1047 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1048 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1049 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1050 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1051 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1052 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1053 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1054 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1055 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1056 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1057 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1058 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1059 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1060 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1061 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1062 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1063 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1064 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1065 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1066 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1067 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1068 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1069 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1070 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1071 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1072 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1073 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1074 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1075 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1076 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1077 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1078 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1079 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1080 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1081 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1082 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1083 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1084 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1085 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1086 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1087 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1088 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1089 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1090 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1091 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1092 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1093 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1094 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1095 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1096 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1097 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1098 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1099 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1100 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1101 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1102 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1103 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1104 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1105 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1106 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1107 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1108 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1109 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1110 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1111 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1112 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1113 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1114 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1115 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1116 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1117 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1118 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1119 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1120 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1121 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1122 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1123 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1124 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1125 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1126 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1127 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1128 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1129 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1130 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1131 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1132 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1133 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1134 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1135 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1136 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1137 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1138 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1139 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1140 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1141 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1142 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1143 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1144 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1145 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1146 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1147 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1148 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1149 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1150 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1151 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1152 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1153 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1154 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1155 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1156 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1157 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1158 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1159 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1160 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1161 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1162 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1163 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1164 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1165 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1166 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1167 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1168 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1169 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1170 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1171 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1172 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1173 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1174 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1175 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1176 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1177 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1178 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1179 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1180 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1181 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1182 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1183 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1184 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1185 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1186 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1187 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1188 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1189 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1190 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1191 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1192 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1193 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1194 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1195 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1196 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1197 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1198 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1199 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1200 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1201 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1202 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1203 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1204 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1205 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1206 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1207 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1208 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1209 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1210 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1211 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1212 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1213 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1214 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1215 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1216 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1217 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1218 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1219 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1220 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1221 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1222 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1223 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1224 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1225 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1226 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1227 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1228 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1229 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1230 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1231 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1232 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1233 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1234 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1235 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1236 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1237 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1238 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1239 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1240 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1241 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1242 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1243 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1244 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1245 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1246 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1247 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1248 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1249 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1250 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1251 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1252 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1253 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1254 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1255 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1256 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1257 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1258 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1259 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1260 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1261 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1262 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1263 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1264 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1265 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1266 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1267 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1268 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1269 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1270 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1271 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1272 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1273 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1274 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1275 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1276 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1277 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1278 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1279 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1280 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1281 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1282 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1283 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1284 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1285 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1286 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1287 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1288 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1289 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1290 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1291 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1292 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1293 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1294 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1295 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1296 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1297 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1298 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1299 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1300 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1301 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1302 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1303 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1304 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1305 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1306 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1307 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1308 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1309 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1310 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1311 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1312 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1313 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1314 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1315 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1316 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1317 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1318 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1319 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1320 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1321 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1322 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1323 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1324 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1325 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1326 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1327 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1328 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1329 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1330 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1331 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1332 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1333 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1334 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1335 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1336 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1337 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1338 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1339 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1340 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1341 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1342 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1343 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1344 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1345 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1346 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1347 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1348 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1349 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1350 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1351 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1352 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1353 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1354 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1355 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1356 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1357 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1358 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1359 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1360 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1361 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1362 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1363 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1364 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1365 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1366 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1367 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1368 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1369 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1370 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1371 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1372 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1373 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1374 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1375 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1376 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1377 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1378 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1379 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1380 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1381 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1382 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1383 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1384 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1385 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1386 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1387 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1388 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1389 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1390 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1391 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1392 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1393 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1394 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1395 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1396 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1397 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1398 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1399 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1400 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1401 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1402 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1403 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1404 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1405 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1406 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1407 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1408 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1409 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1410 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1411 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1412 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1413 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1414 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1415 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1416 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1417 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1418 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1419 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1420 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1421 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1422 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1423 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1424 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1425 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1426 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1427 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1428 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1429 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1430 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1431 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1432 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1433 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1434 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1435 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1436 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1437 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1438 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1439 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1440 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1441 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1442 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1443 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1444 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1445 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1446 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1447 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1448 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1449 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1450 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1451 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1452 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1453 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1454 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1455 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1456 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1457 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1458 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1459 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1460 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1461 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1462 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1463 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1464 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1465 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1466 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1467 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1468 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1469 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1470 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1471 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1472 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1473 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1474 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1475 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1476 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1477 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1478 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1479 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1480 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1481 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1482 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1483 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1484 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1485 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1486 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1487 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1488 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1489 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1490 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1491 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1492 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1493 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1494 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1495 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1496 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1497 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1498 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1499 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1500 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1501 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1502 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1503 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1504 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1505 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1506 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1507 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1508 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1509 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1510 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1511 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1512 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1513 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1514 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1515 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1516 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1517 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1518 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1519 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1520 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1521 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1522 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1523 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1524 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1525 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1526 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1527 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1528 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1529 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1530 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1531 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1532 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1533 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1534 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1535 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1536 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1537 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1538 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1539 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1540 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1541 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1542 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1543 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1544 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1545 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1546 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1547 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1548 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1549 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1550 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1551 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1552 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1553 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1554 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1555 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1556 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1557 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1558 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1559 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1560 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1561 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1562 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1563 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1564 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1565 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1566 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1567 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1568 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1569 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1570 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1571 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1572 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1573 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1574 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1575 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1576 w_n1200_n1200# a_n50_n50# a_112_1150# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1577 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1578 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1579 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1580 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1581 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1582 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1583 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1584 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1585 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1586 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1587 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1588 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1589 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1590 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1591 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1592 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1593 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1594 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1595 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1596 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1597 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1598 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1599 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1600 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1601 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1602 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1603 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1604 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1605 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1606 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1607 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1608 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1609 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1610 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1611 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1612 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1613 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1614 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1615 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1616 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1617 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1618 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1619 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1620 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1621 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1622 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1623 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1624 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1625 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1626 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1627 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1628 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1629 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1630 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1631 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1632 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1633 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1634 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1635 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1636 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1637 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1638 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1639 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1640 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1641 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1642 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1643 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1644 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1645 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1646 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1647 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1648 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1649 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1650 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1651 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1652 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1653 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1654 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1655 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1656 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1657 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1658 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1659 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1660 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1661 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1662 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1663 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1664 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1665 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1666 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1667 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1668 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1669 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1670 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1671 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1672 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1673 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1674 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1675 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1676 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1677 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1678 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1679 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1680 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1681 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1682 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1683 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1684 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1685 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1686 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1687 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1688 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1689 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1690 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1691 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1692 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1693 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1694 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1695 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1696 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1697 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1698 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1699 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1700 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1701 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1702 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1703 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1704 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1705 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1706 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1707 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1708 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1709 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1710 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1711 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1712 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1713 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1714 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1715 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1716 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1717 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1718 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1719 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1720 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1721 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1722 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1723 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1724 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1725 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1726 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1727 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1728 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1729 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1730 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1731 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1732 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1733 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1734 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1735 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1736 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1737 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1738 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1739 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1740 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1741 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1742 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1743 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1744 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1745 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1746 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1747 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1748 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1749 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1750 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1751 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1752 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1753 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1754 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1755 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1756 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1757 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1758 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1759 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1760 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1761 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1762 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1763 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1764 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1765 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1766 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1767 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1768 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1769 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1770 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1771 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1772 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1773 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1774 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1775 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1776 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1777 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1778 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1779 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1780 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1781 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1782 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1783 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1784 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1785 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1786 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1787 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1788 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1789 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1790 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1791 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1792 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1793 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1794 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1795 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1796 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1797 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1798 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1799 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1800 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1801 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1802 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1803 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1804 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1805 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1806 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1807 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1808 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1809 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1810 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1811 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1812 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1813 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1814 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1815 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1816 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1817 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1818 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1819 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1820 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1821 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1822 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1823 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1824 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1825 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1826 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1827 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1828 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1829 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1830 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1831 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1832 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1833 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1834 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1835 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1836 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1837 a_112_1150# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1838 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1839 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1840 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1841 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1842 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1843 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1844 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1845 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1846 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1847 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1848 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1849 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1850 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1851 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1852 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1853 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1854 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1855 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1856 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1857 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1858 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1859 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1860 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1861 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1862 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1863 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1864 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1865 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1866 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1867 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1868 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1869 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1870 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1871 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1872 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1873 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1874 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1875 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1876 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1877 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1878 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1879 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1880 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1881 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1882 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1883 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1884 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1885 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1886 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1887 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1888 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1889 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1890 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1891 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1892 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1893 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1894 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1895 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1896 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1897 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1898 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1899 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1900 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1901 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1902 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1903 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1904 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1905 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1906 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1907 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1908 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1909 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1910 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1911 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1912 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1913 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1914 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1915 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1916 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1917 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1918 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1919 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1920 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1921 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1922 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1923 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1924 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1925 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1926 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1927 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1928 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1929 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1930 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1931 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1932 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1933 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1934 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1935 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1936 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1937 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1938 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1939 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1940 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1941 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1942 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1943 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1944 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1945 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1946 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1947 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1948 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1949 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1950 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1951 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1952 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1953 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1954 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1955 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1956 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1957 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1958 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1959 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1960 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1961 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1962 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1963 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1964 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1965 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1966 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1967 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1968 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1969 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1970 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1971 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1972 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1973 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1974 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1975 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1976 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1977 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1978 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1979 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1980 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1981 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1982 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1983 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1984 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1985 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1986 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1987 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1988 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1989 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1990 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1991 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1992 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1993 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1994 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1995 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1996 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1997 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1998 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1999 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2000 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2001 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2002 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2003 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2004 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2005 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2006 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2007 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2008 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2009 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2010 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2011 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2012 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2013 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2014 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2015 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2016 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2017 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2018 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2019 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2020 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2021 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2022 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2023 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2024 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2025 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2026 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2027 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2028 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2029 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2030 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2031 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2032 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2033 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2034 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2035 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2036 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2037 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2038 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2039 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2040 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2041 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2042 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2043 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2044 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2045 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2046 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2047 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2048 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2049 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2050 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2051 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2052 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2053 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2054 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2055 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2056 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2057 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2058 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2059 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2060 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2061 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2062 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2063 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2064 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2065 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2066 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2067 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2068 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2069 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2070 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2071 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2072 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2073 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2074 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2075 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2076 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2077 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2078 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2079 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2080 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2081 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2082 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2083 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2084 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2085 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2086 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2087 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2088 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2089 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2090 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2091 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2092 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2093 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2094 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2095 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2096 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2097 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2098 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2099 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2100 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2101 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2102 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2103 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2104 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2105 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2106 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2107 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2108 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2109 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2110 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2111 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2112 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2113 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2114 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2115 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2116 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2117 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2118 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2119 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2120 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2121 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2122 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2123 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2124 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2125 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2126 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2127 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2128 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2129 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2130 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2131 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2132 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2133 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2134 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2135 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2136 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2137 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2138 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2139 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2140 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2141 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2142 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2143 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2144 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2145 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2146 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2147 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2148 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2149 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2150 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2151 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2152 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2153 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2154 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2155 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2156 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2157 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2158 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2159 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2160 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2161 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2162 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2163 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2164 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2165 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2166 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2167 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2168 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2169 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2170 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2171 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2172 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2173 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2174 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2175 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2176 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2177 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2178 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2179 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2180 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2181 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2182 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2183 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2184 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2185 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2186 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2187 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2188 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2189 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2190 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2191 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2192 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2193 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2194 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2195 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2196 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2197 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2198 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2199 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2200 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2201 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2202 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2203 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2204 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2205 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2206 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2207 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2208 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2209 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2210 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2211 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2212 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2213 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2214 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2215 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2216 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2217 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2218 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2219 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2220 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2221 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2222 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2223 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2224 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2225 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2226 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2227 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2228 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2229 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2230 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2231 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2232 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2233 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2234 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2235 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2236 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2237 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2238 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2239 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2240 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2241 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2242 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2243 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2244 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2245 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2246 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2247 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2248 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2249 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2250 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2251 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2252 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2253 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2254 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2255 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2256 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2257 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2258 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2259 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2260 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2261 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2262 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2263 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2264 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2265 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2266 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2267 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2268 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2269 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2270 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2271 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2272 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2273 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2274 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2275 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2276 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2277 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2278 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2279 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2280 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2281 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2282 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2283 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2284 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2285 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2286 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2287 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2288 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2289 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2290 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2291 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2292 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2293 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2294 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2295 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2296 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2297 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2298 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2299 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2300 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2301 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2302 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2303 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2304 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2305 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2306 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2307 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2308 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2309 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2310 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2311 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2312 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2313 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2314 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2315 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2316 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2317 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2318 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2319 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2320 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2321 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2322 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2323 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2324 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2325 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2326 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2327 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2328 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2329 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2330 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2331 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2332 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2333 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2334 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2335 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2336 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2337 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2338 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2339 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2340 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2341 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2342 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2343 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2344 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2345 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2346 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2347 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2348 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2349 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2350 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2351 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2352 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2353 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2354 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2355 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2356 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2357 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2358 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2359 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2360 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2361 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2362 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2363 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2364 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2365 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2366 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2367 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2368 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2369 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2370 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2371 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2372 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2373 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2374 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2375 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2376 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2377 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2378 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2379 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2380 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2381 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2382 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2383 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2384 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2385 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2386 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2387 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2388 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2389 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2390 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2391 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2392 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2393 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2394 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2395 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2396 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2397 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2398 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2399 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2400 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2401 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2402 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2403 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2404 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2405 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2406 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2407 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2408 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2409 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2410 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2411 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2412 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2413 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2414 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2415 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2416 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2417 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2418 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2419 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2420 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2421 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2422 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2423 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2424 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2425 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2426 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2427 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2428 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2429 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2430 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2431 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2432 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2433 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2434 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2435 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2436 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2437 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2438 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2439 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2440 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2441 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2442 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2443 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2444 a_112_1150# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2445 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2446 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2447 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2448 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2449 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2450 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2451 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2452 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2453 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2454 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2455 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2456 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2457 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2458 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2459 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2460 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2461 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2462 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2463 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2464 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2465 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2466 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2467 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2468 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2469 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2470 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2471 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2472 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2473 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2474 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2475 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2476 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2477 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2478 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2479 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2480 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2481 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2482 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2483 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2484 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2485 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2486 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2487 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2488 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2489 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2490 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2491 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2492 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2493 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2494 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2495 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2496 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2497 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2498 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2499 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2500 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2501 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2502 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2503 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2504 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2505 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2506 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2507 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2508 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2509 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2510 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2511 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2512 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2513 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2514 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2515 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2516 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2517 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2518 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2519 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
.ends

.subckt pmos_waffle_48x48 w_n1200_n1200# a_n50_n50# a_112_3350# a_112_1150#
X0 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=6.26247e+15p pd=4.24392e+10u as=1.56918e+16p ps=3.81907e+10u w=4.38e+06u l=500000u
X1 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X5 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X6 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X7 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X8 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X9 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X10 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X11 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X12 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X13 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X14 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X15 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X16 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X17 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X18 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X19 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X20 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X21 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X22 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X23 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X24 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X25 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X26 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X27 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X28 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X29 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X30 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X31 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X32 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X33 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X34 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X35 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X36 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X37 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X38 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X39 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X40 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X41 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X42 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X43 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X44 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X45 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X46 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X47 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X48 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X49 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X50 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X51 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X52 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X53 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X54 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X55 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X56 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X57 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X58 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X59 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X60 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X61 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X62 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X63 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X64 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X65 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X66 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X67 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X68 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X69 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X70 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X71 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X72 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X73 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X74 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X75 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X76 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X77 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X78 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X79 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X80 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X81 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X82 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X83 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X84 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X85 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X86 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X87 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X88 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X89 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X90 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X91 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X92 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X93 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X94 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X95 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X96 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X97 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X98 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X99 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X100 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X101 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X102 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X103 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X104 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X105 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X106 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X107 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X108 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X109 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X110 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X111 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X112 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X113 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X114 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X115 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X116 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X117 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X118 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X119 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X120 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X121 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X122 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X123 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X124 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X125 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X126 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X127 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X128 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X129 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X130 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X131 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X132 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X133 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X134 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X135 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X136 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X137 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X138 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X139 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X140 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X141 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X142 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X143 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X144 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X145 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X146 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X147 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X148 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X149 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X150 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X151 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X152 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X153 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X154 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X155 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X156 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X157 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X158 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X159 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X160 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X161 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X162 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X163 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X164 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X165 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X166 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X167 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X168 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X169 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X170 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X171 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X172 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X173 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X174 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X175 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X176 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X177 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X178 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X179 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X180 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X181 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X182 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X183 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X184 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X185 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X186 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X187 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X188 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X189 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X190 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X191 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X192 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X193 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X194 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X195 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X196 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X197 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X198 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X199 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X200 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X201 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X202 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X203 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X204 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X205 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X206 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X207 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X208 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X209 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X210 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X211 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X212 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X213 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X214 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X215 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X216 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X217 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X218 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X219 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X220 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X221 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X222 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X223 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X224 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X225 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X226 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X227 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X228 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X229 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X230 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X231 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X232 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X233 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X234 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X235 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X236 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X237 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X238 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X239 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X240 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X241 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X242 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X243 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X244 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X245 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X246 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X247 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X248 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X249 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X250 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X251 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X252 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X253 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X254 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X255 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X256 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X257 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X258 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X259 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X260 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X261 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X262 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X263 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X264 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X265 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X266 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X267 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X268 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X269 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X270 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X271 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X272 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X273 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X274 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X275 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X276 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X277 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X278 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X279 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X280 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X281 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X282 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X283 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X284 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X285 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X286 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X287 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X288 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X289 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X290 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X291 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X292 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X293 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X294 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X295 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X296 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X297 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X298 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X299 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X300 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X301 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X302 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X303 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X304 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X305 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X306 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X307 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X308 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X309 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X310 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X311 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X312 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X313 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X314 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X315 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X316 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X317 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X318 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X319 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X320 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X321 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X322 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X323 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X324 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X325 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X326 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X327 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X328 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X329 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X330 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X331 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X332 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X333 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X334 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X335 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X336 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X337 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X338 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X339 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X340 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X341 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X342 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X343 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X344 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X345 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X346 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X347 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X348 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X349 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X350 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X351 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X352 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X353 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X354 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X355 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X356 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X357 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X358 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X359 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X360 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X361 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X362 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X363 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X364 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X365 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X366 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X367 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X368 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X369 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X370 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X371 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X372 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X373 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X374 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X375 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X376 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X377 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X378 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X379 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X380 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X381 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X382 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X383 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X384 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X385 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X386 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X387 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X388 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X389 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X390 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X391 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X392 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X393 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X394 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X395 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X396 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X397 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X398 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X399 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X400 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X401 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X402 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X403 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X404 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X405 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X406 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X407 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X408 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X409 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X410 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X411 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X412 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X413 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X414 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X415 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X416 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X417 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X418 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X419 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X420 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X421 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X422 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X423 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X424 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X425 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X426 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X427 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X428 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X429 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X430 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X431 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X432 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X433 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X434 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X435 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X436 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X437 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X438 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X439 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X440 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X441 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X442 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X443 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X444 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X445 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X446 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X447 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X448 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X449 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X450 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X451 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X452 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X453 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X454 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X455 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X456 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X457 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X458 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X459 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X460 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X461 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X462 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X463 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X464 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X465 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X466 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X467 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X468 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X469 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X470 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X471 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X472 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X473 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X474 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X475 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X476 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X477 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X478 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X479 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X480 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X481 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X482 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X483 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X484 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X485 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X486 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X487 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X488 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X489 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X490 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X491 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X492 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X493 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X494 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X495 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X496 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X497 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X498 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X499 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X500 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X501 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X502 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X503 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X504 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X505 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X506 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X507 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X508 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X509 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X510 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X511 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X512 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X513 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X514 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X515 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X516 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X517 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X518 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X519 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X520 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X521 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X522 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X523 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X524 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X525 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X526 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X527 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X528 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X529 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X530 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X531 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X532 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X533 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X534 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X535 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X536 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X537 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X538 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X539 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X540 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X541 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X542 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X543 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X544 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X545 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X546 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X547 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X548 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X549 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X550 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X551 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X552 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X553 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X554 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X555 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X556 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X557 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X558 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X559 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X560 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X561 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X562 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X563 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X564 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X565 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X566 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X567 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X568 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X569 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X570 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X571 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X572 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X573 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X574 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X575 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X576 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X577 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X578 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X579 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X580 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X581 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X582 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X583 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X584 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X585 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X586 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X587 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X588 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X589 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X590 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X591 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X592 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X593 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X594 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X595 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X596 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X597 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X598 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X599 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X600 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X601 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X602 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X603 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X604 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X605 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X606 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X607 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X608 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X609 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X610 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X611 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X612 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X613 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X614 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X615 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X616 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X617 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X618 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X619 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X620 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X621 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X622 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X623 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X624 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X625 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X626 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X627 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X628 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X629 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X630 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X631 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X632 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X633 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X634 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X635 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X636 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X637 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X638 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X639 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X640 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X641 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X642 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X643 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X644 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X645 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X646 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X647 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X648 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X649 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X650 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X651 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X652 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X653 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X654 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X655 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X656 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X657 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X658 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X659 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X660 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X661 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X662 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X663 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X664 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X665 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X666 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X667 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X668 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X669 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X670 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X671 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X672 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X673 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X674 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X675 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X676 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X677 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X678 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X679 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X680 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X681 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X682 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X683 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X684 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X685 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X686 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X687 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X688 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X689 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X690 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X691 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X692 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X693 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X694 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X695 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X696 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X697 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X698 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X699 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X700 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X701 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X702 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X703 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X704 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X705 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X706 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X707 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X708 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X709 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X710 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X711 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X712 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X713 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X714 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X715 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X716 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X717 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X718 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X719 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X720 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X721 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X722 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X723 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X724 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X725 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X726 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X727 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X728 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X729 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X730 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X731 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X732 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X733 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X734 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X735 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X736 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X737 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X738 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X739 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X740 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X741 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X742 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X743 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X744 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X745 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X746 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X747 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X748 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X749 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X750 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X751 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X752 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X753 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X754 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X755 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X756 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X757 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X758 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X759 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X760 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X761 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X762 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X763 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X764 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X765 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X766 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X767 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X768 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X769 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X770 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X771 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X772 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X773 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X774 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X775 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X776 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X777 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X778 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X779 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X780 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X781 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X782 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X783 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X784 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X785 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X786 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X787 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X788 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X789 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X790 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X791 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X792 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X793 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X794 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X795 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X796 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X797 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X798 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X799 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X800 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X801 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X802 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X803 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X804 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X805 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X806 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X807 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X808 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X809 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X810 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X811 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X812 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X813 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X814 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X815 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X816 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X817 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X818 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X819 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X820 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X821 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X822 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X823 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X824 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X825 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X826 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X827 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X828 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X829 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X830 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X831 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X832 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X833 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X834 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X835 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X836 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X837 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X838 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X839 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X840 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X841 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X842 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X843 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X844 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X845 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X846 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X847 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X848 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X849 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X850 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X851 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X852 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X853 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X854 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X855 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X856 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X857 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X858 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X859 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X860 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X861 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X862 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X863 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X864 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X865 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X866 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X867 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X868 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X869 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X870 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X871 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X872 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X873 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X874 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X875 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X876 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X877 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X878 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X879 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X880 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X881 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X882 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X883 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X884 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X885 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X886 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X887 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X888 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X889 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X890 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X891 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X892 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X893 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X894 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X895 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X896 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X897 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X898 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X899 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X900 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X901 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X902 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X903 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X904 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X905 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X906 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X907 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X908 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X909 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X910 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X911 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X912 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X913 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X914 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X915 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X916 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X917 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X918 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X919 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X920 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X921 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X922 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X923 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X924 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X925 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X926 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X927 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X928 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X929 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X930 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X931 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X932 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X933 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X934 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X935 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X936 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X937 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X938 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X939 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X940 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X941 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X942 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X943 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X944 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X945 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X946 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X947 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X948 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X949 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X950 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X951 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X952 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X953 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X954 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X955 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X956 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X957 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X958 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X959 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X960 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X961 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X962 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X963 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X964 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X965 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X966 w_n1200_n1200# a_n50_n50# a_112_1150# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.1096e+12p ps=5.636e+07u w=4.38e+06u l=500000u
X967 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X968 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X969 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X970 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X971 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X972 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X973 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X974 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X975 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X976 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X977 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X978 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X979 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X980 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X981 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X982 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X983 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X984 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X985 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X986 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X987 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X988 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X989 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X990 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X991 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X992 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X993 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X994 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X995 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X996 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X997 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X998 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X999 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1000 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1001 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1002 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1003 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1004 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1005 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1006 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1007 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1008 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1009 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1010 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1011 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1012 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1013 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1014 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1015 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1016 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1017 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1018 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1019 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1020 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1021 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1022 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1023 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1024 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1025 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1026 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1027 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1028 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1029 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1030 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1031 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1032 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1033 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1034 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1035 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1036 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1037 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1038 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1039 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1040 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1041 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1042 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1043 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1044 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1045 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1046 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1047 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1048 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1049 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1050 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1051 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1052 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1053 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1054 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1055 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1056 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1057 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1058 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1059 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1060 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1061 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1062 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1063 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1064 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1065 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1066 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1067 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1068 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1069 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1070 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1071 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1072 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1073 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1074 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1075 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1076 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1077 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1078 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1079 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1080 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1081 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1082 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1083 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1084 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1085 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1086 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1087 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1088 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1089 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1090 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1091 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1092 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1093 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1094 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1095 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1096 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1097 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1098 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1099 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1100 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1101 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1102 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1103 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1104 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1105 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1106 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1107 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1108 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1109 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1110 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1111 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1112 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1113 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1114 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1115 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1116 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1117 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1118 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1119 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1120 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1121 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1122 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1123 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1124 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1125 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1126 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1127 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1128 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1129 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1130 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1131 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1132 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1133 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1134 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1135 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1136 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1137 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1138 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1139 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1140 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1141 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1142 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1143 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1144 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1145 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1146 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1147 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1148 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1149 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1150 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1151 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1152 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1153 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1154 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1155 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1156 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1157 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1158 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1159 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1160 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1161 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1162 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1163 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1164 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1165 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1166 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1167 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1168 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1169 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1170 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1171 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1172 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1173 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1174 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1175 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1176 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1177 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1178 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1179 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1180 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1181 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1182 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1183 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1184 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1185 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1186 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1187 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1188 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1189 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1190 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1191 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1192 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1193 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1194 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1195 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1196 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1197 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1198 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1199 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1200 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1201 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1202 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1203 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1204 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1205 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1206 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1207 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1208 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1209 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1210 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1211 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1212 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1213 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1214 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1215 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1216 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1217 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1218 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1219 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1220 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1221 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1222 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1223 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1224 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1225 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1226 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1227 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1228 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1229 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1230 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1231 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1232 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1233 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1234 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1235 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1236 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1237 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1238 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1239 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1240 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1241 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1242 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1243 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1244 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1245 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1246 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1247 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1248 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1249 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1250 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1251 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1252 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1253 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1254 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1255 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1256 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1257 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1258 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1259 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1260 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1261 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1262 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1263 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1264 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1265 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1266 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1267 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1268 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1269 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1270 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1271 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1272 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1273 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1274 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1275 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1276 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1277 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1278 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1279 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1280 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1281 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1282 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1283 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1284 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1285 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1286 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1287 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1288 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1289 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1290 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1291 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1292 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1293 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1294 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1295 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1296 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1297 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1298 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1299 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1300 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1301 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1302 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1303 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1304 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1305 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1306 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1307 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1308 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1309 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1310 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1311 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1312 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1313 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1314 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1315 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1316 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1317 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1318 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1319 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1320 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1321 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1322 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1323 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1324 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1325 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1326 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1327 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1328 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1329 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1330 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1331 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1332 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1333 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1334 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1335 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1336 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1337 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1338 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1339 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1340 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1341 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1342 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1343 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1344 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1345 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1346 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1347 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1348 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1349 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1350 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1351 w_n1200_n1200# a_n50_n50# a_112_1150# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1352 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1353 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1354 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1355 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1356 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1357 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1358 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1359 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1360 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1361 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1362 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1363 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1364 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1365 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1366 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1367 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1368 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1369 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1370 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1371 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1372 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1373 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1374 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1375 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1376 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1377 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1378 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1379 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1380 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1381 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1382 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1383 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1384 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1385 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1386 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1387 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1388 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1389 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1390 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1391 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1392 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1393 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1394 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1395 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1396 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1397 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1398 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1399 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1400 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1401 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1402 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1403 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1404 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1405 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1406 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1407 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1408 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1409 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1410 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1411 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1412 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1413 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1414 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1415 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1416 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1417 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1418 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1419 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1420 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1421 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1422 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1423 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1424 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1425 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1426 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1427 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1428 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1429 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1430 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1431 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1432 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1433 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1434 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1435 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1436 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1437 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1438 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1439 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1440 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1441 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1442 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1443 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1444 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1445 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1446 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1447 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1448 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1449 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1450 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1451 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1452 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1453 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1454 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1455 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1456 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1457 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1458 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1459 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1460 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1461 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1462 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1463 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1464 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1465 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1466 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1467 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1468 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1469 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1470 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1471 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1472 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1473 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1474 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1475 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1476 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1477 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1478 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1479 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1480 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1481 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1482 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1483 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1484 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1485 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1486 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1487 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1488 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1489 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1490 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1491 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1492 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1493 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1494 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1495 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1496 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1497 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1498 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1499 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1500 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1501 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1502 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1503 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1504 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1505 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1506 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1507 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1508 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1509 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1510 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1511 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1512 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1513 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1514 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1515 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1516 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1517 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1518 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1519 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1520 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1521 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1522 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1523 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1524 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1525 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1526 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1527 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1528 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1529 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1530 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1531 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1532 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1533 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1534 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1535 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1536 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1537 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1538 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1539 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1540 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1541 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1542 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1543 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1544 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1545 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1546 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1547 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1548 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1549 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1550 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1551 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1552 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1553 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1554 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1555 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1556 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1557 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1558 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1559 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1560 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1561 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1562 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1563 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1564 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1565 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1566 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1567 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1568 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1569 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1570 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1571 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1572 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1573 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1574 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1575 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1576 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1577 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1578 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1579 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1580 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1581 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1582 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1583 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1584 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1585 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1586 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1587 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1588 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1589 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1590 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1591 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1592 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1593 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1594 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1595 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1596 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1597 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1598 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1599 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1600 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1601 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1602 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1603 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1604 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1605 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1606 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1607 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1608 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1609 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1610 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1611 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1612 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1613 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1614 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1615 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1616 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1617 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1618 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1619 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1620 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1621 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1622 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1623 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1624 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1625 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1626 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1627 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1628 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1629 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1630 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1631 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1632 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1633 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1634 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1635 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1636 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1637 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1638 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1639 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1640 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1641 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1642 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1643 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1644 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1645 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1646 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1647 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1648 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1649 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1650 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1651 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1652 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1653 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1654 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1655 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1656 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1657 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1658 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1659 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1660 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1661 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1662 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1663 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1664 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1665 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1666 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1667 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1668 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1669 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1670 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1671 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1672 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1673 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1674 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1675 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1676 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1677 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1678 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1679 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1680 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1681 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1682 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1683 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1684 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1685 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1686 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1687 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1688 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1689 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1690 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1691 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1692 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1693 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1694 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1695 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1696 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1697 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1698 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1699 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1700 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1701 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1702 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1703 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1704 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1705 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1706 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1707 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1708 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1709 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1710 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1711 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1712 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1713 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1714 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1715 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1716 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1717 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1718 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1719 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1720 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1721 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1722 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1723 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1724 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1725 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1726 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1727 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1728 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1729 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1730 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1731 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1732 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1733 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1734 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1735 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1736 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1737 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1738 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1739 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1740 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1741 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1742 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1743 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1744 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1745 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1746 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1747 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1748 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1749 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1750 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1751 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1752 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1753 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1754 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1755 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1756 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1757 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1758 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1759 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1760 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1761 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1762 w_n1200_n1200# a_n50_n50# a_112_1150# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1763 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1764 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1765 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1766 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1767 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1768 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1769 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1770 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1771 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1772 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1773 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1774 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1775 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1776 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1777 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1778 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1779 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1780 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1781 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1782 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1783 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1784 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1785 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1786 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1787 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1788 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1789 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1790 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1791 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1792 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1793 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1794 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1795 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1796 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1797 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1798 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1799 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1800 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1801 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1802 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1803 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1804 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1805 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1806 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1807 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1808 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1809 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1810 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1811 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1812 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1813 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1814 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1815 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1816 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1817 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1818 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1819 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1820 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1821 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1822 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1823 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1824 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1825 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1826 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1827 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1828 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1829 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1830 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1831 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1832 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1833 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1834 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1835 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1836 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1837 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1838 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1839 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1840 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1841 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1842 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1843 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1844 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1845 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1846 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1847 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1848 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1849 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1850 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1851 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1852 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1853 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1854 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1855 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1856 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1857 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1858 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1859 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1860 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1861 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1862 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1863 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1864 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1865 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1866 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1867 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1868 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1869 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1870 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1871 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1872 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1873 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1874 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1875 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1876 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1877 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1878 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1879 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1880 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1881 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1882 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1883 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1884 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1885 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1886 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1887 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1888 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1889 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1890 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1891 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1892 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1893 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1894 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1895 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1896 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1897 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1898 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1899 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1900 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1901 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1902 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1903 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1904 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1905 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1906 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1907 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1908 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1909 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1910 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1911 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1912 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1913 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1914 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1915 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1916 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1917 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1918 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1919 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1920 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1921 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1922 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1923 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1924 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1925 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1926 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1927 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1928 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1929 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1930 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1931 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1932 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1933 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1934 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1935 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1936 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1937 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1938 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1939 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1940 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1941 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1942 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1943 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1944 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1945 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1946 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1947 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1948 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1949 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1950 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1951 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1952 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1953 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1954 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1955 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1956 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1957 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1958 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1959 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1960 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1961 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1962 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1963 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1964 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1965 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1966 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1967 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1968 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1969 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1970 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1971 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1972 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1973 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1974 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1975 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1976 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1977 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1978 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1979 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1980 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1981 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1982 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1983 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1984 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1985 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1986 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1987 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1988 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1989 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1990 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1991 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1992 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1993 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1994 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1995 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1996 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1997 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1998 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1999 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2000 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2001 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2002 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2003 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2004 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2005 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2006 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2007 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2008 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2009 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2010 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2011 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2012 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2013 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2014 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2015 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2016 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2017 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2018 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2019 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2020 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2021 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2022 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2023 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2024 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2025 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2026 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2027 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2028 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2029 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2030 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2031 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2032 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2033 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2034 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2035 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2036 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2037 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2038 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2039 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2040 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2041 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2042 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2043 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2044 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2045 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2046 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2047 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2048 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2049 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2050 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2051 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2052 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2053 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2054 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2055 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2056 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2057 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2058 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2059 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2060 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2061 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2062 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2063 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2064 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2065 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2066 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2067 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2068 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2069 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2070 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2071 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2072 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2073 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2074 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2075 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2076 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2077 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2078 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2079 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2080 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2081 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2082 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2083 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2084 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2085 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2086 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2087 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2088 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2089 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2090 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2091 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2092 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2093 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2094 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2095 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2096 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2097 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2098 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2099 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2100 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2101 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2102 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2103 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2104 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2105 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2106 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2107 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2108 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2109 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2110 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2111 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2112 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2113 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2114 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2115 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2116 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2117 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2118 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2119 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2120 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2121 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2122 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2123 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2124 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2125 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2126 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2127 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2128 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2129 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2130 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2131 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2132 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2133 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2134 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2135 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2136 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2137 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2138 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2139 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2140 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2141 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2142 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2143 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2144 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2145 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2146 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2147 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2148 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2149 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2150 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2151 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2152 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2153 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2154 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2155 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2156 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2157 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2158 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2159 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2160 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2161 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2162 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2163 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2164 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2165 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2166 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2167 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2168 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2169 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2170 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2171 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2172 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2173 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2174 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2175 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2176 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2177 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2178 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2179 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2180 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2181 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2182 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2183 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2184 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2185 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2186 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2187 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2188 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2189 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2190 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2191 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2192 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2193 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2194 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2195 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2196 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2197 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2198 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2199 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2200 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2201 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2202 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2203 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2204 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2205 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2206 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2207 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2208 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2209 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2210 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2211 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2212 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2213 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2214 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2215 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2216 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2217 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2218 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2219 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2220 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2221 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2222 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2223 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2224 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2225 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2226 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2227 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2228 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2229 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2230 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2231 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2232 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2233 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2234 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2235 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2236 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2237 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2238 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2239 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2240 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2241 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2242 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2243 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2244 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2245 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2246 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2247 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2248 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2249 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2250 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2251 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2252 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2253 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2254 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2255 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2256 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2257 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2258 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2259 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2260 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2261 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2262 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2263 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2264 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2265 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2266 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2267 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2268 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2269 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2270 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2271 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2272 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2273 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2274 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2275 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2276 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2277 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2278 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2279 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2280 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2281 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2282 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2283 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2284 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2285 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2286 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2287 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2288 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2289 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2290 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2291 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2292 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2293 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2294 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2295 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2296 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2297 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2298 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2299 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2300 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2301 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2302 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2303 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2304 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2305 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2306 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2307 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2308 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2309 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2310 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2311 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2312 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2313 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2314 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2315 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2316 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2317 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2318 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2319 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2320 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2321 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2322 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2323 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2324 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2325 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2326 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2327 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2328 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2329 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2330 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2331 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2332 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2333 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2334 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2335 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2336 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2337 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2338 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2339 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2340 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2341 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2342 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2343 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2344 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2345 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2346 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2347 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2348 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2349 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2350 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2351 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2352 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2353 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2354 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2355 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2356 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2357 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2358 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2359 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2360 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2361 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2362 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2363 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2364 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2365 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2366 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2367 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2368 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2369 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2370 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2371 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2372 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2373 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2374 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2375 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2376 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2377 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2378 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2379 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2380 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2381 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2382 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2383 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2384 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2385 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2386 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2387 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2388 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2389 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2390 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2391 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2392 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2393 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2394 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2395 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2396 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2397 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2398 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2399 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2400 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2401 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2402 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2403 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2404 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2405 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2406 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2407 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2408 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2409 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2410 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2411 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2412 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2413 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2414 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2415 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2416 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2417 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2418 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2419 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2420 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2421 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2422 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2423 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2424 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2425 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2426 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2427 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2428 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2429 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2430 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2431 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2432 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2433 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2434 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2435 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2436 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2437 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2438 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2439 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2440 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2441 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2442 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2443 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2444 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2445 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2446 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2447 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2448 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2449 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2450 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2451 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2452 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2453 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2454 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2455 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2456 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2457 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2458 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2459 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2460 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2461 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2462 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2463 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2464 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2465 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2466 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2467 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2468 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2469 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2470 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2471 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2472 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2473 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2474 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2475 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2476 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2477 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2478 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2479 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2480 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2481 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2482 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2483 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2484 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2485 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2486 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2487 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2488 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2489 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2490 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2491 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2492 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2493 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2494 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2495 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2496 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2497 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2498 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2499 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2500 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2501 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2502 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2503 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2504 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2505 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2506 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2507 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2508 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2509 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2510 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2511 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2512 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2513 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2514 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2515 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2516 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2517 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2518 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2519 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2520 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2521 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2522 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2523 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2524 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2525 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2526 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2527 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2528 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2529 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2530 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2531 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2532 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2533 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2534 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2535 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2536 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2537 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2538 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2539 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2540 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2541 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2542 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2543 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2544 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2545 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2546 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2547 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2548 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2549 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2550 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2551 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2552 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2553 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2554 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2555 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2556 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2557 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2558 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2559 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2560 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2561 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2562 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2563 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2564 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2565 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2566 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2567 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2568 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2569 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2570 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2571 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2572 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2573 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2574 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2575 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2576 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2577 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2578 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2579 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2580 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2581 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2582 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2583 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2584 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2585 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2586 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2587 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2588 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2589 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2590 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2591 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2592 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2593 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2594 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2595 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2596 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2597 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2598 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2599 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2600 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2601 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2602 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2603 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2604 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2605 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2606 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2607 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2608 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2609 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2610 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2611 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2612 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2613 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2614 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2615 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2616 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2617 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2618 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2619 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2620 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2621 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2622 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2623 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2624 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2625 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2626 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2627 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2628 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2629 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2630 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2631 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2632 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2633 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2634 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2635 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2636 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2637 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2638 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2639 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2640 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2641 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2642 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2643 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2644 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2645 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2646 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2647 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2648 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2649 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2650 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2651 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2652 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2653 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2654 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2655 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2656 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2657 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2658 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2659 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2660 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2661 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2662 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2663 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2664 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2665 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2666 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2667 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2668 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2669 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2670 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2671 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2672 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2673 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2674 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2675 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2676 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2677 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2678 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2679 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2680 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2681 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2682 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2683 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2684 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2685 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2686 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2687 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2688 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2689 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2690 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2691 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2692 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2693 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2694 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2695 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2696 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2697 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2698 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2699 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2700 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2701 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2702 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2703 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2704 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2705 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2706 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2707 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2708 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2709 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2710 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2711 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2712 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2713 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2714 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2715 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2716 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2717 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2718 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2719 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2720 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2721 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2722 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2723 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2724 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2725 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2726 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2727 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2728 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2729 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2730 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2731 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2732 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2733 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2734 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2735 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2736 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2737 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2738 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2739 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2740 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2741 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2742 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2743 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2744 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2745 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2746 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2747 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2748 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2749 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2750 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2751 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2752 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2753 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2754 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2755 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2756 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2757 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2758 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2759 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2760 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2761 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2762 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2763 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2764 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2765 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2766 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2767 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2768 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2769 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2770 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2771 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2772 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2773 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2774 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2775 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2776 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2777 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2778 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2779 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2780 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2781 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2782 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2783 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2784 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2785 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2786 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2787 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2788 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2789 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2790 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2791 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2792 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2793 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2794 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2795 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2796 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2797 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2798 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2799 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2800 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2801 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2802 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2803 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2804 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2805 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2806 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2807 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2808 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2809 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2810 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2811 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2812 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2813 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2814 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2815 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2816 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2817 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2818 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2819 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2820 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2821 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2822 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2823 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2824 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2825 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2826 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2827 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2828 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2829 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2830 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2831 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2832 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2833 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2834 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2835 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2836 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2837 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2838 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2839 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2840 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2841 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2842 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2843 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2844 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2845 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2846 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2847 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2848 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2849 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2850 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2851 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2852 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2853 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2854 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2855 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2856 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2857 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2858 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2859 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2860 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2861 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2862 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2863 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2864 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2865 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2866 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2867 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2868 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2869 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2870 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2871 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2872 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2873 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2874 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2875 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2876 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2877 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2878 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2879 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2880 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2881 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2882 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2883 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2884 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2885 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2886 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2887 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2888 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2889 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2890 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2891 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2892 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2893 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2894 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2895 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2896 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2897 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2898 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2899 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2900 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2901 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2902 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2903 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2904 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2905 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2906 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2907 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2908 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2909 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2910 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2911 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2912 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2913 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2914 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2915 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2916 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2917 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2918 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2919 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2920 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2921 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2922 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2923 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2924 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2925 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2926 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2927 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2928 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2929 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2930 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2931 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2932 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2933 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2934 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2935 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2936 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2937 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2938 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2939 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2940 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2941 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2942 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2943 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2944 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2945 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2946 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2947 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2948 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2949 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2950 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2951 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2952 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2953 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2954 w_n1200_n1200# a_n50_n50# a_112_1150# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2955 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2956 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2957 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2958 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2959 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2960 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2961 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2962 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2963 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2964 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2965 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2966 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2967 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2968 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2969 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2970 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2971 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2972 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2973 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2974 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2975 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2976 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2977 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2978 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2979 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2980 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2981 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2982 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2983 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2984 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2985 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2986 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2987 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2988 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2989 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2990 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2991 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2992 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2993 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2994 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2995 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2996 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2997 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2998 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2999 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3000 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3001 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3002 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3003 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3004 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3005 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3006 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3007 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3008 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3009 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3010 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3011 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3012 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3013 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3014 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3015 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3016 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3017 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3018 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3019 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3020 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3021 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3022 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3023 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3024 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3025 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3026 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3027 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3028 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3029 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3030 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3031 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3032 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3033 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3034 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3035 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3036 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3037 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3038 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3039 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3040 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3041 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3042 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3043 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3044 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3045 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3046 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3047 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3048 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3049 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3050 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3051 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3052 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3053 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3054 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3055 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3056 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3057 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3058 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3059 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3060 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3061 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3062 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3063 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3064 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3065 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3066 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3067 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3068 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3069 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3070 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3071 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3072 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3073 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3074 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3075 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3076 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3077 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3078 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3079 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3080 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3081 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3082 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3083 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3084 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3085 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3086 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3087 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3088 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3089 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3090 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3091 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3092 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3093 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3094 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3095 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3096 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3097 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3098 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3099 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3100 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3101 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3102 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3103 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3104 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3105 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3106 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3107 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3108 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3109 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3110 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3111 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3112 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3113 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3114 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3115 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3116 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3117 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3118 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3119 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3120 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3121 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3122 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3123 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3124 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3125 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3126 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3127 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3128 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3129 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3130 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3131 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3132 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3133 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3134 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3135 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3136 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3137 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3138 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3139 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3140 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3141 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3142 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3143 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3144 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3145 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3146 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3147 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3148 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3149 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3150 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3151 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3152 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3153 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3154 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3155 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3156 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3157 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3158 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3159 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3160 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3161 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3162 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3163 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3164 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3165 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3166 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3167 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3168 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3169 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3170 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3171 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3172 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3173 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3174 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3175 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3176 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3177 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3178 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3179 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3180 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3181 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3182 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3183 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3184 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3185 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3186 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3187 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3188 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3189 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3190 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3191 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3192 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3193 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3194 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3195 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3196 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3197 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3198 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3199 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3200 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3201 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3202 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3203 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3204 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3205 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3206 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3207 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3208 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3209 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3210 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3211 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3212 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3213 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3214 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3215 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3216 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3217 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3218 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3219 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3220 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3221 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3222 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3223 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3224 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3225 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3226 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3227 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3228 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3229 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3230 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3231 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3232 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3233 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3234 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3235 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3236 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3237 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3238 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3239 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3240 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3241 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3242 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3243 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3244 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3245 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3246 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3247 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3248 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3249 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3250 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3251 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3252 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3253 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3254 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3255 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3256 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3257 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3258 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3259 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3260 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3261 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3262 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3263 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3264 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3265 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3266 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3267 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3268 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3269 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3270 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3271 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3272 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3273 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3274 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3275 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3276 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3277 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3278 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3279 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3280 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3281 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3282 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3283 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3284 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3285 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3286 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3287 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3288 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3289 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3290 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3291 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3292 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3293 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3294 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3295 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3296 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3297 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3298 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3299 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3300 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3301 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3302 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3303 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3304 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3305 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3306 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3307 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3308 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3309 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3310 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3311 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3312 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3313 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3314 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3315 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3316 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3317 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3318 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3319 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3320 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3321 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3322 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3323 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3324 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3325 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3326 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3327 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3328 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3329 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3330 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3331 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3332 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3333 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3334 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3335 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3336 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3337 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3338 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3339 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3340 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3341 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3342 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3343 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3344 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3345 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3346 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3347 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3348 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3349 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3350 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3351 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3352 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3353 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3354 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3355 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3356 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3357 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3358 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3359 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3360 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3361 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3362 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3363 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3364 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3365 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3366 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3367 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3368 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3369 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3370 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3371 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3372 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3373 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3374 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3375 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3376 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3377 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3378 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3379 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3380 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3381 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3382 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3383 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3384 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3385 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3386 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3387 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3388 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3389 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3390 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3391 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3392 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3393 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3394 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3395 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3396 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3397 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3398 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3399 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3400 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3401 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3402 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3403 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3404 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3405 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3406 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3407 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3408 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3409 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3410 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3411 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3412 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3413 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3414 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3415 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3416 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3417 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3418 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3419 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3420 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3421 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3422 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3423 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3424 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3425 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3426 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3427 a_112_1150# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3428 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3429 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3430 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3431 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3432 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3433 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3434 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3435 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3436 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3437 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3438 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3439 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3440 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3441 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3442 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3443 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3444 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3445 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3446 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3447 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3448 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3449 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3450 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3451 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3452 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3453 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3454 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3455 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3456 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3457 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3458 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3459 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3460 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3461 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3462 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3463 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3464 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3465 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3466 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3467 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3468 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3469 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3470 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3471 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3472 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3473 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3474 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3475 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3476 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3477 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3478 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3479 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3480 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3481 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3482 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3483 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3484 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3485 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3486 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3487 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3488 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3489 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3490 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3491 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3492 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3493 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3494 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3495 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3496 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3497 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3498 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3499 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3500 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3501 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3502 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3503 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3504 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3505 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3506 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3507 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3508 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3509 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3510 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3511 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3512 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3513 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3514 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3515 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3516 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3517 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3518 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3519 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3520 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3521 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3522 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3523 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3524 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3525 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3526 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3527 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3528 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3529 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3530 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3531 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3532 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3533 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3534 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3535 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3536 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3537 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3538 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3539 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3540 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3541 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3542 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3543 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3544 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3545 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3546 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3547 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3548 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3549 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3550 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3551 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3552 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3553 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3554 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3555 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3556 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3557 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3558 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3559 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3560 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3561 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3562 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3563 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3564 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3565 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3566 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3567 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3568 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3569 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3570 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3571 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3572 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3573 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3574 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3575 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3576 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3577 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3578 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3579 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3580 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3581 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3582 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3583 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3584 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3585 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3586 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3587 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3588 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3589 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3590 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3591 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3592 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3593 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3594 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3595 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3596 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3597 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3598 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3599 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3600 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3601 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3602 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3603 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3604 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3605 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3606 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3607 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3608 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3609 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3610 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3611 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3612 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3613 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3614 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3615 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3616 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3617 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3618 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3619 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3620 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3621 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3622 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3623 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3624 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3625 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3626 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3627 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3628 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3629 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3630 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3631 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3632 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3633 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3634 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3635 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3636 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3637 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3638 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3639 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3640 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3641 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3642 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3643 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3644 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3645 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3646 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3647 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3648 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3649 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3650 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3651 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3652 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3653 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3654 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3655 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3656 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3657 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3658 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3659 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3660 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3661 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3662 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3663 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3664 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3665 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3666 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3667 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3668 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3669 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3670 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3671 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3672 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3673 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3674 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3675 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3676 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3677 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3678 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3679 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3680 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3681 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3682 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3683 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3684 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3685 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3686 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3687 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3688 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3689 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3690 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3691 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3692 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3693 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3694 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3695 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3696 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3697 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3698 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3699 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3700 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3701 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3702 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3703 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3704 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3705 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3706 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3707 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3708 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3709 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3710 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3711 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3712 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3713 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3714 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3715 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3716 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3717 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3718 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3719 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3720 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3721 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3722 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3723 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3724 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3725 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3726 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3727 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3728 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3729 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3730 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3731 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3732 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3733 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3734 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3735 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3736 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3737 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3738 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3739 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3740 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3741 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3742 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3743 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3744 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3745 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3746 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3747 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3748 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3749 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3750 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3751 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3752 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3753 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3754 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3755 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3756 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3757 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3758 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3759 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3760 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3761 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3762 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3763 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3764 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3765 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3766 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3767 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3768 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3769 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3770 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3771 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3772 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3773 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3774 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3775 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3776 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3777 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3778 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3779 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3780 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3781 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3782 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3783 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3784 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3785 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3786 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3787 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3788 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3789 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3790 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3791 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3792 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3793 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3794 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3795 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3796 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3797 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3798 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3799 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3800 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3801 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3802 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3803 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3804 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3805 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3806 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3807 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3808 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3809 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3810 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3811 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3812 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3813 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3814 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3815 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3816 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3817 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3818 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3819 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3820 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3821 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3822 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3823 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3824 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3825 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3826 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3827 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3828 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3829 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3830 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3831 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3832 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3833 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3834 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3835 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3836 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3837 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3838 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3839 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3840 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3841 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3842 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3843 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3844 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3845 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3846 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3847 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3848 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3849 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3850 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3851 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3852 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3853 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3854 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3855 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3856 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3857 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3858 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3859 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3860 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3861 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3862 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3863 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3864 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3865 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3866 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3867 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3868 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3869 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3870 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3871 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3872 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3873 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3874 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3875 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3876 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3877 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3878 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3879 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3880 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3881 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3882 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3883 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3884 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3885 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3886 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3887 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3888 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3889 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3890 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3891 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3892 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3893 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3894 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3895 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3896 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3897 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3898 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3899 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3900 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3901 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3902 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3903 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3904 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3905 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3906 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3907 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3908 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3909 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3910 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3911 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3912 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3913 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3914 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3915 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3916 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3917 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3918 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3919 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3920 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3921 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3922 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3923 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3924 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3925 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3926 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3927 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3928 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3929 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3930 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3931 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3932 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3933 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3934 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3935 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3936 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3937 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3938 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3939 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3940 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3941 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3942 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3943 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3944 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3945 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3946 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3947 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3948 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3949 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3950 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3951 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3952 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3953 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3954 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3955 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3956 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3957 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3958 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3959 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3960 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3961 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3962 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3963 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3964 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3965 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3966 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3967 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3968 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3969 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3970 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3971 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3972 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3973 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3974 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3975 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3976 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3977 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3978 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3979 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3980 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3981 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3982 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3983 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3984 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3985 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3986 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3987 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3988 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3989 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3990 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3991 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3992 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3993 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3994 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3995 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3996 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3997 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3998 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3999 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4000 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4001 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4002 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4003 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4004 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4005 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4006 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4007 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4008 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4009 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4010 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4011 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4012 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4013 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4014 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4015 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4016 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4017 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4018 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4019 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4020 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4021 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4022 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4023 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4024 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4025 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4026 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4027 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4028 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4029 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4030 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4031 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4032 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4033 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4034 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4035 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4036 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4037 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4038 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4039 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4040 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4041 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4042 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4043 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4044 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4045 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4046 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4047 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4048 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4049 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4050 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4051 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4052 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4053 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4054 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4055 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4056 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4057 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4058 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4059 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4060 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4061 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4062 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4063 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4064 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4065 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4066 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4067 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4068 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4069 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4070 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4071 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4072 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4073 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4074 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4075 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4076 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4077 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4078 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4079 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4080 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4081 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4082 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4083 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4084 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4085 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4086 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4087 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4088 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4089 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4090 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4091 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4092 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4093 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4094 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4095 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4096 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4097 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4098 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4099 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4100 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4101 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4102 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4103 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4104 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4105 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4106 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4107 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4108 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4109 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4110 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4111 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4112 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4113 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4114 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4115 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4116 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4117 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4118 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4119 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4120 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4121 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4122 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4123 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4124 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4125 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4126 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4127 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4128 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4129 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4130 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4131 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4132 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4133 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4134 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4135 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4136 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4137 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4138 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4139 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4140 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4141 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4142 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4143 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4144 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4145 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4146 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4147 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4148 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4149 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4150 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4151 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4152 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4153 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4154 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4155 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4156 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4157 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4158 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4159 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4160 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4161 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4162 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4163 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4164 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4165 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4166 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4167 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4168 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4169 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4170 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4171 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4172 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4173 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4174 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4175 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4176 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4177 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4178 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4179 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4180 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4181 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4182 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4183 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4184 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4185 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4186 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4187 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4188 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4189 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4190 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4191 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4192 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4193 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4194 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4195 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4196 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4197 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4198 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4199 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4200 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4201 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4202 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4203 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4204 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4205 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4206 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4207 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4208 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4209 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4210 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4211 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4212 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4213 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4214 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4215 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4216 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4217 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4218 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4219 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4220 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4221 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4222 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4223 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4224 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4225 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4226 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4227 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4228 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4229 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4230 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4231 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4232 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4233 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4234 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4235 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4236 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4237 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4238 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4239 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4240 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4241 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4242 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4243 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4244 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4245 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4246 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4247 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4248 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4249 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4250 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4251 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4252 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4253 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4254 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4255 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4256 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4257 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4258 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4259 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4260 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4261 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4262 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4263 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4264 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4265 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4266 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4267 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4268 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4269 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4270 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4271 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4272 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4273 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4274 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4275 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4276 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4277 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4278 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4279 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4280 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4281 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4282 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4283 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4284 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4285 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4286 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4287 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4288 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4289 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4290 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4291 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4292 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4293 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4294 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4295 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4296 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4297 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4298 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4299 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4300 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4301 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4302 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4303 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4304 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4305 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4306 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4307 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4308 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4309 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4310 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4311 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4312 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4313 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4314 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4315 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4316 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4317 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4318 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4319 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4320 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4321 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4322 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4323 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4324 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4325 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4326 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4327 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4328 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4329 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4330 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4331 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4332 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4333 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4334 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4335 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4336 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4337 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4338 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4339 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4340 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4341 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4342 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4343 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4344 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4345 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4346 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4347 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4348 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4349 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4350 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4351 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4352 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4353 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4354 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4355 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4356 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4357 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4358 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4359 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4360 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4361 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4362 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4363 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4364 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4365 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4366 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4367 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4368 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4369 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4370 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4371 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4372 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4373 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4374 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4375 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4376 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4377 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4378 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4379 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4380 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4381 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4382 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4383 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4384 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4385 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4386 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4387 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4388 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4389 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4390 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4391 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4392 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4393 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4394 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4395 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4396 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4397 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4398 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4399 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4400 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4401 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4402 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4403 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4404 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4405 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4406 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4407 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4408 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4409 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4410 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4411 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4412 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4413 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4414 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4415 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4416 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4417 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4418 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4419 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4420 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4421 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4422 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4423 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4424 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4425 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4426 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4427 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4428 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4429 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4430 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4431 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4432 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4433 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4434 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4435 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4436 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4437 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4438 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4439 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4440 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4441 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4442 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4443 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4444 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4445 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4446 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4447 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4448 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4449 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4450 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4451 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4452 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4453 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4454 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4455 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4456 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4457 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4458 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4459 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4460 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4461 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4462 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4463 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4464 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4465 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4466 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4467 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4468 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4469 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4470 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4471 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4472 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4473 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4474 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4475 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4476 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4477 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4478 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4479 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4480 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4481 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4482 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4483 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4484 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4485 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4486 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4487 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4488 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4489 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4490 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4491 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4492 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4493 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4494 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4495 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4496 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4497 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4498 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4499 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4500 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4501 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4502 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4503 a_112_1150# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4504 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4505 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4506 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4507 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4508 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4509 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4510 w_n1200_n1200# a_n50_n50# a_112_3350# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4511 a_112_3350# a_n50_n50# w_n1200_n1200# w_n1200_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
.ends

.subckt power_stage fc2 VN fc1
Xnmos_waffle_36x36_0 VN s4 fc2 fc2 nmos_waffle_36x36
Xnmos_waffle_36x36_1 fc2 s3 out out nmos_waffle_36x36
Xpmos_waffle_48x48_0 fc1 s2 out out pmos_waffle_48x48
Xpmos_waffle_48x48_1 VP s1 fc1 fc1 pmos_waffle_48x48
.ends

.subckt unit_cap c2_30_30# c1_30_30# m3_0_0#
X0 c1_30_30# m3_0_0# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X1 c2_30_30# c1_30_30# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
.ends

.subckt flying_cap m3_142420_294000# m3_2060_293480#
Xunit_cap_360 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_371 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_382 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_393 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1005 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1049 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1016 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1027 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1038 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1561 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1572 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1583 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1594 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1550 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_190 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1380 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1391 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_915 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_959 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_926 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_937 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_948 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_904 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_701 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_734 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_778 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_40 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_84 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_789 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_51 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_95 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_745 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_62 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_756 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_712 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_73 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_767 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_723 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1924 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1968 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1935 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1946 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1902 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1957 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1913 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_542 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_553 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_520 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_531 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_597 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_564 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_575 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_586 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1209 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1710 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1743 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1787 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1754 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1798 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1765 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1721 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1776 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1732 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_361 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_372 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_383 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_394 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_350 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1006 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1017 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1028 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1039 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1562 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1540 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1551 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1573 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1584 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1595 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_180 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_191 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1370 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1381 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1392 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_916 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_927 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_938 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_949 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_905 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_735 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_41 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_52 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_702 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_713 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_30 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_724 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_779 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_85 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_96 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_746 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_63 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_757 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_74 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_768 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1903 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1925 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1969 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1936 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1947 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1958 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1914 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_543 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_510 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_554 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_565 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_521 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_576 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_532 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_587 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_598 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1700 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1744 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1711 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1722 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1733 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1788 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1755 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1799 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1766 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1777 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_362 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_373 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_384 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_340 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_395 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_351 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1007 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1018 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1029 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1563 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1574 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1530 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1585 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1541 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1596 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1552 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_181 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_192 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_170 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1371 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1382 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1393 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1360 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_917 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_906 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_928 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_939 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1190 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_42 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_86 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_53 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_736 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_747 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_703 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_64 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_20 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_758 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_714 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_75 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_31 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_769 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_725 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_97 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1926 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1937 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1904 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1915 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1948 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1959 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_500 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_544 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_588 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_511 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_555 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_599 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_566 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_522 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_577 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_533 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1701 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1745 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1756 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1712 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1767 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1723 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1778 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1734 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1789 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_363 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_330 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_374 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_385 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_341 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_396 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_352 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1008 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1019 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1553 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1520 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1564 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1575 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1531 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1586 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1542 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1597 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_160 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_182 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_193 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_171 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1372 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1383 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1394 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1350 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1361 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_918 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_929 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_907 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1191 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1180 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_43 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_87 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_726 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_54 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_98 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_737 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_10 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_748 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_704 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_65 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_21 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_759 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_715 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_76 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_32 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1927 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1938 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1949 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1905 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1916 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_501 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_545 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_589 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_512 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_556 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_567 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_523 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_578 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_534 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1746 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1702 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1757 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1713 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1768 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1724 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1779 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1735 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_320 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_331 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_342 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_364 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_375 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_386 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_397 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_353 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1009 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1510 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1554 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1521 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1565 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1576 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1532 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1587 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1543 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1598 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_183 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_194 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_150 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_161 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_172 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1340 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1351 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1362 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1373 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1384 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1395 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_919 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_908 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1192 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1170 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1181 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_11 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_44 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_88 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_727 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_99 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_738 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_55 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_749 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_705 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_66 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_22 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_716 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_77 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_33 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1928 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1939 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1906 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1917 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_502 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_513 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_524 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_535 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_546 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_557 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_568 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_579 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1747 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1703 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1758 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1714 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1769 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1725 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1736 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_321 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_365 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_376 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_332 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_343 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_354 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_310 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_387 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_398 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1511 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1522 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1533 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1544 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1500 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1555 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1599 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1566 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1577 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1588 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_184 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_140 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_195 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_151 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_162 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_173 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1330 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1374 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1341 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1385 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1352 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1363 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1396 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_909 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1193 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1160 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1171 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1182 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_12 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_706 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_23 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_717 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_34 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_45 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_89 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_728 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_739 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_56 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_67 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_78 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1929 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1907 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1918 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_503 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_547 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_514 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_558 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_569 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_525 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_536 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1704 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1715 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1726 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1737 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1748 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1759 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_366 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_322 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_377 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_333 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_388 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_344 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_300 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_399 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_355 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_311 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1512 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1556 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1523 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1567 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1578 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1534 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1545 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1501 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1589 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_130 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_174 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_141 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_185 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_196 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_152 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_163 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1331 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1375 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1342 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1386 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1397 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1353 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1364 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1320 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1194 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1150 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1161 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1172 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1183 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_729 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_46 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_57 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_13 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_707 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_68 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_24 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_718 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_35 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_79 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1908 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1919 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_504 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_548 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_559 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_515 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_526 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_537 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1738 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1705 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1749 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1716 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1727 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_301 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_367 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_312 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_323 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_378 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_334 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_389 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_345 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_356 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_890 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1513 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1557 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1524 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1568 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1579 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1535 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1546 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1502 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_131 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_142 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_120 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_175 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_186 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_197 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_153 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_164 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1310 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1332 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1376 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1387 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1343 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1398 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1354 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1365 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1321 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1140 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1151 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1195 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1162 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1173 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1184 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_36 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_47 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_58 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_14 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_708 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_69 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_25 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_719 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1909 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_505 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_549 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_516 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_527 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_538 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1739 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1706 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1717 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1728 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_313 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_324 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_302 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_368 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_379 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_335 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_346 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_357 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_880 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_891 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1514 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1558 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1525 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1569 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1536 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1547 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1503 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_132 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_176 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_143 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_154 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_110 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_165 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_121 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_187 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_198 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1333 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1344 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1300 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1311 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1322 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1377 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1388 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1399 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1355 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1366 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1141 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1152 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1163 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1174 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1130 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1185 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1196 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_37 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_48 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_59 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_15 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_709 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_26 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_506 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_517 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_528 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_539 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1707 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1718 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1729 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_314 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_358 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_325 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_336 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_347 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_303 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_369 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_870 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_881 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_892 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1515 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1526 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1504 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1559 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1537 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1548 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_133 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_177 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_100 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_144 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_188 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_199 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_155 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_111 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_166 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_122 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1334 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1345 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1301 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1356 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1312 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1367 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1323 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1378 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1389 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1890 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1142 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1186 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1153 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1197 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1164 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1120 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1175 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1131 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_16 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_38 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_49 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_27 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_507 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_518 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_529 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1708 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1719 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_315 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_359 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_326 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_337 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_348 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_304 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_871 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_882 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_893 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_860 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1516 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1527 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1538 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1549 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1505 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_134 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_178 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_145 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_189 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_101 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_156 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_112 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_167 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_123 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_690 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1379 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1324 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1335 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1346 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1302 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1357 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1313 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1368 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1880 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1891 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1110 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1143 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1187 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1154 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1198 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1165 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1121 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1176 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1132 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_39 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_17 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_28 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_508 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_519 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1709 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_316 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_327 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_338 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_349 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_305 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_872 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_883 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_894 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_850 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_861 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1517 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1528 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1539 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1506 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_102 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_113 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_124 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_135 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_179 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_146 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_157 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_168 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_680 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_691 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1325 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1336 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1347 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1303 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1358 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1314 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1369 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1881 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1892 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1870 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1100 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1111 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1122 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1133 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1144 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1188 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1155 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1199 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1166 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1177 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_18 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_29 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_509 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_306 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_317 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_328 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_339 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_840 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_851 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_862 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_873 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_884 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_895 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1507 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1518 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1529 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_136 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_147 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_103 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_158 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_114 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_125 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_169 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_681 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_692 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_670 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1326 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1304 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1315 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1337 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1348 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1359 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1860 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1871 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1882 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1893 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1101 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1145 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1112 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1156 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1167 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1123 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1134 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1189 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1178 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1690 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_19 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_318 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_329 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_307 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_830 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_874 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_885 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_841 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_896 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_852 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_863 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1508 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1519 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_137 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_148 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_104 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_159 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_115 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_126 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_682 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_693 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_660 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_671 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1327 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1338 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1349 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1305 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1316 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1883 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1894 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1850 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1861 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1872 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_490 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1102 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1146 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1157 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1113 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1168 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1124 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1179 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1135 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1691 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1680 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_319 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_308 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_820 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_864 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_831 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_875 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_886 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_842 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_897 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_853 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1509 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_138 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_149 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_105 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_116 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_127 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_683 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_650 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_694 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_661 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_672 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1328 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1339 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1306 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1317 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1884 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1840 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1895 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1851 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1862 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1873 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_480 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_491 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1103 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1147 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1158 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1114 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1169 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1125 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1136 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1692 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1670 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1681 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_309 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_810 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_821 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_865 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_832 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_876 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_887 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_843 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_898 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_854 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_106 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_128 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_139 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_117 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_640 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_651 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_662 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_684 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_695 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_673 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1329 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1307 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1318 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1830 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1885 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1841 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1896 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1852 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1863 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1874 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_470 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_481 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_492 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1104 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1115 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1148 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1159 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1126 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1137 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1660 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1671 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1693 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1682 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1490 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_822 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_833 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_844 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_800 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_811 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_866 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_877 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_888 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_899 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_855 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_129 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_107 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_118 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_0 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_641 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_685 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_652 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_696 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_663 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_674 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_630 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1308 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1319 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1831 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1842 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1853 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1820 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1875 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1886 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1897 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1864 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_460 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_471 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_482 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_493 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1149 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1105 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1116 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1127 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1138 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1650 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1694 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1661 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1672 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1683 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_290 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1480 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1491 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_823 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_867 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_834 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_878 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_845 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_801 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_856 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_812 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_889 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_108 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_119 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_642 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_686 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_697 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_653 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_664 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_620 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_675 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_631 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1309 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1832 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1876 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1843 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1887 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1854 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1810 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1865 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1821 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1898 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_450 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_461 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_472 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_483 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_494 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1106 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1117 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1128 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1139 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1651 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1695 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1662 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1673 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1684 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1640 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_280 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_291 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1470 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1481 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1492 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_824 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_868 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_835 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_879 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_846 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_802 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_857 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_813 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_109 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_2 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_610 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_643 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_687 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_698 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_654 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_665 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_621 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_676 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_632 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1833 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1877 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1800 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1844 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1888 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1899 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1855 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1811 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1866 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1822 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_451 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_462 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_440 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_473 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_484 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_495 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1107 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1118 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1129 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1652 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1696 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1663 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1674 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1630 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1685 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1641 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_270 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_281 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_292 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1471 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1460 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1482 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1493 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1290 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_825 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_869 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_836 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_847 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_803 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_858 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_814 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_3 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_600 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_644 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_611 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_622 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_633 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_688 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_699 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_655 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_666 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_677 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1801 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1812 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1834 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1878 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1845 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1889 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1856 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1867 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1823 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_452 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_463 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_474 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_430 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_485 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_441 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_496 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1108 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1119 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1653 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1620 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1631 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1642 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1697 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1664 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1675 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1686 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_271 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_282 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_293 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_260 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1461 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1472 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1483 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1494 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1450 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1280 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1291 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_826 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_804 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_815 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_837 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_848 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_859 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_4 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_634 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_601 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_645 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_656 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_612 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_667 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_623 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_678 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_689 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1835 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1802 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1813 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1824 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1879 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1846 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1857 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1868 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_453 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_497 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_420 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_464 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_475 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_431 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_486 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_442 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1109 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1654 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1610 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1665 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1621 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1676 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1632 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1687 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1643 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1698 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_272 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_283 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_294 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_250 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_261 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1462 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1473 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1484 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1440 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1495 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1451 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1281 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1292 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1270 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_827 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_838 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_849 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_805 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_816 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_5 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_635 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_602 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_646 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_657 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_613 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_668 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_624 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_679 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1836 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1847 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1803 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1858 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1814 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1869 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1825 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_410 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_454 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_498 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_421 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_465 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_476 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_432 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_487 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_443 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1655 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1699 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1600 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1611 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1666 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1622 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1677 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1633 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1688 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1644 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_240 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_251 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_273 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_284 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_295 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_262 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1463 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1430 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1474 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1485 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1441 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1496 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1452 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1260 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1271 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1282 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1293 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_828 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_839 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_806 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_817 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1090 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_6 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_636 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_603 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_647 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_658 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_614 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_669 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_625 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1837 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1848 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1804 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1859 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1815 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1826 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_411 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_422 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_433 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_444 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_400 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_455 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_499 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_466 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_477 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_488 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1601 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1645 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1612 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1656 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1667 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1623 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1678 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1634 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1689 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_274 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_230 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_285 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_241 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_252 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_263 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_296 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1420 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1431 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1442 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1453 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1464 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1475 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1486 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1497 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1283 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1250 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1294 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1261 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1272 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_818 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_829 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_807 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1080 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1091 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_7 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_604 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_615 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_626 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_637 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_648 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_659 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1838 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1849 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1805 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1816 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1827 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_412 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_456 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_467 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_423 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_434 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_445 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_401 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_478 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_489 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_990 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1602 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1613 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1624 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1635 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1646 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1657 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1668 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1679 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_275 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_220 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_231 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_286 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_242 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_297 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_253 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_264 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1421 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1465 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1432 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1476 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1487 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1443 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1454 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1410 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1498 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1240 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1284 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1295 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1251 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1262 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1273 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_808 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_819 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1070 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1081 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1092 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_8 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_638 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_605 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_649 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_616 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_627 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1806 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1817 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1839 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1828 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_413 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_457 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_468 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_424 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_479 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_435 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_446 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_402 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_980 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_991 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1603 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1647 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1614 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1658 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1669 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1625 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1636 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_221 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_276 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_232 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_287 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_243 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_298 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_254 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_210 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_265 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1422 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1466 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1433 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1477 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1488 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1444 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1400 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1499 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1455 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1411 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1241 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1285 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1296 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1252 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1263 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1274 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1230 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_809 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1060 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1071 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1082 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1093 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_9 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_639 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_606 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_617 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_628 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1829 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1807 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1818 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_458 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_414 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_469 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_425 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_436 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_447 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_403 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_970 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_981 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_992 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1604 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1648 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1615 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1659 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1626 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1637 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_222 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_233 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_200 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_211 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_266 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_277 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_288 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_244 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_299 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_255 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1401 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1423 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1467 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1434 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1478 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1489 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1445 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1456 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1412 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1242 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1253 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1220 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1231 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1286 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1297 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1264 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1275 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1050 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1094 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1061 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1072 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1083 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_607 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_618 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_629 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1808 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1819 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_404 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_415 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_426 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_459 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_437 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_448 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_960 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_971 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_982 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_993 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1605 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1649 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1616 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1627 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1638 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_223 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_267 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_234 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_245 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_201 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_256 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_212 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_278 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_289 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_790 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1424 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1435 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1402 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1413 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1468 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1479 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1446 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1457 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1232 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1243 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1254 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1210 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1265 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1221 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1276 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1287 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1298 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1051 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1095 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1062 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1073 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1084 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1040 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_608 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_619 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1809 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_405 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_416 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_427 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_438 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_449 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_961 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_972 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_983 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_994 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_950 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1606 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1617 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1628 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1639 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_224 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_268 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_235 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_279 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_246 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_202 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_257 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_213 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_780 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_791 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1425 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1469 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1436 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1447 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1403 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1458 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1414 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1970 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1233 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1200 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1244 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1288 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1299 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1255 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1211 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1266 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1222 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1277 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1052 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1096 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1063 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1074 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1030 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1085 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1041 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_609 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_406 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_417 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_428 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_439 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_962 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_973 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_984 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_940 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_995 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_951 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1607 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1618 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1629 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_225 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_269 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_236 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_247 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_203 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_258 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_214 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_781 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_792 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_770 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1426 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1437 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1448 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1404 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1459 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1415 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1971 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1960 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1201 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1234 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1278 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1245 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1289 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1256 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1212 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1267 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1223 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1790 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1020 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1031 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1042 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1053 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1097 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1064 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1075 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1086 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_407 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_418 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_429 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_930 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_963 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_974 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_985 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_941 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_996 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_952 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1608 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1619 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_204 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_215 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_226 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_237 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_248 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_259 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_760 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_771 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_782 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_793 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1416 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1427 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1438 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1449 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1405 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1972 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1950 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1961 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_590 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1202 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1213 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1224 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1235 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1279 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1246 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1257 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1268 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1780 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1791 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1010 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1054 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1065 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1021 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1076 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1032 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1043 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1098 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1087 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_408 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_419 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_920 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_931 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_942 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_953 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_964 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_975 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_986 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_997 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1609 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_227 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_238 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_249 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_205 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_216 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_772 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_783 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_794 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_750 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_761 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1417 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1406 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1428 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1439 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1973 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1940 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1951 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1962 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_591 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_580 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1236 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1203 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1247 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1258 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1214 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1225 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1269 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1792 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1770 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1781 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1011 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1055 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1099 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1066 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1022 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1077 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1033 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1088 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1044 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1000 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_409 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_965 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_910 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_921 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_976 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_932 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_987 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_943 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_954 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_998 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_228 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_239 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_206 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_217 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_90 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_773 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_740 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_784 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_795 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_751 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_762 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1418 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1429 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1407 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1930 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1974 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1941 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1952 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1963 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_592 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_570 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_581 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1237 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1204 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1248 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1259 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1215 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1226 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1793 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1760 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1771 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1782 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1056 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1012 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1067 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1023 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1078 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1034 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1089 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1045 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1001 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1590 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_911 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_922 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_966 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_977 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_933 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_988 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_944 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_900 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_999 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_955 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_229 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_207 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_218 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_91 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_730 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_774 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_741 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_785 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_796 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_752 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_763 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_80 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1419 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1408 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1931 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1975 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1942 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1953 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1964 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1920 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_560 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_571 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_593 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_582 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1238 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1249 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1205 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1216 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1227 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1783 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1750 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1794 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1761 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1772 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_390 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1002 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1013 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1024 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1057 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1068 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1079 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1035 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1046 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1580 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1591 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_912 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_901 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_956 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_923 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_967 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_978 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_934 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_989 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_945 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_208 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_219 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_731 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_742 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_753 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_70 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_720 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_81 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_775 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_786 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_92 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_797 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_764 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1409 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1921 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1910 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1976 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1932 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1943 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1954 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1965 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_550 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_594 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_561 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_572 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_583 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1206 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1239 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1217 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1228 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1740 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1751 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1762 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1784 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1795 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1773 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_380 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_391 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1003 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1014 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1058 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1025 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1036 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1047 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1069 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1570 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1581 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1592 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_913 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_924 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_935 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_902 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_957 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_968 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_979 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_946 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_209 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_732 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_776 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_82 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_743 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_787 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_93 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_60 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_754 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_710 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_71 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_765 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_721 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_798 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1922 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1933 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1944 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1900 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1955 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1911 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1977 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1966 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_551 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_595 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_562 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_573 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_584 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_540 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1207 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1218 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1229 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1741 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1785 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1752 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1796 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1763 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1774 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1730 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_370 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_381 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_392 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1004 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1048 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1015 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1059 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1026 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1037 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1560 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1571 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1582 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1593 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1390 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_914 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_958 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_925 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_969 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_936 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_947 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_903 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_733 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_777 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_83 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_744 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_788 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_50 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_94 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_700 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_61 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_799 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_755 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_711 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_72 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_766 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_722 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1923 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1967 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1934 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1945 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1901 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1956 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1912 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_596 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_552 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_563 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_574 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_530 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_585 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_541 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1208 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1219 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1742 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1786 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1753 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1797 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1764 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1720 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1775 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
Xunit_cap_1731 m3_2060_293480# m3_142420_294000# m3_2060_293480# unit_cap
.ends


* Top level circuit converter

Xpower_stage_0 fc2_read power_stage_0/VN fc1_read power_stage
Xflying_cap_0 fc2_read fc1_read flying_cap
.end

