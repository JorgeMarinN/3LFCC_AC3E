magic
tech sky130A
timestamp 1660314476
<< metal3 >>
rect 1000 3030 2000 3085
rect 0 2000 3030 3030
rect 0 1000 3085 2000
rect 0 0 3030 1000
<< mimcap >>
rect 15 3007 3015 3015
rect 15 23 23 3007
rect 3007 23 3015 3007
rect 15 15 3015 23
<< mimcapcontact >>
rect 23 23 3007 3007
<< metal4 >>
rect 1000 3030 2000 3085
rect 0 3007 3030 3030
rect 0 23 23 3007
rect 3007 2000 3030 3007
rect 3007 1000 3085 2000
rect 3007 23 3030 1000
rect 0 0 3030 23
<< end >>
