magic
tech sky130A
timestamp 1666629347
<< metal4 >>
rect 57929 76784 65539 100320
rect 57929 69306 57995 76784
rect 65473 69306 65539 76784
rect 57929 69240 65539 69306
<< via4 >>
rect 57995 69306 65473 76784
<< metal5 >>
rect 50000 85100 92710 92710
rect 50000 77170 84780 84780
rect 50000 57609 57609 77170
rect 57929 76784 65539 76850
rect 57929 69306 57995 76784
rect 65473 69306 65539 76784
rect 57929 65539 65539 69306
rect 77170 65539 84780 77170
rect 57929 57929 84780 65539
rect 85100 57609 92710 85100
rect 50000 50000 92710 57609
<< end >>
