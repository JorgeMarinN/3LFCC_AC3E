magic
tech sky130A
magscale 1 2
timestamp 1663531380
<< error_s >>
rect -4 4682 2 4692
rect 24 4682 30 4684
<< metal1 >>
rect -2436 8898 -2296 8900
rect -2436 8896 -1800 8898
rect -2436 8808 3274 8896
rect -2436 7738 -2296 8808
rect -1870 8806 3274 8808
rect -2436 7140 -2294 7738
rect -2434 2324 -2294 7140
rect -2256 6472 -2116 6482
rect -2256 6372 -2238 6472
rect -2138 6372 -2116 6472
rect -2256 3648 -2116 6372
rect -2256 3548 -2238 3648
rect -2138 3548 -2116 3648
rect -2256 3538 -2116 3548
rect -2078 2866 -1938 6698
rect -116 6568 -106 6586
rect -122 6486 -106 6568
rect 0 6568 10 6586
rect 0 6486 18 6568
rect -122 4682 18 6486
rect -122 4582 -104 4682
rect 2 4582 18 4682
rect -1874 4034 160 4264
rect -158 4012 160 4034
rect -96 4010 160 4012
rect -1876 3184 -1318 3270
rect -2446 2312 -2254 2324
rect -2446 2252 -2434 2312
rect -2374 2252 -2326 2312
rect -2266 2252 -2254 2312
rect -776 2254 -766 2314
rect -706 2254 -696 2314
rect -630 2254 -620 2314
rect -560 2254 -550 2314
rect -476 2254 -466 2314
rect -406 2254 -396 2314
rect -2446 2242 -2254 2252
rect 20 0 160 4010
<< via1 >>
rect -2238 6372 -2138 6472
rect -2238 3548 -2138 3648
rect -106 6486 0 6586
rect -104 4582 2 4682
rect -2434 2252 -2374 2312
rect -2326 2252 -2266 2312
rect -766 2254 -706 2314
rect -620 2254 -560 2314
rect -466 2254 -406 2314
<< metal2 >>
rect -106 6586 0 6596
rect -272 6492 -106 6572
rect -2238 6472 -2138 6482
rect -106 6476 0 6486
rect -2242 6384 -2238 6462
rect -2138 6384 -1784 6462
rect -2238 6362 -2138 6372
rect -104 4682 2 4692
rect 24 4682 392 4684
rect 2 4584 392 4682
rect 2 4582 66 4584
rect -104 4572 2 4582
rect -1897 3705 -1160 3758
rect -2238 3648 -2138 3658
rect -2138 3568 -1252 3628
rect -2238 3538 -2138 3548
rect -1312 3020 -1252 3568
rect -1220 3102 -1160 3705
rect -1220 3068 -1124 3102
rect -1312 2986 -1040 3020
rect -2446 2312 -2254 2324
rect -766 2314 -706 2324
rect -2446 2252 -2434 2312
rect -2374 2252 -2326 2312
rect -2266 2254 -766 2312
rect -620 2314 -560 2324
rect -706 2254 -620 2312
rect -466 2314 -406 2324
rect -560 2254 -466 2312
rect -406 2254 -322 2312
rect -2266 2252 -322 2254
rect -2446 2242 -2254 2252
rect -766 2244 -706 2252
rect -620 2244 -560 2252
rect -466 2244 -406 2252
use cruzados  cruzados_0
timestamp 1663527930
transform 1 0 -880 0 -1 2872
box -1226 -3826 870 654
use inv_1_8  inv_1_8_0
timestamp 1663277475
transform 1 0 -1891 0 -1 4111
box -11 19 600 1019
use inv_400  inv_400_0
timestamp 1663461063
transform 1 0 330 0 1 -32158
box -188 32158 3166 41088
use stage_100  stage_100_0
timestamp 1663462081
transform 1 0 -1914 0 1 6686
box -14 -2532 1760 2244
<< labels >>
rlabel metal1 -1876 3184 -1318 3270 1 VDD
rlabel metal1 -1870 8806 3274 8896 1 VH
rlabel metal1 -2256 3648 -2116 6372 1 IN
rlabel metal1 20 0 160 4264 1 GND
rlabel space 3274 4278 3460 4378 1 OUT
rlabel space 142 0 3496 8930 1 OUT
<< end >>
