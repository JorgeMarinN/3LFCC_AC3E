magic
tech sky130A
timestamp 1668297044
<< metal5 >>
rect 27000 13500 27500 14000
rect 27000 13000 28000 13500
rect 27000 12000 28500 13000
rect 3500 11500 6000 12000
rect 7500 11500 10000 12000
rect 10500 11500 12000 12000
rect 14500 11500 17000 12000
rect 18500 11500 21000 12000
rect 21500 11500 22000 12000
rect 26500 11500 28500 12000
rect 4000 11000 5500 11500
rect 8000 11000 9500 11500
rect 11000 11000 12500 11500
rect 15000 11000 16500 11500
rect 18000 11000 19000 11500
rect 20500 11000 22000 11500
rect 26000 11000 28000 11500
rect 4500 6500 5500 11000
rect 8500 6500 9000 11000
rect 11500 10000 13000 11000
rect 11500 6500 12000 10000
rect 12500 9500 13500 10000
rect 12500 9000 14000 9500
rect 13000 8500 14000 9000
rect 13500 8000 14500 8500
rect 14000 7500 15000 8000
rect 15500 7500 16000 11000
rect 17500 10000 18500 11000
rect 21000 10500 22000 11000
rect 25500 10500 27500 11000
rect 17500 9500 19000 10000
rect 21500 9500 22000 10500
rect 25000 10000 27000 10500
rect 24500 9500 28000 10000
rect 18000 9000 19500 9500
rect 24500 9000 27500 9500
rect 18500 8500 21000 9000
rect 24000 8900 25200 9000
rect 24000 8700 25000 8900
rect 24000 8600 24900 8700
rect 24000 8500 24800 8600
rect 25500 8500 27000 9000
rect 19500 8000 21500 8500
rect 24000 8400 24600 8500
rect 25100 8400 26000 8500
rect 24000 8200 24500 8400
rect 24000 8100 24400 8200
rect 24000 8000 24300 8100
rect 25000 8000 26000 8400
rect 20500 7500 22000 8000
rect 24600 7900 26500 8000
rect 24500 7500 26500 7900
rect 14000 7000 16000 7500
rect 14500 6500 16000 7000
rect 5000 6000 5500 6500
rect 8000 6000 9000 6500
rect 11000 6000 12500 6500
rect 15000 6000 16000 6500
rect 5000 5500 8500 6000
rect 10500 5500 13000 6000
rect 15500 5500 16000 6000
rect 17500 6500 18000 7500
rect 21000 6500 22000 7500
rect 24000 7000 26000 7500
rect 23500 6500 25500 7000
rect 17500 6000 18500 6500
rect 20500 6000 21500 6500
rect 17500 5500 21000 6000
rect 23500 5500 25000 6500
rect 24000 4700 24500 5500
rect 24000 4500 24700 4700
rect 24300 4300 25000 4500
rect 24500 4000 25000 4300
rect 24500 3500 25500 4000
rect 25000 3000 25500 3500
<< comment >>
rect -100 17000 32100 17100
rect -100 0 0 17000
rect 32000 0 32100 17000
rect -100 -100 32100 0
<< end >>
