magic
tech sky130A
timestamp 1668455399
<< metal5 >>
rect 24900 21800 36600 22000
rect 36900 21800 48600 22000
rect 25100 21700 28000 21800
rect 25200 21600 28000 21700
rect 33500 21700 36400 21800
rect 37100 21700 48400 21800
rect 33500 21600 36300 21700
rect 37200 21600 48300 21700
rect 25300 21500 28000 21600
rect 25400 21300 28000 21500
rect 25500 21000 28000 21300
rect 25500 20900 26600 21000
rect 26900 20900 28000 21000
rect 25500 20800 26500 20900
rect 27000 20800 28000 20900
rect 25500 20700 26400 20800
rect 27100 20700 28000 20800
rect 28200 21500 29300 21600
rect 32200 21500 33300 21600
rect 28200 21400 29400 21500
rect 32100 21400 33300 21500
rect 28200 21300 29500 21400
rect 32000 21300 33300 21400
rect 28200 21200 29600 21300
rect 31900 21200 33300 21300
rect 28200 21100 29700 21200
rect 31800 21100 33300 21200
rect 28200 21000 29800 21100
rect 31700 21000 33300 21100
rect 28200 20900 29900 21000
rect 31600 20900 33300 21000
rect 28200 20800 30000 20900
rect 31500 20800 33300 20900
rect 28200 20700 30100 20800
rect 31400 20700 33300 20800
rect 33500 21500 36200 21600
rect 37300 21500 48200 21600
rect 33500 21300 36100 21500
rect 37400 21300 39100 21500
rect 39400 21300 42600 21500
rect 42900 21300 46100 21500
rect 46400 21300 48100 21500
rect 33500 21000 36000 21300
rect 33500 20900 34600 21000
rect 34900 20900 36000 21000
rect 33500 20800 34500 20900
rect 35000 20800 36000 20900
rect 33500 20700 34400 20800
rect 35100 20700 36000 20800
rect 25500 20600 26300 20700
rect 27200 20600 28000 20700
rect 28300 20600 30200 20700
rect 31300 20600 33200 20700
rect 33500 20600 34300 20700
rect 35200 20600 36000 20700
rect 25500 20500 26200 20600
rect 27300 20500 28000 20600
rect 28400 20500 30300 20600
rect 31200 20500 33100 20600
rect 33500 20500 34200 20600
rect 35300 20500 36000 20600
rect 25500 20400 26100 20500
rect 27400 20400 28000 20500
rect 28500 20400 30400 20500
rect 31100 20400 33000 20500
rect 33500 20400 34100 20500
rect 35400 20400 36000 20500
rect 25500 20000 26000 20400
rect 27500 20000 28000 20400
rect 28600 20300 30500 20400
rect 31000 20300 32900 20400
rect 28700 20200 30600 20300
rect 30900 20200 32800 20300
rect 28800 20100 32700 20200
rect 28900 20000 32600 20100
rect 33500 20000 34000 20400
rect 35500 20000 36000 20400
rect 25500 19800 26100 20000
rect 27400 19800 28000 20000
rect 29000 19900 32500 20000
rect 29100 19800 32400 19900
rect 33500 19800 34100 20000
rect 35400 19800 36000 20000
rect 25500 19700 26200 19800
rect 27300 19700 28000 19800
rect 29200 19700 32300 19800
rect 33500 19700 34200 19800
rect 35300 19700 36000 19800
rect 25500 19600 26300 19700
rect 27200 19600 28000 19700
rect 29300 19600 32200 19700
rect 33500 19600 34300 19700
rect 35200 19600 36000 19700
rect 25500 19500 26500 19600
rect 27000 19500 28000 19600
rect 29400 19500 32100 19600
rect 33500 19500 34500 19600
rect 35000 19500 36000 19600
rect 25500 18500 28000 19500
rect 29500 19300 32000 19500
rect 29400 19200 32100 19300
rect 29300 19100 32200 19200
rect 29200 19000 32300 19100
rect 29100 18900 32400 19000
rect 29000 18800 32500 18900
rect 28900 18700 32600 18800
rect 28800 18600 32700 18700
rect 28700 18500 30600 18600
rect 30900 18500 32800 18600
rect 33500 18500 36000 19500
rect 25500 18400 26600 18500
rect 26900 18400 28000 18500
rect 28600 18400 30500 18500
rect 31000 18400 32900 18500
rect 33500 18400 34600 18500
rect 34900 18400 36000 18500
rect 25500 18300 26500 18400
rect 27000 18300 28000 18400
rect 28500 18300 30400 18400
rect 31100 18300 33000 18400
rect 33500 18300 34500 18400
rect 35000 18300 36000 18400
rect 25500 18200 26400 18300
rect 27100 18200 28000 18300
rect 28400 18200 30300 18300
rect 31200 18200 33100 18300
rect 33500 18200 34400 18300
rect 35100 18200 36000 18300
rect 25500 18100 26300 18200
rect 27200 18100 28000 18200
rect 28300 18100 30200 18200
rect 31300 18100 33200 18200
rect 33500 18100 34300 18200
rect 35200 18100 36000 18200
rect 25500 18000 26200 18100
rect 27300 18000 28000 18100
rect 25500 17900 26100 18000
rect 27400 17900 28000 18000
rect 25500 17500 26000 17900
rect 27500 17500 28000 17900
rect 25500 17300 26100 17500
rect 27400 17300 28000 17500
rect 25500 17200 26200 17300
rect 27300 17200 28000 17300
rect 25500 17100 26300 17200
rect 27200 17100 28000 17200
rect 28200 18000 30100 18100
rect 31400 18000 33300 18100
rect 28200 17900 30000 18000
rect 31500 17900 33300 18000
rect 28200 17800 29900 17900
rect 31600 17800 33300 17900
rect 28200 17700 29800 17800
rect 31700 17700 33300 17800
rect 28200 17600 29700 17700
rect 31800 17600 33300 17700
rect 28200 17500 29600 17600
rect 31900 17500 33300 17600
rect 28200 17400 29500 17500
rect 32000 17400 33300 17500
rect 28200 17300 29400 17400
rect 32100 17300 33300 17400
rect 28200 17200 29300 17300
rect 32200 17200 33300 17300
rect 28200 17100 29200 17200
rect 32300 17100 33300 17200
rect 33500 18000 34200 18100
rect 35300 18000 36000 18100
rect 33500 17900 34100 18000
rect 35400 17900 36000 18000
rect 33500 17500 34000 17900
rect 35500 17500 36000 17900
rect 33500 17300 34100 17500
rect 35400 17300 36000 17500
rect 33500 17200 34200 17300
rect 35300 17200 36000 17300
rect 33500 17100 34300 17200
rect 35200 17100 36000 17200
rect 25500 17000 26500 17100
rect 27000 17000 28000 17100
rect 25500 16900 28000 17000
rect 33500 17000 34500 17100
rect 35000 17000 36000 17100
rect 33500 16900 36000 17000
rect 25500 16700 36000 16900
rect 25500 16000 28000 16700
rect 25500 15900 26600 16000
rect 26900 15900 28000 16000
rect 25500 15800 26500 15900
rect 27000 15800 28000 15900
rect 25500 15700 26400 15800
rect 27100 15700 28000 15800
rect 25500 15600 26300 15700
rect 27200 15600 28000 15700
rect 25500 15500 26200 15600
rect 27300 15500 28000 15600
rect 28270 15500 29170 16000
rect 29330 15500 30230 16000
rect 25500 15400 26100 15500
rect 27400 15400 28000 15500
rect 25500 15000 26000 15400
rect 27500 15000 28000 15400
rect 28370 15000 29070 15500
rect 29430 15000 30130 15500
rect 25500 14800 26100 15000
rect 27400 14800 28000 15000
rect 25500 14700 26200 14800
rect 27300 14700 28000 14800
rect 25500 14600 26300 14700
rect 27200 14600 28000 14700
rect 25500 14500 26500 14600
rect 27000 14500 28000 14600
rect 28470 14500 28970 15000
rect 29530 14500 30030 15000
rect 25500 13500 28000 14500
rect 25500 13400 26600 13500
rect 26900 13400 28000 13500
rect 25500 13300 26500 13400
rect 27000 13300 28000 13400
rect 25500 13200 26400 13300
rect 27100 13200 28000 13300
rect 25500 13100 26300 13200
rect 27200 13100 28000 13200
rect 25500 13000 26200 13100
rect 27300 13000 28000 13100
rect 28800 13000 29700 13500
rect 25500 12900 26100 13000
rect 27400 12900 28000 13000
rect 25500 12500 26000 12900
rect 27500 12500 28000 12900
rect 28900 12500 29600 13000
rect 25500 12300 26100 12500
rect 27400 12300 28000 12500
rect 25500 12200 26200 12300
rect 27300 12200 28000 12300
rect 25500 12100 26300 12200
rect 27200 12100 28000 12200
rect 25500 12000 26500 12100
rect 27000 12000 28000 12100
rect 29000 12000 29500 12500
rect 25500 11900 28100 12000
rect 25500 11800 28200 11900
rect 25500 11700 28300 11800
rect 25500 11600 28400 11700
rect 25500 11500 28500 11600
rect 25500 11400 28600 11500
rect 25500 11300 28700 11400
rect 25500 11200 28800 11300
rect 25500 11100 28900 11200
rect 25500 11000 29000 11100
rect 30600 11000 30900 16700
rect 32100 16000 32500 16100
rect 33500 16000 36000 16700
rect 31700 15900 32700 16000
rect 33500 15900 34600 16000
rect 34900 15900 36000 16000
rect 31500 15700 32900 15900
rect 33500 15800 34500 15900
rect 35000 15800 36000 15900
rect 33500 15700 34400 15800
rect 35100 15700 36000 15800
rect 31400 15500 33100 15700
rect 33500 15600 34300 15700
rect 35200 15600 36000 15700
rect 33500 15500 34200 15600
rect 35300 15500 36000 15600
rect 31260 14500 33200 15500
rect 33500 15400 34100 15500
rect 35400 15400 36000 15500
rect 33500 15000 34000 15400
rect 35500 15000 36000 15400
rect 33500 14800 34100 15000
rect 35400 14800 36000 15000
rect 33500 14700 34200 14800
rect 35300 14700 36000 14800
rect 33500 14600 34300 14700
rect 35200 14600 36000 14700
rect 33500 14500 34500 14600
rect 35000 14500 36000 14600
rect 31300 14400 33100 14500
rect 31400 14300 33100 14400
rect 31400 14200 33000 14300
rect 31500 14000 33000 14200
rect 31700 13900 32700 14000
rect 31800 13800 32600 13900
rect 32100 13160 32400 13800
rect 32090 13010 32400 13160
rect 32080 12730 32400 13010
rect 32070 12540 32400 12730
rect 32060 12490 32400 12540
rect 33500 13500 36000 14500
rect 33500 13400 34600 13500
rect 34900 13400 36000 13500
rect 33500 13300 34500 13400
rect 35000 13300 36000 13400
rect 33500 13200 34400 13300
rect 35100 13200 36000 13300
rect 33500 13100 34300 13200
rect 35200 13100 36000 13200
rect 33500 13000 34200 13100
rect 35300 13000 36000 13100
rect 33500 12900 34100 13000
rect 35400 12900 36000 13000
rect 33500 12500 34000 12900
rect 35500 12500 36000 12900
rect 32060 12400 32410 12490
rect 32040 12370 32410 12400
rect 32010 12340 32420 12370
rect 32000 12300 32440 12340
rect 33500 12300 34100 12500
rect 35400 12300 36000 12500
rect 31900 12260 32500 12300
rect 31840 12250 32500 12260
rect 31840 12240 32570 12250
rect 31840 12230 32600 12240
rect 31800 12220 32630 12230
rect 31770 12210 32630 12220
rect 31760 12200 32630 12210
rect 33500 12200 34200 12300
rect 35300 12200 36000 12300
rect 31740 12190 32700 12200
rect 31720 12180 32700 12190
rect 31700 12170 32700 12180
rect 31690 12140 32700 12170
rect 31690 12130 32740 12140
rect 31640 12100 32740 12130
rect 33500 12100 34300 12200
rect 35200 12100 36000 12200
rect 31600 12080 32800 12100
rect 31600 12060 32280 12080
rect 32450 12070 32800 12080
rect 31580 12040 31840 12060
rect 31560 12030 31840 12040
rect 31550 12000 31840 12030
rect 31550 11930 31800 12000
rect 32050 11950 32280 12060
rect 32490 12040 32800 12070
rect 32490 12030 32840 12040
rect 32520 12020 32840 12030
rect 32520 12000 32880 12020
rect 33500 12000 34500 12100
rect 35000 12000 36000 12100
rect 32570 11980 32910 12000
rect 31550 11900 31760 11930
rect 32050 11900 32260 11950
rect 32600 11900 32940 11980
rect 33400 11900 36000 12000
rect 31550 11880 31740 11900
rect 31550 11870 31720 11880
rect 32000 11840 32260 11900
rect 32670 11880 32940 11900
rect 32710 11860 32940 11880
rect 32740 11840 32940 11860
rect 31970 11800 32260 11840
rect 32770 11820 32940 11840
rect 33300 11800 36000 11900
rect 31930 11790 32260 11800
rect 31930 11780 32240 11790
rect 31930 11770 32230 11780
rect 31900 11760 32230 11770
rect 31900 11700 32200 11760
rect 33200 11700 36000 11800
rect 31900 11680 32140 11700
rect 31900 11600 32100 11680
rect 33100 11600 36000 11700
rect 33000 11500 36000 11600
rect 32900 11400 36000 11500
rect 32800 11300 36000 11400
rect 32700 11200 36000 11300
rect 32600 11100 36000 11200
rect 32500 11000 36000 11100
rect 25500 10500 36000 11000
rect 25500 10400 28600 10500
rect 28900 10400 32600 10500
rect 32900 10400 36000 10500
rect 25500 10300 28500 10400
rect 29000 10300 32500 10400
rect 33000 10300 36000 10400
rect 25500 10200 28400 10300
rect 29100 10200 32400 10300
rect 33100 10200 36000 10300
rect 25500 10100 28300 10200
rect 29200 10100 32300 10200
rect 33200 10100 36000 10200
rect 25500 10000 28200 10100
rect 29300 10000 32200 10100
rect 33300 10000 36000 10100
rect 37500 21100 39000 21300
rect 37500 20800 38400 21100
rect 38700 21000 39000 21100
rect 39500 21100 42500 21300
rect 39500 21000 39800 21100
rect 40100 20800 41900 21100
rect 42200 21000 42500 21100
rect 43000 21100 46000 21300
rect 43000 21000 43300 21100
rect 43600 20800 45400 21100
rect 45700 21000 46000 21100
rect 46500 21100 48000 21300
rect 46500 21000 46800 21100
rect 47100 20800 48000 21100
rect 37500 20500 38500 20800
rect 40000 20500 42000 20800
rect 43500 20500 45500 20800
rect 47000 20500 48000 20800
rect 37500 20400 38200 20500
rect 40300 20400 41700 20500
rect 43800 20400 45200 20500
rect 47300 20400 48000 20500
rect 37500 20100 38000 20400
rect 40500 20100 41500 20400
rect 44000 20100 45000 20400
rect 47500 20100 48000 20400
rect 37500 20000 38200 20100
rect 40300 20000 41700 20100
rect 43800 20000 45200 20100
rect 47300 20000 48000 20100
rect 37500 19700 38500 20000
rect 40000 19700 42000 20000
rect 43500 19700 45500 20000
rect 47000 19700 48000 20000
rect 37500 19400 38400 19700
rect 38700 19400 39000 19500
rect 37500 19200 39000 19400
rect 39500 19400 39800 19500
rect 40100 19400 41900 19700
rect 42200 19400 42500 19500
rect 39500 19200 42500 19400
rect 43000 19400 43300 19500
rect 43600 19400 45400 19700
rect 45700 19400 46000 19500
rect 43000 19200 46000 19400
rect 46500 19400 46800 19500
rect 47100 19400 48000 19700
rect 46500 19200 48000 19400
rect 37500 19000 39100 19200
rect 39400 19000 42600 19200
rect 42900 19000 46100 19200
rect 46400 19000 48000 19200
rect 37500 18500 48000 19000
rect 37500 10400 38000 18500
rect 39600 17310 39760 17320
rect 39600 17300 39810 17310
rect 39600 17290 39860 17300
rect 39600 17280 39920 17290
rect 39600 17270 39960 17280
rect 39600 17260 40020 17270
rect 39600 17250 40100 17260
rect 39600 17240 40140 17250
rect 39600 17230 40170 17240
rect 39600 17220 40210 17230
rect 39600 17210 40250 17220
rect 39600 17200 40280 17210
rect 39600 17180 40300 17200
rect 39600 17160 40350 17180
rect 39680 17150 40370 17160
rect 39740 17140 40370 17150
rect 39780 17130 40370 17140
rect 39820 17120 40390 17130
rect 39880 17110 40390 17120
rect 39940 17100 40390 17110
rect 40000 17080 41630 17100
rect 44040 17080 44900 17100
rect 40000 17050 41960 17080
rect 43640 17070 44900 17080
rect 43640 17060 44950 17070
rect 43640 17050 45010 17060
rect 40000 17020 42200 17050
rect 43500 17030 45030 17050
rect 43500 17020 45070 17030
rect 40000 17000 42430 17020
rect 43070 17000 45130 17020
rect 40000 16980 45200 17000
rect 40000 16960 45230 16980
rect 40000 16940 45300 16960
rect 39900 16930 45300 16940
rect 39800 16910 45340 16930
rect 39750 16900 45340 16910
rect 39750 16890 45400 16900
rect 39700 16870 45400 16890
rect 39660 16860 45400 16870
rect 39660 16840 45440 16860
rect 39660 16830 45470 16840
rect 39640 16800 45470 16830
rect 39620 16780 45500 16800
rect 39600 16750 45500 16780
rect 39600 16740 45510 16750
rect 39590 16710 45510 16740
rect 39550 16700 45510 16710
rect 39540 16670 45510 16700
rect 39500 16650 45510 16670
rect 39500 16600 45530 16650
rect 39470 16590 43500 16600
rect 39430 16560 43500 16590
rect 43730 16560 45530 16600
rect 39420 16540 43500 16560
rect 39400 16470 43500 16540
rect 43800 16520 45530 16560
rect 43840 16500 45530 16520
rect 43900 16480 45530 16500
rect 39380 16400 43500 16470
rect 43940 16460 45530 16480
rect 44000 16420 45530 16460
rect 44030 16400 45530 16420
rect 39380 16390 43680 16400
rect 39380 16360 43700 16390
rect 44080 16380 45180 16400
rect 44120 16360 45180 16380
rect 39380 16340 43760 16360
rect 44170 16340 45180 16360
rect 39380 16300 43800 16340
rect 44200 16330 45180 16340
rect 45340 16360 45530 16400
rect 44200 16300 45150 16330
rect 39380 16280 43870 16300
rect 44290 16280 45130 16300
rect 39400 16250 43900 16280
rect 44340 16260 45120 16280
rect 44340 16250 45080 16260
rect 39400 16240 43940 16250
rect 39420 16230 43940 16240
rect 44370 16240 45080 16250
rect 44370 16230 45060 16240
rect 39420 16200 43980 16230
rect 44400 16210 45040 16230
rect 44400 16200 45000 16210
rect 45340 16200 45520 16360
rect 39460 16180 44020 16200
rect 44430 16190 44990 16200
rect 44430 16180 44950 16190
rect 39460 16170 44060 16180
rect 39500 16160 39940 16170
rect 40130 16160 44060 16170
rect 44460 16170 44950 16180
rect 45320 16170 45510 16200
rect 44460 16160 44930 16170
rect 39500 16150 39850 16160
rect 40130 16150 44080 16160
rect 44500 16150 44930 16160
rect 39550 16140 39800 16150
rect 40130 16140 44110 16150
rect 39580 16130 39770 16140
rect 40160 16130 44110 16140
rect 44500 16130 44900 16150
rect 45300 16130 45510 16170
rect 39580 16120 39750 16130
rect 40160 16120 44130 16130
rect 44530 16120 44900 16130
rect 40160 16100 44170 16120
rect 44530 16100 44860 16120
rect 45260 16100 45510 16130
rect 40200 16060 44200 16100
rect 44590 16090 44770 16100
rect 40200 16040 44270 16060
rect 45200 16050 45510 16100
rect 40240 16010 44270 16040
rect 45150 16030 45510 16050
rect 45120 16020 45510 16030
rect 40260 16000 44310 16010
rect 45120 16000 45500 16020
rect 40300 15970 44370 16000
rect 45050 15970 45500 16000
rect 40330 15950 44400 15970
rect 40370 15930 44400 15950
rect 45000 15950 45500 15970
rect 45000 15940 45490 15950
rect 40430 15920 44440 15930
rect 44960 15920 45490 15940
rect 40460 15900 44440 15920
rect 44870 15900 45490 15920
rect 40500 15870 45490 15900
rect 40510 15860 45490 15870
rect 40510 15840 45480 15860
rect 40510 15820 45460 15840
rect 40510 15800 45440 15820
rect 40540 15770 45400 15800
rect 40540 15740 45370 15770
rect 40580 15730 45370 15740
rect 40580 15700 45340 15730
rect 40600 15660 45300 15700
rect 40600 15630 45280 15660
rect 40620 15600 45260 15630
rect 40620 15570 45230 15600
rect 40620 15550 45210 15570
rect 40620 15540 45200 15550
rect 40640 15520 45200 15540
rect 40640 15490 45180 15520
rect 40640 15470 45170 15490
rect 40640 15460 45150 15470
rect 40670 15430 45150 15460
rect 40690 15420 45130 15430
rect 40700 15410 45130 15420
rect 40710 15400 45130 15410
rect 40710 15390 44140 15400
rect 40730 15370 44070 15390
rect 40730 15360 44000 15370
rect 40760 15340 44000 15360
rect 40760 15330 43930 15340
rect 40780 15320 43930 15330
rect 40800 15310 43870 15320
rect 40820 15300 43870 15310
rect 40820 15290 43780 15300
rect 40850 15280 43780 15290
rect 40850 15270 43700 15280
rect 40880 15250 43660 15270
rect 40930 15240 43660 15250
rect 44300 15240 45100 15400
rect 40930 15220 43610 15240
rect 40950 15210 43530 15220
rect 40980 15200 43530 15210
rect 40980 15180 42140 15200
rect 41010 15160 42140 15180
rect 41040 15140 42140 15160
rect 41100 15120 42140 15140
rect 41120 15100 42140 15120
rect 43100 15160 43400 15200
rect 44290 15180 45120 15240
rect 43100 15140 43370 15160
rect 44290 15140 45140 15180
rect 43100 15120 43310 15140
rect 43100 15100 43260 15120
rect 44290 15100 45180 15140
rect 41150 15090 42100 15100
rect 41220 15070 42100 15090
rect 44290 15080 45200 15100
rect 41270 15040 42100 15070
rect 44310 15060 45200 15080
rect 41300 15020 42100 15040
rect 44320 15020 45240 15060
rect 41320 15000 42100 15020
rect 44330 15000 45240 15020
rect 41350 14990 42100 15000
rect 41400 14970 42100 14990
rect 44340 14980 45260 15000
rect 41450 14940 42100 14970
rect 44360 14950 45270 14980
rect 41460 14930 42100 14940
rect 41460 14920 42120 14930
rect 41490 14910 42120 14920
rect 44380 14910 45300 14950
rect 41520 14810 42120 14910
rect 44400 14900 45300 14910
rect 44400 14840 44700 14900
rect 41520 14750 42150 14810
rect 44400 14750 44690 14840
rect 44900 14800 45300 14900
rect 41500 14700 42150 14750
rect 44380 14730 44690 14750
rect 44910 14790 45300 14800
rect 44910 14730 45290 14790
rect 44380 14700 44680 14730
rect 41460 14680 42150 14700
rect 41460 14670 42170 14680
rect 41460 14630 41720 14670
rect 41440 14600 41720 14630
rect 41880 14600 42170 14670
rect 44370 14670 44680 14700
rect 44930 14700 45290 14730
rect 44930 14670 45280 14700
rect 44370 14640 44660 14670
rect 44350 14610 44650 14640
rect 44930 14610 45260 14670
rect 41440 14580 41700 14600
rect 41400 14520 41700 14580
rect 41400 14500 41660 14520
rect 41900 14510 42200 14600
rect 44350 14580 44630 14610
rect 44330 14560 44620 14580
rect 44940 14560 45230 14610
rect 44330 14550 44600 14560
rect 44330 14530 44590 14550
rect 41370 14440 41660 14500
rect 41940 14450 42200 14510
rect 41340 14400 41660 14440
rect 41950 14400 42200 14450
rect 41340 14380 41600 14400
rect 41300 14350 41600 14380
rect 41300 14300 41550 14350
rect 41270 14250 41500 14300
rect 41200 14200 41500 14250
rect 42000 14250 42200 14400
rect 44320 14510 44590 14530
rect 44970 14520 45230 14560
rect 44320 14460 44570 14510
rect 44970 14500 45200 14520
rect 45000 14480 45200 14500
rect 44320 14400 44550 14460
rect 45000 14420 45190 14480
rect 44320 14370 44540 14400
rect 44330 14300 44540 14370
rect 42000 14200 42220 14250
rect 44330 14220 44530 14300
rect 45000 14260 45180 14420
rect 45000 14230 45190 14260
rect 44330 14210 44500 14220
rect 44300 14200 44500 14210
rect 45000 14200 45200 14230
rect 41150 14160 41460 14200
rect 41950 14160 42220 14200
rect 44270 14180 44500 14200
rect 44950 14180 45200 14200
rect 44250 14160 44500 14180
rect 44930 14170 45200 14180
rect 41100 14100 41460 14160
rect 41100 14000 41400 14100
rect 41900 14050 42220 14160
rect 41900 14000 42200 14050
rect 44200 14030 44500 14160
rect 44900 14070 45200 14170
rect 44900 14030 45180 14070
rect 44200 14000 44460 14030
rect 44900 14010 45090 14030
rect 44930 14000 45090 14010
rect 39600 13310 39760 13320
rect 39600 13300 39810 13310
rect 39600 13290 39860 13300
rect 39600 13280 39920 13290
rect 39600 13270 39960 13280
rect 39600 13260 40020 13270
rect 39600 13250 40100 13260
rect 39600 13240 40140 13250
rect 39600 13230 40170 13240
rect 39600 13220 40210 13230
rect 39600 13210 40250 13220
rect 39600 13200 40280 13210
rect 39600 13180 40300 13200
rect 39600 13160 40350 13180
rect 39680 13150 40370 13160
rect 39740 13140 40370 13150
rect 39780 13130 40370 13140
rect 39820 13120 40390 13130
rect 39880 13110 40390 13120
rect 39940 13100 40390 13110
rect 40000 13080 41630 13100
rect 44040 13080 44900 13100
rect 40000 13050 41960 13080
rect 43640 13070 44900 13080
rect 43640 13060 44950 13070
rect 43640 13050 45010 13060
rect 40000 13020 42200 13050
rect 43500 13030 45030 13050
rect 43500 13020 45070 13030
rect 40000 13000 42430 13020
rect 43070 13000 45130 13020
rect 40000 12980 45200 13000
rect 40000 12960 45230 12980
rect 40000 12940 45300 12960
rect 39900 12930 45300 12940
rect 39800 12910 45340 12930
rect 39750 12900 45340 12910
rect 39750 12890 45400 12900
rect 39700 12870 45400 12890
rect 39660 12860 45400 12870
rect 39660 12840 45440 12860
rect 39660 12830 45470 12840
rect 39640 12800 45470 12830
rect 39620 12780 45500 12800
rect 39600 12750 45500 12780
rect 39600 12740 45510 12750
rect 39590 12710 45510 12740
rect 39550 12700 45510 12710
rect 39540 12670 45510 12700
rect 39500 12650 45510 12670
rect 39500 12600 45530 12650
rect 39470 12590 43500 12600
rect 39430 12560 43500 12590
rect 43730 12560 45530 12600
rect 39420 12540 43500 12560
rect 39400 12470 43500 12540
rect 43800 12520 45530 12560
rect 43840 12500 45530 12520
rect 43900 12480 45530 12500
rect 39380 12400 43500 12470
rect 43940 12460 45530 12480
rect 44000 12420 45530 12460
rect 44030 12400 45530 12420
rect 39380 12390 43680 12400
rect 39380 12360 43700 12390
rect 44080 12380 45180 12400
rect 44120 12360 45180 12380
rect 39380 12340 43760 12360
rect 44170 12340 45180 12360
rect 39380 12300 43800 12340
rect 44200 12330 45180 12340
rect 45340 12360 45530 12400
rect 44200 12300 45150 12330
rect 39380 12280 43870 12300
rect 44290 12280 45130 12300
rect 39400 12250 43900 12280
rect 44340 12260 45120 12280
rect 44340 12250 45080 12260
rect 39400 12240 43940 12250
rect 39420 12230 43940 12240
rect 44370 12240 45080 12250
rect 44370 12230 45060 12240
rect 39420 12200 43980 12230
rect 44400 12210 45040 12230
rect 44400 12200 45000 12210
rect 45340 12200 45520 12360
rect 39460 12180 44020 12200
rect 44430 12190 44990 12200
rect 44430 12180 44950 12190
rect 39460 12170 44060 12180
rect 39500 12160 39940 12170
rect 40130 12160 44060 12170
rect 44460 12170 44950 12180
rect 45320 12170 45510 12200
rect 44460 12160 44930 12170
rect 39500 12150 39850 12160
rect 40130 12150 44080 12160
rect 44500 12150 44930 12160
rect 39550 12140 39800 12150
rect 40130 12140 44110 12150
rect 39580 12130 39770 12140
rect 40160 12130 44110 12140
rect 44500 12130 44900 12150
rect 45300 12130 45510 12170
rect 39580 12120 39750 12130
rect 40160 12120 44130 12130
rect 44530 12120 44900 12130
rect 40160 12100 44170 12120
rect 44530 12100 44860 12120
rect 45260 12100 45510 12130
rect 40200 12060 44200 12100
rect 44590 12090 44770 12100
rect 40200 12040 44270 12060
rect 45200 12050 45510 12100
rect 40240 12010 44270 12040
rect 45150 12030 45510 12050
rect 45120 12020 45510 12030
rect 40260 12000 44310 12010
rect 45120 12000 45500 12020
rect 40300 11970 44370 12000
rect 45050 11970 45500 12000
rect 40330 11950 44400 11970
rect 40370 11930 44400 11950
rect 45000 11950 45500 11970
rect 45000 11940 45490 11950
rect 40430 11920 44440 11930
rect 44960 11920 45490 11940
rect 40460 11900 44440 11920
rect 44870 11900 45490 11920
rect 40500 11870 45490 11900
rect 40510 11860 45490 11870
rect 40510 11840 45480 11860
rect 40510 11820 45460 11840
rect 40510 11800 45440 11820
rect 40540 11770 45400 11800
rect 40540 11740 45370 11770
rect 40580 11730 45370 11740
rect 40580 11700 45340 11730
rect 40600 11660 45300 11700
rect 40600 11630 45280 11660
rect 40620 11600 45260 11630
rect 40620 11570 45230 11600
rect 40620 11550 45210 11570
rect 40620 11540 45200 11550
rect 40640 11520 45200 11540
rect 40640 11490 45180 11520
rect 40640 11470 45170 11490
rect 40640 11460 45150 11470
rect 40670 11430 45150 11460
rect 40690 11420 45130 11430
rect 40700 11410 45130 11420
rect 40710 11400 45130 11410
rect 40710 11390 44140 11400
rect 40730 11370 44070 11390
rect 40730 11360 44000 11370
rect 40760 11340 44000 11360
rect 40760 11330 43930 11340
rect 40780 11320 43930 11330
rect 40800 11310 43870 11320
rect 40820 11300 43870 11310
rect 40820 11290 43780 11300
rect 40850 11280 43780 11290
rect 40850 11270 43700 11280
rect 40880 11250 43660 11270
rect 40930 11240 43660 11250
rect 44300 11240 45100 11400
rect 40930 11220 43610 11240
rect 40950 11210 43530 11220
rect 40980 11200 43530 11210
rect 40980 11180 42140 11200
rect 41010 11160 42140 11180
rect 41040 11140 42140 11160
rect 41100 11120 42140 11140
rect 41120 11100 42140 11120
rect 43100 11160 43400 11200
rect 44290 11180 45120 11240
rect 43100 11140 43370 11160
rect 44290 11140 45140 11180
rect 43100 11120 43310 11140
rect 43100 11100 43260 11120
rect 44290 11100 45180 11140
rect 41150 11090 42100 11100
rect 41220 11070 42100 11090
rect 44290 11080 45200 11100
rect 41270 11040 42100 11070
rect 44310 11060 45200 11080
rect 41300 11020 42100 11040
rect 44320 11020 45240 11060
rect 41320 11000 42100 11020
rect 44330 11000 45240 11020
rect 41350 10990 42100 11000
rect 41400 10970 42100 10990
rect 44340 10980 45260 11000
rect 41450 10940 42100 10970
rect 44360 10950 45270 10980
rect 41460 10930 42100 10940
rect 41460 10920 42120 10930
rect 41490 10910 42120 10920
rect 44380 10910 45300 10950
rect 41520 10810 42120 10910
rect 44400 10900 45300 10910
rect 44400 10840 44700 10900
rect 41520 10750 42150 10810
rect 44400 10750 44690 10840
rect 44900 10800 45300 10900
rect 41500 10700 42150 10750
rect 44380 10730 44690 10750
rect 44910 10790 45300 10800
rect 44910 10730 45290 10790
rect 44380 10700 44680 10730
rect 41460 10680 42150 10700
rect 41460 10670 42170 10680
rect 41460 10630 41720 10670
rect 41440 10600 41720 10630
rect 41880 10600 42170 10670
rect 44370 10670 44680 10700
rect 44930 10700 45290 10730
rect 44930 10670 45280 10700
rect 44370 10640 44660 10670
rect 44350 10610 44650 10640
rect 44930 10610 45260 10670
rect 41440 10580 41700 10600
rect 41400 10520 41700 10580
rect 41400 10500 41660 10520
rect 41900 10510 42200 10600
rect 44350 10580 44630 10610
rect 44330 10560 44620 10580
rect 44940 10560 45230 10610
rect 44330 10550 44600 10560
rect 44330 10530 44590 10550
rect 41370 10440 41660 10500
rect 41940 10450 42200 10510
rect 41340 10400 41660 10440
rect 41950 10400 42200 10450
rect 37500 10300 38100 10400
rect 41340 10380 41600 10400
rect 41300 10350 41600 10380
rect 41300 10300 41550 10350
rect 37500 10200 38200 10300
rect 41270 10250 41500 10300
rect 41200 10200 41500 10250
rect 42000 10250 42200 10400
rect 44320 10510 44590 10530
rect 44970 10520 45230 10560
rect 44320 10460 44570 10510
rect 44970 10500 45200 10520
rect 45000 10480 45200 10500
rect 44320 10400 44550 10460
rect 45000 10420 45190 10480
rect 44320 10370 44540 10400
rect 44330 10300 44540 10370
rect 42000 10200 42220 10250
rect 44330 10220 44530 10300
rect 45000 10260 45180 10420
rect 47500 10400 48000 18500
rect 47400 10300 48000 10400
rect 45000 10230 45190 10260
rect 44330 10210 44500 10220
rect 44300 10200 44500 10210
rect 45000 10200 45200 10230
rect 47300 10200 48000 10300
rect 37500 10100 38300 10200
rect 41150 10160 41460 10200
rect 41950 10160 42220 10200
rect 44270 10180 44500 10200
rect 44950 10180 45200 10200
rect 44250 10160 44500 10180
rect 44930 10170 45200 10180
rect 41100 10100 41460 10160
rect 37500 10000 38400 10100
rect 41100 10000 41400 10100
rect 41900 10050 42220 10160
rect 41900 10000 42200 10050
rect 44200 10030 44500 10160
rect 44900 10070 45200 10170
rect 47200 10100 48000 10200
rect 44900 10030 45180 10070
rect 44200 10000 44460 10030
rect 44900 10010 45090 10030
rect 44930 10000 45090 10010
rect 47100 10000 48000 10100
rect 25600 9900 28100 10000
rect 29400 9900 32100 10000
rect 33400 9900 35900 10000
rect 37600 9900 38500 10000
rect 47000 9900 47900 10000
rect 25700 9800 28000 9900
rect 25800 9700 28000 9800
rect 25900 9600 28000 9700
rect 26000 9500 28000 9600
rect 29500 9500 32000 9900
rect 33500 9800 35800 9900
rect 37700 9800 38600 9900
rect 46900 9800 47800 9900
rect 33500 9700 35700 9800
rect 37800 9700 38700 9800
rect 46800 9700 47700 9800
rect 33500 9600 35600 9700
rect 37900 9600 38800 9700
rect 46700 9600 47600 9700
rect 33500 9500 35500 9600
rect 38000 9500 38900 9600
rect 46600 9500 47500 9600
rect 26100 9400 28100 9500
rect 26200 9300 28100 9400
rect 29400 9300 32100 9500
rect 33400 9400 35400 9500
rect 38100 9400 39000 9500
rect 46500 9400 47400 9500
rect 33400 9300 35300 9400
rect 38200 9300 39100 9400
rect 46400 9300 47300 9400
rect 26300 9200 28200 9300
rect 29300 9200 32200 9300
rect 33300 9200 35200 9300
rect 38300 9200 39200 9300
rect 46300 9200 47200 9300
rect 26400 9100 28300 9200
rect 29200 9100 32300 9200
rect 33200 9100 35100 9200
rect 38400 9100 39300 9200
rect 46200 9100 47100 9200
rect 26500 9000 28500 9100
rect 29000 9000 32500 9100
rect 33000 9000 35000 9100
rect 38500 9000 39400 9100
rect 46100 9000 47000 9100
rect 26600 8900 34900 9000
rect 38600 8900 46900 9000
rect 26700 8800 34800 8900
rect 38700 8800 46800 8900
rect 26800 8700 34700 8800
rect 38800 8700 46700 8800
rect 26900 8600 34600 8700
rect 38900 8600 46600 8700
rect 27000 8500 34500 8600
rect 39000 8500 46500 8600
rect 30200 8400 31300 8500
rect 42200 8400 43300 8500
rect 30400 8300 31100 8400
rect 42400 8300 43100 8400
rect 30500 8200 31000 8300
rect 42500 8200 43000 8300
rect 30600 8000 30900 8200
rect 42600 8000 42900 8200
rect 35100 7990 37600 8000
rect 35080 7980 37620 7990
rect 35060 7970 37640 7980
rect 35050 7960 37650 7970
rect 35040 7950 37660 7960
rect 35030 7940 37670 7950
rect 35020 7920 37680 7940
rect 35010 7900 37690 7920
rect 35000 7800 37700 7900
rect 35000 7000 35500 7800
rect 25600 6990 35500 7000
rect 25580 6980 35500 6990
rect 25560 6970 35500 6980
rect 25550 6960 35500 6970
rect 25540 6950 35500 6960
rect 25530 6940 35500 6950
rect 25520 6920 35500 6940
rect 25510 6900 35500 6920
rect 25500 6800 35500 6900
rect 25500 6000 25700 6800
rect 24800 5800 25700 6000
rect 24800 4000 25000 5800
rect 25500 5000 25700 5800
rect 26200 6300 26900 6500
rect 27200 6450 27360 6500
rect 27820 6450 27980 6500
rect 27200 6420 27370 6450
rect 27810 6420 27980 6450
rect 27200 6390 27380 6420
rect 27800 6390 27980 6420
rect 27200 6360 27390 6390
rect 27790 6360 27980 6390
rect 27200 6330 27400 6360
rect 27780 6330 27980 6360
rect 27200 6300 27410 6330
rect 27770 6300 27980 6330
rect 26200 6000 26400 6300
rect 27200 6290 27420 6300
rect 27210 6270 27420 6290
rect 27760 6280 27980 6300
rect 27760 6270 27970 6280
rect 27210 6260 27430 6270
rect 27220 6240 27430 6260
rect 27750 6250 27970 6270
rect 27750 6240 27960 6250
rect 27220 6230 27440 6240
rect 27230 6210 27440 6230
rect 27740 6220 27960 6240
rect 27740 6210 27950 6220
rect 27230 6200 27450 6210
rect 27240 6180 27450 6200
rect 27730 6190 27950 6210
rect 27730 6180 27940 6190
rect 27240 6170 27460 6180
rect 27250 6150 27460 6170
rect 27720 6160 27940 6180
rect 27720 6150 27930 6160
rect 27250 6140 27470 6150
rect 27260 6120 27470 6140
rect 27710 6130 27930 6150
rect 27710 6120 27920 6130
rect 27260 6100 27480 6120
rect 27270 6090 27480 6100
rect 27700 6100 27920 6120
rect 27700 6090 27910 6100
rect 27270 6080 27490 6090
rect 27280 6060 27490 6080
rect 27690 6070 27910 6090
rect 27690 6060 27900 6070
rect 27280 6050 27500 6060
rect 27290 6030 27500 6050
rect 27680 6040 27900 6060
rect 27680 6030 27890 6040
rect 27290 6020 27510 6030
rect 27300 6000 27510 6020
rect 27670 6010 27890 6030
rect 27670 6000 27880 6010
rect 26200 5800 26800 6000
rect 27300 5800 27880 6000
rect 26200 5500 26400 5800
rect 27300 5790 27510 5800
rect 27290 5770 27510 5790
rect 27670 5790 27880 5800
rect 27670 5770 27890 5790
rect 27290 5760 27500 5770
rect 27280 5740 27500 5760
rect 27680 5760 27890 5770
rect 27680 5740 27900 5760
rect 27280 5730 27490 5740
rect 27270 5710 27490 5730
rect 27690 5730 27900 5740
rect 27690 5710 27910 5730
rect 27270 5700 27480 5710
rect 27260 5680 27480 5700
rect 27700 5700 27910 5710
rect 27700 5680 27920 5700
rect 27260 5670 27470 5680
rect 27250 5650 27470 5670
rect 27710 5670 27920 5680
rect 27710 5650 27930 5670
rect 27250 5640 27460 5650
rect 27240 5620 27460 5640
rect 27720 5640 27930 5650
rect 27720 5620 27940 5640
rect 27240 5610 27450 5620
rect 27230 5590 27450 5610
rect 27730 5610 27940 5620
rect 27730 5590 27950 5610
rect 27230 5580 27440 5590
rect 27220 5560 27440 5580
rect 27740 5580 27950 5590
rect 27740 5560 27960 5580
rect 27220 5550 27430 5560
rect 27210 5530 27430 5550
rect 27750 5550 27960 5560
rect 27750 5530 27970 5550
rect 27210 5520 27420 5530
rect 27200 5500 27420 5520
rect 27760 5520 27970 5530
rect 28700 5540 28900 6500
rect 29400 5540 29600 6500
rect 28700 5520 28910 5540
rect 29390 5520 29600 5540
rect 27760 5500 27980 5520
rect 26200 5300 26900 5500
rect 27200 5470 27410 5500
rect 27770 5470 27980 5500
rect 28700 5510 28920 5520
rect 29380 5510 29600 5520
rect 28700 5500 28930 5510
rect 29370 5500 29600 5510
rect 28700 5490 29600 5500
rect 29900 6450 30140 6500
rect 30860 6450 31100 6500
rect 29900 6400 30180 6450
rect 30820 6400 31100 6450
rect 29900 6350 30220 6400
rect 30780 6350 31100 6400
rect 29900 6300 30260 6350
rect 30740 6300 31100 6350
rect 29900 6250 30300 6300
rect 30700 6250 31100 6300
rect 29900 6200 30340 6250
rect 30660 6200 31100 6250
rect 29900 6150 30380 6200
rect 30620 6150 31100 6200
rect 29900 6100 30420 6150
rect 30580 6100 31100 6150
rect 29900 6020 31100 6100
rect 27200 5440 27400 5470
rect 27780 5440 27980 5470
rect 28710 5450 29590 5490
rect 27200 5410 27390 5440
rect 27790 5410 27980 5440
rect 28720 5420 29580 5450
rect 27200 5380 27380 5410
rect 27800 5380 27980 5410
rect 28730 5400 29570 5420
rect 28740 5380 29560 5400
rect 27200 5350 27370 5380
rect 27810 5350 27980 5380
rect 28750 5370 29550 5380
rect 28760 5360 29540 5370
rect 28770 5350 29530 5360
rect 27200 5300 27360 5350
rect 27820 5300 27980 5350
rect 28780 5340 29520 5350
rect 28800 5330 29500 5340
rect 28820 5320 29480 5330
rect 28850 5310 29450 5320
rect 28890 5300 29410 5310
rect 29900 5300 30100 6020
rect 30260 5970 30740 6020
rect 30300 5920 30700 5970
rect 30340 5870 30660 5920
rect 30380 5820 30620 5870
rect 30420 5770 30580 5820
rect 30900 5300 31100 6020
rect 31400 6490 32060 6500
rect 32500 6490 33160 6500
rect 31400 6480 32090 6490
rect 32500 6480 33190 6490
rect 31400 6470 32110 6480
rect 32500 6470 33210 6480
rect 33960 6470 34360 6500
rect 31400 6460 32120 6470
rect 32500 6460 33220 6470
rect 31400 6450 32130 6460
rect 32500 6450 33230 6460
rect 31400 6440 32140 6450
rect 32500 6440 33240 6450
rect 33950 6440 34370 6470
rect 31400 6430 32150 6440
rect 32500 6430 33250 6440
rect 31400 6420 32160 6430
rect 32500 6420 33260 6430
rect 31400 6410 32170 6420
rect 32500 6410 33270 6420
rect 33940 6410 34380 6440
rect 31400 6390 32180 6410
rect 32500 6390 33280 6410
rect 31400 6370 32190 6390
rect 32500 6370 33290 6390
rect 33930 6380 34390 6410
rect 31400 6300 32200 6370
rect 31400 6000 31600 6300
rect 31970 6290 32200 6300
rect 31980 6280 32200 6290
rect 31990 6270 32200 6280
rect 32000 6250 32200 6270
rect 32010 6050 32200 6250
rect 32000 6030 32200 6050
rect 31990 6020 32200 6030
rect 31980 6010 32200 6020
rect 32500 6300 33300 6370
rect 33920 6350 34400 6380
rect 33910 6320 34410 6350
rect 31970 6000 32190 6010
rect 32500 6000 32700 6300
rect 33070 6290 33300 6300
rect 33900 6290 34080 6320
rect 33080 6280 33300 6290
rect 33090 6270 33300 6280
rect 33100 6250 33300 6270
rect 33890 6260 34080 6290
rect 34240 6290 34420 6320
rect 34240 6260 34430 6290
rect 33110 6050 33300 6250
rect 33880 6230 34060 6260
rect 33870 6200 34060 6230
rect 34260 6230 34440 6260
rect 34260 6200 34450 6230
rect 33860 6170 34040 6200
rect 33850 6140 34040 6170
rect 34280 6170 34460 6200
rect 34280 6140 34470 6170
rect 33840 6110 34020 6140
rect 33830 6080 34020 6110
rect 34300 6110 34480 6140
rect 34300 6080 34490 6110
rect 33820 6050 34000 6080
rect 33100 6030 33300 6050
rect 33090 6020 33300 6030
rect 33810 6020 34000 6050
rect 33080 6010 33300 6020
rect 33070 6000 33300 6010
rect 31400 5990 32180 6000
rect 32500 5990 33290 6000
rect 33800 5990 34000 6020
rect 31400 5820 32160 5990
rect 32500 5980 33280 5990
rect 32500 5970 33270 5980
rect 32500 5960 33260 5970
rect 33790 5960 34000 5990
rect 32500 5950 33250 5960
rect 31400 5810 32180 5820
rect 31400 5800 32190 5810
rect 32500 5800 33240 5950
rect 33780 5930 34000 5960
rect 33770 5900 34000 5930
rect 34320 6050 34500 6080
rect 34320 6020 34510 6050
rect 34320 5990 34520 6020
rect 35000 6000 35500 6800
rect 35700 6300 35900 7600
rect 36100 7560 36380 7600
rect 36100 7510 36420 7560
rect 36100 7460 36460 7510
rect 36100 7410 36500 7460
rect 36100 7360 36540 7410
rect 36100 7310 36580 7360
rect 36100 7260 36620 7310
rect 36100 7210 36660 7260
rect 36100 7160 36700 7210
rect 36100 7110 36740 7160
rect 36100 7100 36780 7110
rect 36100 6300 36300 7100
rect 36460 7060 36780 7100
rect 36460 7050 36820 7060
rect 36500 7010 36820 7050
rect 36500 7000 36860 7010
rect 36540 6960 36860 7000
rect 36540 6950 36900 6960
rect 36580 6910 36900 6950
rect 36580 6900 36940 6910
rect 36620 6860 36940 6900
rect 37100 6860 37300 7600
rect 36620 6850 37300 6860
rect 36660 6800 37300 6850
rect 36700 6750 37300 6800
rect 36740 6700 37300 6750
rect 36780 6650 37300 6700
rect 36820 6600 37300 6650
rect 36860 6550 37300 6600
rect 36900 6500 37300 6550
rect 36940 6450 37300 6500
rect 36980 6400 37300 6450
rect 37020 6350 37300 6400
rect 37060 6300 37300 6350
rect 37500 7500 37700 7800
rect 37500 7000 38000 7500
rect 37500 6990 47900 7000
rect 37500 6980 47920 6990
rect 37500 6970 47940 6980
rect 37500 6960 47950 6970
rect 37500 6950 47960 6960
rect 37500 6940 47970 6950
rect 37500 6920 47980 6940
rect 37500 6900 47990 6920
rect 37500 6800 48000 6900
rect 37500 6000 38000 6800
rect 40100 6460 40700 6500
rect 41300 6460 41700 6500
rect 40100 6400 40760 6460
rect 41240 6400 41760 6460
rect 34320 5960 34530 5990
rect 34320 5930 34540 5960
rect 34320 5900 34550 5930
rect 33760 5870 34560 5900
rect 33750 5840 34570 5870
rect 33740 5810 34580 5840
rect 31400 5500 31600 5800
rect 31970 5790 32200 5800
rect 31980 5780 32200 5790
rect 31990 5770 32200 5780
rect 32000 5750 32200 5770
rect 32010 5550 32200 5750
rect 32000 5530 32200 5550
rect 31990 5520 32200 5530
rect 31980 5510 32200 5520
rect 31970 5500 32200 5510
rect 31400 5440 32200 5500
rect 31400 5410 32190 5440
rect 31400 5390 32180 5410
rect 31400 5380 32170 5390
rect 31400 5370 32160 5380
rect 31400 5360 32150 5370
rect 31400 5350 32140 5360
rect 31400 5340 32130 5350
rect 31400 5330 32120 5340
rect 31400 5320 32110 5330
rect 31400 5310 32090 5320
rect 31400 5300 32060 5310
rect 32500 5300 32700 5800
rect 33040 5790 33240 5800
rect 33050 5780 33250 5790
rect 33730 5780 34590 5810
rect 33060 5760 33250 5780
rect 33070 5750 33250 5760
rect 33720 5750 34600 5780
rect 33070 5730 33260 5750
rect 33080 5710 33260 5730
rect 33710 5720 34610 5750
rect 33080 5690 33270 5710
rect 33700 5700 34620 5720
rect 33700 5690 33880 5700
rect 33090 5670 33270 5690
rect 33090 5650 33280 5670
rect 33690 5660 33880 5690
rect 34440 5690 34620 5700
rect 34440 5660 34630 5690
rect 33100 5630 33280 5650
rect 33680 5630 33860 5660
rect 33100 5610 33290 5630
rect 33110 5590 33290 5610
rect 33670 5600 33860 5630
rect 34460 5630 34640 5660
rect 34460 5600 34650 5630
rect 33110 5300 33300 5590
rect 33660 5570 33840 5600
rect 33650 5540 33840 5570
rect 34480 5570 34660 5600
rect 34480 5540 34670 5570
rect 33640 5510 33820 5540
rect 33630 5480 33820 5510
rect 34500 5510 34680 5540
rect 34500 5480 34690 5510
rect 35000 5500 38000 6000
rect 40000 6300 40800 6400
rect 41200 6360 41800 6400
rect 41140 6300 41860 6360
rect 40000 6230 40300 6300
rect 40000 6070 40200 6230
rect 40600 6200 40800 6300
rect 41100 6200 41400 6300
rect 41600 6200 41900 6300
rect 40000 6000 40300 6070
rect 40000 5900 40700 6000
rect 40100 5800 40800 5900
rect 40500 5730 40800 5800
rect 40000 5500 40200 5600
rect 40600 5570 40800 5730
rect 40500 5500 40800 5570
rect 41100 5600 41300 6200
rect 41700 5600 41900 6200
rect 41100 5500 41400 5600
rect 41600 5500 41900 5600
rect 42200 5500 42400 6500
rect 43200 6300 43900 6500
rect 44200 6450 44440 6500
rect 45160 6450 45400 6500
rect 44200 6400 44480 6450
rect 45120 6400 45400 6450
rect 44200 6350 44520 6400
rect 45080 6350 45400 6400
rect 44200 6300 44560 6350
rect 45040 6300 45400 6350
rect 43200 6000 43400 6300
rect 44200 6250 44600 6300
rect 45000 6250 45400 6300
rect 44200 6200 44640 6250
rect 44960 6200 45400 6250
rect 44200 6150 44680 6200
rect 44920 6150 45400 6200
rect 44200 6100 44720 6150
rect 44880 6100 45400 6150
rect 44200 6020 45400 6100
rect 43200 5800 43800 6000
rect 43200 5500 43400 5800
rect 33620 5460 33800 5480
rect 33600 5420 33800 5460
rect 34520 5460 34700 5480
rect 34520 5420 34720 5460
rect 33600 5360 33780 5420
rect 34540 5360 34720 5420
rect 33600 5300 33760 5360
rect 34560 5300 34720 5360
rect 35500 5000 36000 5500
rect 25500 4500 36000 5000
rect 37500 5000 37700 5500
rect 40000 5400 40800 5500
rect 41140 5440 41860 5500
rect 41200 5400 41800 5440
rect 40040 5340 40700 5400
rect 41240 5340 41760 5400
rect 40100 5300 40700 5340
rect 41300 5300 41700 5340
rect 42200 5300 42900 5500
rect 43200 5300 43900 5500
rect 44200 5300 44400 6020
rect 44560 5970 45040 6020
rect 44600 5920 45000 5970
rect 44640 5870 44960 5920
rect 44680 5820 44920 5870
rect 44720 5770 44880 5820
rect 45200 5300 45400 6020
rect 47500 6000 48000 6800
rect 47500 5800 49000 6000
rect 47500 5000 48000 5800
rect 37500 4500 48000 5000
rect 26000 4000 26500 4500
rect 24800 3900 26500 4000
rect 47300 4000 47500 4500
rect 48500 4000 49000 5800
rect 47300 3900 49000 4000
rect 24800 3880 26490 3900
rect 47310 3880 49000 3900
rect 24800 3860 26480 3880
rect 47320 3860 49000 3880
rect 24800 3850 26470 3860
rect 47330 3850 49000 3860
rect 24800 3840 26460 3850
rect 47340 3840 49000 3850
rect 24800 3830 26450 3840
rect 47350 3830 49000 3840
rect 24800 3820 26440 3830
rect 47370 3820 49000 3830
rect 24800 3810 26420 3820
rect 47380 3810 49000 3820
rect 24800 3800 26400 3810
rect 47400 3800 49000 3810
<< comment >>
rect -100 26000 49100 26100
rect -100 0 0 26000
rect 49000 0 49100 26000
rect -100 -100 49100 0
<< end >>
