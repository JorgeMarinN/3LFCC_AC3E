* NGSPICE file created from level_shifter.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_g5v0d10v5_PPR2BY a_n1077_n2026# a_129_n2000# a_503_n2026#
+ a_n445_n2026# a_603_n2000# a_1135_n2026# a_n919_n2026# a_n1551_n2026# a_1235_n2000#
+ a_345_n2026# a_n287_n2026# a_819_n2026# a_n1393_n2026# a_919_n2000# a_445_n2000#
+ a_187_n2026# a_n761_n2026# a_1077_n2000# a_1451_n2026# a_1551_n2000# a_287_n2000#
+ a_661_n2026# a_1293_n2026# a_761_n2000# a_n29_n2000# a_1393_n2000# a_977_n2026#
+ a_n1135_n2000# a_n503_n2000# a_n1609_n2000# a_n345_n2000# a_n819_n2000# a_n1451_n2000#
+ a_n187_n2000# a_n661_n2000# a_n1293_n2000# a_n977_n2000# a_29_n2026# a_n129_n2026#
+ a_n1235_n2026# a_n603_n2026# VSUBS
X0 a_129_n2000# a_29_n2026# a_n29_n2000# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=5.8e+12p pd=4.058e+07u as=5.8e+12p ps=4.058e+07u w=2e+07u l=500000u
X1 a_445_n2000# a_345_n2026# a_287_n2000# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=5.8e+12p pd=4.058e+07u as=5.8e+12p ps=4.058e+07u w=2e+07u l=500000u
X2 a_919_n2000# a_819_n2026# a_761_n2000# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=5.8e+12p pd=4.058e+07u as=5.8e+12p ps=4.058e+07u w=2e+07u l=500000u
X3 a_n1451_n2000# a_n1551_n2026# a_n1609_n2000# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=5.8e+12p pd=4.058e+07u as=5.8e+12p ps=4.058e+07u w=2e+07u l=500000u
X4 a_1077_n2000# a_977_n2026# a_919_n2000# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=5.8e+12p pd=4.058e+07u as=0p ps=0u w=2e+07u l=500000u
X5 a_n345_n2000# a_n445_n2026# a_n503_n2000# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=5.8e+12p pd=4.058e+07u as=5.8e+12p ps=4.058e+07u w=2e+07u l=500000u
X6 a_n819_n2000# a_n919_n2026# a_n977_n2000# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=5.8e+12p pd=4.058e+07u as=5.8e+12p ps=4.058e+07u w=2e+07u l=500000u
X7 a_n977_n2000# a_n1077_n2026# a_n1135_n2000# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=5.8e+12p ps=4.058e+07u w=2e+07u l=500000u
X8 a_1235_n2000# a_1135_n2026# a_1077_n2000# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=5.8e+12p pd=4.058e+07u as=0p ps=0u w=2e+07u l=500000u
X9 a_603_n2000# a_503_n2026# a_445_n2000# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=5.8e+12p pd=4.058e+07u as=0p ps=0u w=2e+07u l=500000u
X10 a_1393_n2000# a_1293_n2026# a_1235_n2000# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=5.8e+12p pd=4.058e+07u as=0p ps=0u w=2e+07u l=500000u
X11 a_761_n2000# a_661_n2026# a_603_n2000# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X12 a_n503_n2000# a_n603_n2026# a_n661_n2000# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=5.8e+12p ps=4.058e+07u w=2e+07u l=500000u
X13 a_287_n2000# a_187_n2026# a_129_n2000# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X14 a_n661_n2000# a_n761_n2026# a_n819_n2000# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X15 a_n1135_n2000# a_n1235_n2026# a_n1293_n2000# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=5.8e+12p ps=4.058e+07u w=2e+07u l=500000u
X16 a_n1293_n2000# a_n1393_n2026# a_n1451_n2000# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X17 a_n29_n2000# a_n129_n2026# a_n187_n2000# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=5.8e+12p ps=4.058e+07u w=2e+07u l=500000u
X18 a_1551_n2000# a_1451_n2026# a_1393_n2000# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=5.8e+12p pd=4.058e+07u as=0p ps=0u w=2e+07u l=500000u
X19 a_n187_n2000# a_n287_n2026# a_n345_n2000# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_VJVCZ4 a_n1077_n2026# a_129_n2000# a_503_n2026#
+ a_n445_n2026# a_603_n2000# a_1135_n2026# a_n919_n2026# a_n1551_n2026# a_1235_n2000#
+ a_345_n2026# a_n287_n2026# a_819_n2026# a_n1393_n2026# a_919_n2000# a_445_n2000#
+ a_187_n2026# a_n761_n2026# a_1077_n2000# a_1451_n2026# a_1551_n2000# a_287_n2000#
+ a_661_n2026# a_1293_n2026# a_761_n2000# a_n29_n2000# a_1393_n2000# a_977_n2026#
+ a_n1135_n2000# a_n503_n2000# a_n1609_n2000# a_n345_n2000# a_n819_n2000# a_n1451_n2000#
+ a_n187_n2000# a_n661_n2000# a_n1293_n2000# a_n977_n2000# a_29_n2026# a_n129_n2026#
+ a_n1235_n2026# a_n603_n2026# w_n1645_n2062#
X0 a_n187_n2000# a_n287_n2026# a_n345_n2000# w_n1645_n2062# sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+12p pd=4.058e+07u as=5.8e+12p ps=4.058e+07u w=2e+07u l=500000u
X1 a_129_n2000# a_29_n2026# a_n29_n2000# w_n1645_n2062# sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+12p pd=4.058e+07u as=5.8e+12p ps=4.058e+07u w=2e+07u l=500000u
X2 a_445_n2000# a_345_n2026# a_287_n2000# w_n1645_n2062# sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+12p pd=4.058e+07u as=5.8e+12p ps=4.058e+07u w=2e+07u l=500000u
X3 a_919_n2000# a_819_n2026# a_761_n2000# w_n1645_n2062# sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+12p pd=4.058e+07u as=5.8e+12p ps=4.058e+07u w=2e+07u l=500000u
X4 a_n1451_n2000# a_n1551_n2026# a_n1609_n2000# w_n1645_n2062# sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+12p pd=4.058e+07u as=5.8e+12p ps=4.058e+07u w=2e+07u l=500000u
X5 a_1077_n2000# a_977_n2026# a_919_n2000# w_n1645_n2062# sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+12p pd=4.058e+07u as=0p ps=0u w=2e+07u l=500000u
X6 a_n345_n2000# a_n445_n2026# a_n503_n2000# w_n1645_n2062# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=5.8e+12p ps=4.058e+07u w=2e+07u l=500000u
X7 a_n977_n2000# a_n1077_n2026# a_n1135_n2000# w_n1645_n2062# sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+12p pd=4.058e+07u as=5.8e+12p ps=4.058e+07u w=2e+07u l=500000u
X8 a_n819_n2000# a_n919_n2026# a_n977_n2000# w_n1645_n2062# sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+12p pd=4.058e+07u as=0p ps=0u w=2e+07u l=500000u
X9 a_1235_n2000# a_1135_n2026# a_1077_n2000# w_n1645_n2062# sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+12p pd=4.058e+07u as=0p ps=0u w=2e+07u l=500000u
X10 a_603_n2000# a_503_n2026# a_445_n2000# w_n1645_n2062# sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+12p pd=4.058e+07u as=0p ps=0u w=2e+07u l=500000u
X11 a_1393_n2000# a_1293_n2026# a_1235_n2000# w_n1645_n2062# sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+12p pd=4.058e+07u as=0p ps=0u w=2e+07u l=500000u
X12 a_761_n2000# a_661_n2026# a_603_n2000# w_n1645_n2062# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X13 a_n503_n2000# a_n603_n2026# a_n661_n2000# w_n1645_n2062# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=5.8e+12p ps=4.058e+07u w=2e+07u l=500000u
X14 a_287_n2000# a_187_n2026# a_129_n2000# w_n1645_n2062# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X15 a_n661_n2000# a_n761_n2026# a_n819_n2000# w_n1645_n2062# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X16 a_n1135_n2000# a_n1235_n2026# a_n1293_n2000# w_n1645_n2062# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=5.8e+12p ps=4.058e+07u w=2e+07u l=500000u
X17 a_n1293_n2000# a_n1393_n2026# a_n1451_n2000# w_n1645_n2062# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X18 a_n29_n2000# a_n129_n2026# a_n187_n2000# w_n1645_n2062# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X19 a_1551_n2000# a_1451_n2026# a_1393_n2000# w_n1645_n2062# sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+12p pd=4.058e+07u as=0p ps=0u w=2e+07u l=500000u
.ends

.subckt inv_400 a_n166_32166# w_n304_36844# cont_poly_min_9/VSUBS IN
Xsky130_fd_pr__nfet_g5v0d10v5_PPR2BY_0 IN OUT IN IN cont_poly_min_9/VSUBS IN IN IN
+ cont_poly_min_9/VSUBS IN IN IN IN cont_poly_min_9/VSUBS OUT IN IN OUT IN cont_poly_min_9/VSUBS
+ cont_poly_min_9/VSUBS IN IN OUT cont_poly_min_9/VSUBS OUT IN OUT OUT cont_poly_min_9/VSUBS
+ cont_poly_min_9/VSUBS OUT OUT OUT cont_poly_min_9/VSUBS cont_poly_min_9/VSUBS cont_poly_min_9/VSUBS
+ IN IN IN IN cont_poly_min_9/VSUBS sky130_fd_pr__nfet_g5v0d10v5_PPR2BY
Xsky130_fd_pr__pfet_g5v0d10v5_VJVCZ4_0 IN OUT IN IN w_n304_36844# IN IN IN w_n304_36844#
+ IN IN IN IN w_n304_36844# OUT IN IN OUT IN w_n304_36844# w_n304_36844# IN IN OUT
+ w_n304_36844# OUT IN OUT OUT w_n304_36844# w_n304_36844# OUT OUT OUT w_n304_36844#
+ w_n304_36844# w_n304_36844# IN IN IN IN w_n304_36844# sky130_fd_pr__pfet_g5v0d10v5_VJVCZ4
.ends

.subckt sky130_fd_pr__nfet_01v8_RBMM6F a_207_n100# a_n207_n126# a_81_n126# a_15_n100#
+ a_n177_n100# a_111_n100# a_n15_n126# a_n111_n126# a_n81_n100# a_177_n126# a_n269_n100#
+ VSUBS
X0 a_207_n100# a_177_n126# a_111_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X1 a_15_n100# a_n15_n126# a_n81_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X2 a_111_n100# a_81_n126# a_15_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_n81_n100# a_n111_n126# a_n177_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X4 a_n177_n100# a_n207_n126# a_n269_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_5S5LDE a_207_n100# a_177_n131# a_81_n126# a_15_n100#
+ a_n177_n100# a_111_n100# a_n111_n126# a_n207_n131# w_n305_n200# a_n81_n100# a_n15_n131#
+ a_n269_n100#
X0 a_207_n100# a_177_n131# a_111_n100# w_n305_n200# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X1 a_15_n100# a_n15_n131# a_n81_n100# w_n305_n200# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X2 a_111_n100# a_81_n126# a_15_n100# w_n305_n200# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_n81_n100# a_n111_n126# a_n177_n100# w_n305_n200# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X4 a_n177_n100# a_n207_n131# a_n269_n100# w_n305_n200# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
.ends

.subckt inv_1_8 OUT VDD IN GND
Xsky130_fd_pr__nfet_01v8_RBMM6F_0 OUT IN IN OUT OUT GND IN IN GND IN GND GND sky130_fd_pr__nfet_01v8_RBMM6F
Xsky130_fd_pr__pfet_01v8_5S5LDE_0 OUT IN IN OUT OUT VDD IN IN VDD VDD IN VDD sky130_fd_pr__pfet_01v8_5S5LDE
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_PVZBWB a_n503_n1000# a_n345_n1000# a_n819_n1000#
+ a_n187_n1000# a_n661_n1000# a_29_n1026# a_n129_n1026# a_n603_n1026# a_129_n1000#
+ a_503_n1026# a_n445_n1026# a_603_n1000# a_345_n1026# a_n287_n1026# a_445_n1000#
+ a_n761_n1026# a_187_n1026# a_287_n1000# a_661_n1026# a_761_n1000# a_n29_n1000# VSUBS
X0 a_445_n1000# a_345_n1026# a_287_n1000# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+12p pd=2.058e+07u as=2.9e+12p ps=2.058e+07u w=1e+07u l=500000u
X1 a_n503_n1000# a_n603_n1026# a_n661_n1000# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+12p pd=2.058e+07u as=2.9e+12p ps=2.058e+07u w=1e+07u l=500000u
X2 a_n29_n1000# a_n129_n1026# a_n187_n1000# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+12p pd=2.058e+07u as=2.9e+12p ps=2.058e+07u w=1e+07u l=500000u
X3 a_603_n1000# a_503_n1026# a_445_n1000# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+12p pd=2.058e+07u as=0p ps=0u w=1e+07u l=500000u
X4 a_n661_n1000# a_n761_n1026# a_n819_n1000# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=2.9e+12p ps=2.058e+07u w=1e+07u l=500000u
X5 a_n187_n1000# a_n287_n1026# a_n345_n1000# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=2.9e+12p ps=2.058e+07u w=1e+07u l=500000u
X6 a_761_n1000# a_661_n1026# a_603_n1000# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+12p pd=2.058e+07u as=0p ps=0u w=1e+07u l=500000u
X7 a_287_n1000# a_187_n1026# a_129_n1000# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=2.9e+12p ps=2.058e+07u w=1e+07u l=500000u
X8 a_n345_n1000# a_n445_n1026# a_n503_n1000# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+07u l=500000u
X9 a_129_n1000# a_29_n1026# a_n29_n1000# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+07u l=500000u
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_VEZS85 a_n503_n1000# a_n345_n1000# a_n819_n1000#
+ a_n187_n1000# a_n661_n1000# a_29_n1026# a_n129_n1026# a_n603_n1026# a_129_n1000#
+ a_503_n1026# a_n445_n1026# w_n855_n1062# a_603_n1000# a_345_n1026# a_n287_n1026#
+ a_445_n1000# a_n761_n1026# a_187_n1026# a_287_n1000# a_661_n1026# a_761_n1000# a_n29_n1000#
X0 a_129_n1000# a_29_n1026# a_n29_n1000# w_n855_n1062# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+12p pd=2.058e+07u as=2.9e+12p ps=2.058e+07u w=1e+07u l=500000u
X1 a_445_n1000# a_345_n1026# a_287_n1000# w_n855_n1062# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+12p pd=2.058e+07u as=2.9e+12p ps=2.058e+07u w=1e+07u l=500000u
X2 a_n503_n1000# a_n603_n1026# a_n661_n1000# w_n855_n1062# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+12p pd=2.058e+07u as=2.9e+12p ps=2.058e+07u w=1e+07u l=500000u
X3 a_n29_n1000# a_n129_n1026# a_n187_n1000# w_n855_n1062# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+12p ps=2.058e+07u w=1e+07u l=500000u
X4 a_603_n1000# a_503_n1026# a_445_n1000# w_n855_n1062# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+12p pd=2.058e+07u as=0p ps=0u w=1e+07u l=500000u
X5 a_n661_n1000# a_n761_n1026# a_n819_n1000# w_n855_n1062# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+12p ps=2.058e+07u w=1e+07u l=500000u
X6 a_n187_n1000# a_n287_n1026# a_n345_n1000# w_n855_n1062# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+12p ps=2.058e+07u w=1e+07u l=500000u
X7 a_761_n1000# a_661_n1026# a_603_n1000# w_n855_n1062# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+12p pd=2.058e+07u as=0p ps=0u w=1e+07u l=500000u
X8 a_287_n1000# a_187_n1026# a_129_n1000# w_n855_n1062# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+07u l=500000u
X9 a_n345_n1000# a_n445_n1026# a_n503_n1000# w_n855_n1062# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+07u l=500000u
.ends

.subckt stage_100 OUT B a_924_n78# VH GND
Xsky130_fd_pr__nfet_g5v0d10v5_PVZBWB_0 GND OUT GND GND OUT B B B GND B B OUT B B GND
+ B B OUT B GND OUT GND sky130_fd_pr__nfet_g5v0d10v5_PVZBWB
Xsky130_fd_pr__pfet_g5v0d10v5_VEZS85_0 VH OUT VH VH OUT a_924_n78# a_924_n78# a_924_n78#
+ VH a_924_n78# a_924_n78# VH OUT a_924_n78# a_924_n78# VH a_924_n78# a_924_n78# OUT
+ a_924_n78# VH OUT sky130_fd_pr__pfet_g5v0d10v5_VEZS85
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_BUUKVD a_n108_n164# a_n50_n261# a_50_n164# w_n144_n264#
X0 a_50_n164# a_n50_n261# a_n108_n164# w_n144_n264# sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_C7Z2GC a_208_n400# a_108_n426# a_n208_n426# a_50_n400#
+ a_n50_n426# a_n108_n400# a_n266_n400# VSUBS
X0 a_50_n400# a_n50_n426# a_n108_n400# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X1 a_n108_n400# a_n208_n426# a_n266_n400# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X2 a_208_n400# a_108_n426# a_50_n400# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4e+06u l=500000u
.ends

.subckt cruzados OUT cont_poly_min_6/VSUBS VH IN2 IN1
Xsky130_fd_pr__pfet_g5v0d10v5_BUUKVD_0 VH m1_108_n44# OUT VH sky130_fd_pr__pfet_g5v0d10v5_BUUKVD
Xsky130_fd_pr__pfet_g5v0d10v5_BUUKVD_1 VH OUT m1_108_n44# VH sky130_fd_pr__pfet_g5v0d10v5_BUUKVD
Xsky130_fd_pr__nfet_g5v0d10v5_C7Z2GC_0 OUT IN1 IN1 cont_poly_min_6/VSUBS IN1 OUT cont_poly_min_6/VSUBS
+ cont_poly_min_6/VSUBS sky130_fd_pr__nfet_g5v0d10v5_C7Z2GC
Xsky130_fd_pr__nfet_g5v0d10v5_C7Z2GC_1 m1_108_n44# IN2 IN2 cont_poly_min_6/VSUBS IN2
+ m1_108_n44# cont_poly_min_6/VSUBS cont_poly_min_6/VSUBS sky130_fd_pr__nfet_g5v0d10v5_C7Z2GC
.ends


* Top level circuit level_shifter

Xinv_400_0 GND VH GND inv_400_0/IN inv_400
Xinv_1_8_0 inv_1_8_0/OUT VDD IN GND inv_1_8
Xstage_100_0 inv_400_0/IN IN cruzados_0/OUT VH GND stage_100
Xcruzados_0 cruzados_0/OUT GND VH IN inv_1_8_0/OUT cruzados
.end

