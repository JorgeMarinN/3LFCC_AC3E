magic
tech sky130A
magscale 1 2
timestamp 1663277475
<< nwell >>
rect -10 839 600 1019
<< psubdiff >>
rect 71 29 95 68
rect 510 29 534 68
<< nsubdiff >>
rect 33 850 100 884
rect 489 850 560 884
<< psubdiffcont >>
rect 95 29 510 68
<< nsubdiffcont >>
rect 100 850 489 884
<< poly >>
rect 88 292 118 603
rect 184 286 214 613
rect 280 287 310 614
rect 376 285 406 612
rect 472 286 502 613
<< viali >>
rect 27 884 562 885
rect 27 850 100 884
rect 100 850 489 884
rect 489 850 562 884
rect 27 849 562 850
rect 30 68 552 71
rect 30 29 95 68
rect 95 29 510 68
rect 510 29 552 68
rect 30 25 552 29
<< metal1 >>
rect 15 885 574 891
rect 15 849 27 885
rect 562 849 574 885
rect 15 843 574 849
rect 38 776 72 843
rect 230 776 264 843
rect 422 775 456 843
rect 35 494 45 546
rect 97 494 107 546
rect 136 406 166 621
rect 211 495 221 547
rect 273 495 283 547
rect 328 406 358 622
rect 404 497 414 549
rect 466 497 476 549
rect 520 407 550 622
rect 116 354 126 406
rect 178 354 188 406
rect 308 354 318 406
rect 370 354 380 406
rect 499 355 509 407
rect 561 355 571 407
rect 136 294 166 354
rect 328 286 358 354
rect 520 286 550 355
rect 38 77 72 132
rect 230 77 264 132
rect 422 77 456 133
rect 18 71 564 77
rect 18 25 30 71
rect 552 25 564 71
rect 18 19 564 25
<< via1 >>
rect 45 494 97 546
rect 221 495 273 547
rect 414 497 466 549
rect 126 354 178 406
rect 318 354 370 406
rect 509 355 561 407
<< metal2 >>
rect 45 546 97 556
rect -10 507 45 535
rect 221 547 273 557
rect 97 507 221 535
rect 45 484 97 494
rect 414 549 466 559
rect 273 507 414 535
rect 221 485 273 495
rect 466 507 600 535
rect 414 487 466 497
rect 126 406 178 416
rect -11 367 126 395
rect 318 406 370 416
rect 178 367 318 395
rect 126 344 178 354
rect 509 407 561 417
rect 370 367 509 395
rect 318 344 370 354
rect 561 367 600 395
rect 509 345 561 355
use cont_poly_min  cont_poly_min_0
timestamp 1663264347
transform 1 0 71 0 1 444
box -33 33 33 99
use cont_poly_min  cont_poly_min_1
timestamp 1663264347
transform 1 0 247 0 1 444
box -33 33 33 99
use cont_poly_min  cont_poly_min_2
timestamp 1663264347
transform 1 0 439 0 1 447
box -33 33 33 99
use sky130_fd_pr__nfet_01v8_RBMM6F  sky130_fd_pr__nfet_01v8_RBMM6F_0
timestamp 1663264347
transform 1 0 295 0 1 226
box -269 -126 269 126
use sky130_fd_pr__pfet_01v8_5S5LDE  sky130_fd_pr__pfet_01v8_5S5LDE_0
timestamp 1663269594
transform 1 0 295 0 1 677
box -305 -200 305 200
<< labels >>
rlabel metal1 18 19 564 25 1 GND
rlabel metal2 561 367 600 395 1 OUT
rlabel metal2 -10 507 45 535 1 IN
rlabel metal1 15 885 574 891 1 VDD
<< end >>
