magic
tech sky130A
timestamp 1667693123
<< metal1 >>
rect 1000 166980 68990 167000
rect 1000 166020 1020 166980
rect 68970 166020 68990 166980
rect 1000 165720 68990 166020
rect -590 165700 68990 165720
rect -590 143730 -570 165700
rect 9390 164000 68990 165700
rect 71000 166980 136000 167000
rect 71000 166020 71200 166980
rect 135960 166020 136000 166980
rect 71000 164000 136000 166020
rect 9390 161000 9410 164000
rect 22000 161000 25000 164000
rect 9390 158000 25000 161000
rect 9390 155000 9410 158000
rect 36000 155000 39000 164000
rect 9390 152000 39000 155000
rect 9390 149000 9410 152000
rect 51000 149000 54000 164000
rect 9390 146000 54000 149000
rect 9390 143730 9410 146000
rect -590 143710 9410 143730
rect 71000 122000 74000 164000
rect 1000 121060 74000 122000
rect -590 121040 74000 121060
rect -590 99070 -570 121040
rect 9390 119000 74000 121040
rect 9390 118000 9410 119000
rect 82000 118000 85000 164000
rect 9390 115000 85000 118000
rect 9390 114000 9410 115000
rect 93000 114000 96000 164000
rect 9390 111000 96000 114000
rect 9390 110000 9410 111000
rect 104000 110000 107000 164000
rect 9390 107000 107000 110000
rect 9390 106000 9410 107000
rect 115000 106000 118000 164000
rect 9390 103000 118000 106000
rect 9390 102000 9410 103000
rect 126000 102000 129000 164000
rect 9390 99070 129000 102000
rect -590 99050 129000 99070
rect 9000 99000 129000 99050
<< via1 >>
rect 1020 166020 68970 166980
rect -570 143730 9390 165700
rect 71200 166020 135960 166980
rect -570 99070 9390 121040
<< metal2 >>
rect 1000 166980 68990 167000
rect 1000 166020 1020 166980
rect 68970 166020 68990 166980
rect 1000 165720 68990 166020
rect -590 165700 68990 165720
rect -590 143730 -570 165700
rect 9390 164000 68990 165700
rect 71000 166980 136000 167000
rect 71000 166020 71200 166980
rect 135960 166020 136000 166980
rect 71000 164000 136000 166020
rect 9390 161000 9410 164000
rect 22000 161000 25000 164000
rect 9390 158000 25000 161000
rect 9390 155000 9410 158000
rect 36000 155000 39000 164000
rect 9390 152000 39000 155000
rect 9390 149000 9410 152000
rect 51000 149000 54000 164000
rect 9390 146000 54000 149000
rect 9390 143730 9410 146000
rect -590 143710 9410 143730
rect 71000 122000 74000 164000
rect 1000 121060 74000 122000
rect -590 121040 74000 121060
rect -590 99070 -570 121040
rect 9390 119000 74000 121040
rect 9390 118000 9410 119000
rect 82000 118000 85000 164000
rect 9390 115000 85000 118000
rect 9390 114000 9410 115000
rect 93000 114000 96000 164000
rect 9390 111000 96000 114000
rect 9390 110000 9410 111000
rect 104000 110000 107000 164000
rect 9390 107000 107000 110000
rect 9390 106000 9410 107000
rect 115000 106000 118000 164000
rect 9390 103000 118000 106000
rect 9390 102000 9410 103000
rect 126000 102000 129000 164000
rect 9390 99070 129000 102000
rect -590 99050 129000 99070
rect 9000 99000 129000 99050
<< via2 >>
rect 1020 166020 68970 166980
rect -570 143730 9390 165700
rect 71200 166020 135960 166980
rect -570 99070 9390 121040
<< metal3 >>
rect 71180 167030 135980 168000
rect 1000 166980 68990 167000
rect 1000 166020 1020 166980
rect 68970 166020 68990 166980
rect 1000 165880 68990 166020
rect 71180 166020 71200 167030
rect 135960 166020 135980 167030
rect 71180 166000 135980 166020
rect 1000 165720 2000 165880
rect 4190 165720 5190 165880
rect 7380 165720 8380 165880
rect -590 165700 9410 165720
rect -590 143730 -570 165700
rect 9390 164690 9410 165700
rect 9390 163690 9570 164690
rect 9390 161500 9410 163690
rect 9390 160500 9570 161500
rect 9390 158310 9410 160500
rect 9390 157310 9570 158310
rect 9390 155120 9410 157310
rect 9390 154120 9570 155120
rect 9390 151930 9410 154120
rect 9390 150930 9570 151930
rect 9390 148740 9410 150930
rect 9390 147740 9570 148740
rect 9390 145550 9410 147740
rect 9390 144550 9570 145550
rect 9390 143730 9410 144550
rect -590 143710 9410 143730
rect 1000 143550 2000 143710
rect 4190 143550 5190 143710
rect 7380 143550 8380 143710
rect -590 121040 9410 121060
rect -590 99070 -570 121040
rect 9390 99070 9410 121040
rect -590 99050 9410 99070
<< via3 >>
rect 1020 166020 68970 166980
rect 71200 166980 135960 167030
rect 71200 166070 135960 166980
rect -570 143730 9390 165700
rect -570 99070 9390 121040
<< metal4 >>
rect 1000 166980 68990 168000
rect 1000 166020 1020 166980
rect 68970 166020 68990 166980
rect 1000 166000 68990 166020
rect 71180 167030 135980 167050
rect 71180 166070 71200 167030
rect 135960 166070 135980 167030
rect 71180 165880 135980 166070
rect -590 165700 9410 165720
rect -590 143730 -570 165700
rect 9390 143730 9410 165700
rect -590 143710 9410 143730
rect 1000 121060 2000 121220
rect 4190 121060 5190 121220
rect 7380 121060 8380 121220
rect -590 121040 9410 121060
rect -590 99070 -570 121040
rect 9390 120030 9410 121040
rect 9390 119030 9570 120030
rect 9390 116840 9410 119030
rect 9390 115840 9570 116840
rect 9390 113650 9410 115840
rect 9390 112650 9570 113650
rect 9390 110460 9410 112650
rect 9390 109460 9570 110460
rect 9390 107270 9410 109460
rect 9390 106270 9570 107270
rect 9390 104080 9410 106270
rect 9390 103080 9570 104080
rect 9390 100890 9410 103080
rect 9390 99890 9570 100890
rect 9390 99070 9410 99890
rect -590 99050 9410 99070
rect 1000 98890 2000 99050
rect 4190 98890 5190 99050
rect 7380 98890 8380 99050
<< via4 >>
rect 1020 166020 68970 166980
rect 71200 166070 135960 167030
rect -570 143730 9390 165700
rect -570 99070 9390 121040
<< metal5 >>
rect 71180 167030 135980 168000
rect 1000 166980 68990 167000
rect 1000 166020 1020 166980
rect 68970 166020 68990 166980
rect 71180 166070 71200 167030
rect 135960 166070 135980 167030
rect 71180 166050 135980 166070
rect 1000 165880 68990 166020
rect 1000 165720 2000 165880
rect 4190 165720 5190 165880
rect 7380 165720 8380 165880
rect -590 165700 9410 165720
rect -590 143730 -570 165700
rect 9390 164690 9410 165700
rect 9390 163690 9570 164690
rect 9390 161500 9410 163690
rect 9390 160500 9570 161500
rect 9390 158310 9410 160500
rect 9390 157310 9570 158310
rect 9390 155120 9410 157310
rect 9390 154120 9570 155120
rect 9390 151930 9410 154120
rect 9390 150930 9570 151930
rect 9390 148740 9410 150930
rect 9390 147740 9570 148740
rect 9390 145550 9410 147740
rect 9390 144550 9570 145550
rect 9390 143730 9410 144550
rect -590 143710 9410 143730
rect 1000 143550 2000 143710
rect 4190 143550 5190 143710
rect 7380 143550 8380 143710
rect -590 121040 9410 121060
rect -590 99070 -570 121040
rect 9390 99070 9410 121040
rect -590 99050 9410 99070
use unit_cap  unit_cap_0
timestamp 1662145021
transform 1 0 0 0 1 0
box 0 0 3190 3190
use unit_cap  unit_cap_1
timestamp 1662145021
transform 1 0 0 0 1 3190
box 0 0 3190 3190
use unit_cap  unit_cap_2
timestamp 1662145021
transform 1 0 0 0 1 6380
box 0 0 3190 3190
use unit_cap  unit_cap_3
timestamp 1662145021
transform 1 0 0 0 1 9570
box 0 0 3190 3190
use unit_cap  unit_cap_4
timestamp 1662145021
transform 1 0 0 0 1 12760
box 0 0 3190 3190
use unit_cap  unit_cap_5
timestamp 1662145021
transform 1 0 0 0 1 15950
box 0 0 3190 3190
use unit_cap  unit_cap_6
timestamp 1662145021
transform 1 0 0 0 1 19140
box 0 0 3190 3190
use unit_cap  unit_cap_7
timestamp 1662145021
transform 1 0 0 0 1 22330
box 0 0 3190 3190
use unit_cap  unit_cap_8
timestamp 1662145021
transform 1 0 0 0 1 25520
box 0 0 3190 3190
use unit_cap  unit_cap_9
timestamp 1662145021
transform 1 0 0 0 1 28710
box 0 0 3190 3190
use unit_cap  unit_cap_10
timestamp 1662145021
transform 1 0 0 0 1 31900
box 0 0 3190 3190
use unit_cap  unit_cap_11
timestamp 1662145021
transform 1 0 0 0 1 35090
box 0 0 3190 3190
use unit_cap  unit_cap_12
timestamp 1662145021
transform 1 0 0 0 1 38280
box 0 0 3190 3190
use unit_cap  unit_cap_13
timestamp 1662145021
transform 1 0 0 0 1 41470
box 0 0 3190 3190
use unit_cap  unit_cap_14
timestamp 1662145021
transform 1 0 0 0 1 44660
box 0 0 3190 3190
use unit_cap  unit_cap_15
timestamp 1662145021
transform 1 0 0 0 1 47850
box 0 0 3190 3190
use unit_cap  unit_cap_16
timestamp 1662145021
transform 1 0 0 0 1 51040
box 0 0 3190 3190
use unit_cap  unit_cap_17
timestamp 1662145021
transform 1 0 0 0 1 54230
box 0 0 3190 3190
use unit_cap  unit_cap_18
timestamp 1662145021
transform 1 0 0 0 1 57420
box 0 0 3190 3190
use unit_cap  unit_cap_19
timestamp 1662145021
transform 1 0 0 0 1 60610
box 0 0 3190 3190
use unit_cap  unit_cap_20
timestamp 1662145021
transform 1 0 0 0 1 63800
box 0 0 3190 3190
use unit_cap  unit_cap_21
timestamp 1662145021
transform 1 0 0 0 1 66990
box 0 0 3190 3190
use unit_cap  unit_cap_22
timestamp 1662145021
transform 1 0 0 0 1 70180
box 0 0 3190 3190
use unit_cap  unit_cap_23
timestamp 1662145021
transform 1 0 0 0 1 73370
box 0 0 3190 3190
use unit_cap  unit_cap_24
timestamp 1662145021
transform 1 0 0 0 1 76560
box 0 0 3190 3190
use unit_cap  unit_cap_25
timestamp 1662145021
transform 1 0 0 0 1 79750
box 0 0 3190 3190
use unit_cap  unit_cap_26
timestamp 1662145021
transform 1 0 0 0 1 82940
box 0 0 3190 3190
use unit_cap  unit_cap_27
timestamp 1662145021
transform 1 0 0 0 1 86130
box 0 0 3190 3190
use unit_cap  unit_cap_28
timestamp 1662145021
transform 1 0 0 0 1 89320
box 0 0 3190 3190
use unit_cap  unit_cap_29
timestamp 1662145021
transform 1 0 0 0 1 92510
box 0 0 3190 3190
use unit_cap  unit_cap_30
timestamp 1662145021
transform 1 0 0 0 1 95700
box 0 0 3190 3190
use unit_cap  unit_cap_38
timestamp 1662145021
transform 1 0 0 0 1 121220
box 0 0 3190 3190
use unit_cap  unit_cap_39
timestamp 1662145021
transform 1 0 0 0 1 124410
box 0 0 3190 3190
use unit_cap  unit_cap_40
timestamp 1662145021
transform 1 0 0 0 1 127600
box 0 0 3190 3190
use unit_cap  unit_cap_41
timestamp 1662145021
transform 1 0 0 0 1 130790
box 0 0 3190 3190
use unit_cap  unit_cap_42
timestamp 1662145021
transform 1 0 0 0 1 133980
box 0 0 3190 3190
use unit_cap  unit_cap_43
timestamp 1662145021
transform 1 0 0 0 1 137170
box 0 0 3190 3190
use unit_cap  unit_cap_44
timestamp 1662145021
transform 1 0 0 0 1 140360
box 0 0 3190 3190
use unit_cap  unit_cap_52
timestamp 1662145021
transform 1 0 3190 0 1 0
box 0 0 3190 3190
use unit_cap  unit_cap_53
timestamp 1662145021
transform 1 0 3190 0 1 3190
box 0 0 3190 3190
use unit_cap  unit_cap_54
timestamp 1662145021
transform 1 0 3190 0 1 6380
box 0 0 3190 3190
use unit_cap  unit_cap_55
timestamp 1662145021
transform 1 0 3190 0 1 9570
box 0 0 3190 3190
use unit_cap  unit_cap_56
timestamp 1662145021
transform 1 0 3190 0 1 12760
box 0 0 3190 3190
use unit_cap  unit_cap_57
timestamp 1662145021
transform 1 0 3190 0 1 15950
box 0 0 3190 3190
use unit_cap  unit_cap_58
timestamp 1662145021
transform 1 0 3190 0 1 19140
box 0 0 3190 3190
use unit_cap  unit_cap_59
timestamp 1662145021
transform 1 0 3190 0 1 22330
box 0 0 3190 3190
use unit_cap  unit_cap_60
timestamp 1662145021
transform 1 0 3190 0 1 25520
box 0 0 3190 3190
use unit_cap  unit_cap_61
timestamp 1662145021
transform 1 0 3190 0 1 28710
box 0 0 3190 3190
use unit_cap  unit_cap_62
timestamp 1662145021
transform 1 0 3190 0 1 31900
box 0 0 3190 3190
use unit_cap  unit_cap_63
timestamp 1662145021
transform 1 0 3190 0 1 35090
box 0 0 3190 3190
use unit_cap  unit_cap_64
timestamp 1662145021
transform 1 0 3190 0 1 38280
box 0 0 3190 3190
use unit_cap  unit_cap_65
timestamp 1662145021
transform 1 0 3190 0 1 41470
box 0 0 3190 3190
use unit_cap  unit_cap_66
timestamp 1662145021
transform 1 0 3190 0 1 44660
box 0 0 3190 3190
use unit_cap  unit_cap_67
timestamp 1662145021
transform 1 0 3190 0 1 47850
box 0 0 3190 3190
use unit_cap  unit_cap_68
timestamp 1662145021
transform 1 0 3190 0 1 51040
box 0 0 3190 3190
use unit_cap  unit_cap_69
timestamp 1662145021
transform 1 0 3190 0 1 54230
box 0 0 3190 3190
use unit_cap  unit_cap_70
timestamp 1662145021
transform 1 0 3190 0 1 57420
box 0 0 3190 3190
use unit_cap  unit_cap_71
timestamp 1662145021
transform 1 0 3190 0 1 60610
box 0 0 3190 3190
use unit_cap  unit_cap_72
timestamp 1662145021
transform 1 0 3190 0 1 63800
box 0 0 3190 3190
use unit_cap  unit_cap_73
timestamp 1662145021
transform 1 0 3190 0 1 66990
box 0 0 3190 3190
use unit_cap  unit_cap_74
timestamp 1662145021
transform 1 0 3190 0 1 70180
box 0 0 3190 3190
use unit_cap  unit_cap_75
timestamp 1662145021
transform 1 0 3190 0 1 73370
box 0 0 3190 3190
use unit_cap  unit_cap_76
timestamp 1662145021
transform 1 0 3190 0 1 76560
box 0 0 3190 3190
use unit_cap  unit_cap_77
timestamp 1662145021
transform 1 0 3190 0 1 79750
box 0 0 3190 3190
use unit_cap  unit_cap_78
timestamp 1662145021
transform 1 0 3190 0 1 82940
box 0 0 3190 3190
use unit_cap  unit_cap_79
timestamp 1662145021
transform 1 0 3190 0 1 86130
box 0 0 3190 3190
use unit_cap  unit_cap_80
timestamp 1662145021
transform 1 0 3190 0 1 89320
box 0 0 3190 3190
use unit_cap  unit_cap_81
timestamp 1662145021
transform 1 0 3190 0 1 92510
box 0 0 3190 3190
use unit_cap  unit_cap_82
timestamp 1662145021
transform 1 0 3190 0 1 95700
box 0 0 3190 3190
use unit_cap  unit_cap_90
timestamp 1662145021
transform 1 0 3190 0 1 121220
box 0 0 3190 3190
use unit_cap  unit_cap_91
timestamp 1662145021
transform 1 0 3190 0 1 124410
box 0 0 3190 3190
use unit_cap  unit_cap_92
timestamp 1662145021
transform 1 0 3190 0 1 127600
box 0 0 3190 3190
use unit_cap  unit_cap_93
timestamp 1662145021
transform 1 0 3190 0 1 130790
box 0 0 3190 3190
use unit_cap  unit_cap_94
timestamp 1662145021
transform 1 0 3190 0 1 133980
box 0 0 3190 3190
use unit_cap  unit_cap_95
timestamp 1662145021
transform 1 0 3190 0 1 137170
box 0 0 3190 3190
use unit_cap  unit_cap_96
timestamp 1662145021
transform 1 0 3190 0 1 140360
box 0 0 3190 3190
use unit_cap  unit_cap_104
timestamp 1662145021
transform 1 0 6380 0 1 0
box 0 0 3190 3190
use unit_cap  unit_cap_105
timestamp 1662145021
transform 1 0 6380 0 1 3190
box 0 0 3190 3190
use unit_cap  unit_cap_106
timestamp 1662145021
transform 1 0 6380 0 1 6380
box 0 0 3190 3190
use unit_cap  unit_cap_107
timestamp 1662145021
transform 1 0 6380 0 1 9570
box 0 0 3190 3190
use unit_cap  unit_cap_108
timestamp 1662145021
transform 1 0 6380 0 1 12760
box 0 0 3190 3190
use unit_cap  unit_cap_109
timestamp 1662145021
transform 1 0 6380 0 1 15950
box 0 0 3190 3190
use unit_cap  unit_cap_110
timestamp 1662145021
transform 1 0 6380 0 1 19140
box 0 0 3190 3190
use unit_cap  unit_cap_111
timestamp 1662145021
transform 1 0 6380 0 1 22330
box 0 0 3190 3190
use unit_cap  unit_cap_112
timestamp 1662145021
transform 1 0 6380 0 1 25520
box 0 0 3190 3190
use unit_cap  unit_cap_113
timestamp 1662145021
transform 1 0 6380 0 1 28710
box 0 0 3190 3190
use unit_cap  unit_cap_114
timestamp 1662145021
transform 1 0 6380 0 1 31900
box 0 0 3190 3190
use unit_cap  unit_cap_115
timestamp 1662145021
transform 1 0 6380 0 1 35090
box 0 0 3190 3190
use unit_cap  unit_cap_116
timestamp 1662145021
transform 1 0 6380 0 1 38280
box 0 0 3190 3190
use unit_cap  unit_cap_117
timestamp 1662145021
transform 1 0 6380 0 1 41470
box 0 0 3190 3190
use unit_cap  unit_cap_118
timestamp 1662145021
transform 1 0 6380 0 1 44660
box 0 0 3190 3190
use unit_cap  unit_cap_119
timestamp 1662145021
transform 1 0 6380 0 1 47850
box 0 0 3190 3190
use unit_cap  unit_cap_120
timestamp 1662145021
transform 1 0 6380 0 1 51040
box 0 0 3190 3190
use unit_cap  unit_cap_121
timestamp 1662145021
transform 1 0 6380 0 1 54230
box 0 0 3190 3190
use unit_cap  unit_cap_122
timestamp 1662145021
transform 1 0 6380 0 1 57420
box 0 0 3190 3190
use unit_cap  unit_cap_123
timestamp 1662145021
transform 1 0 6380 0 1 60610
box 0 0 3190 3190
use unit_cap  unit_cap_124
timestamp 1662145021
transform 1 0 6380 0 1 63800
box 0 0 3190 3190
use unit_cap  unit_cap_125
timestamp 1662145021
transform 1 0 6380 0 1 66990
box 0 0 3190 3190
use unit_cap  unit_cap_126
timestamp 1662145021
transform 1 0 6380 0 1 70180
box 0 0 3190 3190
use unit_cap  unit_cap_127
timestamp 1662145021
transform 1 0 6380 0 1 73370
box 0 0 3190 3190
use unit_cap  unit_cap_128
timestamp 1662145021
transform 1 0 6380 0 1 76560
box 0 0 3190 3190
use unit_cap  unit_cap_129
timestamp 1662145021
transform 1 0 6380 0 1 79750
box 0 0 3190 3190
use unit_cap  unit_cap_130
timestamp 1662145021
transform 1 0 6380 0 1 82940
box 0 0 3190 3190
use unit_cap  unit_cap_131
timestamp 1662145021
transform 1 0 6380 0 1 86130
box 0 0 3190 3190
use unit_cap  unit_cap_132
timestamp 1662145021
transform 1 0 6380 0 1 89320
box 0 0 3190 3190
use unit_cap  unit_cap_133
timestamp 1662145021
transform 1 0 6380 0 1 92510
box 0 0 3190 3190
use unit_cap  unit_cap_134
timestamp 1662145021
transform 1 0 6380 0 1 95700
box 0 0 3190 3190
use unit_cap  unit_cap_142
timestamp 1662145021
transform 1 0 6380 0 1 121220
box 0 0 3190 3190
use unit_cap  unit_cap_143
timestamp 1662145021
transform 1 0 6380 0 1 124410
box 0 0 3190 3190
use unit_cap  unit_cap_144
timestamp 1662145021
transform 1 0 6380 0 1 127600
box 0 0 3190 3190
use unit_cap  unit_cap_145
timestamp 1662145021
transform 1 0 6380 0 1 130790
box 0 0 3190 3190
use unit_cap  unit_cap_146
timestamp 1662145021
transform 1 0 6380 0 1 133980
box 0 0 3190 3190
use unit_cap  unit_cap_147
timestamp 1662145021
transform 1 0 6380 0 1 137170
box 0 0 3190 3190
use unit_cap  unit_cap_148
timestamp 1662145021
transform 1 0 6380 0 1 140360
box 0 0 3190 3190
use unit_cap  unit_cap_156
timestamp 1662145021
transform 1 0 9570 0 1 0
box 0 0 3190 3190
use unit_cap  unit_cap_157
timestamp 1662145021
transform 1 0 9570 0 1 3190
box 0 0 3190 3190
use unit_cap  unit_cap_158
timestamp 1662145021
transform 1 0 9570 0 1 6380
box 0 0 3190 3190
use unit_cap  unit_cap_159
timestamp 1662145021
transform 1 0 9570 0 1 9570
box 0 0 3190 3190
use unit_cap  unit_cap_160
timestamp 1662145021
transform 1 0 9570 0 1 12760
box 0 0 3190 3190
use unit_cap  unit_cap_161
timestamp 1662145021
transform 1 0 9570 0 1 15950
box 0 0 3190 3190
use unit_cap  unit_cap_162
timestamp 1662145021
transform 1 0 9570 0 1 19140
box 0 0 3190 3190
use unit_cap  unit_cap_163
timestamp 1662145021
transform 1 0 9570 0 1 22330
box 0 0 3190 3190
use unit_cap  unit_cap_164
timestamp 1662145021
transform 1 0 9570 0 1 25520
box 0 0 3190 3190
use unit_cap  unit_cap_165
timestamp 1662145021
transform 1 0 9570 0 1 28710
box 0 0 3190 3190
use unit_cap  unit_cap_166
timestamp 1662145021
transform 1 0 9570 0 1 31900
box 0 0 3190 3190
use unit_cap  unit_cap_167
timestamp 1662145021
transform 1 0 9570 0 1 35090
box 0 0 3190 3190
use unit_cap  unit_cap_168
timestamp 1662145021
transform 1 0 9570 0 1 38280
box 0 0 3190 3190
use unit_cap  unit_cap_169
timestamp 1662145021
transform 1 0 9570 0 1 41470
box 0 0 3190 3190
use unit_cap  unit_cap_170
timestamp 1662145021
transform 1 0 9570 0 1 44660
box 0 0 3190 3190
use unit_cap  unit_cap_171
timestamp 1662145021
transform 1 0 9570 0 1 47850
box 0 0 3190 3190
use unit_cap  unit_cap_172
timestamp 1662145021
transform 1 0 9570 0 1 51040
box 0 0 3190 3190
use unit_cap  unit_cap_173
timestamp 1662145021
transform 1 0 9570 0 1 54230
box 0 0 3190 3190
use unit_cap  unit_cap_174
timestamp 1662145021
transform 1 0 9570 0 1 57420
box 0 0 3190 3190
use unit_cap  unit_cap_175
timestamp 1662145021
transform 1 0 9570 0 1 60610
box 0 0 3190 3190
use unit_cap  unit_cap_176
timestamp 1662145021
transform 1 0 9570 0 1 63800
box 0 0 3190 3190
use unit_cap  unit_cap_177
timestamp 1662145021
transform 1 0 9570 0 1 66990
box 0 0 3190 3190
use unit_cap  unit_cap_178
timestamp 1662145021
transform 1 0 9570 0 1 70180
box 0 0 3190 3190
use unit_cap  unit_cap_179
timestamp 1662145021
transform 1 0 9570 0 1 73370
box 0 0 3190 3190
use unit_cap  unit_cap_180
timestamp 1662145021
transform 1 0 9570 0 1 76560
box 0 0 3190 3190
use unit_cap  unit_cap_181
timestamp 1662145021
transform 1 0 9570 0 1 79750
box 0 0 3190 3190
use unit_cap  unit_cap_182
timestamp 1662145021
transform 1 0 9570 0 1 82940
box 0 0 3190 3190
use unit_cap  unit_cap_183
timestamp 1662145021
transform 1 0 9570 0 1 86130
box 0 0 3190 3190
use unit_cap  unit_cap_184
timestamp 1662145021
transform 1 0 9570 0 1 89320
box 0 0 3190 3190
use unit_cap  unit_cap_185
timestamp 1662145021
transform 1 0 9570 0 1 92510
box 0 0 3190 3190
use unit_cap  unit_cap_186
timestamp 1662145021
transform 1 0 9570 0 1 95700
box 0 0 3190 3190
use unit_cap  unit_cap_187
timestamp 1662145021
transform 1 0 9570 0 1 98890
box 0 0 3190 3190
use unit_cap  unit_cap_188
timestamp 1662145021
transform 1 0 9570 0 1 102080
box 0 0 3190 3190
use unit_cap  unit_cap_189
timestamp 1662145021
transform 1 0 9570 0 1 105270
box 0 0 3190 3190
use unit_cap  unit_cap_190
timestamp 1662145021
transform 1 0 9570 0 1 108460
box 0 0 3190 3190
use unit_cap  unit_cap_191
timestamp 1662145021
transform 1 0 9570 0 1 111650
box 0 0 3190 3190
use unit_cap  unit_cap_192
timestamp 1662145021
transform 1 0 9570 0 1 114840
box 0 0 3190 3190
use unit_cap  unit_cap_193
timestamp 1662145021
transform 1 0 9570 0 1 118030
box 0 0 3190 3190
use unit_cap  unit_cap_194
timestamp 1662145021
transform 1 0 9570 0 1 121220
box 0 0 3190 3190
use unit_cap  unit_cap_195
timestamp 1662145021
transform 1 0 9570 0 1 124410
box 0 0 3190 3190
use unit_cap  unit_cap_196
timestamp 1662145021
transform 1 0 9570 0 1 127600
box 0 0 3190 3190
use unit_cap  unit_cap_197
timestamp 1662145021
transform 1 0 9570 0 1 130790
box 0 0 3190 3190
use unit_cap  unit_cap_198
timestamp 1662145021
transform 1 0 9570 0 1 133980
box 0 0 3190 3190
use unit_cap  unit_cap_199
timestamp 1662145021
transform 1 0 9570 0 1 137170
box 0 0 3190 3190
use unit_cap  unit_cap_200
timestamp 1662145021
transform 1 0 9570 0 1 140360
box 0 0 3190 3190
use unit_cap  unit_cap_201
timestamp 1662145021
transform 1 0 9570 0 1 143550
box 0 0 3190 3190
use unit_cap  unit_cap_202
timestamp 1662145021
transform 1 0 9570 0 1 146740
box 0 0 3190 3190
use unit_cap  unit_cap_203
timestamp 1662145021
transform 1 0 9570 0 1 149930
box 0 0 3190 3190
use unit_cap  unit_cap_204
timestamp 1662145021
transform 1 0 9570 0 1 153120
box 0 0 3190 3190
use unit_cap  unit_cap_205
timestamp 1662145021
transform 1 0 9570 0 1 156310
box 0 0 3190 3190
use unit_cap  unit_cap_206
timestamp 1662145021
transform 1 0 9570 0 1 159500
box 0 0 3190 3190
use unit_cap  unit_cap_207
timestamp 1662145021
transform 1 0 9570 0 1 162690
box 0 0 3190 3190
use unit_cap  unit_cap_208
timestamp 1662145021
transform 1 0 12760 0 1 0
box 0 0 3190 3190
use unit_cap  unit_cap_209
timestamp 1662145021
transform 1 0 12760 0 1 3190
box 0 0 3190 3190
use unit_cap  unit_cap_210
timestamp 1662145021
transform 1 0 12760 0 1 6380
box 0 0 3190 3190
use unit_cap  unit_cap_211
timestamp 1662145021
transform 1 0 12760 0 1 9570
box 0 0 3190 3190
use unit_cap  unit_cap_212
timestamp 1662145021
transform 1 0 12760 0 1 12760
box 0 0 3190 3190
use unit_cap  unit_cap_213
timestamp 1662145021
transform 1 0 12760 0 1 15950
box 0 0 3190 3190
use unit_cap  unit_cap_214
timestamp 1662145021
transform 1 0 12760 0 1 19140
box 0 0 3190 3190
use unit_cap  unit_cap_215
timestamp 1662145021
transform 1 0 12760 0 1 22330
box 0 0 3190 3190
use unit_cap  unit_cap_216
timestamp 1662145021
transform 1 0 12760 0 1 25520
box 0 0 3190 3190
use unit_cap  unit_cap_217
timestamp 1662145021
transform 1 0 12760 0 1 28710
box 0 0 3190 3190
use unit_cap  unit_cap_218
timestamp 1662145021
transform 1 0 12760 0 1 31900
box 0 0 3190 3190
use unit_cap  unit_cap_219
timestamp 1662145021
transform 1 0 12760 0 1 35090
box 0 0 3190 3190
use unit_cap  unit_cap_220
timestamp 1662145021
transform 1 0 12760 0 1 38280
box 0 0 3190 3190
use unit_cap  unit_cap_221
timestamp 1662145021
transform 1 0 12760 0 1 41470
box 0 0 3190 3190
use unit_cap  unit_cap_222
timestamp 1662145021
transform 1 0 12760 0 1 44660
box 0 0 3190 3190
use unit_cap  unit_cap_223
timestamp 1662145021
transform 1 0 12760 0 1 47850
box 0 0 3190 3190
use unit_cap  unit_cap_224
timestamp 1662145021
transform 1 0 12760 0 1 51040
box 0 0 3190 3190
use unit_cap  unit_cap_225
timestamp 1662145021
transform 1 0 12760 0 1 54230
box 0 0 3190 3190
use unit_cap  unit_cap_226
timestamp 1662145021
transform 1 0 12760 0 1 57420
box 0 0 3190 3190
use unit_cap  unit_cap_227
timestamp 1662145021
transform 1 0 12760 0 1 60610
box 0 0 3190 3190
use unit_cap  unit_cap_228
timestamp 1662145021
transform 1 0 12760 0 1 63800
box 0 0 3190 3190
use unit_cap  unit_cap_229
timestamp 1662145021
transform 1 0 12760 0 1 66990
box 0 0 3190 3190
use unit_cap  unit_cap_230
timestamp 1662145021
transform 1 0 12760 0 1 70180
box 0 0 3190 3190
use unit_cap  unit_cap_231
timestamp 1662145021
transform 1 0 12760 0 1 73370
box 0 0 3190 3190
use unit_cap  unit_cap_232
timestamp 1662145021
transform 1 0 12760 0 1 76560
box 0 0 3190 3190
use unit_cap  unit_cap_233
timestamp 1662145021
transform 1 0 12760 0 1 79750
box 0 0 3190 3190
use unit_cap  unit_cap_234
timestamp 1662145021
transform 1 0 12760 0 1 82940
box 0 0 3190 3190
use unit_cap  unit_cap_235
timestamp 1662145021
transform 1 0 12760 0 1 86130
box 0 0 3190 3190
use unit_cap  unit_cap_236
timestamp 1662145021
transform 1 0 12760 0 1 89320
box 0 0 3190 3190
use unit_cap  unit_cap_237
timestamp 1662145021
transform 1 0 12760 0 1 92510
box 0 0 3190 3190
use unit_cap  unit_cap_238
timestamp 1662145021
transform 1 0 12760 0 1 95700
box 0 0 3190 3190
use unit_cap  unit_cap_239
timestamp 1662145021
transform 1 0 12760 0 1 98890
box 0 0 3190 3190
use unit_cap  unit_cap_240
timestamp 1662145021
transform 1 0 12760 0 1 102080
box 0 0 3190 3190
use unit_cap  unit_cap_241
timestamp 1662145021
transform 1 0 12760 0 1 105270
box 0 0 3190 3190
use unit_cap  unit_cap_242
timestamp 1662145021
transform 1 0 12760 0 1 108460
box 0 0 3190 3190
use unit_cap  unit_cap_243
timestamp 1662145021
transform 1 0 12760 0 1 111650
box 0 0 3190 3190
use unit_cap  unit_cap_244
timestamp 1662145021
transform 1 0 12760 0 1 114840
box 0 0 3190 3190
use unit_cap  unit_cap_245
timestamp 1662145021
transform 1 0 12760 0 1 118030
box 0 0 3190 3190
use unit_cap  unit_cap_246
timestamp 1662145021
transform 1 0 12760 0 1 121220
box 0 0 3190 3190
use unit_cap  unit_cap_247
timestamp 1662145021
transform 1 0 12760 0 1 124410
box 0 0 3190 3190
use unit_cap  unit_cap_248
timestamp 1662145021
transform 1 0 12760 0 1 127600
box 0 0 3190 3190
use unit_cap  unit_cap_249
timestamp 1662145021
transform 1 0 12760 0 1 130790
box 0 0 3190 3190
use unit_cap  unit_cap_250
timestamp 1662145021
transform 1 0 12760 0 1 133980
box 0 0 3190 3190
use unit_cap  unit_cap_251
timestamp 1662145021
transform 1 0 12760 0 1 137170
box 0 0 3190 3190
use unit_cap  unit_cap_252
timestamp 1662145021
transform 1 0 12760 0 1 140360
box 0 0 3190 3190
use unit_cap  unit_cap_253
timestamp 1662145021
transform 1 0 12760 0 1 143550
box 0 0 3190 3190
use unit_cap  unit_cap_254
timestamp 1662145021
transform 1 0 12760 0 1 146740
box 0 0 3190 3190
use unit_cap  unit_cap_255
timestamp 1662145021
transform 1 0 12760 0 1 149930
box 0 0 3190 3190
use unit_cap  unit_cap_256
timestamp 1662145021
transform 1 0 12760 0 1 153120
box 0 0 3190 3190
use unit_cap  unit_cap_257
timestamp 1662145021
transform 1 0 12760 0 1 156310
box 0 0 3190 3190
use unit_cap  unit_cap_258
timestamp 1662145021
transform 1 0 12760 0 1 159500
box 0 0 3190 3190
use unit_cap  unit_cap_259
timestamp 1662145021
transform 1 0 12760 0 1 162690
box 0 0 3190 3190
use unit_cap  unit_cap_260
timestamp 1662145021
transform 1 0 15950 0 1 0
box 0 0 3190 3190
use unit_cap  unit_cap_261
timestamp 1662145021
transform 1 0 15950 0 1 3190
box 0 0 3190 3190
use unit_cap  unit_cap_262
timestamp 1662145021
transform 1 0 15950 0 1 6380
box 0 0 3190 3190
use unit_cap  unit_cap_263
timestamp 1662145021
transform 1 0 15950 0 1 9570
box 0 0 3190 3190
use unit_cap  unit_cap_264
timestamp 1662145021
transform 1 0 15950 0 1 12760
box 0 0 3190 3190
use unit_cap  unit_cap_265
timestamp 1662145021
transform 1 0 15950 0 1 15950
box 0 0 3190 3190
use unit_cap  unit_cap_266
timestamp 1662145021
transform 1 0 15950 0 1 19140
box 0 0 3190 3190
use unit_cap  unit_cap_267
timestamp 1662145021
transform 1 0 15950 0 1 22330
box 0 0 3190 3190
use unit_cap  unit_cap_268
timestamp 1662145021
transform 1 0 15950 0 1 25520
box 0 0 3190 3190
use unit_cap  unit_cap_269
timestamp 1662145021
transform 1 0 15950 0 1 28710
box 0 0 3190 3190
use unit_cap  unit_cap_270
timestamp 1662145021
transform 1 0 15950 0 1 31900
box 0 0 3190 3190
use unit_cap  unit_cap_271
timestamp 1662145021
transform 1 0 15950 0 1 35090
box 0 0 3190 3190
use unit_cap  unit_cap_272
timestamp 1662145021
transform 1 0 15950 0 1 38280
box 0 0 3190 3190
use unit_cap  unit_cap_273
timestamp 1662145021
transform 1 0 15950 0 1 41470
box 0 0 3190 3190
use unit_cap  unit_cap_274
timestamp 1662145021
transform 1 0 15950 0 1 44660
box 0 0 3190 3190
use unit_cap  unit_cap_275
timestamp 1662145021
transform 1 0 15950 0 1 47850
box 0 0 3190 3190
use unit_cap  unit_cap_276
timestamp 1662145021
transform 1 0 15950 0 1 51040
box 0 0 3190 3190
use unit_cap  unit_cap_277
timestamp 1662145021
transform 1 0 15950 0 1 54230
box 0 0 3190 3190
use unit_cap  unit_cap_278
timestamp 1662145021
transform 1 0 15950 0 1 57420
box 0 0 3190 3190
use unit_cap  unit_cap_279
timestamp 1662145021
transform 1 0 15950 0 1 60610
box 0 0 3190 3190
use unit_cap  unit_cap_280
timestamp 1662145021
transform 1 0 15950 0 1 63800
box 0 0 3190 3190
use unit_cap  unit_cap_281
timestamp 1662145021
transform 1 0 15950 0 1 66990
box 0 0 3190 3190
use unit_cap  unit_cap_282
timestamp 1662145021
transform 1 0 15950 0 1 70180
box 0 0 3190 3190
use unit_cap  unit_cap_283
timestamp 1662145021
transform 1 0 15950 0 1 73370
box 0 0 3190 3190
use unit_cap  unit_cap_284
timestamp 1662145021
transform 1 0 15950 0 1 76560
box 0 0 3190 3190
use unit_cap  unit_cap_285
timestamp 1662145021
transform 1 0 15950 0 1 79750
box 0 0 3190 3190
use unit_cap  unit_cap_286
timestamp 1662145021
transform 1 0 15950 0 1 82940
box 0 0 3190 3190
use unit_cap  unit_cap_287
timestamp 1662145021
transform 1 0 15950 0 1 86130
box 0 0 3190 3190
use unit_cap  unit_cap_288
timestamp 1662145021
transform 1 0 15950 0 1 89320
box 0 0 3190 3190
use unit_cap  unit_cap_289
timestamp 1662145021
transform 1 0 15950 0 1 92510
box 0 0 3190 3190
use unit_cap  unit_cap_290
timestamp 1662145021
transform 1 0 15950 0 1 95700
box 0 0 3190 3190
use unit_cap  unit_cap_291
timestamp 1662145021
transform 1 0 15950 0 1 98890
box 0 0 3190 3190
use unit_cap  unit_cap_292
timestamp 1662145021
transform 1 0 15950 0 1 102080
box 0 0 3190 3190
use unit_cap  unit_cap_293
timestamp 1662145021
transform 1 0 15950 0 1 105270
box 0 0 3190 3190
use unit_cap  unit_cap_294
timestamp 1662145021
transform 1 0 15950 0 1 108460
box 0 0 3190 3190
use unit_cap  unit_cap_295
timestamp 1662145021
transform 1 0 15950 0 1 111650
box 0 0 3190 3190
use unit_cap  unit_cap_296
timestamp 1662145021
transform 1 0 15950 0 1 114840
box 0 0 3190 3190
use unit_cap  unit_cap_297
timestamp 1662145021
transform 1 0 15950 0 1 118030
box 0 0 3190 3190
use unit_cap  unit_cap_298
timestamp 1662145021
transform 1 0 15950 0 1 121220
box 0 0 3190 3190
use unit_cap  unit_cap_299
timestamp 1662145021
transform 1 0 15950 0 1 124410
box 0 0 3190 3190
use unit_cap  unit_cap_300
timestamp 1662145021
transform 1 0 15950 0 1 127600
box 0 0 3190 3190
use unit_cap  unit_cap_301
timestamp 1662145021
transform 1 0 15950 0 1 130790
box 0 0 3190 3190
use unit_cap  unit_cap_302
timestamp 1662145021
transform 1 0 15950 0 1 133980
box 0 0 3190 3190
use unit_cap  unit_cap_303
timestamp 1662145021
transform 1 0 15950 0 1 137170
box 0 0 3190 3190
use unit_cap  unit_cap_304
timestamp 1662145021
transform 1 0 15950 0 1 140360
box 0 0 3190 3190
use unit_cap  unit_cap_305
timestamp 1662145021
transform 1 0 15950 0 1 143550
box 0 0 3190 3190
use unit_cap  unit_cap_306
timestamp 1662145021
transform 1 0 15950 0 1 146740
box 0 0 3190 3190
use unit_cap  unit_cap_307
timestamp 1662145021
transform 1 0 15950 0 1 149930
box 0 0 3190 3190
use unit_cap  unit_cap_308
timestamp 1662145021
transform 1 0 15950 0 1 153120
box 0 0 3190 3190
use unit_cap  unit_cap_309
timestamp 1662145021
transform 1 0 15950 0 1 156310
box 0 0 3190 3190
use unit_cap  unit_cap_310
timestamp 1662145021
transform 1 0 15950 0 1 159500
box 0 0 3190 3190
use unit_cap  unit_cap_311
timestamp 1662145021
transform 1 0 15950 0 1 162690
box 0 0 3190 3190
use unit_cap  unit_cap_312
timestamp 1662145021
transform 1 0 19140 0 1 0
box 0 0 3190 3190
use unit_cap  unit_cap_313
timestamp 1662145021
transform 1 0 19140 0 1 3190
box 0 0 3190 3190
use unit_cap  unit_cap_314
timestamp 1662145021
transform 1 0 19140 0 1 6380
box 0 0 3190 3190
use unit_cap  unit_cap_315
timestamp 1662145021
transform 1 0 19140 0 1 9570
box 0 0 3190 3190
use unit_cap  unit_cap_316
timestamp 1662145021
transform 1 0 19140 0 1 12760
box 0 0 3190 3190
use unit_cap  unit_cap_317
timestamp 1662145021
transform 1 0 19140 0 1 15950
box 0 0 3190 3190
use unit_cap  unit_cap_318
timestamp 1662145021
transform 1 0 19140 0 1 19140
box 0 0 3190 3190
use unit_cap  unit_cap_319
timestamp 1662145021
transform 1 0 19140 0 1 22330
box 0 0 3190 3190
use unit_cap  unit_cap_320
timestamp 1662145021
transform 1 0 19140 0 1 25520
box 0 0 3190 3190
use unit_cap  unit_cap_321
timestamp 1662145021
transform 1 0 19140 0 1 28710
box 0 0 3190 3190
use unit_cap  unit_cap_322
timestamp 1662145021
transform 1 0 19140 0 1 31900
box 0 0 3190 3190
use unit_cap  unit_cap_323
timestamp 1662145021
transform 1 0 19140 0 1 35090
box 0 0 3190 3190
use unit_cap  unit_cap_324
timestamp 1662145021
transform 1 0 19140 0 1 38280
box 0 0 3190 3190
use unit_cap  unit_cap_325
timestamp 1662145021
transform 1 0 19140 0 1 41470
box 0 0 3190 3190
use unit_cap  unit_cap_326
timestamp 1662145021
transform 1 0 19140 0 1 44660
box 0 0 3190 3190
use unit_cap  unit_cap_327
timestamp 1662145021
transform 1 0 19140 0 1 47850
box 0 0 3190 3190
use unit_cap  unit_cap_328
timestamp 1662145021
transform 1 0 19140 0 1 51040
box 0 0 3190 3190
use unit_cap  unit_cap_329
timestamp 1662145021
transform 1 0 19140 0 1 54230
box 0 0 3190 3190
use unit_cap  unit_cap_330
timestamp 1662145021
transform 1 0 19140 0 1 57420
box 0 0 3190 3190
use unit_cap  unit_cap_331
timestamp 1662145021
transform 1 0 19140 0 1 60610
box 0 0 3190 3190
use unit_cap  unit_cap_332
timestamp 1662145021
transform 1 0 19140 0 1 63800
box 0 0 3190 3190
use unit_cap  unit_cap_333
timestamp 1662145021
transform 1 0 19140 0 1 66990
box 0 0 3190 3190
use unit_cap  unit_cap_334
timestamp 1662145021
transform 1 0 19140 0 1 70180
box 0 0 3190 3190
use unit_cap  unit_cap_335
timestamp 1662145021
transform 1 0 19140 0 1 73370
box 0 0 3190 3190
use unit_cap  unit_cap_336
timestamp 1662145021
transform 1 0 19140 0 1 76560
box 0 0 3190 3190
use unit_cap  unit_cap_337
timestamp 1662145021
transform 1 0 19140 0 1 79750
box 0 0 3190 3190
use unit_cap  unit_cap_338
timestamp 1662145021
transform 1 0 19140 0 1 82940
box 0 0 3190 3190
use unit_cap  unit_cap_339
timestamp 1662145021
transform 1 0 19140 0 1 86130
box 0 0 3190 3190
use unit_cap  unit_cap_340
timestamp 1662145021
transform 1 0 19140 0 1 89320
box 0 0 3190 3190
use unit_cap  unit_cap_341
timestamp 1662145021
transform 1 0 19140 0 1 92510
box 0 0 3190 3190
use unit_cap  unit_cap_342
timestamp 1662145021
transform 1 0 19140 0 1 95700
box 0 0 3190 3190
use unit_cap  unit_cap_343
timestamp 1662145021
transform 1 0 19140 0 1 98890
box 0 0 3190 3190
use unit_cap  unit_cap_344
timestamp 1662145021
transform 1 0 19140 0 1 102080
box 0 0 3190 3190
use unit_cap  unit_cap_345
timestamp 1662145021
transform 1 0 19140 0 1 105270
box 0 0 3190 3190
use unit_cap  unit_cap_346
timestamp 1662145021
transform 1 0 19140 0 1 108460
box 0 0 3190 3190
use unit_cap  unit_cap_347
timestamp 1662145021
transform 1 0 19140 0 1 111650
box 0 0 3190 3190
use unit_cap  unit_cap_348
timestamp 1662145021
transform 1 0 19140 0 1 114840
box 0 0 3190 3190
use unit_cap  unit_cap_349
timestamp 1662145021
transform 1 0 19140 0 1 118030
box 0 0 3190 3190
use unit_cap  unit_cap_350
timestamp 1662145021
transform 1 0 19140 0 1 121220
box 0 0 3190 3190
use unit_cap  unit_cap_351
timestamp 1662145021
transform 1 0 19140 0 1 124410
box 0 0 3190 3190
use unit_cap  unit_cap_352
timestamp 1662145021
transform 1 0 19140 0 1 127600
box 0 0 3190 3190
use unit_cap  unit_cap_353
timestamp 1662145021
transform 1 0 19140 0 1 130790
box 0 0 3190 3190
use unit_cap  unit_cap_354
timestamp 1662145021
transform 1 0 19140 0 1 133980
box 0 0 3190 3190
use unit_cap  unit_cap_355
timestamp 1662145021
transform 1 0 19140 0 1 137170
box 0 0 3190 3190
use unit_cap  unit_cap_356
timestamp 1662145021
transform 1 0 19140 0 1 140360
box 0 0 3190 3190
use unit_cap  unit_cap_357
timestamp 1662145021
transform 1 0 19140 0 1 143550
box 0 0 3190 3190
use unit_cap  unit_cap_358
timestamp 1662145021
transform 1 0 19140 0 1 146740
box 0 0 3190 3190
use unit_cap  unit_cap_359
timestamp 1662145021
transform 1 0 19140 0 1 149930
box 0 0 3190 3190
use unit_cap  unit_cap_360
timestamp 1662145021
transform 1 0 19140 0 1 153120
box 0 0 3190 3190
use unit_cap  unit_cap_361
timestamp 1662145021
transform 1 0 19140 0 1 156310
box 0 0 3190 3190
use unit_cap  unit_cap_362
timestamp 1662145021
transform 1 0 19140 0 1 159500
box 0 0 3190 3190
use unit_cap  unit_cap_363
timestamp 1662145021
transform 1 0 19140 0 1 162690
box 0 0 3190 3190
use unit_cap  unit_cap_364
timestamp 1662145021
transform 1 0 22330 0 1 0
box 0 0 3190 3190
use unit_cap  unit_cap_365
timestamp 1662145021
transform 1 0 22330 0 1 3190
box 0 0 3190 3190
use unit_cap  unit_cap_366
timestamp 1662145021
transform 1 0 22330 0 1 6380
box 0 0 3190 3190
use unit_cap  unit_cap_367
timestamp 1662145021
transform 1 0 22330 0 1 9570
box 0 0 3190 3190
use unit_cap  unit_cap_368
timestamp 1662145021
transform 1 0 22330 0 1 12760
box 0 0 3190 3190
use unit_cap  unit_cap_369
timestamp 1662145021
transform 1 0 22330 0 1 15950
box 0 0 3190 3190
use unit_cap  unit_cap_370
timestamp 1662145021
transform 1 0 22330 0 1 19140
box 0 0 3190 3190
use unit_cap  unit_cap_371
timestamp 1662145021
transform 1 0 22330 0 1 22330
box 0 0 3190 3190
use unit_cap  unit_cap_372
timestamp 1662145021
transform 1 0 22330 0 1 25520
box 0 0 3190 3190
use unit_cap  unit_cap_373
timestamp 1662145021
transform 1 0 22330 0 1 28710
box 0 0 3190 3190
use unit_cap  unit_cap_374
timestamp 1662145021
transform 1 0 22330 0 1 31900
box 0 0 3190 3190
use unit_cap  unit_cap_375
timestamp 1662145021
transform 1 0 22330 0 1 35090
box 0 0 3190 3190
use unit_cap  unit_cap_376
timestamp 1662145021
transform 1 0 22330 0 1 38280
box 0 0 3190 3190
use unit_cap  unit_cap_377
timestamp 1662145021
transform 1 0 22330 0 1 41470
box 0 0 3190 3190
use unit_cap  unit_cap_378
timestamp 1662145021
transform 1 0 22330 0 1 44660
box 0 0 3190 3190
use unit_cap  unit_cap_379
timestamp 1662145021
transform 1 0 22330 0 1 47850
box 0 0 3190 3190
use unit_cap  unit_cap_380
timestamp 1662145021
transform 1 0 22330 0 1 51040
box 0 0 3190 3190
use unit_cap  unit_cap_381
timestamp 1662145021
transform 1 0 22330 0 1 54230
box 0 0 3190 3190
use unit_cap  unit_cap_382
timestamp 1662145021
transform 1 0 22330 0 1 57420
box 0 0 3190 3190
use unit_cap  unit_cap_383
timestamp 1662145021
transform 1 0 22330 0 1 60610
box 0 0 3190 3190
use unit_cap  unit_cap_384
timestamp 1662145021
transform 1 0 22330 0 1 63800
box 0 0 3190 3190
use unit_cap  unit_cap_385
timestamp 1662145021
transform 1 0 22330 0 1 66990
box 0 0 3190 3190
use unit_cap  unit_cap_386
timestamp 1662145021
transform 1 0 22330 0 1 70180
box 0 0 3190 3190
use unit_cap  unit_cap_387
timestamp 1662145021
transform 1 0 22330 0 1 73370
box 0 0 3190 3190
use unit_cap  unit_cap_388
timestamp 1662145021
transform 1 0 22330 0 1 76560
box 0 0 3190 3190
use unit_cap  unit_cap_389
timestamp 1662145021
transform 1 0 22330 0 1 79750
box 0 0 3190 3190
use unit_cap  unit_cap_390
timestamp 1662145021
transform 1 0 22330 0 1 82940
box 0 0 3190 3190
use unit_cap  unit_cap_391
timestamp 1662145021
transform 1 0 22330 0 1 86130
box 0 0 3190 3190
use unit_cap  unit_cap_392
timestamp 1662145021
transform 1 0 22330 0 1 89320
box 0 0 3190 3190
use unit_cap  unit_cap_393
timestamp 1662145021
transform 1 0 22330 0 1 92510
box 0 0 3190 3190
use unit_cap  unit_cap_394
timestamp 1662145021
transform 1 0 22330 0 1 95700
box 0 0 3190 3190
use unit_cap  unit_cap_395
timestamp 1662145021
transform 1 0 22330 0 1 98890
box 0 0 3190 3190
use unit_cap  unit_cap_396
timestamp 1662145021
transform 1 0 22330 0 1 102080
box 0 0 3190 3190
use unit_cap  unit_cap_397
timestamp 1662145021
transform 1 0 22330 0 1 105270
box 0 0 3190 3190
use unit_cap  unit_cap_398
timestamp 1662145021
transform 1 0 22330 0 1 108460
box 0 0 3190 3190
use unit_cap  unit_cap_399
timestamp 1662145021
transform 1 0 22330 0 1 111650
box 0 0 3190 3190
use unit_cap  unit_cap_400
timestamp 1662145021
transform 1 0 22330 0 1 114840
box 0 0 3190 3190
use unit_cap  unit_cap_401
timestamp 1662145021
transform 1 0 22330 0 1 118030
box 0 0 3190 3190
use unit_cap  unit_cap_402
timestamp 1662145021
transform 1 0 22330 0 1 121220
box 0 0 3190 3190
use unit_cap  unit_cap_403
timestamp 1662145021
transform 1 0 22330 0 1 124410
box 0 0 3190 3190
use unit_cap  unit_cap_404
timestamp 1662145021
transform 1 0 22330 0 1 127600
box 0 0 3190 3190
use unit_cap  unit_cap_405
timestamp 1662145021
transform 1 0 22330 0 1 130790
box 0 0 3190 3190
use unit_cap  unit_cap_406
timestamp 1662145021
transform 1 0 22330 0 1 133980
box 0 0 3190 3190
use unit_cap  unit_cap_407
timestamp 1662145021
transform 1 0 22330 0 1 137170
box 0 0 3190 3190
use unit_cap  unit_cap_408
timestamp 1662145021
transform 1 0 22330 0 1 140360
box 0 0 3190 3190
use unit_cap  unit_cap_409
timestamp 1662145021
transform 1 0 22330 0 1 143550
box 0 0 3190 3190
use unit_cap  unit_cap_410
timestamp 1662145021
transform 1 0 22330 0 1 146740
box 0 0 3190 3190
use unit_cap  unit_cap_411
timestamp 1662145021
transform 1 0 22330 0 1 149930
box 0 0 3190 3190
use unit_cap  unit_cap_412
timestamp 1662145021
transform 1 0 22330 0 1 153120
box 0 0 3190 3190
use unit_cap  unit_cap_413
timestamp 1662145021
transform 1 0 22330 0 1 156310
box 0 0 3190 3190
use unit_cap  unit_cap_414
timestamp 1662145021
transform 1 0 22330 0 1 159500
box 0 0 3190 3190
use unit_cap  unit_cap_415
timestamp 1662145021
transform 1 0 22330 0 1 162690
box 0 0 3190 3190
use unit_cap  unit_cap_416
timestamp 1662145021
transform 1 0 25520 0 1 0
box 0 0 3190 3190
use unit_cap  unit_cap_417
timestamp 1662145021
transform 1 0 25520 0 1 3190
box 0 0 3190 3190
use unit_cap  unit_cap_418
timestamp 1662145021
transform 1 0 25520 0 1 6380
box 0 0 3190 3190
use unit_cap  unit_cap_419
timestamp 1662145021
transform 1 0 25520 0 1 9570
box 0 0 3190 3190
use unit_cap  unit_cap_420
timestamp 1662145021
transform 1 0 25520 0 1 12760
box 0 0 3190 3190
use unit_cap  unit_cap_421
timestamp 1662145021
transform 1 0 25520 0 1 15950
box 0 0 3190 3190
use unit_cap  unit_cap_422
timestamp 1662145021
transform 1 0 25520 0 1 19140
box 0 0 3190 3190
use unit_cap  unit_cap_423
timestamp 1662145021
transform 1 0 25520 0 1 22330
box 0 0 3190 3190
use unit_cap  unit_cap_424
timestamp 1662145021
transform 1 0 25520 0 1 25520
box 0 0 3190 3190
use unit_cap  unit_cap_425
timestamp 1662145021
transform 1 0 25520 0 1 28710
box 0 0 3190 3190
use unit_cap  unit_cap_426
timestamp 1662145021
transform 1 0 25520 0 1 31900
box 0 0 3190 3190
use unit_cap  unit_cap_427
timestamp 1662145021
transform 1 0 25520 0 1 35090
box 0 0 3190 3190
use unit_cap  unit_cap_428
timestamp 1662145021
transform 1 0 25520 0 1 38280
box 0 0 3190 3190
use unit_cap  unit_cap_429
timestamp 1662145021
transform 1 0 25520 0 1 41470
box 0 0 3190 3190
use unit_cap  unit_cap_430
timestamp 1662145021
transform 1 0 25520 0 1 44660
box 0 0 3190 3190
use unit_cap  unit_cap_431
timestamp 1662145021
transform 1 0 25520 0 1 47850
box 0 0 3190 3190
use unit_cap  unit_cap_432
timestamp 1662145021
transform 1 0 25520 0 1 51040
box 0 0 3190 3190
use unit_cap  unit_cap_433
timestamp 1662145021
transform 1 0 25520 0 1 54230
box 0 0 3190 3190
use unit_cap  unit_cap_434
timestamp 1662145021
transform 1 0 25520 0 1 57420
box 0 0 3190 3190
use unit_cap  unit_cap_435
timestamp 1662145021
transform 1 0 25520 0 1 60610
box 0 0 3190 3190
use unit_cap  unit_cap_436
timestamp 1662145021
transform 1 0 25520 0 1 63800
box 0 0 3190 3190
use unit_cap  unit_cap_437
timestamp 1662145021
transform 1 0 25520 0 1 66990
box 0 0 3190 3190
use unit_cap  unit_cap_438
timestamp 1662145021
transform 1 0 25520 0 1 70180
box 0 0 3190 3190
use unit_cap  unit_cap_439
timestamp 1662145021
transform 1 0 25520 0 1 73370
box 0 0 3190 3190
use unit_cap  unit_cap_440
timestamp 1662145021
transform 1 0 25520 0 1 76560
box 0 0 3190 3190
use unit_cap  unit_cap_441
timestamp 1662145021
transform 1 0 25520 0 1 79750
box 0 0 3190 3190
use unit_cap  unit_cap_442
timestamp 1662145021
transform 1 0 25520 0 1 82940
box 0 0 3190 3190
use unit_cap  unit_cap_443
timestamp 1662145021
transform 1 0 25520 0 1 86130
box 0 0 3190 3190
use unit_cap  unit_cap_444
timestamp 1662145021
transform 1 0 25520 0 1 89320
box 0 0 3190 3190
use unit_cap  unit_cap_445
timestamp 1662145021
transform 1 0 25520 0 1 92510
box 0 0 3190 3190
use unit_cap  unit_cap_446
timestamp 1662145021
transform 1 0 25520 0 1 95700
box 0 0 3190 3190
use unit_cap  unit_cap_447
timestamp 1662145021
transform 1 0 25520 0 1 98890
box 0 0 3190 3190
use unit_cap  unit_cap_448
timestamp 1662145021
transform 1 0 25520 0 1 102080
box 0 0 3190 3190
use unit_cap  unit_cap_449
timestamp 1662145021
transform 1 0 25520 0 1 105270
box 0 0 3190 3190
use unit_cap  unit_cap_450
timestamp 1662145021
transform 1 0 25520 0 1 108460
box 0 0 3190 3190
use unit_cap  unit_cap_451
timestamp 1662145021
transform 1 0 25520 0 1 111650
box 0 0 3190 3190
use unit_cap  unit_cap_452
timestamp 1662145021
transform 1 0 25520 0 1 114840
box 0 0 3190 3190
use unit_cap  unit_cap_453
timestamp 1662145021
transform 1 0 25520 0 1 118030
box 0 0 3190 3190
use unit_cap  unit_cap_454
timestamp 1662145021
transform 1 0 25520 0 1 121220
box 0 0 3190 3190
use unit_cap  unit_cap_455
timestamp 1662145021
transform 1 0 25520 0 1 124410
box 0 0 3190 3190
use unit_cap  unit_cap_456
timestamp 1662145021
transform 1 0 25520 0 1 127600
box 0 0 3190 3190
use unit_cap  unit_cap_457
timestamp 1662145021
transform 1 0 25520 0 1 130790
box 0 0 3190 3190
use unit_cap  unit_cap_458
timestamp 1662145021
transform 1 0 25520 0 1 133980
box 0 0 3190 3190
use unit_cap  unit_cap_459
timestamp 1662145021
transform 1 0 25520 0 1 137170
box 0 0 3190 3190
use unit_cap  unit_cap_460
timestamp 1662145021
transform 1 0 25520 0 1 140360
box 0 0 3190 3190
use unit_cap  unit_cap_461
timestamp 1662145021
transform 1 0 25520 0 1 143550
box 0 0 3190 3190
use unit_cap  unit_cap_462
timestamp 1662145021
transform 1 0 25520 0 1 146740
box 0 0 3190 3190
use unit_cap  unit_cap_463
timestamp 1662145021
transform 1 0 25520 0 1 149930
box 0 0 3190 3190
use unit_cap  unit_cap_464
timestamp 1662145021
transform 1 0 25520 0 1 153120
box 0 0 3190 3190
use unit_cap  unit_cap_465
timestamp 1662145021
transform 1 0 25520 0 1 156310
box 0 0 3190 3190
use unit_cap  unit_cap_466
timestamp 1662145021
transform 1 0 25520 0 1 159500
box 0 0 3190 3190
use unit_cap  unit_cap_467
timestamp 1662145021
transform 1 0 25520 0 1 162690
box 0 0 3190 3190
use unit_cap  unit_cap_468
timestamp 1662145021
transform 1 0 28710 0 1 0
box 0 0 3190 3190
use unit_cap  unit_cap_469
timestamp 1662145021
transform 1 0 28710 0 1 3190
box 0 0 3190 3190
use unit_cap  unit_cap_470
timestamp 1662145021
transform 1 0 28710 0 1 6380
box 0 0 3190 3190
use unit_cap  unit_cap_471
timestamp 1662145021
transform 1 0 28710 0 1 9570
box 0 0 3190 3190
use unit_cap  unit_cap_472
timestamp 1662145021
transform 1 0 28710 0 1 12760
box 0 0 3190 3190
use unit_cap  unit_cap_473
timestamp 1662145021
transform 1 0 28710 0 1 15950
box 0 0 3190 3190
use unit_cap  unit_cap_474
timestamp 1662145021
transform 1 0 28710 0 1 19140
box 0 0 3190 3190
use unit_cap  unit_cap_475
timestamp 1662145021
transform 1 0 28710 0 1 22330
box 0 0 3190 3190
use unit_cap  unit_cap_476
timestamp 1662145021
transform 1 0 28710 0 1 25520
box 0 0 3190 3190
use unit_cap  unit_cap_477
timestamp 1662145021
transform 1 0 28710 0 1 28710
box 0 0 3190 3190
use unit_cap  unit_cap_478
timestamp 1662145021
transform 1 0 28710 0 1 31900
box 0 0 3190 3190
use unit_cap  unit_cap_479
timestamp 1662145021
transform 1 0 28710 0 1 35090
box 0 0 3190 3190
use unit_cap  unit_cap_480
timestamp 1662145021
transform 1 0 28710 0 1 38280
box 0 0 3190 3190
use unit_cap  unit_cap_481
timestamp 1662145021
transform 1 0 28710 0 1 41470
box 0 0 3190 3190
use unit_cap  unit_cap_482
timestamp 1662145021
transform 1 0 28710 0 1 44660
box 0 0 3190 3190
use unit_cap  unit_cap_483
timestamp 1662145021
transform 1 0 28710 0 1 47850
box 0 0 3190 3190
use unit_cap  unit_cap_484
timestamp 1662145021
transform 1 0 28710 0 1 51040
box 0 0 3190 3190
use unit_cap  unit_cap_485
timestamp 1662145021
transform 1 0 28710 0 1 54230
box 0 0 3190 3190
use unit_cap  unit_cap_486
timestamp 1662145021
transform 1 0 28710 0 1 57420
box 0 0 3190 3190
use unit_cap  unit_cap_487
timestamp 1662145021
transform 1 0 28710 0 1 60610
box 0 0 3190 3190
use unit_cap  unit_cap_488
timestamp 1662145021
transform 1 0 28710 0 1 63800
box 0 0 3190 3190
use unit_cap  unit_cap_489
timestamp 1662145021
transform 1 0 28710 0 1 66990
box 0 0 3190 3190
use unit_cap  unit_cap_490
timestamp 1662145021
transform 1 0 28710 0 1 70180
box 0 0 3190 3190
use unit_cap  unit_cap_491
timestamp 1662145021
transform 1 0 28710 0 1 73370
box 0 0 3190 3190
use unit_cap  unit_cap_492
timestamp 1662145021
transform 1 0 28710 0 1 76560
box 0 0 3190 3190
use unit_cap  unit_cap_493
timestamp 1662145021
transform 1 0 28710 0 1 79750
box 0 0 3190 3190
use unit_cap  unit_cap_494
timestamp 1662145021
transform 1 0 28710 0 1 82940
box 0 0 3190 3190
use unit_cap  unit_cap_495
timestamp 1662145021
transform 1 0 28710 0 1 86130
box 0 0 3190 3190
use unit_cap  unit_cap_496
timestamp 1662145021
transform 1 0 28710 0 1 89320
box 0 0 3190 3190
use unit_cap  unit_cap_497
timestamp 1662145021
transform 1 0 28710 0 1 92510
box 0 0 3190 3190
use unit_cap  unit_cap_498
timestamp 1662145021
transform 1 0 28710 0 1 95700
box 0 0 3190 3190
use unit_cap  unit_cap_499
timestamp 1662145021
transform 1 0 28710 0 1 98890
box 0 0 3190 3190
use unit_cap  unit_cap_500
timestamp 1662145021
transform 1 0 28710 0 1 102080
box 0 0 3190 3190
use unit_cap  unit_cap_501
timestamp 1662145021
transform 1 0 28710 0 1 105270
box 0 0 3190 3190
use unit_cap  unit_cap_502
timestamp 1662145021
transform 1 0 28710 0 1 108460
box 0 0 3190 3190
use unit_cap  unit_cap_503
timestamp 1662145021
transform 1 0 28710 0 1 111650
box 0 0 3190 3190
use unit_cap  unit_cap_504
timestamp 1662145021
transform 1 0 28710 0 1 114840
box 0 0 3190 3190
use unit_cap  unit_cap_505
timestamp 1662145021
transform 1 0 28710 0 1 118030
box 0 0 3190 3190
use unit_cap  unit_cap_506
timestamp 1662145021
transform 1 0 28710 0 1 121220
box 0 0 3190 3190
use unit_cap  unit_cap_507
timestamp 1662145021
transform 1 0 28710 0 1 124410
box 0 0 3190 3190
use unit_cap  unit_cap_508
timestamp 1662145021
transform 1 0 28710 0 1 127600
box 0 0 3190 3190
use unit_cap  unit_cap_509
timestamp 1662145021
transform 1 0 28710 0 1 130790
box 0 0 3190 3190
use unit_cap  unit_cap_510
timestamp 1662145021
transform 1 0 28710 0 1 133980
box 0 0 3190 3190
use unit_cap  unit_cap_511
timestamp 1662145021
transform 1 0 28710 0 1 137170
box 0 0 3190 3190
use unit_cap  unit_cap_512
timestamp 1662145021
transform 1 0 28710 0 1 140360
box 0 0 3190 3190
use unit_cap  unit_cap_513
timestamp 1662145021
transform 1 0 28710 0 1 143550
box 0 0 3190 3190
use unit_cap  unit_cap_514
timestamp 1662145021
transform 1 0 28710 0 1 146740
box 0 0 3190 3190
use unit_cap  unit_cap_515
timestamp 1662145021
transform 1 0 28710 0 1 149930
box 0 0 3190 3190
use unit_cap  unit_cap_516
timestamp 1662145021
transform 1 0 28710 0 1 153120
box 0 0 3190 3190
use unit_cap  unit_cap_517
timestamp 1662145021
transform 1 0 28710 0 1 156310
box 0 0 3190 3190
use unit_cap  unit_cap_518
timestamp 1662145021
transform 1 0 28710 0 1 159500
box 0 0 3190 3190
use unit_cap  unit_cap_519
timestamp 1662145021
transform 1 0 28710 0 1 162690
box 0 0 3190 3190
use unit_cap  unit_cap_520
timestamp 1662145021
transform 1 0 31900 0 1 0
box 0 0 3190 3190
use unit_cap  unit_cap_521
timestamp 1662145021
transform 1 0 31900 0 1 3190
box 0 0 3190 3190
use unit_cap  unit_cap_522
timestamp 1662145021
transform 1 0 31900 0 1 6380
box 0 0 3190 3190
use unit_cap  unit_cap_523
timestamp 1662145021
transform 1 0 31900 0 1 9570
box 0 0 3190 3190
use unit_cap  unit_cap_524
timestamp 1662145021
transform 1 0 31900 0 1 12760
box 0 0 3190 3190
use unit_cap  unit_cap_525
timestamp 1662145021
transform 1 0 31900 0 1 15950
box 0 0 3190 3190
use unit_cap  unit_cap_526
timestamp 1662145021
transform 1 0 31900 0 1 19140
box 0 0 3190 3190
use unit_cap  unit_cap_527
timestamp 1662145021
transform 1 0 31900 0 1 22330
box 0 0 3190 3190
use unit_cap  unit_cap_528
timestamp 1662145021
transform 1 0 31900 0 1 25520
box 0 0 3190 3190
use unit_cap  unit_cap_529
timestamp 1662145021
transform 1 0 31900 0 1 28710
box 0 0 3190 3190
use unit_cap  unit_cap_530
timestamp 1662145021
transform 1 0 31900 0 1 31900
box 0 0 3190 3190
use unit_cap  unit_cap_531
timestamp 1662145021
transform 1 0 31900 0 1 35090
box 0 0 3190 3190
use unit_cap  unit_cap_532
timestamp 1662145021
transform 1 0 31900 0 1 38280
box 0 0 3190 3190
use unit_cap  unit_cap_533
timestamp 1662145021
transform 1 0 31900 0 1 41470
box 0 0 3190 3190
use unit_cap  unit_cap_534
timestamp 1662145021
transform 1 0 31900 0 1 44660
box 0 0 3190 3190
use unit_cap  unit_cap_535
timestamp 1662145021
transform 1 0 31900 0 1 47850
box 0 0 3190 3190
use unit_cap  unit_cap_536
timestamp 1662145021
transform 1 0 31900 0 1 51040
box 0 0 3190 3190
use unit_cap  unit_cap_537
timestamp 1662145021
transform 1 0 31900 0 1 54230
box 0 0 3190 3190
use unit_cap  unit_cap_538
timestamp 1662145021
transform 1 0 31900 0 1 57420
box 0 0 3190 3190
use unit_cap  unit_cap_539
timestamp 1662145021
transform 1 0 31900 0 1 60610
box 0 0 3190 3190
use unit_cap  unit_cap_540
timestamp 1662145021
transform 1 0 31900 0 1 63800
box 0 0 3190 3190
use unit_cap  unit_cap_541
timestamp 1662145021
transform 1 0 31900 0 1 66990
box 0 0 3190 3190
use unit_cap  unit_cap_542
timestamp 1662145021
transform 1 0 31900 0 1 70180
box 0 0 3190 3190
use unit_cap  unit_cap_543
timestamp 1662145021
transform 1 0 31900 0 1 73370
box 0 0 3190 3190
use unit_cap  unit_cap_544
timestamp 1662145021
transform 1 0 31900 0 1 76560
box 0 0 3190 3190
use unit_cap  unit_cap_545
timestamp 1662145021
transform 1 0 31900 0 1 79750
box 0 0 3190 3190
use unit_cap  unit_cap_546
timestamp 1662145021
transform 1 0 31900 0 1 82940
box 0 0 3190 3190
use unit_cap  unit_cap_547
timestamp 1662145021
transform 1 0 31900 0 1 86130
box 0 0 3190 3190
use unit_cap  unit_cap_548
timestamp 1662145021
transform 1 0 31900 0 1 89320
box 0 0 3190 3190
use unit_cap  unit_cap_549
timestamp 1662145021
transform 1 0 31900 0 1 92510
box 0 0 3190 3190
use unit_cap  unit_cap_550
timestamp 1662145021
transform 1 0 31900 0 1 95700
box 0 0 3190 3190
use unit_cap  unit_cap_551
timestamp 1662145021
transform 1 0 31900 0 1 98890
box 0 0 3190 3190
use unit_cap  unit_cap_552
timestamp 1662145021
transform 1 0 31900 0 1 102080
box 0 0 3190 3190
use unit_cap  unit_cap_553
timestamp 1662145021
transform 1 0 31900 0 1 105270
box 0 0 3190 3190
use unit_cap  unit_cap_554
timestamp 1662145021
transform 1 0 31900 0 1 108460
box 0 0 3190 3190
use unit_cap  unit_cap_555
timestamp 1662145021
transform 1 0 31900 0 1 111650
box 0 0 3190 3190
use unit_cap  unit_cap_556
timestamp 1662145021
transform 1 0 31900 0 1 114840
box 0 0 3190 3190
use unit_cap  unit_cap_557
timestamp 1662145021
transform 1 0 31900 0 1 118030
box 0 0 3190 3190
use unit_cap  unit_cap_558
timestamp 1662145021
transform 1 0 31900 0 1 121220
box 0 0 3190 3190
use unit_cap  unit_cap_559
timestamp 1662145021
transform 1 0 31900 0 1 124410
box 0 0 3190 3190
use unit_cap  unit_cap_560
timestamp 1662145021
transform 1 0 31900 0 1 127600
box 0 0 3190 3190
use unit_cap  unit_cap_561
timestamp 1662145021
transform 1 0 31900 0 1 130790
box 0 0 3190 3190
use unit_cap  unit_cap_562
timestamp 1662145021
transform 1 0 31900 0 1 133980
box 0 0 3190 3190
use unit_cap  unit_cap_563
timestamp 1662145021
transform 1 0 31900 0 1 137170
box 0 0 3190 3190
use unit_cap  unit_cap_564
timestamp 1662145021
transform 1 0 31900 0 1 140360
box 0 0 3190 3190
use unit_cap  unit_cap_565
timestamp 1662145021
transform 1 0 31900 0 1 143550
box 0 0 3190 3190
use unit_cap  unit_cap_566
timestamp 1662145021
transform 1 0 31900 0 1 146740
box 0 0 3190 3190
use unit_cap  unit_cap_567
timestamp 1662145021
transform 1 0 31900 0 1 149930
box 0 0 3190 3190
use unit_cap  unit_cap_568
timestamp 1662145021
transform 1 0 31900 0 1 153120
box 0 0 3190 3190
use unit_cap  unit_cap_569
timestamp 1662145021
transform 1 0 31900 0 1 156310
box 0 0 3190 3190
use unit_cap  unit_cap_570
timestamp 1662145021
transform 1 0 31900 0 1 159500
box 0 0 3190 3190
use unit_cap  unit_cap_571
timestamp 1662145021
transform 1 0 31900 0 1 162690
box 0 0 3190 3190
use unit_cap  unit_cap_572
timestamp 1662145021
transform 1 0 35090 0 1 0
box 0 0 3190 3190
use unit_cap  unit_cap_573
timestamp 1662145021
transform 1 0 35090 0 1 3190
box 0 0 3190 3190
use unit_cap  unit_cap_574
timestamp 1662145021
transform 1 0 35090 0 1 6380
box 0 0 3190 3190
use unit_cap  unit_cap_575
timestamp 1662145021
transform 1 0 35090 0 1 9570
box 0 0 3190 3190
use unit_cap  unit_cap_576
timestamp 1662145021
transform 1 0 35090 0 1 12760
box 0 0 3190 3190
use unit_cap  unit_cap_577
timestamp 1662145021
transform 1 0 35090 0 1 15950
box 0 0 3190 3190
use unit_cap  unit_cap_578
timestamp 1662145021
transform 1 0 35090 0 1 19140
box 0 0 3190 3190
use unit_cap  unit_cap_579
timestamp 1662145021
transform 1 0 35090 0 1 22330
box 0 0 3190 3190
use unit_cap  unit_cap_580
timestamp 1662145021
transform 1 0 35090 0 1 25520
box 0 0 3190 3190
use unit_cap  unit_cap_581
timestamp 1662145021
transform 1 0 35090 0 1 28710
box 0 0 3190 3190
use unit_cap  unit_cap_582
timestamp 1662145021
transform 1 0 35090 0 1 31900
box 0 0 3190 3190
use unit_cap  unit_cap_583
timestamp 1662145021
transform 1 0 35090 0 1 35090
box 0 0 3190 3190
use unit_cap  unit_cap_584
timestamp 1662145021
transform 1 0 35090 0 1 38280
box 0 0 3190 3190
use unit_cap  unit_cap_585
timestamp 1662145021
transform 1 0 35090 0 1 41470
box 0 0 3190 3190
use unit_cap  unit_cap_586
timestamp 1662145021
transform 1 0 35090 0 1 44660
box 0 0 3190 3190
use unit_cap  unit_cap_587
timestamp 1662145021
transform 1 0 35090 0 1 47850
box 0 0 3190 3190
use unit_cap  unit_cap_588
timestamp 1662145021
transform 1 0 35090 0 1 51040
box 0 0 3190 3190
use unit_cap  unit_cap_589
timestamp 1662145021
transform 1 0 35090 0 1 54230
box 0 0 3190 3190
use unit_cap  unit_cap_590
timestamp 1662145021
transform 1 0 35090 0 1 57420
box 0 0 3190 3190
use unit_cap  unit_cap_591
timestamp 1662145021
transform 1 0 35090 0 1 60610
box 0 0 3190 3190
use unit_cap  unit_cap_592
timestamp 1662145021
transform 1 0 35090 0 1 63800
box 0 0 3190 3190
use unit_cap  unit_cap_593
timestamp 1662145021
transform 1 0 35090 0 1 66990
box 0 0 3190 3190
use unit_cap  unit_cap_594
timestamp 1662145021
transform 1 0 35090 0 1 70180
box 0 0 3190 3190
use unit_cap  unit_cap_595
timestamp 1662145021
transform 1 0 35090 0 1 73370
box 0 0 3190 3190
use unit_cap  unit_cap_596
timestamp 1662145021
transform 1 0 35090 0 1 76560
box 0 0 3190 3190
use unit_cap  unit_cap_597
timestamp 1662145021
transform 1 0 35090 0 1 79750
box 0 0 3190 3190
use unit_cap  unit_cap_598
timestamp 1662145021
transform 1 0 35090 0 1 82940
box 0 0 3190 3190
use unit_cap  unit_cap_599
timestamp 1662145021
transform 1 0 35090 0 1 86130
box 0 0 3190 3190
use unit_cap  unit_cap_600
timestamp 1662145021
transform 1 0 35090 0 1 89320
box 0 0 3190 3190
use unit_cap  unit_cap_601
timestamp 1662145021
transform 1 0 35090 0 1 92510
box 0 0 3190 3190
use unit_cap  unit_cap_602
timestamp 1662145021
transform 1 0 35090 0 1 95700
box 0 0 3190 3190
use unit_cap  unit_cap_603
timestamp 1662145021
transform 1 0 35090 0 1 98890
box 0 0 3190 3190
use unit_cap  unit_cap_604
timestamp 1662145021
transform 1 0 35090 0 1 102080
box 0 0 3190 3190
use unit_cap  unit_cap_605
timestamp 1662145021
transform 1 0 35090 0 1 105270
box 0 0 3190 3190
use unit_cap  unit_cap_606
timestamp 1662145021
transform 1 0 35090 0 1 108460
box 0 0 3190 3190
use unit_cap  unit_cap_607
timestamp 1662145021
transform 1 0 35090 0 1 111650
box 0 0 3190 3190
use unit_cap  unit_cap_608
timestamp 1662145021
transform 1 0 35090 0 1 114840
box 0 0 3190 3190
use unit_cap  unit_cap_609
timestamp 1662145021
transform 1 0 35090 0 1 118030
box 0 0 3190 3190
use unit_cap  unit_cap_610
timestamp 1662145021
transform 1 0 35090 0 1 121220
box 0 0 3190 3190
use unit_cap  unit_cap_611
timestamp 1662145021
transform 1 0 35090 0 1 124410
box 0 0 3190 3190
use unit_cap  unit_cap_612
timestamp 1662145021
transform 1 0 35090 0 1 127600
box 0 0 3190 3190
use unit_cap  unit_cap_613
timestamp 1662145021
transform 1 0 35090 0 1 130790
box 0 0 3190 3190
use unit_cap  unit_cap_614
timestamp 1662145021
transform 1 0 35090 0 1 133980
box 0 0 3190 3190
use unit_cap  unit_cap_615
timestamp 1662145021
transform 1 0 35090 0 1 137170
box 0 0 3190 3190
use unit_cap  unit_cap_616
timestamp 1662145021
transform 1 0 35090 0 1 140360
box 0 0 3190 3190
use unit_cap  unit_cap_617
timestamp 1662145021
transform 1 0 35090 0 1 143550
box 0 0 3190 3190
use unit_cap  unit_cap_618
timestamp 1662145021
transform 1 0 35090 0 1 146740
box 0 0 3190 3190
use unit_cap  unit_cap_619
timestamp 1662145021
transform 1 0 35090 0 1 149930
box 0 0 3190 3190
use unit_cap  unit_cap_620
timestamp 1662145021
transform 1 0 35090 0 1 153120
box 0 0 3190 3190
use unit_cap  unit_cap_621
timestamp 1662145021
transform 1 0 35090 0 1 156310
box 0 0 3190 3190
use unit_cap  unit_cap_622
timestamp 1662145021
transform 1 0 35090 0 1 159500
box 0 0 3190 3190
use unit_cap  unit_cap_623
timestamp 1662145021
transform 1 0 35090 0 1 162690
box 0 0 3190 3190
use unit_cap  unit_cap_624
timestamp 1662145021
transform 1 0 38280 0 1 0
box 0 0 3190 3190
use unit_cap  unit_cap_625
timestamp 1662145021
transform 1 0 38280 0 1 3190
box 0 0 3190 3190
use unit_cap  unit_cap_626
timestamp 1662145021
transform 1 0 38280 0 1 6380
box 0 0 3190 3190
use unit_cap  unit_cap_627
timestamp 1662145021
transform 1 0 38280 0 1 9570
box 0 0 3190 3190
use unit_cap  unit_cap_628
timestamp 1662145021
transform 1 0 38280 0 1 12760
box 0 0 3190 3190
use unit_cap  unit_cap_629
timestamp 1662145021
transform 1 0 38280 0 1 15950
box 0 0 3190 3190
use unit_cap  unit_cap_630
timestamp 1662145021
transform 1 0 38280 0 1 19140
box 0 0 3190 3190
use unit_cap  unit_cap_631
timestamp 1662145021
transform 1 0 38280 0 1 22330
box 0 0 3190 3190
use unit_cap  unit_cap_632
timestamp 1662145021
transform 1 0 38280 0 1 25520
box 0 0 3190 3190
use unit_cap  unit_cap_633
timestamp 1662145021
transform 1 0 38280 0 1 28710
box 0 0 3190 3190
use unit_cap  unit_cap_634
timestamp 1662145021
transform 1 0 38280 0 1 31900
box 0 0 3190 3190
use unit_cap  unit_cap_635
timestamp 1662145021
transform 1 0 38280 0 1 35090
box 0 0 3190 3190
use unit_cap  unit_cap_636
timestamp 1662145021
transform 1 0 38280 0 1 38280
box 0 0 3190 3190
use unit_cap  unit_cap_637
timestamp 1662145021
transform 1 0 38280 0 1 41470
box 0 0 3190 3190
use unit_cap  unit_cap_638
timestamp 1662145021
transform 1 0 38280 0 1 44660
box 0 0 3190 3190
use unit_cap  unit_cap_639
timestamp 1662145021
transform 1 0 38280 0 1 47850
box 0 0 3190 3190
use unit_cap  unit_cap_640
timestamp 1662145021
transform 1 0 38280 0 1 51040
box 0 0 3190 3190
use unit_cap  unit_cap_641
timestamp 1662145021
transform 1 0 38280 0 1 54230
box 0 0 3190 3190
use unit_cap  unit_cap_642
timestamp 1662145021
transform 1 0 38280 0 1 57420
box 0 0 3190 3190
use unit_cap  unit_cap_643
timestamp 1662145021
transform 1 0 38280 0 1 60610
box 0 0 3190 3190
use unit_cap  unit_cap_644
timestamp 1662145021
transform 1 0 38280 0 1 63800
box 0 0 3190 3190
use unit_cap  unit_cap_645
timestamp 1662145021
transform 1 0 38280 0 1 66990
box 0 0 3190 3190
use unit_cap  unit_cap_646
timestamp 1662145021
transform 1 0 38280 0 1 70180
box 0 0 3190 3190
use unit_cap  unit_cap_647
timestamp 1662145021
transform 1 0 38280 0 1 73370
box 0 0 3190 3190
use unit_cap  unit_cap_648
timestamp 1662145021
transform 1 0 38280 0 1 76560
box 0 0 3190 3190
use unit_cap  unit_cap_649
timestamp 1662145021
transform 1 0 38280 0 1 79750
box 0 0 3190 3190
use unit_cap  unit_cap_650
timestamp 1662145021
transform 1 0 38280 0 1 82940
box 0 0 3190 3190
use unit_cap  unit_cap_651
timestamp 1662145021
transform 1 0 38280 0 1 86130
box 0 0 3190 3190
use unit_cap  unit_cap_652
timestamp 1662145021
transform 1 0 38280 0 1 89320
box 0 0 3190 3190
use unit_cap  unit_cap_653
timestamp 1662145021
transform 1 0 38280 0 1 92510
box 0 0 3190 3190
use unit_cap  unit_cap_654
timestamp 1662145021
transform 1 0 38280 0 1 95700
box 0 0 3190 3190
use unit_cap  unit_cap_655
timestamp 1662145021
transform 1 0 38280 0 1 98890
box 0 0 3190 3190
use unit_cap  unit_cap_656
timestamp 1662145021
transform 1 0 38280 0 1 102080
box 0 0 3190 3190
use unit_cap  unit_cap_657
timestamp 1662145021
transform 1 0 38280 0 1 105270
box 0 0 3190 3190
use unit_cap  unit_cap_658
timestamp 1662145021
transform 1 0 38280 0 1 108460
box 0 0 3190 3190
use unit_cap  unit_cap_659
timestamp 1662145021
transform 1 0 38280 0 1 111650
box 0 0 3190 3190
use unit_cap  unit_cap_660
timestamp 1662145021
transform 1 0 38280 0 1 114840
box 0 0 3190 3190
use unit_cap  unit_cap_661
timestamp 1662145021
transform 1 0 38280 0 1 118030
box 0 0 3190 3190
use unit_cap  unit_cap_662
timestamp 1662145021
transform 1 0 38280 0 1 121220
box 0 0 3190 3190
use unit_cap  unit_cap_663
timestamp 1662145021
transform 1 0 38280 0 1 124410
box 0 0 3190 3190
use unit_cap  unit_cap_664
timestamp 1662145021
transform 1 0 38280 0 1 127600
box 0 0 3190 3190
use unit_cap  unit_cap_665
timestamp 1662145021
transform 1 0 38280 0 1 130790
box 0 0 3190 3190
use unit_cap  unit_cap_666
timestamp 1662145021
transform 1 0 38280 0 1 133980
box 0 0 3190 3190
use unit_cap  unit_cap_667
timestamp 1662145021
transform 1 0 38280 0 1 137170
box 0 0 3190 3190
use unit_cap  unit_cap_668
timestamp 1662145021
transform 1 0 38280 0 1 140360
box 0 0 3190 3190
use unit_cap  unit_cap_669
timestamp 1662145021
transform 1 0 38280 0 1 143550
box 0 0 3190 3190
use unit_cap  unit_cap_670
timestamp 1662145021
transform 1 0 38280 0 1 146740
box 0 0 3190 3190
use unit_cap  unit_cap_671
timestamp 1662145021
transform 1 0 38280 0 1 149930
box 0 0 3190 3190
use unit_cap  unit_cap_672
timestamp 1662145021
transform 1 0 38280 0 1 153120
box 0 0 3190 3190
use unit_cap  unit_cap_673
timestamp 1662145021
transform 1 0 38280 0 1 156310
box 0 0 3190 3190
use unit_cap  unit_cap_674
timestamp 1662145021
transform 1 0 38280 0 1 159500
box 0 0 3190 3190
use unit_cap  unit_cap_675
timestamp 1662145021
transform 1 0 38280 0 1 162690
box 0 0 3190 3190
use unit_cap  unit_cap_676
timestamp 1662145021
transform 1 0 41470 0 1 0
box 0 0 3190 3190
use unit_cap  unit_cap_677
timestamp 1662145021
transform 1 0 41470 0 1 3190
box 0 0 3190 3190
use unit_cap  unit_cap_678
timestamp 1662145021
transform 1 0 41470 0 1 6380
box 0 0 3190 3190
use unit_cap  unit_cap_679
timestamp 1662145021
transform 1 0 41470 0 1 9570
box 0 0 3190 3190
use unit_cap  unit_cap_680
timestamp 1662145021
transform 1 0 41470 0 1 12760
box 0 0 3190 3190
use unit_cap  unit_cap_681
timestamp 1662145021
transform 1 0 41470 0 1 15950
box 0 0 3190 3190
use unit_cap  unit_cap_682
timestamp 1662145021
transform 1 0 41470 0 1 19140
box 0 0 3190 3190
use unit_cap  unit_cap_683
timestamp 1662145021
transform 1 0 41470 0 1 22330
box 0 0 3190 3190
use unit_cap  unit_cap_684
timestamp 1662145021
transform 1 0 41470 0 1 25520
box 0 0 3190 3190
use unit_cap  unit_cap_685
timestamp 1662145021
transform 1 0 41470 0 1 28710
box 0 0 3190 3190
use unit_cap  unit_cap_686
timestamp 1662145021
transform 1 0 41470 0 1 31900
box 0 0 3190 3190
use unit_cap  unit_cap_687
timestamp 1662145021
transform 1 0 41470 0 1 35090
box 0 0 3190 3190
use unit_cap  unit_cap_688
timestamp 1662145021
transform 1 0 41470 0 1 38280
box 0 0 3190 3190
use unit_cap  unit_cap_689
timestamp 1662145021
transform 1 0 41470 0 1 41470
box 0 0 3190 3190
use unit_cap  unit_cap_690
timestamp 1662145021
transform 1 0 41470 0 1 44660
box 0 0 3190 3190
use unit_cap  unit_cap_691
timestamp 1662145021
transform 1 0 41470 0 1 47850
box 0 0 3190 3190
use unit_cap  unit_cap_692
timestamp 1662145021
transform 1 0 41470 0 1 51040
box 0 0 3190 3190
use unit_cap  unit_cap_693
timestamp 1662145021
transform 1 0 41470 0 1 54230
box 0 0 3190 3190
use unit_cap  unit_cap_694
timestamp 1662145021
transform 1 0 41470 0 1 57420
box 0 0 3190 3190
use unit_cap  unit_cap_695
timestamp 1662145021
transform 1 0 41470 0 1 60610
box 0 0 3190 3190
use unit_cap  unit_cap_696
timestamp 1662145021
transform 1 0 41470 0 1 63800
box 0 0 3190 3190
use unit_cap  unit_cap_697
timestamp 1662145021
transform 1 0 41470 0 1 66990
box 0 0 3190 3190
use unit_cap  unit_cap_698
timestamp 1662145021
transform 1 0 41470 0 1 70180
box 0 0 3190 3190
use unit_cap  unit_cap_699
timestamp 1662145021
transform 1 0 41470 0 1 73370
box 0 0 3190 3190
use unit_cap  unit_cap_700
timestamp 1662145021
transform 1 0 41470 0 1 76560
box 0 0 3190 3190
use unit_cap  unit_cap_701
timestamp 1662145021
transform 1 0 41470 0 1 79750
box 0 0 3190 3190
use unit_cap  unit_cap_702
timestamp 1662145021
transform 1 0 41470 0 1 82940
box 0 0 3190 3190
use unit_cap  unit_cap_703
timestamp 1662145021
transform 1 0 41470 0 1 86130
box 0 0 3190 3190
use unit_cap  unit_cap_704
timestamp 1662145021
transform 1 0 41470 0 1 89320
box 0 0 3190 3190
use unit_cap  unit_cap_705
timestamp 1662145021
transform 1 0 41470 0 1 92510
box 0 0 3190 3190
use unit_cap  unit_cap_706
timestamp 1662145021
transform 1 0 41470 0 1 95700
box 0 0 3190 3190
use unit_cap  unit_cap_707
timestamp 1662145021
transform 1 0 41470 0 1 98890
box 0 0 3190 3190
use unit_cap  unit_cap_708
timestamp 1662145021
transform 1 0 41470 0 1 102080
box 0 0 3190 3190
use unit_cap  unit_cap_709
timestamp 1662145021
transform 1 0 41470 0 1 105270
box 0 0 3190 3190
use unit_cap  unit_cap_710
timestamp 1662145021
transform 1 0 41470 0 1 108460
box 0 0 3190 3190
use unit_cap  unit_cap_711
timestamp 1662145021
transform 1 0 41470 0 1 111650
box 0 0 3190 3190
use unit_cap  unit_cap_712
timestamp 1662145021
transform 1 0 41470 0 1 114840
box 0 0 3190 3190
use unit_cap  unit_cap_713
timestamp 1662145021
transform 1 0 41470 0 1 118030
box 0 0 3190 3190
use unit_cap  unit_cap_714
timestamp 1662145021
transform 1 0 41470 0 1 121220
box 0 0 3190 3190
use unit_cap  unit_cap_715
timestamp 1662145021
transform 1 0 41470 0 1 124410
box 0 0 3190 3190
use unit_cap  unit_cap_716
timestamp 1662145021
transform 1 0 41470 0 1 127600
box 0 0 3190 3190
use unit_cap  unit_cap_717
timestamp 1662145021
transform 1 0 41470 0 1 130790
box 0 0 3190 3190
use unit_cap  unit_cap_718
timestamp 1662145021
transform 1 0 41470 0 1 133980
box 0 0 3190 3190
use unit_cap  unit_cap_719
timestamp 1662145021
transform 1 0 41470 0 1 137170
box 0 0 3190 3190
use unit_cap  unit_cap_720
timestamp 1662145021
transform 1 0 41470 0 1 140360
box 0 0 3190 3190
use unit_cap  unit_cap_721
timestamp 1662145021
transform 1 0 41470 0 1 143550
box 0 0 3190 3190
use unit_cap  unit_cap_722
timestamp 1662145021
transform 1 0 41470 0 1 146740
box 0 0 3190 3190
use unit_cap  unit_cap_723
timestamp 1662145021
transform 1 0 41470 0 1 149930
box 0 0 3190 3190
use unit_cap  unit_cap_724
timestamp 1662145021
transform 1 0 41470 0 1 153120
box 0 0 3190 3190
use unit_cap  unit_cap_725
timestamp 1662145021
transform 1 0 41470 0 1 156310
box 0 0 3190 3190
use unit_cap  unit_cap_726
timestamp 1662145021
transform 1 0 41470 0 1 159500
box 0 0 3190 3190
use unit_cap  unit_cap_727
timestamp 1662145021
transform 1 0 41470 0 1 162690
box 0 0 3190 3190
use unit_cap  unit_cap_728
timestamp 1662145021
transform 1 0 44660 0 1 0
box 0 0 3190 3190
use unit_cap  unit_cap_729
timestamp 1662145021
transform 1 0 44660 0 1 3190
box 0 0 3190 3190
use unit_cap  unit_cap_730
timestamp 1662145021
transform 1 0 44660 0 1 6380
box 0 0 3190 3190
use unit_cap  unit_cap_731
timestamp 1662145021
transform 1 0 44660 0 1 9570
box 0 0 3190 3190
use unit_cap  unit_cap_732
timestamp 1662145021
transform 1 0 44660 0 1 12760
box 0 0 3190 3190
use unit_cap  unit_cap_733
timestamp 1662145021
transform 1 0 44660 0 1 15950
box 0 0 3190 3190
use unit_cap  unit_cap_734
timestamp 1662145021
transform 1 0 44660 0 1 19140
box 0 0 3190 3190
use unit_cap  unit_cap_735
timestamp 1662145021
transform 1 0 44660 0 1 22330
box 0 0 3190 3190
use unit_cap  unit_cap_736
timestamp 1662145021
transform 1 0 44660 0 1 25520
box 0 0 3190 3190
use unit_cap  unit_cap_737
timestamp 1662145021
transform 1 0 44660 0 1 28710
box 0 0 3190 3190
use unit_cap  unit_cap_738
timestamp 1662145021
transform 1 0 44660 0 1 31900
box 0 0 3190 3190
use unit_cap  unit_cap_739
timestamp 1662145021
transform 1 0 44660 0 1 35090
box 0 0 3190 3190
use unit_cap  unit_cap_740
timestamp 1662145021
transform 1 0 44660 0 1 38280
box 0 0 3190 3190
use unit_cap  unit_cap_741
timestamp 1662145021
transform 1 0 44660 0 1 41470
box 0 0 3190 3190
use unit_cap  unit_cap_742
timestamp 1662145021
transform 1 0 44660 0 1 44660
box 0 0 3190 3190
use unit_cap  unit_cap_743
timestamp 1662145021
transform 1 0 44660 0 1 47850
box 0 0 3190 3190
use unit_cap  unit_cap_744
timestamp 1662145021
transform 1 0 44660 0 1 51040
box 0 0 3190 3190
use unit_cap  unit_cap_745
timestamp 1662145021
transform 1 0 44660 0 1 54230
box 0 0 3190 3190
use unit_cap  unit_cap_746
timestamp 1662145021
transform 1 0 44660 0 1 57420
box 0 0 3190 3190
use unit_cap  unit_cap_747
timestamp 1662145021
transform 1 0 44660 0 1 60610
box 0 0 3190 3190
use unit_cap  unit_cap_748
timestamp 1662145021
transform 1 0 44660 0 1 63800
box 0 0 3190 3190
use unit_cap  unit_cap_749
timestamp 1662145021
transform 1 0 44660 0 1 66990
box 0 0 3190 3190
use unit_cap  unit_cap_750
timestamp 1662145021
transform 1 0 44660 0 1 70180
box 0 0 3190 3190
use unit_cap  unit_cap_751
timestamp 1662145021
transform 1 0 44660 0 1 73370
box 0 0 3190 3190
use unit_cap  unit_cap_752
timestamp 1662145021
transform 1 0 44660 0 1 76560
box 0 0 3190 3190
use unit_cap  unit_cap_753
timestamp 1662145021
transform 1 0 44660 0 1 79750
box 0 0 3190 3190
use unit_cap  unit_cap_754
timestamp 1662145021
transform 1 0 44660 0 1 82940
box 0 0 3190 3190
use unit_cap  unit_cap_755
timestamp 1662145021
transform 1 0 44660 0 1 86130
box 0 0 3190 3190
use unit_cap  unit_cap_756
timestamp 1662145021
transform 1 0 44660 0 1 89320
box 0 0 3190 3190
use unit_cap  unit_cap_757
timestamp 1662145021
transform 1 0 44660 0 1 92510
box 0 0 3190 3190
use unit_cap  unit_cap_758
timestamp 1662145021
transform 1 0 44660 0 1 95700
box 0 0 3190 3190
use unit_cap  unit_cap_759
timestamp 1662145021
transform 1 0 44660 0 1 98890
box 0 0 3190 3190
use unit_cap  unit_cap_760
timestamp 1662145021
transform 1 0 44660 0 1 102080
box 0 0 3190 3190
use unit_cap  unit_cap_761
timestamp 1662145021
transform 1 0 44660 0 1 105270
box 0 0 3190 3190
use unit_cap  unit_cap_762
timestamp 1662145021
transform 1 0 44660 0 1 108460
box 0 0 3190 3190
use unit_cap  unit_cap_763
timestamp 1662145021
transform 1 0 44660 0 1 111650
box 0 0 3190 3190
use unit_cap  unit_cap_764
timestamp 1662145021
transform 1 0 44660 0 1 114840
box 0 0 3190 3190
use unit_cap  unit_cap_765
timestamp 1662145021
transform 1 0 44660 0 1 118030
box 0 0 3190 3190
use unit_cap  unit_cap_766
timestamp 1662145021
transform 1 0 44660 0 1 121220
box 0 0 3190 3190
use unit_cap  unit_cap_767
timestamp 1662145021
transform 1 0 44660 0 1 124410
box 0 0 3190 3190
use unit_cap  unit_cap_768
timestamp 1662145021
transform 1 0 44660 0 1 127600
box 0 0 3190 3190
use unit_cap  unit_cap_769
timestamp 1662145021
transform 1 0 44660 0 1 130790
box 0 0 3190 3190
use unit_cap  unit_cap_770
timestamp 1662145021
transform 1 0 44660 0 1 133980
box 0 0 3190 3190
use unit_cap  unit_cap_771
timestamp 1662145021
transform 1 0 44660 0 1 137170
box 0 0 3190 3190
use unit_cap  unit_cap_772
timestamp 1662145021
transform 1 0 44660 0 1 140360
box 0 0 3190 3190
use unit_cap  unit_cap_773
timestamp 1662145021
transform 1 0 44660 0 1 143550
box 0 0 3190 3190
use unit_cap  unit_cap_774
timestamp 1662145021
transform 1 0 44660 0 1 146740
box 0 0 3190 3190
use unit_cap  unit_cap_775
timestamp 1662145021
transform 1 0 44660 0 1 149930
box 0 0 3190 3190
use unit_cap  unit_cap_776
timestamp 1662145021
transform 1 0 44660 0 1 153120
box 0 0 3190 3190
use unit_cap  unit_cap_777
timestamp 1662145021
transform 1 0 44660 0 1 156310
box 0 0 3190 3190
use unit_cap  unit_cap_778
timestamp 1662145021
transform 1 0 44660 0 1 159500
box 0 0 3190 3190
use unit_cap  unit_cap_779
timestamp 1662145021
transform 1 0 44660 0 1 162690
box 0 0 3190 3190
use unit_cap  unit_cap_780
timestamp 1662145021
transform 1 0 47850 0 1 0
box 0 0 3190 3190
use unit_cap  unit_cap_781
timestamp 1662145021
transform 1 0 47850 0 1 3190
box 0 0 3190 3190
use unit_cap  unit_cap_782
timestamp 1662145021
transform 1 0 47850 0 1 6380
box 0 0 3190 3190
use unit_cap  unit_cap_783
timestamp 1662145021
transform 1 0 47850 0 1 9570
box 0 0 3190 3190
use unit_cap  unit_cap_784
timestamp 1662145021
transform 1 0 47850 0 1 12760
box 0 0 3190 3190
use unit_cap  unit_cap_785
timestamp 1662145021
transform 1 0 47850 0 1 15950
box 0 0 3190 3190
use unit_cap  unit_cap_786
timestamp 1662145021
transform 1 0 47850 0 1 19140
box 0 0 3190 3190
use unit_cap  unit_cap_787
timestamp 1662145021
transform 1 0 47850 0 1 22330
box 0 0 3190 3190
use unit_cap  unit_cap_788
timestamp 1662145021
transform 1 0 47850 0 1 25520
box 0 0 3190 3190
use unit_cap  unit_cap_789
timestamp 1662145021
transform 1 0 47850 0 1 28710
box 0 0 3190 3190
use unit_cap  unit_cap_790
timestamp 1662145021
transform 1 0 47850 0 1 31900
box 0 0 3190 3190
use unit_cap  unit_cap_791
timestamp 1662145021
transform 1 0 47850 0 1 35090
box 0 0 3190 3190
use unit_cap  unit_cap_792
timestamp 1662145021
transform 1 0 47850 0 1 38280
box 0 0 3190 3190
use unit_cap  unit_cap_793
timestamp 1662145021
transform 1 0 47850 0 1 41470
box 0 0 3190 3190
use unit_cap  unit_cap_794
timestamp 1662145021
transform 1 0 47850 0 1 44660
box 0 0 3190 3190
use unit_cap  unit_cap_795
timestamp 1662145021
transform 1 0 47850 0 1 47850
box 0 0 3190 3190
use unit_cap  unit_cap_796
timestamp 1662145021
transform 1 0 47850 0 1 51040
box 0 0 3190 3190
use unit_cap  unit_cap_797
timestamp 1662145021
transform 1 0 47850 0 1 54230
box 0 0 3190 3190
use unit_cap  unit_cap_798
timestamp 1662145021
transform 1 0 47850 0 1 57420
box 0 0 3190 3190
use unit_cap  unit_cap_799
timestamp 1662145021
transform 1 0 47850 0 1 60610
box 0 0 3190 3190
use unit_cap  unit_cap_800
timestamp 1662145021
transform 1 0 47850 0 1 63800
box 0 0 3190 3190
use unit_cap  unit_cap_801
timestamp 1662145021
transform 1 0 47850 0 1 66990
box 0 0 3190 3190
use unit_cap  unit_cap_802
timestamp 1662145021
transform 1 0 47850 0 1 70180
box 0 0 3190 3190
use unit_cap  unit_cap_803
timestamp 1662145021
transform 1 0 47850 0 1 73370
box 0 0 3190 3190
use unit_cap  unit_cap_804
timestamp 1662145021
transform 1 0 47850 0 1 76560
box 0 0 3190 3190
use unit_cap  unit_cap_805
timestamp 1662145021
transform 1 0 47850 0 1 79750
box 0 0 3190 3190
use unit_cap  unit_cap_806
timestamp 1662145021
transform 1 0 47850 0 1 82940
box 0 0 3190 3190
use unit_cap  unit_cap_807
timestamp 1662145021
transform 1 0 47850 0 1 86130
box 0 0 3190 3190
use unit_cap  unit_cap_808
timestamp 1662145021
transform 1 0 47850 0 1 89320
box 0 0 3190 3190
use unit_cap  unit_cap_809
timestamp 1662145021
transform 1 0 47850 0 1 92510
box 0 0 3190 3190
use unit_cap  unit_cap_810
timestamp 1662145021
transform 1 0 47850 0 1 95700
box 0 0 3190 3190
use unit_cap  unit_cap_811
timestamp 1662145021
transform 1 0 47850 0 1 98890
box 0 0 3190 3190
use unit_cap  unit_cap_812
timestamp 1662145021
transform 1 0 47850 0 1 102080
box 0 0 3190 3190
use unit_cap  unit_cap_813
timestamp 1662145021
transform 1 0 47850 0 1 105270
box 0 0 3190 3190
use unit_cap  unit_cap_814
timestamp 1662145021
transform 1 0 47850 0 1 108460
box 0 0 3190 3190
use unit_cap  unit_cap_815
timestamp 1662145021
transform 1 0 47850 0 1 111650
box 0 0 3190 3190
use unit_cap  unit_cap_816
timestamp 1662145021
transform 1 0 47850 0 1 114840
box 0 0 3190 3190
use unit_cap  unit_cap_817
timestamp 1662145021
transform 1 0 47850 0 1 118030
box 0 0 3190 3190
use unit_cap  unit_cap_818
timestamp 1662145021
transform 1 0 47850 0 1 121220
box 0 0 3190 3190
use unit_cap  unit_cap_819
timestamp 1662145021
transform 1 0 47850 0 1 124410
box 0 0 3190 3190
use unit_cap  unit_cap_820
timestamp 1662145021
transform 1 0 47850 0 1 127600
box 0 0 3190 3190
use unit_cap  unit_cap_821
timestamp 1662145021
transform 1 0 47850 0 1 130790
box 0 0 3190 3190
use unit_cap  unit_cap_822
timestamp 1662145021
transform 1 0 47850 0 1 133980
box 0 0 3190 3190
use unit_cap  unit_cap_823
timestamp 1662145021
transform 1 0 47850 0 1 137170
box 0 0 3190 3190
use unit_cap  unit_cap_824
timestamp 1662145021
transform 1 0 47850 0 1 140360
box 0 0 3190 3190
use unit_cap  unit_cap_825
timestamp 1662145021
transform 1 0 47850 0 1 143550
box 0 0 3190 3190
use unit_cap  unit_cap_826
timestamp 1662145021
transform 1 0 47850 0 1 146740
box 0 0 3190 3190
use unit_cap  unit_cap_827
timestamp 1662145021
transform 1 0 47850 0 1 149930
box 0 0 3190 3190
use unit_cap  unit_cap_828
timestamp 1662145021
transform 1 0 47850 0 1 153120
box 0 0 3190 3190
use unit_cap  unit_cap_829
timestamp 1662145021
transform 1 0 47850 0 1 156310
box 0 0 3190 3190
use unit_cap  unit_cap_830
timestamp 1662145021
transform 1 0 47850 0 1 159500
box 0 0 3190 3190
use unit_cap  unit_cap_831
timestamp 1662145021
transform 1 0 47850 0 1 162690
box 0 0 3190 3190
use unit_cap  unit_cap_832
timestamp 1662145021
transform 1 0 51040 0 1 0
box 0 0 3190 3190
use unit_cap  unit_cap_833
timestamp 1662145021
transform 1 0 51040 0 1 3190
box 0 0 3190 3190
use unit_cap  unit_cap_834
timestamp 1662145021
transform 1 0 51040 0 1 6380
box 0 0 3190 3190
use unit_cap  unit_cap_835
timestamp 1662145021
transform 1 0 51040 0 1 9570
box 0 0 3190 3190
use unit_cap  unit_cap_836
timestamp 1662145021
transform 1 0 51040 0 1 12760
box 0 0 3190 3190
use unit_cap  unit_cap_837
timestamp 1662145021
transform 1 0 51040 0 1 15950
box 0 0 3190 3190
use unit_cap  unit_cap_838
timestamp 1662145021
transform 1 0 51040 0 1 19140
box 0 0 3190 3190
use unit_cap  unit_cap_839
timestamp 1662145021
transform 1 0 51040 0 1 22330
box 0 0 3190 3190
use unit_cap  unit_cap_840
timestamp 1662145021
transform 1 0 51040 0 1 25520
box 0 0 3190 3190
use unit_cap  unit_cap_841
timestamp 1662145021
transform 1 0 51040 0 1 28710
box 0 0 3190 3190
use unit_cap  unit_cap_842
timestamp 1662145021
transform 1 0 51040 0 1 31900
box 0 0 3190 3190
use unit_cap  unit_cap_843
timestamp 1662145021
transform 1 0 51040 0 1 35090
box 0 0 3190 3190
use unit_cap  unit_cap_844
timestamp 1662145021
transform 1 0 51040 0 1 38280
box 0 0 3190 3190
use unit_cap  unit_cap_845
timestamp 1662145021
transform 1 0 51040 0 1 41470
box 0 0 3190 3190
use unit_cap  unit_cap_846
timestamp 1662145021
transform 1 0 51040 0 1 44660
box 0 0 3190 3190
use unit_cap  unit_cap_847
timestamp 1662145021
transform 1 0 51040 0 1 47850
box 0 0 3190 3190
use unit_cap  unit_cap_848
timestamp 1662145021
transform 1 0 51040 0 1 51040
box 0 0 3190 3190
use unit_cap  unit_cap_849
timestamp 1662145021
transform 1 0 51040 0 1 54230
box 0 0 3190 3190
use unit_cap  unit_cap_850
timestamp 1662145021
transform 1 0 51040 0 1 57420
box 0 0 3190 3190
use unit_cap  unit_cap_851
timestamp 1662145021
transform 1 0 51040 0 1 60610
box 0 0 3190 3190
use unit_cap  unit_cap_852
timestamp 1662145021
transform 1 0 51040 0 1 63800
box 0 0 3190 3190
use unit_cap  unit_cap_853
timestamp 1662145021
transform 1 0 51040 0 1 66990
box 0 0 3190 3190
use unit_cap  unit_cap_854
timestamp 1662145021
transform 1 0 51040 0 1 70180
box 0 0 3190 3190
use unit_cap  unit_cap_855
timestamp 1662145021
transform 1 0 51040 0 1 73370
box 0 0 3190 3190
use unit_cap  unit_cap_856
timestamp 1662145021
transform 1 0 51040 0 1 76560
box 0 0 3190 3190
use unit_cap  unit_cap_857
timestamp 1662145021
transform 1 0 51040 0 1 79750
box 0 0 3190 3190
use unit_cap  unit_cap_858
timestamp 1662145021
transform 1 0 51040 0 1 82940
box 0 0 3190 3190
use unit_cap  unit_cap_859
timestamp 1662145021
transform 1 0 51040 0 1 86130
box 0 0 3190 3190
use unit_cap  unit_cap_860
timestamp 1662145021
transform 1 0 51040 0 1 89320
box 0 0 3190 3190
use unit_cap  unit_cap_861
timestamp 1662145021
transform 1 0 51040 0 1 92510
box 0 0 3190 3190
use unit_cap  unit_cap_862
timestamp 1662145021
transform 1 0 51040 0 1 95700
box 0 0 3190 3190
use unit_cap  unit_cap_863
timestamp 1662145021
transform 1 0 51040 0 1 98890
box 0 0 3190 3190
use unit_cap  unit_cap_864
timestamp 1662145021
transform 1 0 51040 0 1 102080
box 0 0 3190 3190
use unit_cap  unit_cap_865
timestamp 1662145021
transform 1 0 51040 0 1 105270
box 0 0 3190 3190
use unit_cap  unit_cap_866
timestamp 1662145021
transform 1 0 51040 0 1 108460
box 0 0 3190 3190
use unit_cap  unit_cap_867
timestamp 1662145021
transform 1 0 51040 0 1 111650
box 0 0 3190 3190
use unit_cap  unit_cap_868
timestamp 1662145021
transform 1 0 51040 0 1 114840
box 0 0 3190 3190
use unit_cap  unit_cap_869
timestamp 1662145021
transform 1 0 51040 0 1 118030
box 0 0 3190 3190
use unit_cap  unit_cap_870
timestamp 1662145021
transform 1 0 51040 0 1 121220
box 0 0 3190 3190
use unit_cap  unit_cap_871
timestamp 1662145021
transform 1 0 51040 0 1 124410
box 0 0 3190 3190
use unit_cap  unit_cap_872
timestamp 1662145021
transform 1 0 51040 0 1 127600
box 0 0 3190 3190
use unit_cap  unit_cap_873
timestamp 1662145021
transform 1 0 51040 0 1 130790
box 0 0 3190 3190
use unit_cap  unit_cap_874
timestamp 1662145021
transform 1 0 51040 0 1 133980
box 0 0 3190 3190
use unit_cap  unit_cap_875
timestamp 1662145021
transform 1 0 51040 0 1 137170
box 0 0 3190 3190
use unit_cap  unit_cap_876
timestamp 1662145021
transform 1 0 51040 0 1 140360
box 0 0 3190 3190
use unit_cap  unit_cap_877
timestamp 1662145021
transform 1 0 51040 0 1 143550
box 0 0 3190 3190
use unit_cap  unit_cap_878
timestamp 1662145021
transform 1 0 51040 0 1 146740
box 0 0 3190 3190
use unit_cap  unit_cap_879
timestamp 1662145021
transform 1 0 51040 0 1 149930
box 0 0 3190 3190
use unit_cap  unit_cap_880
timestamp 1662145021
transform 1 0 51040 0 1 153120
box 0 0 3190 3190
use unit_cap  unit_cap_881
timestamp 1662145021
transform 1 0 51040 0 1 156310
box 0 0 3190 3190
use unit_cap  unit_cap_882
timestamp 1662145021
transform 1 0 51040 0 1 159500
box 0 0 3190 3190
use unit_cap  unit_cap_883
timestamp 1662145021
transform 1 0 51040 0 1 162690
box 0 0 3190 3190
use unit_cap  unit_cap_884
timestamp 1662145021
transform 1 0 54230 0 1 0
box 0 0 3190 3190
use unit_cap  unit_cap_885
timestamp 1662145021
transform 1 0 54230 0 1 3190
box 0 0 3190 3190
use unit_cap  unit_cap_886
timestamp 1662145021
transform 1 0 54230 0 1 6380
box 0 0 3190 3190
use unit_cap  unit_cap_887
timestamp 1662145021
transform 1 0 54230 0 1 9570
box 0 0 3190 3190
use unit_cap  unit_cap_888
timestamp 1662145021
transform 1 0 54230 0 1 12760
box 0 0 3190 3190
use unit_cap  unit_cap_889
timestamp 1662145021
transform 1 0 54230 0 1 15950
box 0 0 3190 3190
use unit_cap  unit_cap_890
timestamp 1662145021
transform 1 0 54230 0 1 19140
box 0 0 3190 3190
use unit_cap  unit_cap_891
timestamp 1662145021
transform 1 0 54230 0 1 22330
box 0 0 3190 3190
use unit_cap  unit_cap_892
timestamp 1662145021
transform 1 0 54230 0 1 25520
box 0 0 3190 3190
use unit_cap  unit_cap_893
timestamp 1662145021
transform 1 0 54230 0 1 28710
box 0 0 3190 3190
use unit_cap  unit_cap_894
timestamp 1662145021
transform 1 0 54230 0 1 31900
box 0 0 3190 3190
use unit_cap  unit_cap_895
timestamp 1662145021
transform 1 0 54230 0 1 35090
box 0 0 3190 3190
use unit_cap  unit_cap_896
timestamp 1662145021
transform 1 0 54230 0 1 38280
box 0 0 3190 3190
use unit_cap  unit_cap_897
timestamp 1662145021
transform 1 0 54230 0 1 41470
box 0 0 3190 3190
use unit_cap  unit_cap_898
timestamp 1662145021
transform 1 0 54230 0 1 44660
box 0 0 3190 3190
use unit_cap  unit_cap_899
timestamp 1662145021
transform 1 0 54230 0 1 47850
box 0 0 3190 3190
use unit_cap  unit_cap_900
timestamp 1662145021
transform 1 0 54230 0 1 51040
box 0 0 3190 3190
use unit_cap  unit_cap_901
timestamp 1662145021
transform 1 0 54230 0 1 54230
box 0 0 3190 3190
use unit_cap  unit_cap_902
timestamp 1662145021
transform 1 0 54230 0 1 57420
box 0 0 3190 3190
use unit_cap  unit_cap_903
timestamp 1662145021
transform 1 0 54230 0 1 60610
box 0 0 3190 3190
use unit_cap  unit_cap_904
timestamp 1662145021
transform 1 0 54230 0 1 63800
box 0 0 3190 3190
use unit_cap  unit_cap_905
timestamp 1662145021
transform 1 0 54230 0 1 66990
box 0 0 3190 3190
use unit_cap  unit_cap_906
timestamp 1662145021
transform 1 0 54230 0 1 70180
box 0 0 3190 3190
use unit_cap  unit_cap_907
timestamp 1662145021
transform 1 0 54230 0 1 73370
box 0 0 3190 3190
use unit_cap  unit_cap_908
timestamp 1662145021
transform 1 0 54230 0 1 76560
box 0 0 3190 3190
use unit_cap  unit_cap_909
timestamp 1662145021
transform 1 0 54230 0 1 79750
box 0 0 3190 3190
use unit_cap  unit_cap_910
timestamp 1662145021
transform 1 0 54230 0 1 82940
box 0 0 3190 3190
use unit_cap  unit_cap_911
timestamp 1662145021
transform 1 0 54230 0 1 86130
box 0 0 3190 3190
use unit_cap  unit_cap_912
timestamp 1662145021
transform 1 0 54230 0 1 89320
box 0 0 3190 3190
use unit_cap  unit_cap_913
timestamp 1662145021
transform 1 0 54230 0 1 92510
box 0 0 3190 3190
use unit_cap  unit_cap_914
timestamp 1662145021
transform 1 0 54230 0 1 95700
box 0 0 3190 3190
use unit_cap  unit_cap_915
timestamp 1662145021
transform 1 0 54230 0 1 98890
box 0 0 3190 3190
use unit_cap  unit_cap_916
timestamp 1662145021
transform 1 0 54230 0 1 102080
box 0 0 3190 3190
use unit_cap  unit_cap_917
timestamp 1662145021
transform 1 0 54230 0 1 105270
box 0 0 3190 3190
use unit_cap  unit_cap_918
timestamp 1662145021
transform 1 0 54230 0 1 108460
box 0 0 3190 3190
use unit_cap  unit_cap_919
timestamp 1662145021
transform 1 0 54230 0 1 111650
box 0 0 3190 3190
use unit_cap  unit_cap_920
timestamp 1662145021
transform 1 0 54230 0 1 114840
box 0 0 3190 3190
use unit_cap  unit_cap_921
timestamp 1662145021
transform 1 0 54230 0 1 118030
box 0 0 3190 3190
use unit_cap  unit_cap_922
timestamp 1662145021
transform 1 0 54230 0 1 121220
box 0 0 3190 3190
use unit_cap  unit_cap_923
timestamp 1662145021
transform 1 0 54230 0 1 124410
box 0 0 3190 3190
use unit_cap  unit_cap_924
timestamp 1662145021
transform 1 0 54230 0 1 127600
box 0 0 3190 3190
use unit_cap  unit_cap_925
timestamp 1662145021
transform 1 0 54230 0 1 130790
box 0 0 3190 3190
use unit_cap  unit_cap_926
timestamp 1662145021
transform 1 0 54230 0 1 133980
box 0 0 3190 3190
use unit_cap  unit_cap_927
timestamp 1662145021
transform 1 0 54230 0 1 137170
box 0 0 3190 3190
use unit_cap  unit_cap_928
timestamp 1662145021
transform 1 0 54230 0 1 140360
box 0 0 3190 3190
use unit_cap  unit_cap_929
timestamp 1662145021
transform 1 0 54230 0 1 143550
box 0 0 3190 3190
use unit_cap  unit_cap_930
timestamp 1662145021
transform 1 0 54230 0 1 146740
box 0 0 3190 3190
use unit_cap  unit_cap_931
timestamp 1662145021
transform 1 0 54230 0 1 149930
box 0 0 3190 3190
use unit_cap  unit_cap_932
timestamp 1662145021
transform 1 0 54230 0 1 153120
box 0 0 3190 3190
use unit_cap  unit_cap_933
timestamp 1662145021
transform 1 0 54230 0 1 156310
box 0 0 3190 3190
use unit_cap  unit_cap_934
timestamp 1662145021
transform 1 0 54230 0 1 159500
box 0 0 3190 3190
use unit_cap  unit_cap_935
timestamp 1662145021
transform 1 0 54230 0 1 162690
box 0 0 3190 3190
use unit_cap  unit_cap_936
timestamp 1662145021
transform 1 0 57420 0 1 0
box 0 0 3190 3190
use unit_cap  unit_cap_937
timestamp 1662145021
transform 1 0 57420 0 1 3190
box 0 0 3190 3190
use unit_cap  unit_cap_938
timestamp 1662145021
transform 1 0 57420 0 1 6380
box 0 0 3190 3190
use unit_cap  unit_cap_939
timestamp 1662145021
transform 1 0 57420 0 1 9570
box 0 0 3190 3190
use unit_cap  unit_cap_940
timestamp 1662145021
transform 1 0 57420 0 1 12760
box 0 0 3190 3190
use unit_cap  unit_cap_941
timestamp 1662145021
transform 1 0 57420 0 1 15950
box 0 0 3190 3190
use unit_cap  unit_cap_942
timestamp 1662145021
transform 1 0 57420 0 1 19140
box 0 0 3190 3190
use unit_cap  unit_cap_943
timestamp 1662145021
transform 1 0 57420 0 1 22330
box 0 0 3190 3190
use unit_cap  unit_cap_944
timestamp 1662145021
transform 1 0 57420 0 1 25520
box 0 0 3190 3190
use unit_cap  unit_cap_945
timestamp 1662145021
transform 1 0 57420 0 1 28710
box 0 0 3190 3190
use unit_cap  unit_cap_946
timestamp 1662145021
transform 1 0 57420 0 1 31900
box 0 0 3190 3190
use unit_cap  unit_cap_947
timestamp 1662145021
transform 1 0 57420 0 1 35090
box 0 0 3190 3190
use unit_cap  unit_cap_948
timestamp 1662145021
transform 1 0 57420 0 1 38280
box 0 0 3190 3190
use unit_cap  unit_cap_949
timestamp 1662145021
transform 1 0 57420 0 1 41470
box 0 0 3190 3190
use unit_cap  unit_cap_950
timestamp 1662145021
transform 1 0 57420 0 1 44660
box 0 0 3190 3190
use unit_cap  unit_cap_951
timestamp 1662145021
transform 1 0 57420 0 1 47850
box 0 0 3190 3190
use unit_cap  unit_cap_952
timestamp 1662145021
transform 1 0 57420 0 1 51040
box 0 0 3190 3190
use unit_cap  unit_cap_953
timestamp 1662145021
transform 1 0 57420 0 1 54230
box 0 0 3190 3190
use unit_cap  unit_cap_954
timestamp 1662145021
transform 1 0 57420 0 1 57420
box 0 0 3190 3190
use unit_cap  unit_cap_955
timestamp 1662145021
transform 1 0 57420 0 1 60610
box 0 0 3190 3190
use unit_cap  unit_cap_956
timestamp 1662145021
transform 1 0 57420 0 1 63800
box 0 0 3190 3190
use unit_cap  unit_cap_957
timestamp 1662145021
transform 1 0 57420 0 1 66990
box 0 0 3190 3190
use unit_cap  unit_cap_958
timestamp 1662145021
transform 1 0 57420 0 1 70180
box 0 0 3190 3190
use unit_cap  unit_cap_959
timestamp 1662145021
transform 1 0 57420 0 1 73370
box 0 0 3190 3190
use unit_cap  unit_cap_960
timestamp 1662145021
transform 1 0 57420 0 1 76560
box 0 0 3190 3190
use unit_cap  unit_cap_961
timestamp 1662145021
transform 1 0 57420 0 1 79750
box 0 0 3190 3190
use unit_cap  unit_cap_962
timestamp 1662145021
transform 1 0 57420 0 1 82940
box 0 0 3190 3190
use unit_cap  unit_cap_963
timestamp 1662145021
transform 1 0 57420 0 1 86130
box 0 0 3190 3190
use unit_cap  unit_cap_964
timestamp 1662145021
transform 1 0 57420 0 1 89320
box 0 0 3190 3190
use unit_cap  unit_cap_965
timestamp 1662145021
transform 1 0 57420 0 1 92510
box 0 0 3190 3190
use unit_cap  unit_cap_966
timestamp 1662145021
transform 1 0 57420 0 1 95700
box 0 0 3190 3190
use unit_cap  unit_cap_967
timestamp 1662145021
transform 1 0 57420 0 1 98890
box 0 0 3190 3190
use unit_cap  unit_cap_968
timestamp 1662145021
transform 1 0 57420 0 1 102080
box 0 0 3190 3190
use unit_cap  unit_cap_969
timestamp 1662145021
transform 1 0 57420 0 1 105270
box 0 0 3190 3190
use unit_cap  unit_cap_970
timestamp 1662145021
transform 1 0 57420 0 1 108460
box 0 0 3190 3190
use unit_cap  unit_cap_971
timestamp 1662145021
transform 1 0 57420 0 1 111650
box 0 0 3190 3190
use unit_cap  unit_cap_972
timestamp 1662145021
transform 1 0 57420 0 1 114840
box 0 0 3190 3190
use unit_cap  unit_cap_973
timestamp 1662145021
transform 1 0 57420 0 1 118030
box 0 0 3190 3190
use unit_cap  unit_cap_974
timestamp 1662145021
transform 1 0 57420 0 1 121220
box 0 0 3190 3190
use unit_cap  unit_cap_975
timestamp 1662145021
transform 1 0 57420 0 1 124410
box 0 0 3190 3190
use unit_cap  unit_cap_976
timestamp 1662145021
transform 1 0 57420 0 1 127600
box 0 0 3190 3190
use unit_cap  unit_cap_977
timestamp 1662145021
transform 1 0 57420 0 1 130790
box 0 0 3190 3190
use unit_cap  unit_cap_978
timestamp 1662145021
transform 1 0 57420 0 1 133980
box 0 0 3190 3190
use unit_cap  unit_cap_979
timestamp 1662145021
transform 1 0 57420 0 1 137170
box 0 0 3190 3190
use unit_cap  unit_cap_980
timestamp 1662145021
transform 1 0 57420 0 1 140360
box 0 0 3190 3190
use unit_cap  unit_cap_981
timestamp 1662145021
transform 1 0 57420 0 1 143550
box 0 0 3190 3190
use unit_cap  unit_cap_982
timestamp 1662145021
transform 1 0 57420 0 1 146740
box 0 0 3190 3190
use unit_cap  unit_cap_983
timestamp 1662145021
transform 1 0 57420 0 1 149930
box 0 0 3190 3190
use unit_cap  unit_cap_984
timestamp 1662145021
transform 1 0 57420 0 1 153120
box 0 0 3190 3190
use unit_cap  unit_cap_985
timestamp 1662145021
transform 1 0 57420 0 1 156310
box 0 0 3190 3190
use unit_cap  unit_cap_986
timestamp 1662145021
transform 1 0 57420 0 1 159500
box 0 0 3190 3190
use unit_cap  unit_cap_987
timestamp 1662145021
transform 1 0 57420 0 1 162690
box 0 0 3190 3190
use unit_cap  unit_cap_988
timestamp 1662145021
transform 1 0 60610 0 1 0
box 0 0 3190 3190
use unit_cap  unit_cap_989
timestamp 1662145021
transform 1 0 60610 0 1 3190
box 0 0 3190 3190
use unit_cap  unit_cap_990
timestamp 1662145021
transform 1 0 60610 0 1 6380
box 0 0 3190 3190
use unit_cap  unit_cap_991
timestamp 1662145021
transform 1 0 60610 0 1 9570
box 0 0 3190 3190
use unit_cap  unit_cap_992
timestamp 1662145021
transform 1 0 60610 0 1 12760
box 0 0 3190 3190
use unit_cap  unit_cap_993
timestamp 1662145021
transform 1 0 60610 0 1 15950
box 0 0 3190 3190
use unit_cap  unit_cap_994
timestamp 1662145021
transform 1 0 60610 0 1 19140
box 0 0 3190 3190
use unit_cap  unit_cap_995
timestamp 1662145021
transform 1 0 60610 0 1 22330
box 0 0 3190 3190
use unit_cap  unit_cap_996
timestamp 1662145021
transform 1 0 60610 0 1 25520
box 0 0 3190 3190
use unit_cap  unit_cap_997
timestamp 1662145021
transform 1 0 60610 0 1 28710
box 0 0 3190 3190
use unit_cap  unit_cap_998
timestamp 1662145021
transform 1 0 60610 0 1 31900
box 0 0 3190 3190
use unit_cap  unit_cap_999
timestamp 1662145021
transform 1 0 60610 0 1 35090
box 0 0 3190 3190
use unit_cap  unit_cap_1000
timestamp 1662145021
transform 1 0 60610 0 1 38280
box 0 0 3190 3190
use unit_cap  unit_cap_1001
timestamp 1662145021
transform 1 0 60610 0 1 41470
box 0 0 3190 3190
use unit_cap  unit_cap_1002
timestamp 1662145021
transform 1 0 60610 0 1 44660
box 0 0 3190 3190
use unit_cap  unit_cap_1003
timestamp 1662145021
transform 1 0 60610 0 1 47850
box 0 0 3190 3190
use unit_cap  unit_cap_1004
timestamp 1662145021
transform 1 0 60610 0 1 51040
box 0 0 3190 3190
use unit_cap  unit_cap_1005
timestamp 1662145021
transform 1 0 60610 0 1 54230
box 0 0 3190 3190
use unit_cap  unit_cap_1006
timestamp 1662145021
transform 1 0 60610 0 1 57420
box 0 0 3190 3190
use unit_cap  unit_cap_1007
timestamp 1662145021
transform 1 0 60610 0 1 60610
box 0 0 3190 3190
use unit_cap  unit_cap_1008
timestamp 1662145021
transform 1 0 60610 0 1 63800
box 0 0 3190 3190
use unit_cap  unit_cap_1009
timestamp 1662145021
transform 1 0 60610 0 1 66990
box 0 0 3190 3190
use unit_cap  unit_cap_1010
timestamp 1662145021
transform 1 0 60610 0 1 70180
box 0 0 3190 3190
use unit_cap  unit_cap_1011
timestamp 1662145021
transform 1 0 60610 0 1 73370
box 0 0 3190 3190
use unit_cap  unit_cap_1012
timestamp 1662145021
transform 1 0 60610 0 1 76560
box 0 0 3190 3190
use unit_cap  unit_cap_1013
timestamp 1662145021
transform 1 0 60610 0 1 79750
box 0 0 3190 3190
use unit_cap  unit_cap_1014
timestamp 1662145021
transform 1 0 60610 0 1 82940
box 0 0 3190 3190
use unit_cap  unit_cap_1015
timestamp 1662145021
transform 1 0 60610 0 1 86130
box 0 0 3190 3190
use unit_cap  unit_cap_1016
timestamp 1662145021
transform 1 0 60610 0 1 89320
box 0 0 3190 3190
use unit_cap  unit_cap_1017
timestamp 1662145021
transform 1 0 60610 0 1 92510
box 0 0 3190 3190
use unit_cap  unit_cap_1018
timestamp 1662145021
transform 1 0 60610 0 1 95700
box 0 0 3190 3190
use unit_cap  unit_cap_1019
timestamp 1662145021
transform 1 0 60610 0 1 98890
box 0 0 3190 3190
use unit_cap  unit_cap_1020
timestamp 1662145021
transform 1 0 60610 0 1 102080
box 0 0 3190 3190
use unit_cap  unit_cap_1021
timestamp 1662145021
transform 1 0 60610 0 1 105270
box 0 0 3190 3190
use unit_cap  unit_cap_1022
timestamp 1662145021
transform 1 0 60610 0 1 108460
box 0 0 3190 3190
use unit_cap  unit_cap_1023
timestamp 1662145021
transform 1 0 60610 0 1 111650
box 0 0 3190 3190
use unit_cap  unit_cap_1024
timestamp 1662145021
transform 1 0 60610 0 1 114840
box 0 0 3190 3190
use unit_cap  unit_cap_1025
timestamp 1662145021
transform 1 0 60610 0 1 118030
box 0 0 3190 3190
use unit_cap  unit_cap_1026
timestamp 1662145021
transform 1 0 60610 0 1 121220
box 0 0 3190 3190
use unit_cap  unit_cap_1027
timestamp 1662145021
transform 1 0 60610 0 1 124410
box 0 0 3190 3190
use unit_cap  unit_cap_1028
timestamp 1662145021
transform 1 0 60610 0 1 127600
box 0 0 3190 3190
use unit_cap  unit_cap_1029
timestamp 1662145021
transform 1 0 60610 0 1 130790
box 0 0 3190 3190
use unit_cap  unit_cap_1030
timestamp 1662145021
transform 1 0 60610 0 1 133980
box 0 0 3190 3190
use unit_cap  unit_cap_1031
timestamp 1662145021
transform 1 0 60610 0 1 137170
box 0 0 3190 3190
use unit_cap  unit_cap_1032
timestamp 1662145021
transform 1 0 60610 0 1 140360
box 0 0 3190 3190
use unit_cap  unit_cap_1033
timestamp 1662145021
transform 1 0 60610 0 1 143550
box 0 0 3190 3190
use unit_cap  unit_cap_1034
timestamp 1662145021
transform 1 0 60610 0 1 146740
box 0 0 3190 3190
use unit_cap  unit_cap_1035
timestamp 1662145021
transform 1 0 60610 0 1 149930
box 0 0 3190 3190
use unit_cap  unit_cap_1036
timestamp 1662145021
transform 1 0 60610 0 1 153120
box 0 0 3190 3190
use unit_cap  unit_cap_1037
timestamp 1662145021
transform 1 0 60610 0 1 156310
box 0 0 3190 3190
use unit_cap  unit_cap_1038
timestamp 1662145021
transform 1 0 60610 0 1 159500
box 0 0 3190 3190
use unit_cap  unit_cap_1039
timestamp 1662145021
transform 1 0 60610 0 1 162690
box 0 0 3190 3190
use unit_cap  unit_cap_1040
timestamp 1662145021
transform 1 0 63800 0 1 0
box 0 0 3190 3190
use unit_cap  unit_cap_1041
timestamp 1662145021
transform 1 0 63800 0 1 3190
box 0 0 3190 3190
use unit_cap  unit_cap_1042
timestamp 1662145021
transform 1 0 63800 0 1 6380
box 0 0 3190 3190
use unit_cap  unit_cap_1043
timestamp 1662145021
transform 1 0 63800 0 1 9570
box 0 0 3190 3190
use unit_cap  unit_cap_1044
timestamp 1662145021
transform 1 0 63800 0 1 12760
box 0 0 3190 3190
use unit_cap  unit_cap_1045
timestamp 1662145021
transform 1 0 63800 0 1 15950
box 0 0 3190 3190
use unit_cap  unit_cap_1046
timestamp 1662145021
transform 1 0 63800 0 1 19140
box 0 0 3190 3190
use unit_cap  unit_cap_1047
timestamp 1662145021
transform 1 0 63800 0 1 22330
box 0 0 3190 3190
use unit_cap  unit_cap_1048
timestamp 1662145021
transform 1 0 63800 0 1 25520
box 0 0 3190 3190
use unit_cap  unit_cap_1049
timestamp 1662145021
transform 1 0 63800 0 1 28710
box 0 0 3190 3190
use unit_cap  unit_cap_1050
timestamp 1662145021
transform 1 0 63800 0 1 31900
box 0 0 3190 3190
use unit_cap  unit_cap_1051
timestamp 1662145021
transform 1 0 63800 0 1 35090
box 0 0 3190 3190
use unit_cap  unit_cap_1052
timestamp 1662145021
transform 1 0 63800 0 1 38280
box 0 0 3190 3190
use unit_cap  unit_cap_1053
timestamp 1662145021
transform 1 0 63800 0 1 41470
box 0 0 3190 3190
use unit_cap  unit_cap_1054
timestamp 1662145021
transform 1 0 63800 0 1 44660
box 0 0 3190 3190
use unit_cap  unit_cap_1055
timestamp 1662145021
transform 1 0 63800 0 1 47850
box 0 0 3190 3190
use unit_cap  unit_cap_1056
timestamp 1662145021
transform 1 0 63800 0 1 51040
box 0 0 3190 3190
use unit_cap  unit_cap_1057
timestamp 1662145021
transform 1 0 63800 0 1 54230
box 0 0 3190 3190
use unit_cap  unit_cap_1058
timestamp 1662145021
transform 1 0 63800 0 1 57420
box 0 0 3190 3190
use unit_cap  unit_cap_1059
timestamp 1662145021
transform 1 0 63800 0 1 60610
box 0 0 3190 3190
use unit_cap  unit_cap_1060
timestamp 1662145021
transform 1 0 63800 0 1 63800
box 0 0 3190 3190
use unit_cap  unit_cap_1061
timestamp 1662145021
transform 1 0 63800 0 1 66990
box 0 0 3190 3190
use unit_cap  unit_cap_1062
timestamp 1662145021
transform 1 0 63800 0 1 70180
box 0 0 3190 3190
use unit_cap  unit_cap_1063
timestamp 1662145021
transform 1 0 63800 0 1 73370
box 0 0 3190 3190
use unit_cap  unit_cap_1064
timestamp 1662145021
transform 1 0 63800 0 1 76560
box 0 0 3190 3190
use unit_cap  unit_cap_1065
timestamp 1662145021
transform 1 0 63800 0 1 79750
box 0 0 3190 3190
use unit_cap  unit_cap_1066
timestamp 1662145021
transform 1 0 63800 0 1 82940
box 0 0 3190 3190
use unit_cap  unit_cap_1067
timestamp 1662145021
transform 1 0 63800 0 1 86130
box 0 0 3190 3190
use unit_cap  unit_cap_1068
timestamp 1662145021
transform 1 0 63800 0 1 89320
box 0 0 3190 3190
use unit_cap  unit_cap_1069
timestamp 1662145021
transform 1 0 63800 0 1 92510
box 0 0 3190 3190
use unit_cap  unit_cap_1070
timestamp 1662145021
transform 1 0 63800 0 1 95700
box 0 0 3190 3190
use unit_cap  unit_cap_1071
timestamp 1662145021
transform 1 0 63800 0 1 98890
box 0 0 3190 3190
use unit_cap  unit_cap_1072
timestamp 1662145021
transform 1 0 63800 0 1 102080
box 0 0 3190 3190
use unit_cap  unit_cap_1073
timestamp 1662145021
transform 1 0 63800 0 1 105270
box 0 0 3190 3190
use unit_cap  unit_cap_1074
timestamp 1662145021
transform 1 0 63800 0 1 108460
box 0 0 3190 3190
use unit_cap  unit_cap_1075
timestamp 1662145021
transform 1 0 63800 0 1 111650
box 0 0 3190 3190
use unit_cap  unit_cap_1076
timestamp 1662145021
transform 1 0 63800 0 1 114840
box 0 0 3190 3190
use unit_cap  unit_cap_1077
timestamp 1662145021
transform 1 0 63800 0 1 118030
box 0 0 3190 3190
use unit_cap  unit_cap_1078
timestamp 1662145021
transform 1 0 63800 0 1 121220
box 0 0 3190 3190
use unit_cap  unit_cap_1079
timestamp 1662145021
transform 1 0 63800 0 1 124410
box 0 0 3190 3190
use unit_cap  unit_cap_1080
timestamp 1662145021
transform 1 0 63800 0 1 127600
box 0 0 3190 3190
use unit_cap  unit_cap_1081
timestamp 1662145021
transform 1 0 63800 0 1 130790
box 0 0 3190 3190
use unit_cap  unit_cap_1082
timestamp 1662145021
transform 1 0 63800 0 1 133980
box 0 0 3190 3190
use unit_cap  unit_cap_1083
timestamp 1662145021
transform 1 0 63800 0 1 137170
box 0 0 3190 3190
use unit_cap  unit_cap_1084
timestamp 1662145021
transform 1 0 63800 0 1 140360
box 0 0 3190 3190
use unit_cap  unit_cap_1085
timestamp 1662145021
transform 1 0 63800 0 1 143550
box 0 0 3190 3190
use unit_cap  unit_cap_1086
timestamp 1662145021
transform 1 0 63800 0 1 146740
box 0 0 3190 3190
use unit_cap  unit_cap_1087
timestamp 1662145021
transform 1 0 63800 0 1 149930
box 0 0 3190 3190
use unit_cap  unit_cap_1088
timestamp 1662145021
transform 1 0 63800 0 1 153120
box 0 0 3190 3190
use unit_cap  unit_cap_1089
timestamp 1662145021
transform 1 0 63800 0 1 156310
box 0 0 3190 3190
use unit_cap  unit_cap_1090
timestamp 1662145021
transform 1 0 63800 0 1 159500
box 0 0 3190 3190
use unit_cap  unit_cap_1091
timestamp 1662145021
transform 1 0 63800 0 1 162690
box 0 0 3190 3190
use unit_cap  unit_cap_1092
timestamp 1662145021
transform 1 0 66990 0 1 0
box 0 0 3190 3190
use unit_cap  unit_cap_1093
timestamp 1662145021
transform 1 0 66990 0 1 3190
box 0 0 3190 3190
use unit_cap  unit_cap_1094
timestamp 1662145021
transform 1 0 66990 0 1 6380
box 0 0 3190 3190
use unit_cap  unit_cap_1095
timestamp 1662145021
transform 1 0 66990 0 1 9570
box 0 0 3190 3190
use unit_cap  unit_cap_1096
timestamp 1662145021
transform 1 0 66990 0 1 12760
box 0 0 3190 3190
use unit_cap  unit_cap_1097
timestamp 1662145021
transform 1 0 66990 0 1 15950
box 0 0 3190 3190
use unit_cap  unit_cap_1098
timestamp 1662145021
transform 1 0 66990 0 1 19140
box 0 0 3190 3190
use unit_cap  unit_cap_1099
timestamp 1662145021
transform 1 0 66990 0 1 22330
box 0 0 3190 3190
use unit_cap  unit_cap_1100
timestamp 1662145021
transform 1 0 66990 0 1 25520
box 0 0 3190 3190
use unit_cap  unit_cap_1101
timestamp 1662145021
transform 1 0 66990 0 1 28710
box 0 0 3190 3190
use unit_cap  unit_cap_1102
timestamp 1662145021
transform 1 0 66990 0 1 31900
box 0 0 3190 3190
use unit_cap  unit_cap_1103
timestamp 1662145021
transform 1 0 66990 0 1 35090
box 0 0 3190 3190
use unit_cap  unit_cap_1104
timestamp 1662145021
transform 1 0 66990 0 1 38280
box 0 0 3190 3190
use unit_cap  unit_cap_1105
timestamp 1662145021
transform 1 0 66990 0 1 41470
box 0 0 3190 3190
use unit_cap  unit_cap_1106
timestamp 1662145021
transform 1 0 66990 0 1 44660
box 0 0 3190 3190
use unit_cap  unit_cap_1107
timestamp 1662145021
transform 1 0 66990 0 1 47850
box 0 0 3190 3190
use unit_cap  unit_cap_1108
timestamp 1662145021
transform 1 0 66990 0 1 51040
box 0 0 3190 3190
use unit_cap  unit_cap_1109
timestamp 1662145021
transform 1 0 66990 0 1 54230
box 0 0 3190 3190
use unit_cap  unit_cap_1110
timestamp 1662145021
transform 1 0 66990 0 1 57420
box 0 0 3190 3190
use unit_cap  unit_cap_1111
timestamp 1662145021
transform 1 0 66990 0 1 60610
box 0 0 3190 3190
use unit_cap  unit_cap_1112
timestamp 1662145021
transform 1 0 66990 0 1 63800
box 0 0 3190 3190
use unit_cap  unit_cap_1113
timestamp 1662145021
transform 1 0 66990 0 1 66990
box 0 0 3190 3190
use unit_cap  unit_cap_1114
timestamp 1662145021
transform 1 0 66990 0 1 70180
box 0 0 3190 3190
use unit_cap  unit_cap_1115
timestamp 1662145021
transform 1 0 66990 0 1 73370
box 0 0 3190 3190
use unit_cap  unit_cap_1116
timestamp 1662145021
transform 1 0 66990 0 1 76560
box 0 0 3190 3190
use unit_cap  unit_cap_1117
timestamp 1662145021
transform 1 0 66990 0 1 79750
box 0 0 3190 3190
use unit_cap  unit_cap_1118
timestamp 1662145021
transform 1 0 66990 0 1 82940
box 0 0 3190 3190
use unit_cap  unit_cap_1119
timestamp 1662145021
transform 1 0 66990 0 1 86130
box 0 0 3190 3190
use unit_cap  unit_cap_1120
timestamp 1662145021
transform 1 0 66990 0 1 89320
box 0 0 3190 3190
use unit_cap  unit_cap_1121
timestamp 1662145021
transform 1 0 66990 0 1 92510
box 0 0 3190 3190
use unit_cap  unit_cap_1122
timestamp 1662145021
transform 1 0 66990 0 1 95700
box 0 0 3190 3190
use unit_cap  unit_cap_1123
timestamp 1662145021
transform 1 0 66990 0 1 98890
box 0 0 3190 3190
use unit_cap  unit_cap_1124
timestamp 1662145021
transform 1 0 66990 0 1 102080
box 0 0 3190 3190
use unit_cap  unit_cap_1125
timestamp 1662145021
transform 1 0 66990 0 1 105270
box 0 0 3190 3190
use unit_cap  unit_cap_1126
timestamp 1662145021
transform 1 0 66990 0 1 108460
box 0 0 3190 3190
use unit_cap  unit_cap_1127
timestamp 1662145021
transform 1 0 66990 0 1 111650
box 0 0 3190 3190
use unit_cap  unit_cap_1128
timestamp 1662145021
transform 1 0 66990 0 1 114840
box 0 0 3190 3190
use unit_cap  unit_cap_1129
timestamp 1662145021
transform 1 0 66990 0 1 118030
box 0 0 3190 3190
use unit_cap  unit_cap_1130
timestamp 1662145021
transform 1 0 66990 0 1 121220
box 0 0 3190 3190
use unit_cap  unit_cap_1131
timestamp 1662145021
transform 1 0 66990 0 1 124410
box 0 0 3190 3190
use unit_cap  unit_cap_1132
timestamp 1662145021
transform 1 0 66990 0 1 127600
box 0 0 3190 3190
use unit_cap  unit_cap_1133
timestamp 1662145021
transform 1 0 66990 0 1 130790
box 0 0 3190 3190
use unit_cap  unit_cap_1134
timestamp 1662145021
transform 1 0 66990 0 1 133980
box 0 0 3190 3190
use unit_cap  unit_cap_1135
timestamp 1662145021
transform 1 0 66990 0 1 137170
box 0 0 3190 3190
use unit_cap  unit_cap_1136
timestamp 1662145021
transform 1 0 66990 0 1 140360
box 0 0 3190 3190
use unit_cap  unit_cap_1137
timestamp 1662145021
transform 1 0 66990 0 1 143550
box 0 0 3190 3190
use unit_cap  unit_cap_1138
timestamp 1662145021
transform 1 0 66990 0 1 146740
box 0 0 3190 3190
use unit_cap  unit_cap_1139
timestamp 1662145021
transform 1 0 66990 0 1 149930
box 0 0 3190 3190
use unit_cap  unit_cap_1140
timestamp 1662145021
transform 1 0 66990 0 1 153120
box 0 0 3190 3190
use unit_cap  unit_cap_1141
timestamp 1662145021
transform 1 0 66990 0 1 156310
box 0 0 3190 3190
use unit_cap  unit_cap_1142
timestamp 1662145021
transform 1 0 66990 0 1 159500
box 0 0 3190 3190
use unit_cap  unit_cap_1143
timestamp 1662145021
transform 1 0 66990 0 1 162690
box 0 0 3190 3190
use unit_cap  unit_cap_1144
timestamp 1662145021
transform 1 0 70180 0 1 0
box 0 0 3190 3190
use unit_cap  unit_cap_1145
timestamp 1662145021
transform 1 0 70180 0 1 3190
box 0 0 3190 3190
use unit_cap  unit_cap_1146
timestamp 1662145021
transform 1 0 70180 0 1 6380
box 0 0 3190 3190
use unit_cap  unit_cap_1147
timestamp 1662145021
transform 1 0 70180 0 1 9570
box 0 0 3190 3190
use unit_cap  unit_cap_1148
timestamp 1662145021
transform 1 0 70180 0 1 12760
box 0 0 3190 3190
use unit_cap  unit_cap_1149
timestamp 1662145021
transform 1 0 70180 0 1 15950
box 0 0 3190 3190
use unit_cap  unit_cap_1150
timestamp 1662145021
transform 1 0 70180 0 1 19140
box 0 0 3190 3190
use unit_cap  unit_cap_1151
timestamp 1662145021
transform 1 0 70180 0 1 22330
box 0 0 3190 3190
use unit_cap  unit_cap_1152
timestamp 1662145021
transform 1 0 70180 0 1 25520
box 0 0 3190 3190
use unit_cap  unit_cap_1153
timestamp 1662145021
transform 1 0 70180 0 1 28710
box 0 0 3190 3190
use unit_cap  unit_cap_1154
timestamp 1662145021
transform 1 0 70180 0 1 31900
box 0 0 3190 3190
use unit_cap  unit_cap_1155
timestamp 1662145021
transform 1 0 70180 0 1 35090
box 0 0 3190 3190
use unit_cap  unit_cap_1156
timestamp 1662145021
transform 1 0 70180 0 1 38280
box 0 0 3190 3190
use unit_cap  unit_cap_1157
timestamp 1662145021
transform 1 0 70180 0 1 41470
box 0 0 3190 3190
use unit_cap  unit_cap_1158
timestamp 1662145021
transform 1 0 70180 0 1 44660
box 0 0 3190 3190
use unit_cap  unit_cap_1159
timestamp 1662145021
transform 1 0 70180 0 1 47850
box 0 0 3190 3190
use unit_cap  unit_cap_1160
timestamp 1662145021
transform 1 0 70180 0 1 51040
box 0 0 3190 3190
use unit_cap  unit_cap_1161
timestamp 1662145021
transform 1 0 70180 0 1 54230
box 0 0 3190 3190
use unit_cap  unit_cap_1162
timestamp 1662145021
transform 1 0 70180 0 1 57420
box 0 0 3190 3190
use unit_cap  unit_cap_1163
timestamp 1662145021
transform 1 0 70180 0 1 60610
box 0 0 3190 3190
use unit_cap  unit_cap_1164
timestamp 1662145021
transform 1 0 70180 0 1 63800
box 0 0 3190 3190
use unit_cap  unit_cap_1165
timestamp 1662145021
transform 1 0 70180 0 1 66990
box 0 0 3190 3190
use unit_cap  unit_cap_1166
timestamp 1662145021
transform 1 0 70180 0 1 70180
box 0 0 3190 3190
use unit_cap  unit_cap_1167
timestamp 1662145021
transform 1 0 70180 0 1 73370
box 0 0 3190 3190
use unit_cap  unit_cap_1168
timestamp 1662145021
transform 1 0 70180 0 1 76560
box 0 0 3190 3190
use unit_cap  unit_cap_1169
timestamp 1662145021
transform 1 0 70180 0 1 79750
box 0 0 3190 3190
use unit_cap  unit_cap_1170
timestamp 1662145021
transform 1 0 70180 0 1 82940
box 0 0 3190 3190
use unit_cap  unit_cap_1171
timestamp 1662145021
transform 1 0 70180 0 1 86130
box 0 0 3190 3190
use unit_cap  unit_cap_1172
timestamp 1662145021
transform 1 0 70180 0 1 89320
box 0 0 3190 3190
use unit_cap  unit_cap_1173
timestamp 1662145021
transform 1 0 70180 0 1 92510
box 0 0 3190 3190
use unit_cap  unit_cap_1174
timestamp 1662145021
transform 1 0 70180 0 1 95700
box 0 0 3190 3190
use unit_cap  unit_cap_1175
timestamp 1662145021
transform 1 0 70180 0 1 98890
box 0 0 3190 3190
use unit_cap  unit_cap_1176
timestamp 1662145021
transform 1 0 70180 0 1 102080
box 0 0 3190 3190
use unit_cap  unit_cap_1177
timestamp 1662145021
transform 1 0 70180 0 1 105270
box 0 0 3190 3190
use unit_cap  unit_cap_1178
timestamp 1662145021
transform 1 0 70180 0 1 108460
box 0 0 3190 3190
use unit_cap  unit_cap_1179
timestamp 1662145021
transform 1 0 70180 0 1 111650
box 0 0 3190 3190
use unit_cap  unit_cap_1180
timestamp 1662145021
transform 1 0 70180 0 1 114840
box 0 0 3190 3190
use unit_cap  unit_cap_1181
timestamp 1662145021
transform 1 0 70180 0 1 118030
box 0 0 3190 3190
use unit_cap  unit_cap_1182
timestamp 1662145021
transform 1 0 70180 0 1 121220
box 0 0 3190 3190
use unit_cap  unit_cap_1183
timestamp 1662145021
transform 1 0 70180 0 1 124410
box 0 0 3190 3190
use unit_cap  unit_cap_1184
timestamp 1662145021
transform 1 0 70180 0 1 127600
box 0 0 3190 3190
use unit_cap  unit_cap_1185
timestamp 1662145021
transform 1 0 70180 0 1 130790
box 0 0 3190 3190
use unit_cap  unit_cap_1186
timestamp 1662145021
transform 1 0 70180 0 1 133980
box 0 0 3190 3190
use unit_cap  unit_cap_1187
timestamp 1662145021
transform 1 0 70180 0 1 137170
box 0 0 3190 3190
use unit_cap  unit_cap_1188
timestamp 1662145021
transform 1 0 70180 0 1 140360
box 0 0 3190 3190
use unit_cap  unit_cap_1189
timestamp 1662145021
transform 1 0 70180 0 1 143550
box 0 0 3190 3190
use unit_cap  unit_cap_1190
timestamp 1662145021
transform 1 0 70180 0 1 146740
box 0 0 3190 3190
use unit_cap  unit_cap_1191
timestamp 1662145021
transform 1 0 70180 0 1 149930
box 0 0 3190 3190
use unit_cap  unit_cap_1192
timestamp 1662145021
transform 1 0 70180 0 1 153120
box 0 0 3190 3190
use unit_cap  unit_cap_1193
timestamp 1662145021
transform 1 0 70180 0 1 156310
box 0 0 3190 3190
use unit_cap  unit_cap_1194
timestamp 1662145021
transform 1 0 70180 0 1 159500
box 0 0 3190 3190
use unit_cap  unit_cap_1195
timestamp 1662145021
transform 1 0 70180 0 1 162690
box 0 0 3190 3190
use unit_cap  unit_cap_1196
timestamp 1662145021
transform 1 0 73370 0 1 0
box 0 0 3190 3190
use unit_cap  unit_cap_1197
timestamp 1662145021
transform 1 0 73370 0 1 3190
box 0 0 3190 3190
use unit_cap  unit_cap_1198
timestamp 1662145021
transform 1 0 73370 0 1 6380
box 0 0 3190 3190
use unit_cap  unit_cap_1199
timestamp 1662145021
transform 1 0 73370 0 1 9570
box 0 0 3190 3190
use unit_cap  unit_cap_1200
timestamp 1662145021
transform 1 0 73370 0 1 12760
box 0 0 3190 3190
use unit_cap  unit_cap_1201
timestamp 1662145021
transform 1 0 73370 0 1 15950
box 0 0 3190 3190
use unit_cap  unit_cap_1202
timestamp 1662145021
transform 1 0 73370 0 1 19140
box 0 0 3190 3190
use unit_cap  unit_cap_1203
timestamp 1662145021
transform 1 0 73370 0 1 22330
box 0 0 3190 3190
use unit_cap  unit_cap_1204
timestamp 1662145021
transform 1 0 73370 0 1 25520
box 0 0 3190 3190
use unit_cap  unit_cap_1205
timestamp 1662145021
transform 1 0 73370 0 1 28710
box 0 0 3190 3190
use unit_cap  unit_cap_1206
timestamp 1662145021
transform 1 0 73370 0 1 31900
box 0 0 3190 3190
use unit_cap  unit_cap_1207
timestamp 1662145021
transform 1 0 73370 0 1 35090
box 0 0 3190 3190
use unit_cap  unit_cap_1208
timestamp 1662145021
transform 1 0 73370 0 1 38280
box 0 0 3190 3190
use unit_cap  unit_cap_1209
timestamp 1662145021
transform 1 0 73370 0 1 41470
box 0 0 3190 3190
use unit_cap  unit_cap_1210
timestamp 1662145021
transform 1 0 73370 0 1 44660
box 0 0 3190 3190
use unit_cap  unit_cap_1211
timestamp 1662145021
transform 1 0 73370 0 1 47850
box 0 0 3190 3190
use unit_cap  unit_cap_1212
timestamp 1662145021
transform 1 0 73370 0 1 51040
box 0 0 3190 3190
use unit_cap  unit_cap_1213
timestamp 1662145021
transform 1 0 73370 0 1 54230
box 0 0 3190 3190
use unit_cap  unit_cap_1214
timestamp 1662145021
transform 1 0 73370 0 1 57420
box 0 0 3190 3190
use unit_cap  unit_cap_1215
timestamp 1662145021
transform 1 0 73370 0 1 60610
box 0 0 3190 3190
use unit_cap  unit_cap_1216
timestamp 1662145021
transform 1 0 73370 0 1 63800
box 0 0 3190 3190
use unit_cap  unit_cap_1217
timestamp 1662145021
transform 1 0 73370 0 1 66990
box 0 0 3190 3190
use unit_cap  unit_cap_1218
timestamp 1662145021
transform 1 0 73370 0 1 70180
box 0 0 3190 3190
use unit_cap  unit_cap_1219
timestamp 1662145021
transform 1 0 73370 0 1 73370
box 0 0 3190 3190
use unit_cap  unit_cap_1220
timestamp 1662145021
transform 1 0 73370 0 1 76560
box 0 0 3190 3190
use unit_cap  unit_cap_1221
timestamp 1662145021
transform 1 0 73370 0 1 79750
box 0 0 3190 3190
use unit_cap  unit_cap_1222
timestamp 1662145021
transform 1 0 73370 0 1 82940
box 0 0 3190 3190
use unit_cap  unit_cap_1223
timestamp 1662145021
transform 1 0 73370 0 1 86130
box 0 0 3190 3190
use unit_cap  unit_cap_1224
timestamp 1662145021
transform 1 0 73370 0 1 89320
box 0 0 3190 3190
use unit_cap  unit_cap_1225
timestamp 1662145021
transform 1 0 73370 0 1 92510
box 0 0 3190 3190
use unit_cap  unit_cap_1226
timestamp 1662145021
transform 1 0 73370 0 1 95700
box 0 0 3190 3190
use unit_cap  unit_cap_1227
timestamp 1662145021
transform 1 0 73370 0 1 98890
box 0 0 3190 3190
use unit_cap  unit_cap_1228
timestamp 1662145021
transform 1 0 73370 0 1 102080
box 0 0 3190 3190
use unit_cap  unit_cap_1229
timestamp 1662145021
transform 1 0 73370 0 1 105270
box 0 0 3190 3190
use unit_cap  unit_cap_1230
timestamp 1662145021
transform 1 0 73370 0 1 108460
box 0 0 3190 3190
use unit_cap  unit_cap_1231
timestamp 1662145021
transform 1 0 73370 0 1 111650
box 0 0 3190 3190
use unit_cap  unit_cap_1232
timestamp 1662145021
transform 1 0 73370 0 1 114840
box 0 0 3190 3190
use unit_cap  unit_cap_1233
timestamp 1662145021
transform 1 0 73370 0 1 118030
box 0 0 3190 3190
use unit_cap  unit_cap_1234
timestamp 1662145021
transform 1 0 73370 0 1 121220
box 0 0 3190 3190
use unit_cap  unit_cap_1235
timestamp 1662145021
transform 1 0 73370 0 1 124410
box 0 0 3190 3190
use unit_cap  unit_cap_1236
timestamp 1662145021
transform 1 0 73370 0 1 127600
box 0 0 3190 3190
use unit_cap  unit_cap_1237
timestamp 1662145021
transform 1 0 73370 0 1 130790
box 0 0 3190 3190
use unit_cap  unit_cap_1238
timestamp 1662145021
transform 1 0 73370 0 1 133980
box 0 0 3190 3190
use unit_cap  unit_cap_1239
timestamp 1662145021
transform 1 0 73370 0 1 137170
box 0 0 3190 3190
use unit_cap  unit_cap_1240
timestamp 1662145021
transform 1 0 73370 0 1 140360
box 0 0 3190 3190
use unit_cap  unit_cap_1241
timestamp 1662145021
transform 1 0 73370 0 1 143550
box 0 0 3190 3190
use unit_cap  unit_cap_1242
timestamp 1662145021
transform 1 0 73370 0 1 146740
box 0 0 3190 3190
use unit_cap  unit_cap_1243
timestamp 1662145021
transform 1 0 73370 0 1 149930
box 0 0 3190 3190
use unit_cap  unit_cap_1244
timestamp 1662145021
transform 1 0 73370 0 1 153120
box 0 0 3190 3190
use unit_cap  unit_cap_1245
timestamp 1662145021
transform 1 0 73370 0 1 156310
box 0 0 3190 3190
use unit_cap  unit_cap_1246
timestamp 1662145021
transform 1 0 73370 0 1 159500
box 0 0 3190 3190
use unit_cap  unit_cap_1247
timestamp 1662145021
transform 1 0 73370 0 1 162690
box 0 0 3190 3190
use unit_cap  unit_cap_1248
timestamp 1662145021
transform 1 0 76560 0 1 0
box 0 0 3190 3190
use unit_cap  unit_cap_1249
timestamp 1662145021
transform 1 0 76560 0 1 3190
box 0 0 3190 3190
use unit_cap  unit_cap_1250
timestamp 1662145021
transform 1 0 76560 0 1 6380
box 0 0 3190 3190
use unit_cap  unit_cap_1251
timestamp 1662145021
transform 1 0 76560 0 1 9570
box 0 0 3190 3190
use unit_cap  unit_cap_1252
timestamp 1662145021
transform 1 0 76560 0 1 12760
box 0 0 3190 3190
use unit_cap  unit_cap_1253
timestamp 1662145021
transform 1 0 76560 0 1 15950
box 0 0 3190 3190
use unit_cap  unit_cap_1254
timestamp 1662145021
transform 1 0 76560 0 1 19140
box 0 0 3190 3190
use unit_cap  unit_cap_1255
timestamp 1662145021
transform 1 0 76560 0 1 22330
box 0 0 3190 3190
use unit_cap  unit_cap_1256
timestamp 1662145021
transform 1 0 76560 0 1 25520
box 0 0 3190 3190
use unit_cap  unit_cap_1257
timestamp 1662145021
transform 1 0 76560 0 1 28710
box 0 0 3190 3190
use unit_cap  unit_cap_1258
timestamp 1662145021
transform 1 0 76560 0 1 31900
box 0 0 3190 3190
use unit_cap  unit_cap_1259
timestamp 1662145021
transform 1 0 76560 0 1 35090
box 0 0 3190 3190
use unit_cap  unit_cap_1260
timestamp 1662145021
transform 1 0 76560 0 1 38280
box 0 0 3190 3190
use unit_cap  unit_cap_1261
timestamp 1662145021
transform 1 0 76560 0 1 41470
box 0 0 3190 3190
use unit_cap  unit_cap_1262
timestamp 1662145021
transform 1 0 76560 0 1 44660
box 0 0 3190 3190
use unit_cap  unit_cap_1263
timestamp 1662145021
transform 1 0 76560 0 1 47850
box 0 0 3190 3190
use unit_cap  unit_cap_1264
timestamp 1662145021
transform 1 0 76560 0 1 51040
box 0 0 3190 3190
use unit_cap  unit_cap_1265
timestamp 1662145021
transform 1 0 76560 0 1 54230
box 0 0 3190 3190
use unit_cap  unit_cap_1266
timestamp 1662145021
transform 1 0 76560 0 1 57420
box 0 0 3190 3190
use unit_cap  unit_cap_1267
timestamp 1662145021
transform 1 0 76560 0 1 60610
box 0 0 3190 3190
use unit_cap  unit_cap_1268
timestamp 1662145021
transform 1 0 76560 0 1 63800
box 0 0 3190 3190
use unit_cap  unit_cap_1269
timestamp 1662145021
transform 1 0 76560 0 1 66990
box 0 0 3190 3190
use unit_cap  unit_cap_1270
timestamp 1662145021
transform 1 0 76560 0 1 70180
box 0 0 3190 3190
use unit_cap  unit_cap_1271
timestamp 1662145021
transform 1 0 76560 0 1 73370
box 0 0 3190 3190
use unit_cap  unit_cap_1272
timestamp 1662145021
transform 1 0 76560 0 1 76560
box 0 0 3190 3190
use unit_cap  unit_cap_1273
timestamp 1662145021
transform 1 0 76560 0 1 79750
box 0 0 3190 3190
use unit_cap  unit_cap_1274
timestamp 1662145021
transform 1 0 76560 0 1 82940
box 0 0 3190 3190
use unit_cap  unit_cap_1275
timestamp 1662145021
transform 1 0 76560 0 1 86130
box 0 0 3190 3190
use unit_cap  unit_cap_1276
timestamp 1662145021
transform 1 0 76560 0 1 89320
box 0 0 3190 3190
use unit_cap  unit_cap_1277
timestamp 1662145021
transform 1 0 76560 0 1 92510
box 0 0 3190 3190
use unit_cap  unit_cap_1278
timestamp 1662145021
transform 1 0 76560 0 1 95700
box 0 0 3190 3190
use unit_cap  unit_cap_1279
timestamp 1662145021
transform 1 0 76560 0 1 98890
box 0 0 3190 3190
use unit_cap  unit_cap_1280
timestamp 1662145021
transform 1 0 76560 0 1 102080
box 0 0 3190 3190
use unit_cap  unit_cap_1281
timestamp 1662145021
transform 1 0 76560 0 1 105270
box 0 0 3190 3190
use unit_cap  unit_cap_1282
timestamp 1662145021
transform 1 0 76560 0 1 108460
box 0 0 3190 3190
use unit_cap  unit_cap_1283
timestamp 1662145021
transform 1 0 76560 0 1 111650
box 0 0 3190 3190
use unit_cap  unit_cap_1284
timestamp 1662145021
transform 1 0 76560 0 1 114840
box 0 0 3190 3190
use unit_cap  unit_cap_1285
timestamp 1662145021
transform 1 0 76560 0 1 118030
box 0 0 3190 3190
use unit_cap  unit_cap_1286
timestamp 1662145021
transform 1 0 76560 0 1 121220
box 0 0 3190 3190
use unit_cap  unit_cap_1287
timestamp 1662145021
transform 1 0 76560 0 1 124410
box 0 0 3190 3190
use unit_cap  unit_cap_1288
timestamp 1662145021
transform 1 0 76560 0 1 127600
box 0 0 3190 3190
use unit_cap  unit_cap_1289
timestamp 1662145021
transform 1 0 76560 0 1 130790
box 0 0 3190 3190
use unit_cap  unit_cap_1290
timestamp 1662145021
transform 1 0 76560 0 1 133980
box 0 0 3190 3190
use unit_cap  unit_cap_1291
timestamp 1662145021
transform 1 0 76560 0 1 137170
box 0 0 3190 3190
use unit_cap  unit_cap_1292
timestamp 1662145021
transform 1 0 76560 0 1 140360
box 0 0 3190 3190
use unit_cap  unit_cap_1293
timestamp 1662145021
transform 1 0 76560 0 1 143550
box 0 0 3190 3190
use unit_cap  unit_cap_1294
timestamp 1662145021
transform 1 0 76560 0 1 146740
box 0 0 3190 3190
use unit_cap  unit_cap_1295
timestamp 1662145021
transform 1 0 76560 0 1 149930
box 0 0 3190 3190
use unit_cap  unit_cap_1296
timestamp 1662145021
transform 1 0 76560 0 1 153120
box 0 0 3190 3190
use unit_cap  unit_cap_1297
timestamp 1662145021
transform 1 0 76560 0 1 156310
box 0 0 3190 3190
use unit_cap  unit_cap_1298
timestamp 1662145021
transform 1 0 76560 0 1 159500
box 0 0 3190 3190
use unit_cap  unit_cap_1299
timestamp 1662145021
transform 1 0 76560 0 1 162690
box 0 0 3190 3190
use unit_cap  unit_cap_1300
timestamp 1662145021
transform 1 0 79750 0 1 0
box 0 0 3190 3190
use unit_cap  unit_cap_1301
timestamp 1662145021
transform 1 0 79750 0 1 3190
box 0 0 3190 3190
use unit_cap  unit_cap_1302
timestamp 1662145021
transform 1 0 79750 0 1 6380
box 0 0 3190 3190
use unit_cap  unit_cap_1303
timestamp 1662145021
transform 1 0 79750 0 1 9570
box 0 0 3190 3190
use unit_cap  unit_cap_1304
timestamp 1662145021
transform 1 0 79750 0 1 12760
box 0 0 3190 3190
use unit_cap  unit_cap_1305
timestamp 1662145021
transform 1 0 79750 0 1 15950
box 0 0 3190 3190
use unit_cap  unit_cap_1306
timestamp 1662145021
transform 1 0 79750 0 1 19140
box 0 0 3190 3190
use unit_cap  unit_cap_1307
timestamp 1662145021
transform 1 0 79750 0 1 22330
box 0 0 3190 3190
use unit_cap  unit_cap_1308
timestamp 1662145021
transform 1 0 79750 0 1 25520
box 0 0 3190 3190
use unit_cap  unit_cap_1309
timestamp 1662145021
transform 1 0 79750 0 1 28710
box 0 0 3190 3190
use unit_cap  unit_cap_1310
timestamp 1662145021
transform 1 0 79750 0 1 31900
box 0 0 3190 3190
use unit_cap  unit_cap_1311
timestamp 1662145021
transform 1 0 79750 0 1 35090
box 0 0 3190 3190
use unit_cap  unit_cap_1312
timestamp 1662145021
transform 1 0 79750 0 1 38280
box 0 0 3190 3190
use unit_cap  unit_cap_1313
timestamp 1662145021
transform 1 0 79750 0 1 41470
box 0 0 3190 3190
use unit_cap  unit_cap_1314
timestamp 1662145021
transform 1 0 79750 0 1 44660
box 0 0 3190 3190
use unit_cap  unit_cap_1315
timestamp 1662145021
transform 1 0 79750 0 1 47850
box 0 0 3190 3190
use unit_cap  unit_cap_1316
timestamp 1662145021
transform 1 0 79750 0 1 51040
box 0 0 3190 3190
use unit_cap  unit_cap_1317
timestamp 1662145021
transform 1 0 79750 0 1 54230
box 0 0 3190 3190
use unit_cap  unit_cap_1318
timestamp 1662145021
transform 1 0 79750 0 1 57420
box 0 0 3190 3190
use unit_cap  unit_cap_1319
timestamp 1662145021
transform 1 0 79750 0 1 60610
box 0 0 3190 3190
use unit_cap  unit_cap_1320
timestamp 1662145021
transform 1 0 79750 0 1 63800
box 0 0 3190 3190
use unit_cap  unit_cap_1321
timestamp 1662145021
transform 1 0 79750 0 1 66990
box 0 0 3190 3190
use unit_cap  unit_cap_1322
timestamp 1662145021
transform 1 0 79750 0 1 70180
box 0 0 3190 3190
use unit_cap  unit_cap_1323
timestamp 1662145021
transform 1 0 79750 0 1 73370
box 0 0 3190 3190
use unit_cap  unit_cap_1324
timestamp 1662145021
transform 1 0 79750 0 1 76560
box 0 0 3190 3190
use unit_cap  unit_cap_1325
timestamp 1662145021
transform 1 0 79750 0 1 79750
box 0 0 3190 3190
use unit_cap  unit_cap_1326
timestamp 1662145021
transform 1 0 79750 0 1 82940
box 0 0 3190 3190
use unit_cap  unit_cap_1327
timestamp 1662145021
transform 1 0 79750 0 1 86130
box 0 0 3190 3190
use unit_cap  unit_cap_1328
timestamp 1662145021
transform 1 0 79750 0 1 89320
box 0 0 3190 3190
use unit_cap  unit_cap_1329
timestamp 1662145021
transform 1 0 79750 0 1 92510
box 0 0 3190 3190
use unit_cap  unit_cap_1330
timestamp 1662145021
transform 1 0 79750 0 1 95700
box 0 0 3190 3190
use unit_cap  unit_cap_1331
timestamp 1662145021
transform 1 0 79750 0 1 98890
box 0 0 3190 3190
use unit_cap  unit_cap_1332
timestamp 1662145021
transform 1 0 79750 0 1 102080
box 0 0 3190 3190
use unit_cap  unit_cap_1333
timestamp 1662145021
transform 1 0 79750 0 1 105270
box 0 0 3190 3190
use unit_cap  unit_cap_1334
timestamp 1662145021
transform 1 0 79750 0 1 108460
box 0 0 3190 3190
use unit_cap  unit_cap_1335
timestamp 1662145021
transform 1 0 79750 0 1 111650
box 0 0 3190 3190
use unit_cap  unit_cap_1336
timestamp 1662145021
transform 1 0 79750 0 1 114840
box 0 0 3190 3190
use unit_cap  unit_cap_1337
timestamp 1662145021
transform 1 0 79750 0 1 118030
box 0 0 3190 3190
use unit_cap  unit_cap_1338
timestamp 1662145021
transform 1 0 79750 0 1 121220
box 0 0 3190 3190
use unit_cap  unit_cap_1339
timestamp 1662145021
transform 1 0 79750 0 1 124410
box 0 0 3190 3190
use unit_cap  unit_cap_1340
timestamp 1662145021
transform 1 0 79750 0 1 127600
box 0 0 3190 3190
use unit_cap  unit_cap_1341
timestamp 1662145021
transform 1 0 79750 0 1 130790
box 0 0 3190 3190
use unit_cap  unit_cap_1342
timestamp 1662145021
transform 1 0 79750 0 1 133980
box 0 0 3190 3190
use unit_cap  unit_cap_1343
timestamp 1662145021
transform 1 0 79750 0 1 137170
box 0 0 3190 3190
use unit_cap  unit_cap_1344
timestamp 1662145021
transform 1 0 79750 0 1 140360
box 0 0 3190 3190
use unit_cap  unit_cap_1345
timestamp 1662145021
transform 1 0 79750 0 1 143550
box 0 0 3190 3190
use unit_cap  unit_cap_1346
timestamp 1662145021
transform 1 0 79750 0 1 146740
box 0 0 3190 3190
use unit_cap  unit_cap_1347
timestamp 1662145021
transform 1 0 79750 0 1 149930
box 0 0 3190 3190
use unit_cap  unit_cap_1348
timestamp 1662145021
transform 1 0 79750 0 1 153120
box 0 0 3190 3190
use unit_cap  unit_cap_1349
timestamp 1662145021
transform 1 0 79750 0 1 156310
box 0 0 3190 3190
use unit_cap  unit_cap_1350
timestamp 1662145021
transform 1 0 79750 0 1 159500
box 0 0 3190 3190
use unit_cap  unit_cap_1351
timestamp 1662145021
transform 1 0 79750 0 1 162690
box 0 0 3190 3190
use unit_cap  unit_cap_1352
timestamp 1662145021
transform 1 0 82940 0 1 0
box 0 0 3190 3190
use unit_cap  unit_cap_1353
timestamp 1662145021
transform 1 0 82940 0 1 3190
box 0 0 3190 3190
use unit_cap  unit_cap_1354
timestamp 1662145021
transform 1 0 82940 0 1 6380
box 0 0 3190 3190
use unit_cap  unit_cap_1355
timestamp 1662145021
transform 1 0 82940 0 1 9570
box 0 0 3190 3190
use unit_cap  unit_cap_1356
timestamp 1662145021
transform 1 0 82940 0 1 12760
box 0 0 3190 3190
use unit_cap  unit_cap_1357
timestamp 1662145021
transform 1 0 82940 0 1 15950
box 0 0 3190 3190
use unit_cap  unit_cap_1358
timestamp 1662145021
transform 1 0 82940 0 1 19140
box 0 0 3190 3190
use unit_cap  unit_cap_1359
timestamp 1662145021
transform 1 0 82940 0 1 22330
box 0 0 3190 3190
use unit_cap  unit_cap_1360
timestamp 1662145021
transform 1 0 82940 0 1 25520
box 0 0 3190 3190
use unit_cap  unit_cap_1361
timestamp 1662145021
transform 1 0 82940 0 1 28710
box 0 0 3190 3190
use unit_cap  unit_cap_1362
timestamp 1662145021
transform 1 0 82940 0 1 31900
box 0 0 3190 3190
use unit_cap  unit_cap_1363
timestamp 1662145021
transform 1 0 82940 0 1 35090
box 0 0 3190 3190
use unit_cap  unit_cap_1364
timestamp 1662145021
transform 1 0 82940 0 1 38280
box 0 0 3190 3190
use unit_cap  unit_cap_1365
timestamp 1662145021
transform 1 0 82940 0 1 41470
box 0 0 3190 3190
use unit_cap  unit_cap_1366
timestamp 1662145021
transform 1 0 82940 0 1 44660
box 0 0 3190 3190
use unit_cap  unit_cap_1367
timestamp 1662145021
transform 1 0 82940 0 1 47850
box 0 0 3190 3190
use unit_cap  unit_cap_1368
timestamp 1662145021
transform 1 0 82940 0 1 51040
box 0 0 3190 3190
use unit_cap  unit_cap_1369
timestamp 1662145021
transform 1 0 82940 0 1 54230
box 0 0 3190 3190
use unit_cap  unit_cap_1370
timestamp 1662145021
transform 1 0 82940 0 1 57420
box 0 0 3190 3190
use unit_cap  unit_cap_1371
timestamp 1662145021
transform 1 0 82940 0 1 60610
box 0 0 3190 3190
use unit_cap  unit_cap_1372
timestamp 1662145021
transform 1 0 82940 0 1 63800
box 0 0 3190 3190
use unit_cap  unit_cap_1373
timestamp 1662145021
transform 1 0 82940 0 1 66990
box 0 0 3190 3190
use unit_cap  unit_cap_1374
timestamp 1662145021
transform 1 0 82940 0 1 70180
box 0 0 3190 3190
use unit_cap  unit_cap_1375
timestamp 1662145021
transform 1 0 82940 0 1 73370
box 0 0 3190 3190
use unit_cap  unit_cap_1376
timestamp 1662145021
transform 1 0 82940 0 1 76560
box 0 0 3190 3190
use unit_cap  unit_cap_1377
timestamp 1662145021
transform 1 0 82940 0 1 79750
box 0 0 3190 3190
use unit_cap  unit_cap_1378
timestamp 1662145021
transform 1 0 82940 0 1 82940
box 0 0 3190 3190
use unit_cap  unit_cap_1379
timestamp 1662145021
transform 1 0 82940 0 1 86130
box 0 0 3190 3190
use unit_cap  unit_cap_1380
timestamp 1662145021
transform 1 0 82940 0 1 89320
box 0 0 3190 3190
use unit_cap  unit_cap_1381
timestamp 1662145021
transform 1 0 82940 0 1 92510
box 0 0 3190 3190
use unit_cap  unit_cap_1382
timestamp 1662145021
transform 1 0 82940 0 1 95700
box 0 0 3190 3190
use unit_cap  unit_cap_1383
timestamp 1662145021
transform 1 0 82940 0 1 98890
box 0 0 3190 3190
use unit_cap  unit_cap_1384
timestamp 1662145021
transform 1 0 82940 0 1 102080
box 0 0 3190 3190
use unit_cap  unit_cap_1385
timestamp 1662145021
transform 1 0 82940 0 1 105270
box 0 0 3190 3190
use unit_cap  unit_cap_1386
timestamp 1662145021
transform 1 0 82940 0 1 108460
box 0 0 3190 3190
use unit_cap  unit_cap_1387
timestamp 1662145021
transform 1 0 82940 0 1 111650
box 0 0 3190 3190
use unit_cap  unit_cap_1388
timestamp 1662145021
transform 1 0 82940 0 1 114840
box 0 0 3190 3190
use unit_cap  unit_cap_1389
timestamp 1662145021
transform 1 0 82940 0 1 118030
box 0 0 3190 3190
use unit_cap  unit_cap_1390
timestamp 1662145021
transform 1 0 82940 0 1 121220
box 0 0 3190 3190
use unit_cap  unit_cap_1391
timestamp 1662145021
transform 1 0 82940 0 1 124410
box 0 0 3190 3190
use unit_cap  unit_cap_1392
timestamp 1662145021
transform 1 0 82940 0 1 127600
box 0 0 3190 3190
use unit_cap  unit_cap_1393
timestamp 1662145021
transform 1 0 82940 0 1 130790
box 0 0 3190 3190
use unit_cap  unit_cap_1394
timestamp 1662145021
transform 1 0 82940 0 1 133980
box 0 0 3190 3190
use unit_cap  unit_cap_1395
timestamp 1662145021
transform 1 0 82940 0 1 137170
box 0 0 3190 3190
use unit_cap  unit_cap_1396
timestamp 1662145021
transform 1 0 82940 0 1 140360
box 0 0 3190 3190
use unit_cap  unit_cap_1397
timestamp 1662145021
transform 1 0 82940 0 1 143550
box 0 0 3190 3190
use unit_cap  unit_cap_1398
timestamp 1662145021
transform 1 0 82940 0 1 146740
box 0 0 3190 3190
use unit_cap  unit_cap_1399
timestamp 1662145021
transform 1 0 82940 0 1 149930
box 0 0 3190 3190
use unit_cap  unit_cap_1400
timestamp 1662145021
transform 1 0 82940 0 1 153120
box 0 0 3190 3190
use unit_cap  unit_cap_1401
timestamp 1662145021
transform 1 0 82940 0 1 156310
box 0 0 3190 3190
use unit_cap  unit_cap_1402
timestamp 1662145021
transform 1 0 82940 0 1 159500
box 0 0 3190 3190
use unit_cap  unit_cap_1403
timestamp 1662145021
transform 1 0 82940 0 1 162690
box 0 0 3190 3190
use unit_cap  unit_cap_1404
timestamp 1662145021
transform 1 0 86130 0 1 0
box 0 0 3190 3190
use unit_cap  unit_cap_1405
timestamp 1662145021
transform 1 0 86130 0 1 3190
box 0 0 3190 3190
use unit_cap  unit_cap_1406
timestamp 1662145021
transform 1 0 86130 0 1 6380
box 0 0 3190 3190
use unit_cap  unit_cap_1407
timestamp 1662145021
transform 1 0 86130 0 1 9570
box 0 0 3190 3190
use unit_cap  unit_cap_1408
timestamp 1662145021
transform 1 0 86130 0 1 12760
box 0 0 3190 3190
use unit_cap  unit_cap_1409
timestamp 1662145021
transform 1 0 86130 0 1 15950
box 0 0 3190 3190
use unit_cap  unit_cap_1410
timestamp 1662145021
transform 1 0 86130 0 1 19140
box 0 0 3190 3190
use unit_cap  unit_cap_1411
timestamp 1662145021
transform 1 0 86130 0 1 22330
box 0 0 3190 3190
use unit_cap  unit_cap_1412
timestamp 1662145021
transform 1 0 86130 0 1 25520
box 0 0 3190 3190
use unit_cap  unit_cap_1413
timestamp 1662145021
transform 1 0 86130 0 1 28710
box 0 0 3190 3190
use unit_cap  unit_cap_1414
timestamp 1662145021
transform 1 0 86130 0 1 31900
box 0 0 3190 3190
use unit_cap  unit_cap_1415
timestamp 1662145021
transform 1 0 86130 0 1 35090
box 0 0 3190 3190
use unit_cap  unit_cap_1416
timestamp 1662145021
transform 1 0 86130 0 1 38280
box 0 0 3190 3190
use unit_cap  unit_cap_1417
timestamp 1662145021
transform 1 0 86130 0 1 41470
box 0 0 3190 3190
use unit_cap  unit_cap_1418
timestamp 1662145021
transform 1 0 86130 0 1 44660
box 0 0 3190 3190
use unit_cap  unit_cap_1419
timestamp 1662145021
transform 1 0 86130 0 1 47850
box 0 0 3190 3190
use unit_cap  unit_cap_1420
timestamp 1662145021
transform 1 0 86130 0 1 51040
box 0 0 3190 3190
use unit_cap  unit_cap_1421
timestamp 1662145021
transform 1 0 86130 0 1 54230
box 0 0 3190 3190
use unit_cap  unit_cap_1422
timestamp 1662145021
transform 1 0 86130 0 1 57420
box 0 0 3190 3190
use unit_cap  unit_cap_1423
timestamp 1662145021
transform 1 0 86130 0 1 60610
box 0 0 3190 3190
use unit_cap  unit_cap_1424
timestamp 1662145021
transform 1 0 86130 0 1 63800
box 0 0 3190 3190
use unit_cap  unit_cap_1425
timestamp 1662145021
transform 1 0 86130 0 1 66990
box 0 0 3190 3190
use unit_cap  unit_cap_1426
timestamp 1662145021
transform 1 0 86130 0 1 70180
box 0 0 3190 3190
use unit_cap  unit_cap_1427
timestamp 1662145021
transform 1 0 86130 0 1 73370
box 0 0 3190 3190
use unit_cap  unit_cap_1428
timestamp 1662145021
transform 1 0 86130 0 1 76560
box 0 0 3190 3190
use unit_cap  unit_cap_1429
timestamp 1662145021
transform 1 0 86130 0 1 79750
box 0 0 3190 3190
use unit_cap  unit_cap_1430
timestamp 1662145021
transform 1 0 86130 0 1 82940
box 0 0 3190 3190
use unit_cap  unit_cap_1431
timestamp 1662145021
transform 1 0 86130 0 1 86130
box 0 0 3190 3190
use unit_cap  unit_cap_1432
timestamp 1662145021
transform 1 0 86130 0 1 89320
box 0 0 3190 3190
use unit_cap  unit_cap_1433
timestamp 1662145021
transform 1 0 86130 0 1 92510
box 0 0 3190 3190
use unit_cap  unit_cap_1434
timestamp 1662145021
transform 1 0 86130 0 1 95700
box 0 0 3190 3190
use unit_cap  unit_cap_1435
timestamp 1662145021
transform 1 0 86130 0 1 98890
box 0 0 3190 3190
use unit_cap  unit_cap_1436
timestamp 1662145021
transform 1 0 86130 0 1 102080
box 0 0 3190 3190
use unit_cap  unit_cap_1437
timestamp 1662145021
transform 1 0 86130 0 1 105270
box 0 0 3190 3190
use unit_cap  unit_cap_1438
timestamp 1662145021
transform 1 0 86130 0 1 108460
box 0 0 3190 3190
use unit_cap  unit_cap_1439
timestamp 1662145021
transform 1 0 86130 0 1 111650
box 0 0 3190 3190
use unit_cap  unit_cap_1440
timestamp 1662145021
transform 1 0 86130 0 1 114840
box 0 0 3190 3190
use unit_cap  unit_cap_1441
timestamp 1662145021
transform 1 0 86130 0 1 118030
box 0 0 3190 3190
use unit_cap  unit_cap_1442
timestamp 1662145021
transform 1 0 86130 0 1 121220
box 0 0 3190 3190
use unit_cap  unit_cap_1443
timestamp 1662145021
transform 1 0 86130 0 1 124410
box 0 0 3190 3190
use unit_cap  unit_cap_1444
timestamp 1662145021
transform 1 0 86130 0 1 127600
box 0 0 3190 3190
use unit_cap  unit_cap_1445
timestamp 1662145021
transform 1 0 86130 0 1 130790
box 0 0 3190 3190
use unit_cap  unit_cap_1446
timestamp 1662145021
transform 1 0 86130 0 1 133980
box 0 0 3190 3190
use unit_cap  unit_cap_1447
timestamp 1662145021
transform 1 0 86130 0 1 137170
box 0 0 3190 3190
use unit_cap  unit_cap_1448
timestamp 1662145021
transform 1 0 86130 0 1 140360
box 0 0 3190 3190
use unit_cap  unit_cap_1449
timestamp 1662145021
transform 1 0 86130 0 1 143550
box 0 0 3190 3190
use unit_cap  unit_cap_1450
timestamp 1662145021
transform 1 0 86130 0 1 146740
box 0 0 3190 3190
use unit_cap  unit_cap_1451
timestamp 1662145021
transform 1 0 86130 0 1 149930
box 0 0 3190 3190
use unit_cap  unit_cap_1452
timestamp 1662145021
transform 1 0 86130 0 1 153120
box 0 0 3190 3190
use unit_cap  unit_cap_1453
timestamp 1662145021
transform 1 0 86130 0 1 156310
box 0 0 3190 3190
use unit_cap  unit_cap_1454
timestamp 1662145021
transform 1 0 86130 0 1 159500
box 0 0 3190 3190
use unit_cap  unit_cap_1455
timestamp 1662145021
transform 1 0 86130 0 1 162690
box 0 0 3190 3190
use unit_cap  unit_cap_1456
timestamp 1662145021
transform 1 0 89320 0 1 0
box 0 0 3190 3190
use unit_cap  unit_cap_1457
timestamp 1662145021
transform 1 0 89320 0 1 3190
box 0 0 3190 3190
use unit_cap  unit_cap_1458
timestamp 1662145021
transform 1 0 89320 0 1 6380
box 0 0 3190 3190
use unit_cap  unit_cap_1459
timestamp 1662145021
transform 1 0 89320 0 1 9570
box 0 0 3190 3190
use unit_cap  unit_cap_1460
timestamp 1662145021
transform 1 0 89320 0 1 12760
box 0 0 3190 3190
use unit_cap  unit_cap_1461
timestamp 1662145021
transform 1 0 89320 0 1 15950
box 0 0 3190 3190
use unit_cap  unit_cap_1462
timestamp 1662145021
transform 1 0 89320 0 1 19140
box 0 0 3190 3190
use unit_cap  unit_cap_1463
timestamp 1662145021
transform 1 0 89320 0 1 22330
box 0 0 3190 3190
use unit_cap  unit_cap_1464
timestamp 1662145021
transform 1 0 89320 0 1 25520
box 0 0 3190 3190
use unit_cap  unit_cap_1465
timestamp 1662145021
transform 1 0 89320 0 1 28710
box 0 0 3190 3190
use unit_cap  unit_cap_1466
timestamp 1662145021
transform 1 0 89320 0 1 31900
box 0 0 3190 3190
use unit_cap  unit_cap_1467
timestamp 1662145021
transform 1 0 89320 0 1 35090
box 0 0 3190 3190
use unit_cap  unit_cap_1468
timestamp 1662145021
transform 1 0 89320 0 1 38280
box 0 0 3190 3190
use unit_cap  unit_cap_1469
timestamp 1662145021
transform 1 0 89320 0 1 41470
box 0 0 3190 3190
use unit_cap  unit_cap_1470
timestamp 1662145021
transform 1 0 89320 0 1 44660
box 0 0 3190 3190
use unit_cap  unit_cap_1471
timestamp 1662145021
transform 1 0 89320 0 1 47850
box 0 0 3190 3190
use unit_cap  unit_cap_1472
timestamp 1662145021
transform 1 0 89320 0 1 51040
box 0 0 3190 3190
use unit_cap  unit_cap_1473
timestamp 1662145021
transform 1 0 89320 0 1 54230
box 0 0 3190 3190
use unit_cap  unit_cap_1474
timestamp 1662145021
transform 1 0 89320 0 1 57420
box 0 0 3190 3190
use unit_cap  unit_cap_1475
timestamp 1662145021
transform 1 0 89320 0 1 60610
box 0 0 3190 3190
use unit_cap  unit_cap_1476
timestamp 1662145021
transform 1 0 89320 0 1 63800
box 0 0 3190 3190
use unit_cap  unit_cap_1477
timestamp 1662145021
transform 1 0 89320 0 1 66990
box 0 0 3190 3190
use unit_cap  unit_cap_1478
timestamp 1662145021
transform 1 0 89320 0 1 70180
box 0 0 3190 3190
use unit_cap  unit_cap_1479
timestamp 1662145021
transform 1 0 89320 0 1 73370
box 0 0 3190 3190
use unit_cap  unit_cap_1480
timestamp 1662145021
transform 1 0 89320 0 1 76560
box 0 0 3190 3190
use unit_cap  unit_cap_1481
timestamp 1662145021
transform 1 0 89320 0 1 79750
box 0 0 3190 3190
use unit_cap  unit_cap_1482
timestamp 1662145021
transform 1 0 89320 0 1 82940
box 0 0 3190 3190
use unit_cap  unit_cap_1483
timestamp 1662145021
transform 1 0 89320 0 1 86130
box 0 0 3190 3190
use unit_cap  unit_cap_1484
timestamp 1662145021
transform 1 0 89320 0 1 89320
box 0 0 3190 3190
use unit_cap  unit_cap_1485
timestamp 1662145021
transform 1 0 89320 0 1 92510
box 0 0 3190 3190
use unit_cap  unit_cap_1486
timestamp 1662145021
transform 1 0 89320 0 1 95700
box 0 0 3190 3190
use unit_cap  unit_cap_1487
timestamp 1662145021
transform 1 0 89320 0 1 98890
box 0 0 3190 3190
use unit_cap  unit_cap_1488
timestamp 1662145021
transform 1 0 89320 0 1 102080
box 0 0 3190 3190
use unit_cap  unit_cap_1489
timestamp 1662145021
transform 1 0 89320 0 1 105270
box 0 0 3190 3190
use unit_cap  unit_cap_1490
timestamp 1662145021
transform 1 0 89320 0 1 108460
box 0 0 3190 3190
use unit_cap  unit_cap_1491
timestamp 1662145021
transform 1 0 89320 0 1 111650
box 0 0 3190 3190
use unit_cap  unit_cap_1492
timestamp 1662145021
transform 1 0 89320 0 1 114840
box 0 0 3190 3190
use unit_cap  unit_cap_1493
timestamp 1662145021
transform 1 0 89320 0 1 118030
box 0 0 3190 3190
use unit_cap  unit_cap_1494
timestamp 1662145021
transform 1 0 89320 0 1 121220
box 0 0 3190 3190
use unit_cap  unit_cap_1495
timestamp 1662145021
transform 1 0 89320 0 1 124410
box 0 0 3190 3190
use unit_cap  unit_cap_1496
timestamp 1662145021
transform 1 0 89320 0 1 127600
box 0 0 3190 3190
use unit_cap  unit_cap_1497
timestamp 1662145021
transform 1 0 89320 0 1 130790
box 0 0 3190 3190
use unit_cap  unit_cap_1498
timestamp 1662145021
transform 1 0 89320 0 1 133980
box 0 0 3190 3190
use unit_cap  unit_cap_1499
timestamp 1662145021
transform 1 0 89320 0 1 137170
box 0 0 3190 3190
use unit_cap  unit_cap_1500
timestamp 1662145021
transform 1 0 89320 0 1 140360
box 0 0 3190 3190
use unit_cap  unit_cap_1501
timestamp 1662145021
transform 1 0 89320 0 1 143550
box 0 0 3190 3190
use unit_cap  unit_cap_1502
timestamp 1662145021
transform 1 0 89320 0 1 146740
box 0 0 3190 3190
use unit_cap  unit_cap_1503
timestamp 1662145021
transform 1 0 89320 0 1 149930
box 0 0 3190 3190
use unit_cap  unit_cap_1504
timestamp 1662145021
transform 1 0 89320 0 1 153120
box 0 0 3190 3190
use unit_cap  unit_cap_1505
timestamp 1662145021
transform 1 0 89320 0 1 156310
box 0 0 3190 3190
use unit_cap  unit_cap_1506
timestamp 1662145021
transform 1 0 89320 0 1 159500
box 0 0 3190 3190
use unit_cap  unit_cap_1507
timestamp 1662145021
transform 1 0 89320 0 1 162690
box 0 0 3190 3190
use unit_cap  unit_cap_1508
timestamp 1662145021
transform 1 0 92510 0 1 0
box 0 0 3190 3190
use unit_cap  unit_cap_1509
timestamp 1662145021
transform 1 0 92510 0 1 3190
box 0 0 3190 3190
use unit_cap  unit_cap_1510
timestamp 1662145021
transform 1 0 92510 0 1 6380
box 0 0 3190 3190
use unit_cap  unit_cap_1511
timestamp 1662145021
transform 1 0 92510 0 1 9570
box 0 0 3190 3190
use unit_cap  unit_cap_1512
timestamp 1662145021
transform 1 0 92510 0 1 12760
box 0 0 3190 3190
use unit_cap  unit_cap_1513
timestamp 1662145021
transform 1 0 92510 0 1 15950
box 0 0 3190 3190
use unit_cap  unit_cap_1514
timestamp 1662145021
transform 1 0 92510 0 1 19140
box 0 0 3190 3190
use unit_cap  unit_cap_1515
timestamp 1662145021
transform 1 0 92510 0 1 22330
box 0 0 3190 3190
use unit_cap  unit_cap_1516
timestamp 1662145021
transform 1 0 92510 0 1 25520
box 0 0 3190 3190
use unit_cap  unit_cap_1517
timestamp 1662145021
transform 1 0 92510 0 1 28710
box 0 0 3190 3190
use unit_cap  unit_cap_1518
timestamp 1662145021
transform 1 0 92510 0 1 31900
box 0 0 3190 3190
use unit_cap  unit_cap_1519
timestamp 1662145021
transform 1 0 92510 0 1 35090
box 0 0 3190 3190
use unit_cap  unit_cap_1520
timestamp 1662145021
transform 1 0 92510 0 1 38280
box 0 0 3190 3190
use unit_cap  unit_cap_1521
timestamp 1662145021
transform 1 0 92510 0 1 41470
box 0 0 3190 3190
use unit_cap  unit_cap_1522
timestamp 1662145021
transform 1 0 92510 0 1 44660
box 0 0 3190 3190
use unit_cap  unit_cap_1523
timestamp 1662145021
transform 1 0 92510 0 1 47850
box 0 0 3190 3190
use unit_cap  unit_cap_1524
timestamp 1662145021
transform 1 0 92510 0 1 51040
box 0 0 3190 3190
use unit_cap  unit_cap_1525
timestamp 1662145021
transform 1 0 92510 0 1 54230
box 0 0 3190 3190
use unit_cap  unit_cap_1526
timestamp 1662145021
transform 1 0 92510 0 1 57420
box 0 0 3190 3190
use unit_cap  unit_cap_1527
timestamp 1662145021
transform 1 0 92510 0 1 60610
box 0 0 3190 3190
use unit_cap  unit_cap_1528
timestamp 1662145021
transform 1 0 92510 0 1 63800
box 0 0 3190 3190
use unit_cap  unit_cap_1529
timestamp 1662145021
transform 1 0 92510 0 1 66990
box 0 0 3190 3190
use unit_cap  unit_cap_1530
timestamp 1662145021
transform 1 0 92510 0 1 70180
box 0 0 3190 3190
use unit_cap  unit_cap_1531
timestamp 1662145021
transform 1 0 92510 0 1 73370
box 0 0 3190 3190
use unit_cap  unit_cap_1532
timestamp 1662145021
transform 1 0 92510 0 1 76560
box 0 0 3190 3190
use unit_cap  unit_cap_1533
timestamp 1662145021
transform 1 0 92510 0 1 79750
box 0 0 3190 3190
use unit_cap  unit_cap_1534
timestamp 1662145021
transform 1 0 92510 0 1 82940
box 0 0 3190 3190
use unit_cap  unit_cap_1535
timestamp 1662145021
transform 1 0 92510 0 1 86130
box 0 0 3190 3190
use unit_cap  unit_cap_1536
timestamp 1662145021
transform 1 0 92510 0 1 89320
box 0 0 3190 3190
use unit_cap  unit_cap_1537
timestamp 1662145021
transform 1 0 92510 0 1 92510
box 0 0 3190 3190
use unit_cap  unit_cap_1538
timestamp 1662145021
transform 1 0 92510 0 1 95700
box 0 0 3190 3190
use unit_cap  unit_cap_1539
timestamp 1662145021
transform 1 0 92510 0 1 98890
box 0 0 3190 3190
use unit_cap  unit_cap_1540
timestamp 1662145021
transform 1 0 92510 0 1 102080
box 0 0 3190 3190
use unit_cap  unit_cap_1541
timestamp 1662145021
transform 1 0 92510 0 1 105270
box 0 0 3190 3190
use unit_cap  unit_cap_1542
timestamp 1662145021
transform 1 0 92510 0 1 108460
box 0 0 3190 3190
use unit_cap  unit_cap_1543
timestamp 1662145021
transform 1 0 92510 0 1 111650
box 0 0 3190 3190
use unit_cap  unit_cap_1544
timestamp 1662145021
transform 1 0 92510 0 1 114840
box 0 0 3190 3190
use unit_cap  unit_cap_1545
timestamp 1662145021
transform 1 0 92510 0 1 118030
box 0 0 3190 3190
use unit_cap  unit_cap_1546
timestamp 1662145021
transform 1 0 92510 0 1 121220
box 0 0 3190 3190
use unit_cap  unit_cap_1547
timestamp 1662145021
transform 1 0 92510 0 1 124410
box 0 0 3190 3190
use unit_cap  unit_cap_1548
timestamp 1662145021
transform 1 0 92510 0 1 127600
box 0 0 3190 3190
use unit_cap  unit_cap_1549
timestamp 1662145021
transform 1 0 92510 0 1 130790
box 0 0 3190 3190
use unit_cap  unit_cap_1550
timestamp 1662145021
transform 1 0 92510 0 1 133980
box 0 0 3190 3190
use unit_cap  unit_cap_1551
timestamp 1662145021
transform 1 0 92510 0 1 137170
box 0 0 3190 3190
use unit_cap  unit_cap_1552
timestamp 1662145021
transform 1 0 92510 0 1 140360
box 0 0 3190 3190
use unit_cap  unit_cap_1553
timestamp 1662145021
transform 1 0 92510 0 1 143550
box 0 0 3190 3190
use unit_cap  unit_cap_1554
timestamp 1662145021
transform 1 0 92510 0 1 146740
box 0 0 3190 3190
use unit_cap  unit_cap_1555
timestamp 1662145021
transform 1 0 92510 0 1 149930
box 0 0 3190 3190
use unit_cap  unit_cap_1556
timestamp 1662145021
transform 1 0 92510 0 1 153120
box 0 0 3190 3190
use unit_cap  unit_cap_1557
timestamp 1662145021
transform 1 0 92510 0 1 156310
box 0 0 3190 3190
use unit_cap  unit_cap_1558
timestamp 1662145021
transform 1 0 92510 0 1 159500
box 0 0 3190 3190
use unit_cap  unit_cap_1559
timestamp 1662145021
transform 1 0 92510 0 1 162690
box 0 0 3190 3190
use unit_cap  unit_cap_1560
timestamp 1662145021
transform 1 0 95700 0 1 0
box 0 0 3190 3190
use unit_cap  unit_cap_1561
timestamp 1662145021
transform 1 0 95700 0 1 3190
box 0 0 3190 3190
use unit_cap  unit_cap_1562
timestamp 1662145021
transform 1 0 95700 0 1 6380
box 0 0 3190 3190
use unit_cap  unit_cap_1563
timestamp 1662145021
transform 1 0 95700 0 1 9570
box 0 0 3190 3190
use unit_cap  unit_cap_1564
timestamp 1662145021
transform 1 0 95700 0 1 12760
box 0 0 3190 3190
use unit_cap  unit_cap_1565
timestamp 1662145021
transform 1 0 95700 0 1 15950
box 0 0 3190 3190
use unit_cap  unit_cap_1566
timestamp 1662145021
transform 1 0 95700 0 1 19140
box 0 0 3190 3190
use unit_cap  unit_cap_1567
timestamp 1662145021
transform 1 0 95700 0 1 22330
box 0 0 3190 3190
use unit_cap  unit_cap_1568
timestamp 1662145021
transform 1 0 95700 0 1 25520
box 0 0 3190 3190
use unit_cap  unit_cap_1569
timestamp 1662145021
transform 1 0 95700 0 1 28710
box 0 0 3190 3190
use unit_cap  unit_cap_1570
timestamp 1662145021
transform 1 0 95700 0 1 31900
box 0 0 3190 3190
use unit_cap  unit_cap_1571
timestamp 1662145021
transform 1 0 95700 0 1 35090
box 0 0 3190 3190
use unit_cap  unit_cap_1572
timestamp 1662145021
transform 1 0 95700 0 1 38280
box 0 0 3190 3190
use unit_cap  unit_cap_1573
timestamp 1662145021
transform 1 0 95700 0 1 41470
box 0 0 3190 3190
use unit_cap  unit_cap_1574
timestamp 1662145021
transform 1 0 95700 0 1 44660
box 0 0 3190 3190
use unit_cap  unit_cap_1575
timestamp 1662145021
transform 1 0 95700 0 1 47850
box 0 0 3190 3190
use unit_cap  unit_cap_1576
timestamp 1662145021
transform 1 0 95700 0 1 51040
box 0 0 3190 3190
use unit_cap  unit_cap_1577
timestamp 1662145021
transform 1 0 95700 0 1 54230
box 0 0 3190 3190
use unit_cap  unit_cap_1578
timestamp 1662145021
transform 1 0 95700 0 1 57420
box 0 0 3190 3190
use unit_cap  unit_cap_1579
timestamp 1662145021
transform 1 0 95700 0 1 60610
box 0 0 3190 3190
use unit_cap  unit_cap_1580
timestamp 1662145021
transform 1 0 95700 0 1 63800
box 0 0 3190 3190
use unit_cap  unit_cap_1581
timestamp 1662145021
transform 1 0 95700 0 1 66990
box 0 0 3190 3190
use unit_cap  unit_cap_1582
timestamp 1662145021
transform 1 0 95700 0 1 70180
box 0 0 3190 3190
use unit_cap  unit_cap_1583
timestamp 1662145021
transform 1 0 95700 0 1 73370
box 0 0 3190 3190
use unit_cap  unit_cap_1584
timestamp 1662145021
transform 1 0 95700 0 1 76560
box 0 0 3190 3190
use unit_cap  unit_cap_1585
timestamp 1662145021
transform 1 0 95700 0 1 79750
box 0 0 3190 3190
use unit_cap  unit_cap_1586
timestamp 1662145021
transform 1 0 95700 0 1 82940
box 0 0 3190 3190
use unit_cap  unit_cap_1587
timestamp 1662145021
transform 1 0 95700 0 1 86130
box 0 0 3190 3190
use unit_cap  unit_cap_1588
timestamp 1662145021
transform 1 0 95700 0 1 89320
box 0 0 3190 3190
use unit_cap  unit_cap_1589
timestamp 1662145021
transform 1 0 95700 0 1 92510
box 0 0 3190 3190
use unit_cap  unit_cap_1590
timestamp 1662145021
transform 1 0 95700 0 1 95700
box 0 0 3190 3190
use unit_cap  unit_cap_1591
timestamp 1662145021
transform 1 0 95700 0 1 98890
box 0 0 3190 3190
use unit_cap  unit_cap_1592
timestamp 1662145021
transform 1 0 95700 0 1 102080
box 0 0 3190 3190
use unit_cap  unit_cap_1593
timestamp 1662145021
transform 1 0 95700 0 1 105270
box 0 0 3190 3190
use unit_cap  unit_cap_1594
timestamp 1662145021
transform 1 0 95700 0 1 108460
box 0 0 3190 3190
use unit_cap  unit_cap_1595
timestamp 1662145021
transform 1 0 95700 0 1 111650
box 0 0 3190 3190
use unit_cap  unit_cap_1596
timestamp 1662145021
transform 1 0 95700 0 1 114840
box 0 0 3190 3190
use unit_cap  unit_cap_1597
timestamp 1662145021
transform 1 0 95700 0 1 118030
box 0 0 3190 3190
use unit_cap  unit_cap_1598
timestamp 1662145021
transform 1 0 95700 0 1 121220
box 0 0 3190 3190
use unit_cap  unit_cap_1599
timestamp 1662145021
transform 1 0 95700 0 1 124410
box 0 0 3190 3190
use unit_cap  unit_cap_1600
timestamp 1662145021
transform 1 0 95700 0 1 127600
box 0 0 3190 3190
use unit_cap  unit_cap_1601
timestamp 1662145021
transform 1 0 95700 0 1 130790
box 0 0 3190 3190
use unit_cap  unit_cap_1602
timestamp 1662145021
transform 1 0 95700 0 1 133980
box 0 0 3190 3190
use unit_cap  unit_cap_1603
timestamp 1662145021
transform 1 0 95700 0 1 137170
box 0 0 3190 3190
use unit_cap  unit_cap_1604
timestamp 1662145021
transform 1 0 95700 0 1 140360
box 0 0 3190 3190
use unit_cap  unit_cap_1605
timestamp 1662145021
transform 1 0 95700 0 1 143550
box 0 0 3190 3190
use unit_cap  unit_cap_1606
timestamp 1662145021
transform 1 0 95700 0 1 146740
box 0 0 3190 3190
use unit_cap  unit_cap_1607
timestamp 1662145021
transform 1 0 95700 0 1 149930
box 0 0 3190 3190
use unit_cap  unit_cap_1608
timestamp 1662145021
transform 1 0 95700 0 1 153120
box 0 0 3190 3190
use unit_cap  unit_cap_1609
timestamp 1662145021
transform 1 0 95700 0 1 156310
box 0 0 3190 3190
use unit_cap  unit_cap_1610
timestamp 1662145021
transform 1 0 95700 0 1 159500
box 0 0 3190 3190
use unit_cap  unit_cap_1611
timestamp 1662145021
transform 1 0 95700 0 1 162690
box 0 0 3190 3190
use unit_cap  unit_cap_1612
timestamp 1662145021
transform 1 0 98890 0 1 0
box 0 0 3190 3190
use unit_cap  unit_cap_1613
timestamp 1662145021
transform 1 0 98890 0 1 3190
box 0 0 3190 3190
use unit_cap  unit_cap_1614
timestamp 1662145021
transform 1 0 98890 0 1 6380
box 0 0 3190 3190
use unit_cap  unit_cap_1615
timestamp 1662145021
transform 1 0 98890 0 1 9570
box 0 0 3190 3190
use unit_cap  unit_cap_1616
timestamp 1662145021
transform 1 0 98890 0 1 12760
box 0 0 3190 3190
use unit_cap  unit_cap_1617
timestamp 1662145021
transform 1 0 98890 0 1 15950
box 0 0 3190 3190
use unit_cap  unit_cap_1618
timestamp 1662145021
transform 1 0 98890 0 1 19140
box 0 0 3190 3190
use unit_cap  unit_cap_1619
timestamp 1662145021
transform 1 0 98890 0 1 22330
box 0 0 3190 3190
use unit_cap  unit_cap_1620
timestamp 1662145021
transform 1 0 98890 0 1 25520
box 0 0 3190 3190
use unit_cap  unit_cap_1621
timestamp 1662145021
transform 1 0 98890 0 1 28710
box 0 0 3190 3190
use unit_cap  unit_cap_1622
timestamp 1662145021
transform 1 0 98890 0 1 31900
box 0 0 3190 3190
use unit_cap  unit_cap_1623
timestamp 1662145021
transform 1 0 98890 0 1 35090
box 0 0 3190 3190
use unit_cap  unit_cap_1624
timestamp 1662145021
transform 1 0 98890 0 1 38280
box 0 0 3190 3190
use unit_cap  unit_cap_1625
timestamp 1662145021
transform 1 0 98890 0 1 41470
box 0 0 3190 3190
use unit_cap  unit_cap_1626
timestamp 1662145021
transform 1 0 98890 0 1 44660
box 0 0 3190 3190
use unit_cap  unit_cap_1627
timestamp 1662145021
transform 1 0 98890 0 1 47850
box 0 0 3190 3190
use unit_cap  unit_cap_1628
timestamp 1662145021
transform 1 0 98890 0 1 51040
box 0 0 3190 3190
use unit_cap  unit_cap_1629
timestamp 1662145021
transform 1 0 98890 0 1 54230
box 0 0 3190 3190
use unit_cap  unit_cap_1630
timestamp 1662145021
transform 1 0 98890 0 1 57420
box 0 0 3190 3190
use unit_cap  unit_cap_1631
timestamp 1662145021
transform 1 0 98890 0 1 60610
box 0 0 3190 3190
use unit_cap  unit_cap_1632
timestamp 1662145021
transform 1 0 98890 0 1 63800
box 0 0 3190 3190
use unit_cap  unit_cap_1633
timestamp 1662145021
transform 1 0 98890 0 1 66990
box 0 0 3190 3190
use unit_cap  unit_cap_1634
timestamp 1662145021
transform 1 0 98890 0 1 70180
box 0 0 3190 3190
use unit_cap  unit_cap_1635
timestamp 1662145021
transform 1 0 98890 0 1 73370
box 0 0 3190 3190
use unit_cap  unit_cap_1636
timestamp 1662145021
transform 1 0 98890 0 1 76560
box 0 0 3190 3190
use unit_cap  unit_cap_1637
timestamp 1662145021
transform 1 0 98890 0 1 79750
box 0 0 3190 3190
use unit_cap  unit_cap_1638
timestamp 1662145021
transform 1 0 98890 0 1 82940
box 0 0 3190 3190
use unit_cap  unit_cap_1639
timestamp 1662145021
transform 1 0 98890 0 1 86130
box 0 0 3190 3190
use unit_cap  unit_cap_1640
timestamp 1662145021
transform 1 0 98890 0 1 89320
box 0 0 3190 3190
use unit_cap  unit_cap_1641
timestamp 1662145021
transform 1 0 98890 0 1 92510
box 0 0 3190 3190
use unit_cap  unit_cap_1642
timestamp 1662145021
transform 1 0 98890 0 1 95700
box 0 0 3190 3190
use unit_cap  unit_cap_1643
timestamp 1662145021
transform 1 0 98890 0 1 98890
box 0 0 3190 3190
use unit_cap  unit_cap_1644
timestamp 1662145021
transform 1 0 98890 0 1 102080
box 0 0 3190 3190
use unit_cap  unit_cap_1645
timestamp 1662145021
transform 1 0 98890 0 1 105270
box 0 0 3190 3190
use unit_cap  unit_cap_1646
timestamp 1662145021
transform 1 0 98890 0 1 108460
box 0 0 3190 3190
use unit_cap  unit_cap_1647
timestamp 1662145021
transform 1 0 98890 0 1 111650
box 0 0 3190 3190
use unit_cap  unit_cap_1648
timestamp 1662145021
transform 1 0 98890 0 1 114840
box 0 0 3190 3190
use unit_cap  unit_cap_1649
timestamp 1662145021
transform 1 0 98890 0 1 118030
box 0 0 3190 3190
use unit_cap  unit_cap_1650
timestamp 1662145021
transform 1 0 98890 0 1 121220
box 0 0 3190 3190
use unit_cap  unit_cap_1651
timestamp 1662145021
transform 1 0 98890 0 1 124410
box 0 0 3190 3190
use unit_cap  unit_cap_1652
timestamp 1662145021
transform 1 0 98890 0 1 127600
box 0 0 3190 3190
use unit_cap  unit_cap_1653
timestamp 1662145021
transform 1 0 98890 0 1 130790
box 0 0 3190 3190
use unit_cap  unit_cap_1654
timestamp 1662145021
transform 1 0 98890 0 1 133980
box 0 0 3190 3190
use unit_cap  unit_cap_1655
timestamp 1662145021
transform 1 0 98890 0 1 137170
box 0 0 3190 3190
use unit_cap  unit_cap_1656
timestamp 1662145021
transform 1 0 98890 0 1 140360
box 0 0 3190 3190
use unit_cap  unit_cap_1657
timestamp 1662145021
transform 1 0 98890 0 1 143550
box 0 0 3190 3190
use unit_cap  unit_cap_1658
timestamp 1662145021
transform 1 0 98890 0 1 146740
box 0 0 3190 3190
use unit_cap  unit_cap_1659
timestamp 1662145021
transform 1 0 98890 0 1 149930
box 0 0 3190 3190
use unit_cap  unit_cap_1660
timestamp 1662145021
transform 1 0 98890 0 1 153120
box 0 0 3190 3190
use unit_cap  unit_cap_1661
timestamp 1662145021
transform 1 0 98890 0 1 156310
box 0 0 3190 3190
use unit_cap  unit_cap_1662
timestamp 1662145021
transform 1 0 98890 0 1 159500
box 0 0 3190 3190
use unit_cap  unit_cap_1663
timestamp 1662145021
transform 1 0 98890 0 1 162690
box 0 0 3190 3190
use unit_cap  unit_cap_1664
timestamp 1662145021
transform 1 0 102080 0 1 0
box 0 0 3190 3190
use unit_cap  unit_cap_1665
timestamp 1662145021
transform 1 0 102080 0 1 3190
box 0 0 3190 3190
use unit_cap  unit_cap_1666
timestamp 1662145021
transform 1 0 102080 0 1 6380
box 0 0 3190 3190
use unit_cap  unit_cap_1667
timestamp 1662145021
transform 1 0 102080 0 1 9570
box 0 0 3190 3190
use unit_cap  unit_cap_1668
timestamp 1662145021
transform 1 0 102080 0 1 12760
box 0 0 3190 3190
use unit_cap  unit_cap_1669
timestamp 1662145021
transform 1 0 102080 0 1 15950
box 0 0 3190 3190
use unit_cap  unit_cap_1670
timestamp 1662145021
transform 1 0 102080 0 1 19140
box 0 0 3190 3190
use unit_cap  unit_cap_1671
timestamp 1662145021
transform 1 0 102080 0 1 22330
box 0 0 3190 3190
use unit_cap  unit_cap_1672
timestamp 1662145021
transform 1 0 102080 0 1 25520
box 0 0 3190 3190
use unit_cap  unit_cap_1673
timestamp 1662145021
transform 1 0 102080 0 1 28710
box 0 0 3190 3190
use unit_cap  unit_cap_1674
timestamp 1662145021
transform 1 0 102080 0 1 31900
box 0 0 3190 3190
use unit_cap  unit_cap_1675
timestamp 1662145021
transform 1 0 102080 0 1 35090
box 0 0 3190 3190
use unit_cap  unit_cap_1676
timestamp 1662145021
transform 1 0 102080 0 1 38280
box 0 0 3190 3190
use unit_cap  unit_cap_1677
timestamp 1662145021
transform 1 0 102080 0 1 41470
box 0 0 3190 3190
use unit_cap  unit_cap_1678
timestamp 1662145021
transform 1 0 102080 0 1 44660
box 0 0 3190 3190
use unit_cap  unit_cap_1679
timestamp 1662145021
transform 1 0 102080 0 1 47850
box 0 0 3190 3190
use unit_cap  unit_cap_1680
timestamp 1662145021
transform 1 0 102080 0 1 51040
box 0 0 3190 3190
use unit_cap  unit_cap_1681
timestamp 1662145021
transform 1 0 102080 0 1 54230
box 0 0 3190 3190
use unit_cap  unit_cap_1682
timestamp 1662145021
transform 1 0 102080 0 1 57420
box 0 0 3190 3190
use unit_cap  unit_cap_1683
timestamp 1662145021
transform 1 0 102080 0 1 60610
box 0 0 3190 3190
use unit_cap  unit_cap_1684
timestamp 1662145021
transform 1 0 102080 0 1 63800
box 0 0 3190 3190
use unit_cap  unit_cap_1685
timestamp 1662145021
transform 1 0 102080 0 1 66990
box 0 0 3190 3190
use unit_cap  unit_cap_1686
timestamp 1662145021
transform 1 0 102080 0 1 70180
box 0 0 3190 3190
use unit_cap  unit_cap_1687
timestamp 1662145021
transform 1 0 102080 0 1 73370
box 0 0 3190 3190
use unit_cap  unit_cap_1688
timestamp 1662145021
transform 1 0 102080 0 1 76560
box 0 0 3190 3190
use unit_cap  unit_cap_1689
timestamp 1662145021
transform 1 0 102080 0 1 79750
box 0 0 3190 3190
use unit_cap  unit_cap_1690
timestamp 1662145021
transform 1 0 102080 0 1 82940
box 0 0 3190 3190
use unit_cap  unit_cap_1691
timestamp 1662145021
transform 1 0 102080 0 1 86130
box 0 0 3190 3190
use unit_cap  unit_cap_1692
timestamp 1662145021
transform 1 0 102080 0 1 89320
box 0 0 3190 3190
use unit_cap  unit_cap_1693
timestamp 1662145021
transform 1 0 102080 0 1 92510
box 0 0 3190 3190
use unit_cap  unit_cap_1694
timestamp 1662145021
transform 1 0 102080 0 1 95700
box 0 0 3190 3190
use unit_cap  unit_cap_1695
timestamp 1662145021
transform 1 0 102080 0 1 98890
box 0 0 3190 3190
use unit_cap  unit_cap_1696
timestamp 1662145021
transform 1 0 102080 0 1 102080
box 0 0 3190 3190
use unit_cap  unit_cap_1697
timestamp 1662145021
transform 1 0 102080 0 1 105270
box 0 0 3190 3190
use unit_cap  unit_cap_1698
timestamp 1662145021
transform 1 0 102080 0 1 108460
box 0 0 3190 3190
use unit_cap  unit_cap_1699
timestamp 1662145021
transform 1 0 102080 0 1 111650
box 0 0 3190 3190
use unit_cap  unit_cap_1700
timestamp 1662145021
transform 1 0 102080 0 1 114840
box 0 0 3190 3190
use unit_cap  unit_cap_1701
timestamp 1662145021
transform 1 0 102080 0 1 118030
box 0 0 3190 3190
use unit_cap  unit_cap_1702
timestamp 1662145021
transform 1 0 102080 0 1 121220
box 0 0 3190 3190
use unit_cap  unit_cap_1703
timestamp 1662145021
transform 1 0 102080 0 1 124410
box 0 0 3190 3190
use unit_cap  unit_cap_1704
timestamp 1662145021
transform 1 0 102080 0 1 127600
box 0 0 3190 3190
use unit_cap  unit_cap_1705
timestamp 1662145021
transform 1 0 102080 0 1 130790
box 0 0 3190 3190
use unit_cap  unit_cap_1706
timestamp 1662145021
transform 1 0 102080 0 1 133980
box 0 0 3190 3190
use unit_cap  unit_cap_1707
timestamp 1662145021
transform 1 0 102080 0 1 137170
box 0 0 3190 3190
use unit_cap  unit_cap_1708
timestamp 1662145021
transform 1 0 102080 0 1 140360
box 0 0 3190 3190
use unit_cap  unit_cap_1709
timestamp 1662145021
transform 1 0 102080 0 1 143550
box 0 0 3190 3190
use unit_cap  unit_cap_1710
timestamp 1662145021
transform 1 0 102080 0 1 146740
box 0 0 3190 3190
use unit_cap  unit_cap_1711
timestamp 1662145021
transform 1 0 102080 0 1 149930
box 0 0 3190 3190
use unit_cap  unit_cap_1712
timestamp 1662145021
transform 1 0 102080 0 1 153120
box 0 0 3190 3190
use unit_cap  unit_cap_1713
timestamp 1662145021
transform 1 0 102080 0 1 156310
box 0 0 3190 3190
use unit_cap  unit_cap_1714
timestamp 1662145021
transform 1 0 102080 0 1 159500
box 0 0 3190 3190
use unit_cap  unit_cap_1715
timestamp 1662145021
transform 1 0 102080 0 1 162690
box 0 0 3190 3190
use unit_cap  unit_cap_1716
timestamp 1662145021
transform 1 0 105270 0 1 0
box 0 0 3190 3190
use unit_cap  unit_cap_1717
timestamp 1662145021
transform 1 0 105270 0 1 3190
box 0 0 3190 3190
use unit_cap  unit_cap_1718
timestamp 1662145021
transform 1 0 105270 0 1 6380
box 0 0 3190 3190
use unit_cap  unit_cap_1719
timestamp 1662145021
transform 1 0 105270 0 1 9570
box 0 0 3190 3190
use unit_cap  unit_cap_1720
timestamp 1662145021
transform 1 0 105270 0 1 12760
box 0 0 3190 3190
use unit_cap  unit_cap_1721
timestamp 1662145021
transform 1 0 105270 0 1 15950
box 0 0 3190 3190
use unit_cap  unit_cap_1722
timestamp 1662145021
transform 1 0 105270 0 1 19140
box 0 0 3190 3190
use unit_cap  unit_cap_1723
timestamp 1662145021
transform 1 0 105270 0 1 22330
box 0 0 3190 3190
use unit_cap  unit_cap_1724
timestamp 1662145021
transform 1 0 105270 0 1 25520
box 0 0 3190 3190
use unit_cap  unit_cap_1725
timestamp 1662145021
transform 1 0 105270 0 1 28710
box 0 0 3190 3190
use unit_cap  unit_cap_1726
timestamp 1662145021
transform 1 0 105270 0 1 31900
box 0 0 3190 3190
use unit_cap  unit_cap_1727
timestamp 1662145021
transform 1 0 105270 0 1 35090
box 0 0 3190 3190
use unit_cap  unit_cap_1728
timestamp 1662145021
transform 1 0 105270 0 1 38280
box 0 0 3190 3190
use unit_cap  unit_cap_1729
timestamp 1662145021
transform 1 0 105270 0 1 41470
box 0 0 3190 3190
use unit_cap  unit_cap_1730
timestamp 1662145021
transform 1 0 105270 0 1 44660
box 0 0 3190 3190
use unit_cap  unit_cap_1731
timestamp 1662145021
transform 1 0 105270 0 1 47850
box 0 0 3190 3190
use unit_cap  unit_cap_1732
timestamp 1662145021
transform 1 0 105270 0 1 51040
box 0 0 3190 3190
use unit_cap  unit_cap_1733
timestamp 1662145021
transform 1 0 105270 0 1 54230
box 0 0 3190 3190
use unit_cap  unit_cap_1734
timestamp 1662145021
transform 1 0 105270 0 1 57420
box 0 0 3190 3190
use unit_cap  unit_cap_1735
timestamp 1662145021
transform 1 0 105270 0 1 60610
box 0 0 3190 3190
use unit_cap  unit_cap_1736
timestamp 1662145021
transform 1 0 105270 0 1 63800
box 0 0 3190 3190
use unit_cap  unit_cap_1737
timestamp 1662145021
transform 1 0 105270 0 1 66990
box 0 0 3190 3190
use unit_cap  unit_cap_1738
timestamp 1662145021
transform 1 0 105270 0 1 70180
box 0 0 3190 3190
use unit_cap  unit_cap_1739
timestamp 1662145021
transform 1 0 105270 0 1 73370
box 0 0 3190 3190
use unit_cap  unit_cap_1740
timestamp 1662145021
transform 1 0 105270 0 1 76560
box 0 0 3190 3190
use unit_cap  unit_cap_1741
timestamp 1662145021
transform 1 0 105270 0 1 79750
box 0 0 3190 3190
use unit_cap  unit_cap_1742
timestamp 1662145021
transform 1 0 105270 0 1 82940
box 0 0 3190 3190
use unit_cap  unit_cap_1743
timestamp 1662145021
transform 1 0 105270 0 1 86130
box 0 0 3190 3190
use unit_cap  unit_cap_1744
timestamp 1662145021
transform 1 0 105270 0 1 89320
box 0 0 3190 3190
use unit_cap  unit_cap_1745
timestamp 1662145021
transform 1 0 105270 0 1 92510
box 0 0 3190 3190
use unit_cap  unit_cap_1746
timestamp 1662145021
transform 1 0 105270 0 1 95700
box 0 0 3190 3190
use unit_cap  unit_cap_1747
timestamp 1662145021
transform 1 0 105270 0 1 98890
box 0 0 3190 3190
use unit_cap  unit_cap_1748
timestamp 1662145021
transform 1 0 105270 0 1 102080
box 0 0 3190 3190
use unit_cap  unit_cap_1749
timestamp 1662145021
transform 1 0 105270 0 1 105270
box 0 0 3190 3190
use unit_cap  unit_cap_1750
timestamp 1662145021
transform 1 0 105270 0 1 108460
box 0 0 3190 3190
use unit_cap  unit_cap_1751
timestamp 1662145021
transform 1 0 105270 0 1 111650
box 0 0 3190 3190
use unit_cap  unit_cap_1752
timestamp 1662145021
transform 1 0 105270 0 1 114840
box 0 0 3190 3190
use unit_cap  unit_cap_1753
timestamp 1662145021
transform 1 0 105270 0 1 118030
box 0 0 3190 3190
use unit_cap  unit_cap_1754
timestamp 1662145021
transform 1 0 105270 0 1 121220
box 0 0 3190 3190
use unit_cap  unit_cap_1755
timestamp 1662145021
transform 1 0 105270 0 1 124410
box 0 0 3190 3190
use unit_cap  unit_cap_1756
timestamp 1662145021
transform 1 0 105270 0 1 127600
box 0 0 3190 3190
use unit_cap  unit_cap_1757
timestamp 1662145021
transform 1 0 105270 0 1 130790
box 0 0 3190 3190
use unit_cap  unit_cap_1758
timestamp 1662145021
transform 1 0 105270 0 1 133980
box 0 0 3190 3190
use unit_cap  unit_cap_1759
timestamp 1662145021
transform 1 0 105270 0 1 137170
box 0 0 3190 3190
use unit_cap  unit_cap_1760
timestamp 1662145021
transform 1 0 105270 0 1 140360
box 0 0 3190 3190
use unit_cap  unit_cap_1761
timestamp 1662145021
transform 1 0 105270 0 1 143550
box 0 0 3190 3190
use unit_cap  unit_cap_1762
timestamp 1662145021
transform 1 0 105270 0 1 146740
box 0 0 3190 3190
use unit_cap  unit_cap_1763
timestamp 1662145021
transform 1 0 105270 0 1 149930
box 0 0 3190 3190
use unit_cap  unit_cap_1764
timestamp 1662145021
transform 1 0 105270 0 1 153120
box 0 0 3190 3190
use unit_cap  unit_cap_1765
timestamp 1662145021
transform 1 0 105270 0 1 156310
box 0 0 3190 3190
use unit_cap  unit_cap_1766
timestamp 1662145021
transform 1 0 105270 0 1 159500
box 0 0 3190 3190
use unit_cap  unit_cap_1767
timestamp 1662145021
transform 1 0 105270 0 1 162690
box 0 0 3190 3190
use unit_cap  unit_cap_1768
timestamp 1662145021
transform 1 0 108460 0 1 0
box 0 0 3190 3190
use unit_cap  unit_cap_1769
timestamp 1662145021
transform 1 0 108460 0 1 3190
box 0 0 3190 3190
use unit_cap  unit_cap_1770
timestamp 1662145021
transform 1 0 108460 0 1 6380
box 0 0 3190 3190
use unit_cap  unit_cap_1771
timestamp 1662145021
transform 1 0 108460 0 1 9570
box 0 0 3190 3190
use unit_cap  unit_cap_1772
timestamp 1662145021
transform 1 0 108460 0 1 12760
box 0 0 3190 3190
use unit_cap  unit_cap_1773
timestamp 1662145021
transform 1 0 108460 0 1 15950
box 0 0 3190 3190
use unit_cap  unit_cap_1774
timestamp 1662145021
transform 1 0 108460 0 1 19140
box 0 0 3190 3190
use unit_cap  unit_cap_1775
timestamp 1662145021
transform 1 0 108460 0 1 22330
box 0 0 3190 3190
use unit_cap  unit_cap_1776
timestamp 1662145021
transform 1 0 108460 0 1 25520
box 0 0 3190 3190
use unit_cap  unit_cap_1777
timestamp 1662145021
transform 1 0 108460 0 1 28710
box 0 0 3190 3190
use unit_cap  unit_cap_1778
timestamp 1662145021
transform 1 0 108460 0 1 31900
box 0 0 3190 3190
use unit_cap  unit_cap_1779
timestamp 1662145021
transform 1 0 108460 0 1 35090
box 0 0 3190 3190
use unit_cap  unit_cap_1780
timestamp 1662145021
transform 1 0 108460 0 1 38280
box 0 0 3190 3190
use unit_cap  unit_cap_1781
timestamp 1662145021
transform 1 0 108460 0 1 41470
box 0 0 3190 3190
use unit_cap  unit_cap_1782
timestamp 1662145021
transform 1 0 108460 0 1 44660
box 0 0 3190 3190
use unit_cap  unit_cap_1783
timestamp 1662145021
transform 1 0 108460 0 1 47850
box 0 0 3190 3190
use unit_cap  unit_cap_1784
timestamp 1662145021
transform 1 0 108460 0 1 51040
box 0 0 3190 3190
use unit_cap  unit_cap_1785
timestamp 1662145021
transform 1 0 108460 0 1 54230
box 0 0 3190 3190
use unit_cap  unit_cap_1786
timestamp 1662145021
transform 1 0 108460 0 1 57420
box 0 0 3190 3190
use unit_cap  unit_cap_1787
timestamp 1662145021
transform 1 0 108460 0 1 60610
box 0 0 3190 3190
use unit_cap  unit_cap_1788
timestamp 1662145021
transform 1 0 108460 0 1 63800
box 0 0 3190 3190
use unit_cap  unit_cap_1789
timestamp 1662145021
transform 1 0 108460 0 1 66990
box 0 0 3190 3190
use unit_cap  unit_cap_1790
timestamp 1662145021
transform 1 0 108460 0 1 70180
box 0 0 3190 3190
use unit_cap  unit_cap_1791
timestamp 1662145021
transform 1 0 108460 0 1 73370
box 0 0 3190 3190
use unit_cap  unit_cap_1792
timestamp 1662145021
transform 1 0 108460 0 1 76560
box 0 0 3190 3190
use unit_cap  unit_cap_1793
timestamp 1662145021
transform 1 0 108460 0 1 79750
box 0 0 3190 3190
use unit_cap  unit_cap_1794
timestamp 1662145021
transform 1 0 108460 0 1 82940
box 0 0 3190 3190
use unit_cap  unit_cap_1795
timestamp 1662145021
transform 1 0 108460 0 1 86130
box 0 0 3190 3190
use unit_cap  unit_cap_1796
timestamp 1662145021
transform 1 0 108460 0 1 89320
box 0 0 3190 3190
use unit_cap  unit_cap_1797
timestamp 1662145021
transform 1 0 108460 0 1 92510
box 0 0 3190 3190
use unit_cap  unit_cap_1798
timestamp 1662145021
transform 1 0 108460 0 1 95700
box 0 0 3190 3190
use unit_cap  unit_cap_1799
timestamp 1662145021
transform 1 0 108460 0 1 98890
box 0 0 3190 3190
use unit_cap  unit_cap_1800
timestamp 1662145021
transform 1 0 108460 0 1 102080
box 0 0 3190 3190
use unit_cap  unit_cap_1801
timestamp 1662145021
transform 1 0 108460 0 1 105270
box 0 0 3190 3190
use unit_cap  unit_cap_1802
timestamp 1662145021
transform 1 0 108460 0 1 108460
box 0 0 3190 3190
use unit_cap  unit_cap_1803
timestamp 1662145021
transform 1 0 108460 0 1 111650
box 0 0 3190 3190
use unit_cap  unit_cap_1804
timestamp 1662145021
transform 1 0 108460 0 1 114840
box 0 0 3190 3190
use unit_cap  unit_cap_1805
timestamp 1662145021
transform 1 0 108460 0 1 118030
box 0 0 3190 3190
use unit_cap  unit_cap_1806
timestamp 1662145021
transform 1 0 108460 0 1 121220
box 0 0 3190 3190
use unit_cap  unit_cap_1807
timestamp 1662145021
transform 1 0 108460 0 1 124410
box 0 0 3190 3190
use unit_cap  unit_cap_1808
timestamp 1662145021
transform 1 0 108460 0 1 127600
box 0 0 3190 3190
use unit_cap  unit_cap_1809
timestamp 1662145021
transform 1 0 108460 0 1 130790
box 0 0 3190 3190
use unit_cap  unit_cap_1810
timestamp 1662145021
transform 1 0 108460 0 1 133980
box 0 0 3190 3190
use unit_cap  unit_cap_1811
timestamp 1662145021
transform 1 0 108460 0 1 137170
box 0 0 3190 3190
use unit_cap  unit_cap_1812
timestamp 1662145021
transform 1 0 108460 0 1 140360
box 0 0 3190 3190
use unit_cap  unit_cap_1813
timestamp 1662145021
transform 1 0 108460 0 1 143550
box 0 0 3190 3190
use unit_cap  unit_cap_1814
timestamp 1662145021
transform 1 0 108460 0 1 146740
box 0 0 3190 3190
use unit_cap  unit_cap_1815
timestamp 1662145021
transform 1 0 108460 0 1 149930
box 0 0 3190 3190
use unit_cap  unit_cap_1816
timestamp 1662145021
transform 1 0 108460 0 1 153120
box 0 0 3190 3190
use unit_cap  unit_cap_1817
timestamp 1662145021
transform 1 0 108460 0 1 156310
box 0 0 3190 3190
use unit_cap  unit_cap_1818
timestamp 1662145021
transform 1 0 108460 0 1 159500
box 0 0 3190 3190
use unit_cap  unit_cap_1819
timestamp 1662145021
transform 1 0 108460 0 1 162690
box 0 0 3190 3190
use unit_cap  unit_cap_1820
timestamp 1662145021
transform 1 0 111650 0 1 0
box 0 0 3190 3190
use unit_cap  unit_cap_1821
timestamp 1662145021
transform 1 0 111650 0 1 3190
box 0 0 3190 3190
use unit_cap  unit_cap_1822
timestamp 1662145021
transform 1 0 111650 0 1 6380
box 0 0 3190 3190
use unit_cap  unit_cap_1823
timestamp 1662145021
transform 1 0 111650 0 1 9570
box 0 0 3190 3190
use unit_cap  unit_cap_1824
timestamp 1662145021
transform 1 0 111650 0 1 12760
box 0 0 3190 3190
use unit_cap  unit_cap_1825
timestamp 1662145021
transform 1 0 111650 0 1 15950
box 0 0 3190 3190
use unit_cap  unit_cap_1826
timestamp 1662145021
transform 1 0 111650 0 1 19140
box 0 0 3190 3190
use unit_cap  unit_cap_1827
timestamp 1662145021
transform 1 0 111650 0 1 22330
box 0 0 3190 3190
use unit_cap  unit_cap_1828
timestamp 1662145021
transform 1 0 111650 0 1 25520
box 0 0 3190 3190
use unit_cap  unit_cap_1829
timestamp 1662145021
transform 1 0 111650 0 1 28710
box 0 0 3190 3190
use unit_cap  unit_cap_1830
timestamp 1662145021
transform 1 0 111650 0 1 31900
box 0 0 3190 3190
use unit_cap  unit_cap_1831
timestamp 1662145021
transform 1 0 111650 0 1 35090
box 0 0 3190 3190
use unit_cap  unit_cap_1832
timestamp 1662145021
transform 1 0 111650 0 1 38280
box 0 0 3190 3190
use unit_cap  unit_cap_1833
timestamp 1662145021
transform 1 0 111650 0 1 41470
box 0 0 3190 3190
use unit_cap  unit_cap_1834
timestamp 1662145021
transform 1 0 111650 0 1 44660
box 0 0 3190 3190
use unit_cap  unit_cap_1835
timestamp 1662145021
transform 1 0 111650 0 1 47850
box 0 0 3190 3190
use unit_cap  unit_cap_1836
timestamp 1662145021
transform 1 0 111650 0 1 51040
box 0 0 3190 3190
use unit_cap  unit_cap_1837
timestamp 1662145021
transform 1 0 111650 0 1 54230
box 0 0 3190 3190
use unit_cap  unit_cap_1838
timestamp 1662145021
transform 1 0 111650 0 1 57420
box 0 0 3190 3190
use unit_cap  unit_cap_1839
timestamp 1662145021
transform 1 0 111650 0 1 60610
box 0 0 3190 3190
use unit_cap  unit_cap_1840
timestamp 1662145021
transform 1 0 111650 0 1 63800
box 0 0 3190 3190
use unit_cap  unit_cap_1841
timestamp 1662145021
transform 1 0 111650 0 1 66990
box 0 0 3190 3190
use unit_cap  unit_cap_1842
timestamp 1662145021
transform 1 0 111650 0 1 70180
box 0 0 3190 3190
use unit_cap  unit_cap_1843
timestamp 1662145021
transform 1 0 111650 0 1 73370
box 0 0 3190 3190
use unit_cap  unit_cap_1844
timestamp 1662145021
transform 1 0 111650 0 1 76560
box 0 0 3190 3190
use unit_cap  unit_cap_1845
timestamp 1662145021
transform 1 0 111650 0 1 79750
box 0 0 3190 3190
use unit_cap  unit_cap_1846
timestamp 1662145021
transform 1 0 111650 0 1 82940
box 0 0 3190 3190
use unit_cap  unit_cap_1847
timestamp 1662145021
transform 1 0 111650 0 1 86130
box 0 0 3190 3190
use unit_cap  unit_cap_1848
timestamp 1662145021
transform 1 0 111650 0 1 89320
box 0 0 3190 3190
use unit_cap  unit_cap_1849
timestamp 1662145021
transform 1 0 111650 0 1 92510
box 0 0 3190 3190
use unit_cap  unit_cap_1850
timestamp 1662145021
transform 1 0 111650 0 1 95700
box 0 0 3190 3190
use unit_cap  unit_cap_1851
timestamp 1662145021
transform 1 0 111650 0 1 98890
box 0 0 3190 3190
use unit_cap  unit_cap_1852
timestamp 1662145021
transform 1 0 111650 0 1 102080
box 0 0 3190 3190
use unit_cap  unit_cap_1853
timestamp 1662145021
transform 1 0 111650 0 1 105270
box 0 0 3190 3190
use unit_cap  unit_cap_1854
timestamp 1662145021
transform 1 0 111650 0 1 108460
box 0 0 3190 3190
use unit_cap  unit_cap_1855
timestamp 1662145021
transform 1 0 111650 0 1 111650
box 0 0 3190 3190
use unit_cap  unit_cap_1856
timestamp 1662145021
transform 1 0 111650 0 1 114840
box 0 0 3190 3190
use unit_cap  unit_cap_1857
timestamp 1662145021
transform 1 0 111650 0 1 118030
box 0 0 3190 3190
use unit_cap  unit_cap_1858
timestamp 1662145021
transform 1 0 111650 0 1 121220
box 0 0 3190 3190
use unit_cap  unit_cap_1859
timestamp 1662145021
transform 1 0 111650 0 1 124410
box 0 0 3190 3190
use unit_cap  unit_cap_1860
timestamp 1662145021
transform 1 0 111650 0 1 127600
box 0 0 3190 3190
use unit_cap  unit_cap_1861
timestamp 1662145021
transform 1 0 111650 0 1 130790
box 0 0 3190 3190
use unit_cap  unit_cap_1862
timestamp 1662145021
transform 1 0 111650 0 1 133980
box 0 0 3190 3190
use unit_cap  unit_cap_1863
timestamp 1662145021
transform 1 0 111650 0 1 137170
box 0 0 3190 3190
use unit_cap  unit_cap_1864
timestamp 1662145021
transform 1 0 111650 0 1 140360
box 0 0 3190 3190
use unit_cap  unit_cap_1865
timestamp 1662145021
transform 1 0 111650 0 1 143550
box 0 0 3190 3190
use unit_cap  unit_cap_1866
timestamp 1662145021
transform 1 0 111650 0 1 146740
box 0 0 3190 3190
use unit_cap  unit_cap_1867
timestamp 1662145021
transform 1 0 111650 0 1 149930
box 0 0 3190 3190
use unit_cap  unit_cap_1868
timestamp 1662145021
transform 1 0 111650 0 1 153120
box 0 0 3190 3190
use unit_cap  unit_cap_1869
timestamp 1662145021
transform 1 0 111650 0 1 156310
box 0 0 3190 3190
use unit_cap  unit_cap_1870
timestamp 1662145021
transform 1 0 111650 0 1 159500
box 0 0 3190 3190
use unit_cap  unit_cap_1871
timestamp 1662145021
transform 1 0 111650 0 1 162690
box 0 0 3190 3190
use unit_cap  unit_cap_1872
timestamp 1662145021
transform 1 0 114840 0 1 0
box 0 0 3190 3190
use unit_cap  unit_cap_1873
timestamp 1662145021
transform 1 0 114840 0 1 3190
box 0 0 3190 3190
use unit_cap  unit_cap_1874
timestamp 1662145021
transform 1 0 114840 0 1 6380
box 0 0 3190 3190
use unit_cap  unit_cap_1875
timestamp 1662145021
transform 1 0 114840 0 1 9570
box 0 0 3190 3190
use unit_cap  unit_cap_1876
timestamp 1662145021
transform 1 0 114840 0 1 12760
box 0 0 3190 3190
use unit_cap  unit_cap_1877
timestamp 1662145021
transform 1 0 114840 0 1 15950
box 0 0 3190 3190
use unit_cap  unit_cap_1878
timestamp 1662145021
transform 1 0 114840 0 1 19140
box 0 0 3190 3190
use unit_cap  unit_cap_1879
timestamp 1662145021
transform 1 0 114840 0 1 22330
box 0 0 3190 3190
use unit_cap  unit_cap_1880
timestamp 1662145021
transform 1 0 114840 0 1 25520
box 0 0 3190 3190
use unit_cap  unit_cap_1881
timestamp 1662145021
transform 1 0 114840 0 1 28710
box 0 0 3190 3190
use unit_cap  unit_cap_1882
timestamp 1662145021
transform 1 0 114840 0 1 31900
box 0 0 3190 3190
use unit_cap  unit_cap_1883
timestamp 1662145021
transform 1 0 114840 0 1 35090
box 0 0 3190 3190
use unit_cap  unit_cap_1884
timestamp 1662145021
transform 1 0 114840 0 1 38280
box 0 0 3190 3190
use unit_cap  unit_cap_1885
timestamp 1662145021
transform 1 0 114840 0 1 41470
box 0 0 3190 3190
use unit_cap  unit_cap_1886
timestamp 1662145021
transform 1 0 114840 0 1 44660
box 0 0 3190 3190
use unit_cap  unit_cap_1887
timestamp 1662145021
transform 1 0 114840 0 1 47850
box 0 0 3190 3190
use unit_cap  unit_cap_1888
timestamp 1662145021
transform 1 0 114840 0 1 51040
box 0 0 3190 3190
use unit_cap  unit_cap_1889
timestamp 1662145021
transform 1 0 114840 0 1 54230
box 0 0 3190 3190
use unit_cap  unit_cap_1890
timestamp 1662145021
transform 1 0 114840 0 1 57420
box 0 0 3190 3190
use unit_cap  unit_cap_1891
timestamp 1662145021
transform 1 0 114840 0 1 60610
box 0 0 3190 3190
use unit_cap  unit_cap_1892
timestamp 1662145021
transform 1 0 114840 0 1 63800
box 0 0 3190 3190
use unit_cap  unit_cap_1893
timestamp 1662145021
transform 1 0 114840 0 1 66990
box 0 0 3190 3190
use unit_cap  unit_cap_1894
timestamp 1662145021
transform 1 0 114840 0 1 70180
box 0 0 3190 3190
use unit_cap  unit_cap_1895
timestamp 1662145021
transform 1 0 114840 0 1 73370
box 0 0 3190 3190
use unit_cap  unit_cap_1896
timestamp 1662145021
transform 1 0 114840 0 1 76560
box 0 0 3190 3190
use unit_cap  unit_cap_1897
timestamp 1662145021
transform 1 0 114840 0 1 79750
box 0 0 3190 3190
use unit_cap  unit_cap_1898
timestamp 1662145021
transform 1 0 114840 0 1 82940
box 0 0 3190 3190
use unit_cap  unit_cap_1899
timestamp 1662145021
transform 1 0 114840 0 1 86130
box 0 0 3190 3190
use unit_cap  unit_cap_1900
timestamp 1662145021
transform 1 0 114840 0 1 89320
box 0 0 3190 3190
use unit_cap  unit_cap_1901
timestamp 1662145021
transform 1 0 114840 0 1 92510
box 0 0 3190 3190
use unit_cap  unit_cap_1902
timestamp 1662145021
transform 1 0 114840 0 1 95700
box 0 0 3190 3190
use unit_cap  unit_cap_1903
timestamp 1662145021
transform 1 0 114840 0 1 98890
box 0 0 3190 3190
use unit_cap  unit_cap_1904
timestamp 1662145021
transform 1 0 114840 0 1 102080
box 0 0 3190 3190
use unit_cap  unit_cap_1905
timestamp 1662145021
transform 1 0 114840 0 1 105270
box 0 0 3190 3190
use unit_cap  unit_cap_1906
timestamp 1662145021
transform 1 0 114840 0 1 108460
box 0 0 3190 3190
use unit_cap  unit_cap_1907
timestamp 1662145021
transform 1 0 114840 0 1 111650
box 0 0 3190 3190
use unit_cap  unit_cap_1908
timestamp 1662145021
transform 1 0 114840 0 1 114840
box 0 0 3190 3190
use unit_cap  unit_cap_1909
timestamp 1662145021
transform 1 0 114840 0 1 118030
box 0 0 3190 3190
use unit_cap  unit_cap_1910
timestamp 1662145021
transform 1 0 114840 0 1 121220
box 0 0 3190 3190
use unit_cap  unit_cap_1911
timestamp 1662145021
transform 1 0 114840 0 1 124410
box 0 0 3190 3190
use unit_cap  unit_cap_1912
timestamp 1662145021
transform 1 0 114840 0 1 127600
box 0 0 3190 3190
use unit_cap  unit_cap_1913
timestamp 1662145021
transform 1 0 114840 0 1 130790
box 0 0 3190 3190
use unit_cap  unit_cap_1914
timestamp 1662145021
transform 1 0 114840 0 1 133980
box 0 0 3190 3190
use unit_cap  unit_cap_1915
timestamp 1662145021
transform 1 0 114840 0 1 137170
box 0 0 3190 3190
use unit_cap  unit_cap_1916
timestamp 1662145021
transform 1 0 114840 0 1 140360
box 0 0 3190 3190
use unit_cap  unit_cap_1917
timestamp 1662145021
transform 1 0 114840 0 1 143550
box 0 0 3190 3190
use unit_cap  unit_cap_1918
timestamp 1662145021
transform 1 0 114840 0 1 146740
box 0 0 3190 3190
use unit_cap  unit_cap_1919
timestamp 1662145021
transform 1 0 114840 0 1 149930
box 0 0 3190 3190
use unit_cap  unit_cap_1920
timestamp 1662145021
transform 1 0 114840 0 1 153120
box 0 0 3190 3190
use unit_cap  unit_cap_1921
timestamp 1662145021
transform 1 0 114840 0 1 156310
box 0 0 3190 3190
use unit_cap  unit_cap_1922
timestamp 1662145021
transform 1 0 114840 0 1 159500
box 0 0 3190 3190
use unit_cap  unit_cap_1923
timestamp 1662145021
transform 1 0 114840 0 1 162690
box 0 0 3190 3190
use unit_cap  unit_cap_1924
timestamp 1662145021
transform 1 0 118030 0 1 0
box 0 0 3190 3190
use unit_cap  unit_cap_1925
timestamp 1662145021
transform 1 0 118030 0 1 3190
box 0 0 3190 3190
use unit_cap  unit_cap_1926
timestamp 1662145021
transform 1 0 118030 0 1 6380
box 0 0 3190 3190
use unit_cap  unit_cap_1927
timestamp 1662145021
transform 1 0 118030 0 1 9570
box 0 0 3190 3190
use unit_cap  unit_cap_1928
timestamp 1662145021
transform 1 0 118030 0 1 12760
box 0 0 3190 3190
use unit_cap  unit_cap_1929
timestamp 1662145021
transform 1 0 118030 0 1 15950
box 0 0 3190 3190
use unit_cap  unit_cap_1930
timestamp 1662145021
transform 1 0 118030 0 1 19140
box 0 0 3190 3190
use unit_cap  unit_cap_1931
timestamp 1662145021
transform 1 0 118030 0 1 22330
box 0 0 3190 3190
use unit_cap  unit_cap_1932
timestamp 1662145021
transform 1 0 118030 0 1 25520
box 0 0 3190 3190
use unit_cap  unit_cap_1933
timestamp 1662145021
transform 1 0 118030 0 1 28710
box 0 0 3190 3190
use unit_cap  unit_cap_1934
timestamp 1662145021
transform 1 0 118030 0 1 31900
box 0 0 3190 3190
use unit_cap  unit_cap_1935
timestamp 1662145021
transform 1 0 118030 0 1 35090
box 0 0 3190 3190
use unit_cap  unit_cap_1936
timestamp 1662145021
transform 1 0 118030 0 1 38280
box 0 0 3190 3190
use unit_cap  unit_cap_1937
timestamp 1662145021
transform 1 0 118030 0 1 41470
box 0 0 3190 3190
use unit_cap  unit_cap_1938
timestamp 1662145021
transform 1 0 118030 0 1 44660
box 0 0 3190 3190
use unit_cap  unit_cap_1939
timestamp 1662145021
transform 1 0 118030 0 1 47850
box 0 0 3190 3190
use unit_cap  unit_cap_1940
timestamp 1662145021
transform 1 0 118030 0 1 51040
box 0 0 3190 3190
use unit_cap  unit_cap_1941
timestamp 1662145021
transform 1 0 118030 0 1 54230
box 0 0 3190 3190
use unit_cap  unit_cap_1942
timestamp 1662145021
transform 1 0 118030 0 1 57420
box 0 0 3190 3190
use unit_cap  unit_cap_1943
timestamp 1662145021
transform 1 0 118030 0 1 60610
box 0 0 3190 3190
use unit_cap  unit_cap_1944
timestamp 1662145021
transform 1 0 118030 0 1 63800
box 0 0 3190 3190
use unit_cap  unit_cap_1945
timestamp 1662145021
transform 1 0 118030 0 1 66990
box 0 0 3190 3190
use unit_cap  unit_cap_1946
timestamp 1662145021
transform 1 0 118030 0 1 70180
box 0 0 3190 3190
use unit_cap  unit_cap_1947
timestamp 1662145021
transform 1 0 118030 0 1 73370
box 0 0 3190 3190
use unit_cap  unit_cap_1948
timestamp 1662145021
transform 1 0 118030 0 1 76560
box 0 0 3190 3190
use unit_cap  unit_cap_1949
timestamp 1662145021
transform 1 0 118030 0 1 79750
box 0 0 3190 3190
use unit_cap  unit_cap_1950
timestamp 1662145021
transform 1 0 118030 0 1 82940
box 0 0 3190 3190
use unit_cap  unit_cap_1951
timestamp 1662145021
transform 1 0 118030 0 1 86130
box 0 0 3190 3190
use unit_cap  unit_cap_1952
timestamp 1662145021
transform 1 0 118030 0 1 89320
box 0 0 3190 3190
use unit_cap  unit_cap_1953
timestamp 1662145021
transform 1 0 118030 0 1 92510
box 0 0 3190 3190
use unit_cap  unit_cap_1954
timestamp 1662145021
transform 1 0 118030 0 1 95700
box 0 0 3190 3190
use unit_cap  unit_cap_1955
timestamp 1662145021
transform 1 0 118030 0 1 98890
box 0 0 3190 3190
use unit_cap  unit_cap_1956
timestamp 1662145021
transform 1 0 118030 0 1 102080
box 0 0 3190 3190
use unit_cap  unit_cap_1957
timestamp 1662145021
transform 1 0 118030 0 1 105270
box 0 0 3190 3190
use unit_cap  unit_cap_1958
timestamp 1662145021
transform 1 0 118030 0 1 108460
box 0 0 3190 3190
use unit_cap  unit_cap_1959
timestamp 1662145021
transform 1 0 118030 0 1 111650
box 0 0 3190 3190
use unit_cap  unit_cap_1960
timestamp 1662145021
transform 1 0 118030 0 1 114840
box 0 0 3190 3190
use unit_cap  unit_cap_1961
timestamp 1662145021
transform 1 0 118030 0 1 118030
box 0 0 3190 3190
use unit_cap  unit_cap_1962
timestamp 1662145021
transform 1 0 118030 0 1 121220
box 0 0 3190 3190
use unit_cap  unit_cap_1963
timestamp 1662145021
transform 1 0 118030 0 1 124410
box 0 0 3190 3190
use unit_cap  unit_cap_1964
timestamp 1662145021
transform 1 0 118030 0 1 127600
box 0 0 3190 3190
use unit_cap  unit_cap_1965
timestamp 1662145021
transform 1 0 118030 0 1 130790
box 0 0 3190 3190
use unit_cap  unit_cap_1966
timestamp 1662145021
transform 1 0 118030 0 1 133980
box 0 0 3190 3190
use unit_cap  unit_cap_1967
timestamp 1662145021
transform 1 0 118030 0 1 137170
box 0 0 3190 3190
use unit_cap  unit_cap_1968
timestamp 1662145021
transform 1 0 118030 0 1 140360
box 0 0 3190 3190
use unit_cap  unit_cap_1969
timestamp 1662145021
transform 1 0 118030 0 1 143550
box 0 0 3190 3190
use unit_cap  unit_cap_1970
timestamp 1662145021
transform 1 0 118030 0 1 146740
box 0 0 3190 3190
use unit_cap  unit_cap_1971
timestamp 1662145021
transform 1 0 118030 0 1 149930
box 0 0 3190 3190
use unit_cap  unit_cap_1972
timestamp 1662145021
transform 1 0 118030 0 1 153120
box 0 0 3190 3190
use unit_cap  unit_cap_1973
timestamp 1662145021
transform 1 0 118030 0 1 156310
box 0 0 3190 3190
use unit_cap  unit_cap_1974
timestamp 1662145021
transform 1 0 118030 0 1 159500
box 0 0 3190 3190
use unit_cap  unit_cap_1975
timestamp 1662145021
transform 1 0 118030 0 1 162690
box 0 0 3190 3190
use unit_cap  unit_cap_1976
timestamp 1662145021
transform 1 0 121220 0 1 0
box 0 0 3190 3190
use unit_cap  unit_cap_1977
timestamp 1662145021
transform 1 0 121220 0 1 3190
box 0 0 3190 3190
use unit_cap  unit_cap_1978
timestamp 1662145021
transform 1 0 121220 0 1 6380
box 0 0 3190 3190
use unit_cap  unit_cap_1979
timestamp 1662145021
transform 1 0 121220 0 1 9570
box 0 0 3190 3190
use unit_cap  unit_cap_1980
timestamp 1662145021
transform 1 0 121220 0 1 12760
box 0 0 3190 3190
use unit_cap  unit_cap_1981
timestamp 1662145021
transform 1 0 121220 0 1 15950
box 0 0 3190 3190
use unit_cap  unit_cap_1982
timestamp 1662145021
transform 1 0 121220 0 1 19140
box 0 0 3190 3190
use unit_cap  unit_cap_1983
timestamp 1662145021
transform 1 0 121220 0 1 22330
box 0 0 3190 3190
use unit_cap  unit_cap_1984
timestamp 1662145021
transform 1 0 121220 0 1 25520
box 0 0 3190 3190
use unit_cap  unit_cap_1985
timestamp 1662145021
transform 1 0 121220 0 1 28710
box 0 0 3190 3190
use unit_cap  unit_cap_1986
timestamp 1662145021
transform 1 0 121220 0 1 31900
box 0 0 3190 3190
use unit_cap  unit_cap_1987
timestamp 1662145021
transform 1 0 121220 0 1 35090
box 0 0 3190 3190
use unit_cap  unit_cap_1988
timestamp 1662145021
transform 1 0 121220 0 1 38280
box 0 0 3190 3190
use unit_cap  unit_cap_1989
timestamp 1662145021
transform 1 0 121220 0 1 41470
box 0 0 3190 3190
use unit_cap  unit_cap_1990
timestamp 1662145021
transform 1 0 121220 0 1 44660
box 0 0 3190 3190
use unit_cap  unit_cap_1991
timestamp 1662145021
transform 1 0 121220 0 1 47850
box 0 0 3190 3190
use unit_cap  unit_cap_1992
timestamp 1662145021
transform 1 0 121220 0 1 51040
box 0 0 3190 3190
use unit_cap  unit_cap_1993
timestamp 1662145021
transform 1 0 121220 0 1 54230
box 0 0 3190 3190
use unit_cap  unit_cap_1994
timestamp 1662145021
transform 1 0 121220 0 1 57420
box 0 0 3190 3190
use unit_cap  unit_cap_1995
timestamp 1662145021
transform 1 0 121220 0 1 60610
box 0 0 3190 3190
use unit_cap  unit_cap_1996
timestamp 1662145021
transform 1 0 121220 0 1 63800
box 0 0 3190 3190
use unit_cap  unit_cap_1997
timestamp 1662145021
transform 1 0 121220 0 1 66990
box 0 0 3190 3190
use unit_cap  unit_cap_1998
timestamp 1662145021
transform 1 0 121220 0 1 70180
box 0 0 3190 3190
use unit_cap  unit_cap_1999
timestamp 1662145021
transform 1 0 121220 0 1 73370
box 0 0 3190 3190
use unit_cap  unit_cap_2000
timestamp 1662145021
transform 1 0 121220 0 1 76560
box 0 0 3190 3190
use unit_cap  unit_cap_2001
timestamp 1662145021
transform 1 0 121220 0 1 79750
box 0 0 3190 3190
use unit_cap  unit_cap_2002
timestamp 1662145021
transform 1 0 121220 0 1 82940
box 0 0 3190 3190
use unit_cap  unit_cap_2003
timestamp 1662145021
transform 1 0 121220 0 1 86130
box 0 0 3190 3190
use unit_cap  unit_cap_2004
timestamp 1662145021
transform 1 0 121220 0 1 89320
box 0 0 3190 3190
use unit_cap  unit_cap_2005
timestamp 1662145021
transform 1 0 121220 0 1 92510
box 0 0 3190 3190
use unit_cap  unit_cap_2006
timestamp 1662145021
transform 1 0 121220 0 1 95700
box 0 0 3190 3190
use unit_cap  unit_cap_2007
timestamp 1662145021
transform 1 0 121220 0 1 98890
box 0 0 3190 3190
use unit_cap  unit_cap_2008
timestamp 1662145021
transform 1 0 121220 0 1 102080
box 0 0 3190 3190
use unit_cap  unit_cap_2009
timestamp 1662145021
transform 1 0 121220 0 1 105270
box 0 0 3190 3190
use unit_cap  unit_cap_2010
timestamp 1662145021
transform 1 0 121220 0 1 108460
box 0 0 3190 3190
use unit_cap  unit_cap_2011
timestamp 1662145021
transform 1 0 121220 0 1 111650
box 0 0 3190 3190
use unit_cap  unit_cap_2012
timestamp 1662145021
transform 1 0 121220 0 1 114840
box 0 0 3190 3190
use unit_cap  unit_cap_2013
timestamp 1662145021
transform 1 0 121220 0 1 118030
box 0 0 3190 3190
use unit_cap  unit_cap_2014
timestamp 1662145021
transform 1 0 121220 0 1 121220
box 0 0 3190 3190
use unit_cap  unit_cap_2015
timestamp 1662145021
transform 1 0 121220 0 1 124410
box 0 0 3190 3190
use unit_cap  unit_cap_2016
timestamp 1662145021
transform 1 0 121220 0 1 127600
box 0 0 3190 3190
use unit_cap  unit_cap_2017
timestamp 1662145021
transform 1 0 121220 0 1 130790
box 0 0 3190 3190
use unit_cap  unit_cap_2018
timestamp 1662145021
transform 1 0 121220 0 1 133980
box 0 0 3190 3190
use unit_cap  unit_cap_2019
timestamp 1662145021
transform 1 0 121220 0 1 137170
box 0 0 3190 3190
use unit_cap  unit_cap_2020
timestamp 1662145021
transform 1 0 121220 0 1 140360
box 0 0 3190 3190
use unit_cap  unit_cap_2021
timestamp 1662145021
transform 1 0 121220 0 1 143550
box 0 0 3190 3190
use unit_cap  unit_cap_2022
timestamp 1662145021
transform 1 0 121220 0 1 146740
box 0 0 3190 3190
use unit_cap  unit_cap_2023
timestamp 1662145021
transform 1 0 121220 0 1 149930
box 0 0 3190 3190
use unit_cap  unit_cap_2024
timestamp 1662145021
transform 1 0 121220 0 1 153120
box 0 0 3190 3190
use unit_cap  unit_cap_2025
timestamp 1662145021
transform 1 0 121220 0 1 156310
box 0 0 3190 3190
use unit_cap  unit_cap_2026
timestamp 1662145021
transform 1 0 121220 0 1 159500
box 0 0 3190 3190
use unit_cap  unit_cap_2027
timestamp 1662145021
transform 1 0 121220 0 1 162690
box 0 0 3190 3190
use unit_cap  unit_cap_2028
timestamp 1662145021
transform 1 0 124410 0 1 0
box 0 0 3190 3190
use unit_cap  unit_cap_2029
timestamp 1662145021
transform 1 0 124410 0 1 3190
box 0 0 3190 3190
use unit_cap  unit_cap_2030
timestamp 1662145021
transform 1 0 124410 0 1 6380
box 0 0 3190 3190
use unit_cap  unit_cap_2031
timestamp 1662145021
transform 1 0 124410 0 1 9570
box 0 0 3190 3190
use unit_cap  unit_cap_2032
timestamp 1662145021
transform 1 0 124410 0 1 12760
box 0 0 3190 3190
use unit_cap  unit_cap_2033
timestamp 1662145021
transform 1 0 124410 0 1 15950
box 0 0 3190 3190
use unit_cap  unit_cap_2034
timestamp 1662145021
transform 1 0 124410 0 1 19140
box 0 0 3190 3190
use unit_cap  unit_cap_2035
timestamp 1662145021
transform 1 0 124410 0 1 22330
box 0 0 3190 3190
use unit_cap  unit_cap_2036
timestamp 1662145021
transform 1 0 124410 0 1 25520
box 0 0 3190 3190
use unit_cap  unit_cap_2037
timestamp 1662145021
transform 1 0 124410 0 1 28710
box 0 0 3190 3190
use unit_cap  unit_cap_2038
timestamp 1662145021
transform 1 0 124410 0 1 31900
box 0 0 3190 3190
use unit_cap  unit_cap_2039
timestamp 1662145021
transform 1 0 124410 0 1 35090
box 0 0 3190 3190
use unit_cap  unit_cap_2040
timestamp 1662145021
transform 1 0 124410 0 1 38280
box 0 0 3190 3190
use unit_cap  unit_cap_2041
timestamp 1662145021
transform 1 0 124410 0 1 41470
box 0 0 3190 3190
use unit_cap  unit_cap_2042
timestamp 1662145021
transform 1 0 124410 0 1 44660
box 0 0 3190 3190
use unit_cap  unit_cap_2043
timestamp 1662145021
transform 1 0 124410 0 1 47850
box 0 0 3190 3190
use unit_cap  unit_cap_2044
timestamp 1662145021
transform 1 0 124410 0 1 51040
box 0 0 3190 3190
use unit_cap  unit_cap_2045
timestamp 1662145021
transform 1 0 124410 0 1 54230
box 0 0 3190 3190
use unit_cap  unit_cap_2046
timestamp 1662145021
transform 1 0 124410 0 1 57420
box 0 0 3190 3190
use unit_cap  unit_cap_2047
timestamp 1662145021
transform 1 0 124410 0 1 60610
box 0 0 3190 3190
use unit_cap  unit_cap_2048
timestamp 1662145021
transform 1 0 124410 0 1 63800
box 0 0 3190 3190
use unit_cap  unit_cap_2049
timestamp 1662145021
transform 1 0 124410 0 1 66990
box 0 0 3190 3190
use unit_cap  unit_cap_2050
timestamp 1662145021
transform 1 0 124410 0 1 70180
box 0 0 3190 3190
use unit_cap  unit_cap_2051
timestamp 1662145021
transform 1 0 124410 0 1 73370
box 0 0 3190 3190
use unit_cap  unit_cap_2052
timestamp 1662145021
transform 1 0 124410 0 1 76560
box 0 0 3190 3190
use unit_cap  unit_cap_2053
timestamp 1662145021
transform 1 0 124410 0 1 79750
box 0 0 3190 3190
use unit_cap  unit_cap_2054
timestamp 1662145021
transform 1 0 124410 0 1 82940
box 0 0 3190 3190
use unit_cap  unit_cap_2055
timestamp 1662145021
transform 1 0 124410 0 1 86130
box 0 0 3190 3190
use unit_cap  unit_cap_2056
timestamp 1662145021
transform 1 0 124410 0 1 89320
box 0 0 3190 3190
use unit_cap  unit_cap_2057
timestamp 1662145021
transform 1 0 124410 0 1 92510
box 0 0 3190 3190
use unit_cap  unit_cap_2058
timestamp 1662145021
transform 1 0 124410 0 1 95700
box 0 0 3190 3190
use unit_cap  unit_cap_2059
timestamp 1662145021
transform 1 0 124410 0 1 98890
box 0 0 3190 3190
use unit_cap  unit_cap_2060
timestamp 1662145021
transform 1 0 124410 0 1 102080
box 0 0 3190 3190
use unit_cap  unit_cap_2061
timestamp 1662145021
transform 1 0 124410 0 1 105270
box 0 0 3190 3190
use unit_cap  unit_cap_2062
timestamp 1662145021
transform 1 0 124410 0 1 108460
box 0 0 3190 3190
use unit_cap  unit_cap_2063
timestamp 1662145021
transform 1 0 124410 0 1 111650
box 0 0 3190 3190
use unit_cap  unit_cap_2064
timestamp 1662145021
transform 1 0 124410 0 1 114840
box 0 0 3190 3190
use unit_cap  unit_cap_2065
timestamp 1662145021
transform 1 0 124410 0 1 118030
box 0 0 3190 3190
use unit_cap  unit_cap_2066
timestamp 1662145021
transform 1 0 124410 0 1 121220
box 0 0 3190 3190
use unit_cap  unit_cap_2067
timestamp 1662145021
transform 1 0 124410 0 1 124410
box 0 0 3190 3190
use unit_cap  unit_cap_2068
timestamp 1662145021
transform 1 0 124410 0 1 127600
box 0 0 3190 3190
use unit_cap  unit_cap_2069
timestamp 1662145021
transform 1 0 124410 0 1 130790
box 0 0 3190 3190
use unit_cap  unit_cap_2070
timestamp 1662145021
transform 1 0 124410 0 1 133980
box 0 0 3190 3190
use unit_cap  unit_cap_2071
timestamp 1662145021
transform 1 0 124410 0 1 137170
box 0 0 3190 3190
use unit_cap  unit_cap_2072
timestamp 1662145021
transform 1 0 124410 0 1 140360
box 0 0 3190 3190
use unit_cap  unit_cap_2073
timestamp 1662145021
transform 1 0 124410 0 1 143550
box 0 0 3190 3190
use unit_cap  unit_cap_2074
timestamp 1662145021
transform 1 0 124410 0 1 146740
box 0 0 3190 3190
use unit_cap  unit_cap_2075
timestamp 1662145021
transform 1 0 124410 0 1 149930
box 0 0 3190 3190
use unit_cap  unit_cap_2076
timestamp 1662145021
transform 1 0 124410 0 1 153120
box 0 0 3190 3190
use unit_cap  unit_cap_2077
timestamp 1662145021
transform 1 0 124410 0 1 156310
box 0 0 3190 3190
use unit_cap  unit_cap_2078
timestamp 1662145021
transform 1 0 124410 0 1 159500
box 0 0 3190 3190
use unit_cap  unit_cap_2079
timestamp 1662145021
transform 1 0 124410 0 1 162690
box 0 0 3190 3190
use unit_cap  unit_cap_2080
timestamp 1662145021
transform 1 0 127600 0 1 0
box 0 0 3190 3190
use unit_cap  unit_cap_2081
timestamp 1662145021
transform 1 0 127600 0 1 3190
box 0 0 3190 3190
use unit_cap  unit_cap_2082
timestamp 1662145021
transform 1 0 127600 0 1 6380
box 0 0 3190 3190
use unit_cap  unit_cap_2083
timestamp 1662145021
transform 1 0 127600 0 1 9570
box 0 0 3190 3190
use unit_cap  unit_cap_2084
timestamp 1662145021
transform 1 0 127600 0 1 12760
box 0 0 3190 3190
use unit_cap  unit_cap_2085
timestamp 1662145021
transform 1 0 127600 0 1 15950
box 0 0 3190 3190
use unit_cap  unit_cap_2086
timestamp 1662145021
transform 1 0 127600 0 1 19140
box 0 0 3190 3190
use unit_cap  unit_cap_2087
timestamp 1662145021
transform 1 0 127600 0 1 22330
box 0 0 3190 3190
use unit_cap  unit_cap_2088
timestamp 1662145021
transform 1 0 127600 0 1 25520
box 0 0 3190 3190
use unit_cap  unit_cap_2089
timestamp 1662145021
transform 1 0 127600 0 1 28710
box 0 0 3190 3190
use unit_cap  unit_cap_2090
timestamp 1662145021
transform 1 0 127600 0 1 31900
box 0 0 3190 3190
use unit_cap  unit_cap_2091
timestamp 1662145021
transform 1 0 127600 0 1 35090
box 0 0 3190 3190
use unit_cap  unit_cap_2092
timestamp 1662145021
transform 1 0 127600 0 1 38280
box 0 0 3190 3190
use unit_cap  unit_cap_2093
timestamp 1662145021
transform 1 0 127600 0 1 41470
box 0 0 3190 3190
use unit_cap  unit_cap_2094
timestamp 1662145021
transform 1 0 127600 0 1 44660
box 0 0 3190 3190
use unit_cap  unit_cap_2095
timestamp 1662145021
transform 1 0 127600 0 1 47850
box 0 0 3190 3190
use unit_cap  unit_cap_2096
timestamp 1662145021
transform 1 0 127600 0 1 51040
box 0 0 3190 3190
use unit_cap  unit_cap_2097
timestamp 1662145021
transform 1 0 127600 0 1 54230
box 0 0 3190 3190
use unit_cap  unit_cap_2098
timestamp 1662145021
transform 1 0 127600 0 1 57420
box 0 0 3190 3190
use unit_cap  unit_cap_2099
timestamp 1662145021
transform 1 0 127600 0 1 60610
box 0 0 3190 3190
use unit_cap  unit_cap_2100
timestamp 1662145021
transform 1 0 127600 0 1 63800
box 0 0 3190 3190
use unit_cap  unit_cap_2101
timestamp 1662145021
transform 1 0 127600 0 1 66990
box 0 0 3190 3190
use unit_cap  unit_cap_2102
timestamp 1662145021
transform 1 0 127600 0 1 70180
box 0 0 3190 3190
use unit_cap  unit_cap_2103
timestamp 1662145021
transform 1 0 127600 0 1 73370
box 0 0 3190 3190
use unit_cap  unit_cap_2104
timestamp 1662145021
transform 1 0 127600 0 1 76560
box 0 0 3190 3190
use unit_cap  unit_cap_2105
timestamp 1662145021
transform 1 0 127600 0 1 79750
box 0 0 3190 3190
use unit_cap  unit_cap_2106
timestamp 1662145021
transform 1 0 127600 0 1 82940
box 0 0 3190 3190
use unit_cap  unit_cap_2107
timestamp 1662145021
transform 1 0 127600 0 1 86130
box 0 0 3190 3190
use unit_cap  unit_cap_2108
timestamp 1662145021
transform 1 0 127600 0 1 89320
box 0 0 3190 3190
use unit_cap  unit_cap_2109
timestamp 1662145021
transform 1 0 127600 0 1 92510
box 0 0 3190 3190
use unit_cap  unit_cap_2110
timestamp 1662145021
transform 1 0 127600 0 1 95700
box 0 0 3190 3190
use unit_cap  unit_cap_2111
timestamp 1662145021
transform 1 0 127600 0 1 98890
box 0 0 3190 3190
use unit_cap  unit_cap_2112
timestamp 1662145021
transform 1 0 127600 0 1 102080
box 0 0 3190 3190
use unit_cap  unit_cap_2113
timestamp 1662145021
transform 1 0 127600 0 1 105270
box 0 0 3190 3190
use unit_cap  unit_cap_2114
timestamp 1662145021
transform 1 0 127600 0 1 108460
box 0 0 3190 3190
use unit_cap  unit_cap_2115
timestamp 1662145021
transform 1 0 127600 0 1 111650
box 0 0 3190 3190
use unit_cap  unit_cap_2116
timestamp 1662145021
transform 1 0 127600 0 1 114840
box 0 0 3190 3190
use unit_cap  unit_cap_2117
timestamp 1662145021
transform 1 0 127600 0 1 118030
box 0 0 3190 3190
use unit_cap  unit_cap_2118
timestamp 1662145021
transform 1 0 127600 0 1 121220
box 0 0 3190 3190
use unit_cap  unit_cap_2119
timestamp 1662145021
transform 1 0 127600 0 1 124410
box 0 0 3190 3190
use unit_cap  unit_cap_2120
timestamp 1662145021
transform 1 0 127600 0 1 127600
box 0 0 3190 3190
use unit_cap  unit_cap_2121
timestamp 1662145021
transform 1 0 127600 0 1 130790
box 0 0 3190 3190
use unit_cap  unit_cap_2122
timestamp 1662145021
transform 1 0 127600 0 1 133980
box 0 0 3190 3190
use unit_cap  unit_cap_2123
timestamp 1662145021
transform 1 0 127600 0 1 137170
box 0 0 3190 3190
use unit_cap  unit_cap_2124
timestamp 1662145021
transform 1 0 127600 0 1 140360
box 0 0 3190 3190
use unit_cap  unit_cap_2125
timestamp 1662145021
transform 1 0 127600 0 1 143550
box 0 0 3190 3190
use unit_cap  unit_cap_2126
timestamp 1662145021
transform 1 0 127600 0 1 146740
box 0 0 3190 3190
use unit_cap  unit_cap_2127
timestamp 1662145021
transform 1 0 127600 0 1 149930
box 0 0 3190 3190
use unit_cap  unit_cap_2128
timestamp 1662145021
transform 1 0 127600 0 1 153120
box 0 0 3190 3190
use unit_cap  unit_cap_2129
timestamp 1662145021
transform 1 0 127600 0 1 156310
box 0 0 3190 3190
use unit_cap  unit_cap_2130
timestamp 1662145021
transform 1 0 127600 0 1 159500
box 0 0 3190 3190
use unit_cap  unit_cap_2131
timestamp 1662145021
transform 1 0 127600 0 1 162690
box 0 0 3190 3190
use unit_cap  unit_cap_2132
timestamp 1662145021
transform 1 0 130790 0 1 0
box 0 0 3190 3190
use unit_cap  unit_cap_2133
timestamp 1662145021
transform 1 0 130790 0 1 3190
box 0 0 3190 3190
use unit_cap  unit_cap_2134
timestamp 1662145021
transform 1 0 130790 0 1 6380
box 0 0 3190 3190
use unit_cap  unit_cap_2135
timestamp 1662145021
transform 1 0 130790 0 1 9570
box 0 0 3190 3190
use unit_cap  unit_cap_2136
timestamp 1662145021
transform 1 0 130790 0 1 12760
box 0 0 3190 3190
use unit_cap  unit_cap_2137
timestamp 1662145021
transform 1 0 130790 0 1 15950
box 0 0 3190 3190
use unit_cap  unit_cap_2138
timestamp 1662145021
transform 1 0 130790 0 1 19140
box 0 0 3190 3190
use unit_cap  unit_cap_2139
timestamp 1662145021
transform 1 0 130790 0 1 22330
box 0 0 3190 3190
use unit_cap  unit_cap_2140
timestamp 1662145021
transform 1 0 130790 0 1 25520
box 0 0 3190 3190
use unit_cap  unit_cap_2141
timestamp 1662145021
transform 1 0 130790 0 1 28710
box 0 0 3190 3190
use unit_cap  unit_cap_2142
timestamp 1662145021
transform 1 0 130790 0 1 31900
box 0 0 3190 3190
use unit_cap  unit_cap_2143
timestamp 1662145021
transform 1 0 130790 0 1 35090
box 0 0 3190 3190
use unit_cap  unit_cap_2144
timestamp 1662145021
transform 1 0 130790 0 1 38280
box 0 0 3190 3190
use unit_cap  unit_cap_2145
timestamp 1662145021
transform 1 0 130790 0 1 41470
box 0 0 3190 3190
use unit_cap  unit_cap_2146
timestamp 1662145021
transform 1 0 130790 0 1 44660
box 0 0 3190 3190
use unit_cap  unit_cap_2147
timestamp 1662145021
transform 1 0 130790 0 1 47850
box 0 0 3190 3190
use unit_cap  unit_cap_2148
timestamp 1662145021
transform 1 0 130790 0 1 51040
box 0 0 3190 3190
use unit_cap  unit_cap_2149
timestamp 1662145021
transform 1 0 130790 0 1 54230
box 0 0 3190 3190
use unit_cap  unit_cap_2150
timestamp 1662145021
transform 1 0 130790 0 1 57420
box 0 0 3190 3190
use unit_cap  unit_cap_2151
timestamp 1662145021
transform 1 0 130790 0 1 60610
box 0 0 3190 3190
use unit_cap  unit_cap_2152
timestamp 1662145021
transform 1 0 130790 0 1 63800
box 0 0 3190 3190
use unit_cap  unit_cap_2153
timestamp 1662145021
transform 1 0 130790 0 1 66990
box 0 0 3190 3190
use unit_cap  unit_cap_2154
timestamp 1662145021
transform 1 0 130790 0 1 70180
box 0 0 3190 3190
use unit_cap  unit_cap_2155
timestamp 1662145021
transform 1 0 130790 0 1 73370
box 0 0 3190 3190
use unit_cap  unit_cap_2156
timestamp 1662145021
transform 1 0 130790 0 1 76560
box 0 0 3190 3190
use unit_cap  unit_cap_2157
timestamp 1662145021
transform 1 0 130790 0 1 79750
box 0 0 3190 3190
use unit_cap  unit_cap_2158
timestamp 1662145021
transform 1 0 130790 0 1 82940
box 0 0 3190 3190
use unit_cap  unit_cap_2159
timestamp 1662145021
transform 1 0 130790 0 1 86130
box 0 0 3190 3190
use unit_cap  unit_cap_2160
timestamp 1662145021
transform 1 0 130790 0 1 89320
box 0 0 3190 3190
use unit_cap  unit_cap_2161
timestamp 1662145021
transform 1 0 130790 0 1 92510
box 0 0 3190 3190
use unit_cap  unit_cap_2162
timestamp 1662145021
transform 1 0 130790 0 1 95700
box 0 0 3190 3190
use unit_cap  unit_cap_2163
timestamp 1662145021
transform 1 0 130790 0 1 98890
box 0 0 3190 3190
use unit_cap  unit_cap_2164
timestamp 1662145021
transform 1 0 130790 0 1 102080
box 0 0 3190 3190
use unit_cap  unit_cap_2165
timestamp 1662145021
transform 1 0 130790 0 1 105270
box 0 0 3190 3190
use unit_cap  unit_cap_2166
timestamp 1662145021
transform 1 0 130790 0 1 108460
box 0 0 3190 3190
use unit_cap  unit_cap_2167
timestamp 1662145021
transform 1 0 130790 0 1 111650
box 0 0 3190 3190
use unit_cap  unit_cap_2168
timestamp 1662145021
transform 1 0 130790 0 1 114840
box 0 0 3190 3190
use unit_cap  unit_cap_2169
timestamp 1662145021
transform 1 0 130790 0 1 118030
box 0 0 3190 3190
use unit_cap  unit_cap_2170
timestamp 1662145021
transform 1 0 130790 0 1 121220
box 0 0 3190 3190
use unit_cap  unit_cap_2171
timestamp 1662145021
transform 1 0 130790 0 1 124410
box 0 0 3190 3190
use unit_cap  unit_cap_2172
timestamp 1662145021
transform 1 0 130790 0 1 127600
box 0 0 3190 3190
use unit_cap  unit_cap_2173
timestamp 1662145021
transform 1 0 130790 0 1 130790
box 0 0 3190 3190
use unit_cap  unit_cap_2174
timestamp 1662145021
transform 1 0 130790 0 1 133980
box 0 0 3190 3190
use unit_cap  unit_cap_2175
timestamp 1662145021
transform 1 0 130790 0 1 137170
box 0 0 3190 3190
use unit_cap  unit_cap_2176
timestamp 1662145021
transform 1 0 130790 0 1 140360
box 0 0 3190 3190
use unit_cap  unit_cap_2177
timestamp 1662145021
transform 1 0 130790 0 1 143550
box 0 0 3190 3190
use unit_cap  unit_cap_2178
timestamp 1662145021
transform 1 0 130790 0 1 146740
box 0 0 3190 3190
use unit_cap  unit_cap_2179
timestamp 1662145021
transform 1 0 130790 0 1 149930
box 0 0 3190 3190
use unit_cap  unit_cap_2180
timestamp 1662145021
transform 1 0 130790 0 1 153120
box 0 0 3190 3190
use unit_cap  unit_cap_2181
timestamp 1662145021
transform 1 0 130790 0 1 156310
box 0 0 3190 3190
use unit_cap  unit_cap_2182
timestamp 1662145021
transform 1 0 130790 0 1 159500
box 0 0 3190 3190
use unit_cap  unit_cap_2183
timestamp 1662145021
transform 1 0 130790 0 1 162690
box 0 0 3190 3190
use unit_cap  unit_cap_2184
timestamp 1662145021
transform 1 0 133980 0 1 0
box 0 0 3190 3190
use unit_cap  unit_cap_2185
timestamp 1662145021
transform 1 0 133980 0 1 3190
box 0 0 3190 3190
use unit_cap  unit_cap_2186
timestamp 1662145021
transform 1 0 133980 0 1 6380
box 0 0 3190 3190
use unit_cap  unit_cap_2187
timestamp 1662145021
transform 1 0 133980 0 1 9570
box 0 0 3190 3190
use unit_cap  unit_cap_2188
timestamp 1662145021
transform 1 0 133980 0 1 12760
box 0 0 3190 3190
use unit_cap  unit_cap_2189
timestamp 1662145021
transform 1 0 133980 0 1 15950
box 0 0 3190 3190
use unit_cap  unit_cap_2190
timestamp 1662145021
transform 1 0 133980 0 1 19140
box 0 0 3190 3190
use unit_cap  unit_cap_2191
timestamp 1662145021
transform 1 0 133980 0 1 22330
box 0 0 3190 3190
use unit_cap  unit_cap_2192
timestamp 1662145021
transform 1 0 133980 0 1 25520
box 0 0 3190 3190
use unit_cap  unit_cap_2193
timestamp 1662145021
transform 1 0 133980 0 1 28710
box 0 0 3190 3190
use unit_cap  unit_cap_2194
timestamp 1662145021
transform 1 0 133980 0 1 31900
box 0 0 3190 3190
use unit_cap  unit_cap_2195
timestamp 1662145021
transform 1 0 133980 0 1 35090
box 0 0 3190 3190
use unit_cap  unit_cap_2196
timestamp 1662145021
transform 1 0 133980 0 1 38280
box 0 0 3190 3190
use unit_cap  unit_cap_2197
timestamp 1662145021
transform 1 0 133980 0 1 41470
box 0 0 3190 3190
use unit_cap  unit_cap_2198
timestamp 1662145021
transform 1 0 133980 0 1 44660
box 0 0 3190 3190
use unit_cap  unit_cap_2199
timestamp 1662145021
transform 1 0 133980 0 1 47850
box 0 0 3190 3190
use unit_cap  unit_cap_2200
timestamp 1662145021
transform 1 0 133980 0 1 51040
box 0 0 3190 3190
use unit_cap  unit_cap_2201
timestamp 1662145021
transform 1 0 133980 0 1 54230
box 0 0 3190 3190
use unit_cap  unit_cap_2202
timestamp 1662145021
transform 1 0 133980 0 1 57420
box 0 0 3190 3190
use unit_cap  unit_cap_2203
timestamp 1662145021
transform 1 0 133980 0 1 60610
box 0 0 3190 3190
use unit_cap  unit_cap_2204
timestamp 1662145021
transform 1 0 133980 0 1 63800
box 0 0 3190 3190
use unit_cap  unit_cap_2205
timestamp 1662145021
transform 1 0 133980 0 1 66990
box 0 0 3190 3190
use unit_cap  unit_cap_2206
timestamp 1662145021
transform 1 0 133980 0 1 70180
box 0 0 3190 3190
use unit_cap  unit_cap_2207
timestamp 1662145021
transform 1 0 133980 0 1 73370
box 0 0 3190 3190
use unit_cap  unit_cap_2208
timestamp 1662145021
transform 1 0 133980 0 1 76560
box 0 0 3190 3190
use unit_cap  unit_cap_2209
timestamp 1662145021
transform 1 0 133980 0 1 79750
box 0 0 3190 3190
use unit_cap  unit_cap_2210
timestamp 1662145021
transform 1 0 133980 0 1 82940
box 0 0 3190 3190
use unit_cap  unit_cap_2211
timestamp 1662145021
transform 1 0 133980 0 1 86130
box 0 0 3190 3190
use unit_cap  unit_cap_2212
timestamp 1662145021
transform 1 0 133980 0 1 89320
box 0 0 3190 3190
use unit_cap  unit_cap_2213
timestamp 1662145021
transform 1 0 133980 0 1 92510
box 0 0 3190 3190
use unit_cap  unit_cap_2214
timestamp 1662145021
transform 1 0 133980 0 1 95700
box 0 0 3190 3190
use unit_cap  unit_cap_2215
timestamp 1662145021
transform 1 0 133980 0 1 98890
box 0 0 3190 3190
use unit_cap  unit_cap_2216
timestamp 1662145021
transform 1 0 133980 0 1 102080
box 0 0 3190 3190
use unit_cap  unit_cap_2217
timestamp 1662145021
transform 1 0 133980 0 1 105270
box 0 0 3190 3190
use unit_cap  unit_cap_2218
timestamp 1662145021
transform 1 0 133980 0 1 108460
box 0 0 3190 3190
use unit_cap  unit_cap_2219
timestamp 1662145021
transform 1 0 133980 0 1 111650
box 0 0 3190 3190
use unit_cap  unit_cap_2220
timestamp 1662145021
transform 1 0 133980 0 1 114840
box 0 0 3190 3190
use unit_cap  unit_cap_2221
timestamp 1662145021
transform 1 0 133980 0 1 118030
box 0 0 3190 3190
use unit_cap  unit_cap_2222
timestamp 1662145021
transform 1 0 133980 0 1 121220
box 0 0 3190 3190
use unit_cap  unit_cap_2223
timestamp 1662145021
transform 1 0 133980 0 1 124410
box 0 0 3190 3190
use unit_cap  unit_cap_2224
timestamp 1662145021
transform 1 0 133980 0 1 127600
box 0 0 3190 3190
use unit_cap  unit_cap_2225
timestamp 1662145021
transform 1 0 133980 0 1 130790
box 0 0 3190 3190
use unit_cap  unit_cap_2226
timestamp 1662145021
transform 1 0 133980 0 1 133980
box 0 0 3190 3190
use unit_cap  unit_cap_2227
timestamp 1662145021
transform 1 0 133980 0 1 137170
box 0 0 3190 3190
use unit_cap  unit_cap_2228
timestamp 1662145021
transform 1 0 133980 0 1 140360
box 0 0 3190 3190
use unit_cap  unit_cap_2229
timestamp 1662145021
transform 1 0 133980 0 1 143550
box 0 0 3190 3190
use unit_cap  unit_cap_2230
timestamp 1662145021
transform 1 0 133980 0 1 146740
box 0 0 3190 3190
use unit_cap  unit_cap_2231
timestamp 1662145021
transform 1 0 133980 0 1 149930
box 0 0 3190 3190
use unit_cap  unit_cap_2232
timestamp 1662145021
transform 1 0 133980 0 1 153120
box 0 0 3190 3190
use unit_cap  unit_cap_2233
timestamp 1662145021
transform 1 0 133980 0 1 156310
box 0 0 3190 3190
use unit_cap  unit_cap_2234
timestamp 1662145021
transform 1 0 133980 0 1 159500
box 0 0 3190 3190
use unit_cap  unit_cap_2235
timestamp 1662145021
transform 1 0 133980 0 1 162690
box 0 0 3190 3190
<< end >>
