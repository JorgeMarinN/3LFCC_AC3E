magic
tech sky130A
timestamp 1666362992
<< checkpaint >>
rect -1966 39166 139136 209966
rect -1966 -1966 139166 39166
<< metal3 >>
rect 7000 36000 56000 41000
rect 7000 33000 7100 36000
rect 55900 33000 56000 36000
<< via3 >>
rect 7100 33000 55900 36000
rect 69100 33000 129900 36000
<< metal4 >>
rect 69000 36000 130000 41000
rect 69000 33000 69100 36000
rect 129900 33000 130000 36000
<< via4 >>
rect 7100 33000 55900 36000
rect 69100 33000 129900 36000
<< metal5 >>
rect 7000 36000 56000 41000
rect 7000 33000 7100 36000
rect 55900 33000 56000 36000
use flying_cap  flying_cap_0
timestamp 1665353312
transform -1 0 137170 0 -1 208000
box 0 0 137170 168000
use power_stage  power_stage_0
timestamp 1663434482
transform 0 1 0 -1 0 37200
box 0 0 37200 137200
<< end >>
