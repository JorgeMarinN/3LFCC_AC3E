magic
tech sky130A
timestamp 1668294652
<< metal5 >>
rect 19600 27400 20900 27500
rect 19200 27300 21200 27400
rect 18900 27200 21500 27300
rect 18700 27100 21700 27200
rect 18500 27000 21900 27100
rect 18400 26900 22000 27000
rect 18200 26800 22100 26900
rect 18100 26700 22200 26800
rect 17900 26600 22300 26700
rect 17800 26500 22400 26600
rect 17700 26400 22500 26500
rect 17600 26300 22500 26400
rect 17500 26200 22600 26300
rect 17400 26100 22700 26200
rect 17300 26000 22700 26100
rect 17200 25900 22800 26000
rect 17200 25800 22900 25900
rect 17100 25700 22900 25800
rect 17000 25500 23000 25700
rect 16900 25300 23100 25500
rect 16800 25200 23200 25300
rect 16700 25100 23200 25200
rect 16600 24900 23300 25100
rect 16500 24800 23400 24900
rect 16400 24700 23400 24800
rect 16300 24500 23500 24700
rect 16200 24300 23600 24500
rect 16100 24200 23700 24300
rect 16000 24100 23700 24200
rect 16000 24000 23800 24100
rect 15900 23900 19300 24000
rect 19900 23900 23800 24000
rect 15900 23800 19000 23900
rect 20200 23800 23900 23900
rect 15800 23700 18700 23800
rect 20500 23700 23900 23800
rect 15700 23600 18500 23700
rect 20700 23600 24000 23700
rect 15700 23500 18300 23600
rect 20900 23500 24000 23600
rect 15600 23400 18200 23500
rect 21100 23400 24100 23500
rect 15500 23300 18000 23400
rect 21200 23300 24100 23400
rect 15400 23200 17900 23300
rect 21300 23200 24200 23300
rect 15400 23100 17700 23200
rect 21400 23100 24200 23200
rect 15300 23000 17600 23100
rect 21500 23000 24300 23100
rect 15200 22900 17500 23000
rect 21600 22900 24300 23000
rect 15200 22800 17400 22900
rect 21600 22800 24400 22900
rect 15100 22700 17300 22800
rect 21700 22700 24400 22800
rect 15000 22600 17200 22700
rect 21800 22600 24500 22700
rect 15000 22500 17100 22600
rect 21900 22500 24500 22600
rect 2900 22400 4200 22500
rect 14900 22400 17100 22500
rect 2600 22300 4600 22400
rect 14900 22300 17000 22400
rect 22000 22300 24600 22500
rect 2300 22200 4800 22300
rect 14800 22200 16900 22300
rect 22100 22200 24600 22300
rect 2100 22100 5000 22200
rect 14700 22100 16800 22200
rect 22200 22100 24700 22200
rect 1900 22000 3100 22100
rect 3700 22000 5300 22100
rect 14700 22000 16700 22100
rect 1700 21900 2900 22000
rect 4100 21900 5500 22000
rect 14600 21900 16700 22000
rect 22300 22000 24700 22100
rect 22300 21900 24800 22000
rect 1600 21800 2700 21900
rect 4300 21800 5700 21900
rect 14500 21800 16600 21900
rect 22400 21800 24800 21900
rect 1600 21700 2500 21800
rect 4500 21700 5900 21800
rect 14500 21700 16500 21800
rect 22500 21700 24900 21800
rect 1600 21600 2400 21700
rect 4600 21600 6000 21700
rect 14400 21600 16400 21700
rect 22600 21600 24900 21700
rect 1700 21500 2200 21600
rect 4800 21500 6200 21600
rect 14300 21500 16400 21600
rect 4900 21400 6300 21500
rect 14200 21400 16300 21500
rect 22700 21400 25000 21600
rect 5100 21300 6400 21400
rect 5200 21200 6600 21300
rect 14100 21200 16200 21400
rect 22800 21300 25100 21400
rect 22900 21200 25100 21300
rect 5300 21100 6700 21200
rect 14000 21100 16100 21200
rect 5400 21000 6800 21100
rect 5500 20900 6900 21000
rect 13900 20900 16000 21100
rect 23000 21000 25200 21200
rect 23100 20900 25300 21000
rect 5600 20800 7100 20900
rect 13800 20800 15900 20900
rect 23200 20800 25300 20900
rect 5700 20700 7200 20800
rect 13700 20700 15900 20800
rect 23300 20700 25400 20800
rect 5700 20600 7300 20700
rect 13700 20600 15800 20700
rect 23400 20600 25400 20700
rect 5800 20500 7400 20600
rect 13600 20500 15800 20600
rect 5900 20400 7600 20500
rect 6000 20300 7700 20400
rect 13500 20300 15700 20500
rect 23500 20400 25500 20600
rect 23600 20300 25600 20400
rect 6100 20200 7800 20300
rect 13400 20200 15600 20300
rect 23700 20200 25600 20300
rect 6100 20100 7900 20200
rect 13300 20100 15600 20200
rect 23800 20100 25700 20200
rect 6200 20000 8000 20100
rect 13300 20000 15500 20100
rect 23900 20000 25700 20100
rect 6300 19900 8100 20000
rect 13200 19900 15500 20000
rect 24000 19900 25800 20000
rect 6300 19800 8200 19900
rect 13100 19800 15500 19900
rect 24100 19800 25800 19900
rect 6400 19700 8300 19800
rect 13000 19700 15400 19800
rect 24100 19700 25900 19800
rect 6500 19600 8400 19700
rect 12900 19600 15400 19700
rect 24200 19600 25900 19700
rect 6600 19500 8500 19600
rect 6600 19400 8600 19500
rect 12800 19400 15300 19600
rect 24300 19500 26000 19600
rect 24400 19400 26000 19500
rect 6700 19300 8700 19400
rect 12700 19300 15200 19400
rect 6800 19200 8800 19300
rect 12600 19200 15200 19300
rect 24500 19200 26100 19400
rect 6800 19100 8900 19200
rect 12500 19100 15100 19200
rect 24600 19100 26200 19200
rect 6900 19000 9000 19100
rect 12400 19000 15100 19100
rect 24700 19000 26200 19100
rect 7000 18900 9100 19000
rect 7000 18800 9300 18900
rect 12300 18800 15000 19000
rect 24800 18900 26300 19000
rect 24900 18800 26400 18900
rect 7100 18700 9400 18800
rect 12200 18700 14900 18800
rect 25000 18700 26400 18800
rect 7200 18600 9600 18700
rect 12100 18600 14900 18700
rect 25100 18600 26500 18700
rect 7200 18500 9700 18600
rect 12000 18500 14800 18600
rect 25100 18500 26600 18600
rect 7300 18400 9900 18500
rect 11800 18400 14800 18500
rect 25200 18400 26600 18500
rect 7300 18300 10100 18400
rect 11600 18300 14700 18400
rect 25300 18300 26700 18400
rect 7400 18200 10500 18300
rect 11400 18200 14700 18300
rect 25400 18200 26800 18300
rect 7500 18100 14700 18200
rect 25500 18100 26800 18200
rect 7500 18000 14600 18100
rect 25600 18000 26900 18100
rect 7600 17900 14600 18000
rect 25700 17900 27000 18000
rect 7700 17700 14500 17900
rect 25800 17700 27100 17900
rect 7800 17600 14500 17700
rect 25900 17600 27200 17700
rect 7900 17500 14400 17600
rect 26000 17500 27300 17600
rect 8000 17400 14400 17500
rect 26100 17400 27400 17500
rect 8000 17300 14300 17400
rect 26200 17300 27400 17400
rect 8100 17200 14300 17300
rect 26300 17200 27500 17300
rect 8100 17100 14200 17200
rect 26400 17100 27600 17200
rect 8200 17000 14200 17100
rect 26500 17000 27700 17100
rect 8300 16800 14100 17000
rect 26700 16900 27800 17000
rect 26800 16800 28000 16900
rect 8400 16700 14000 16800
rect 26900 16700 28100 16800
rect 8500 16500 13900 16700
rect 27000 16600 28300 16700
rect 27100 16500 28500 16600
rect 29500 16500 29800 16600
rect 8600 16400 13800 16500
rect 27300 16400 28800 16500
rect 29200 16400 29800 16500
rect 8700 16300 13800 16400
rect 27400 16300 29700 16400
rect 8700 16200 13700 16300
rect 27600 16200 29500 16300
rect 8800 16100 13600 16200
rect 27800 16100 29300 16200
rect 8900 16000 13600 16100
rect 28100 16000 29000 16100
rect 8900 15900 13500 16000
rect 9000 15800 13400 15900
rect 9100 15700 13400 15800
rect 9100 15600 13300 15700
rect 9200 15500 13200 15600
rect 9300 15400 13200 15500
rect 9300 15300 13100 15400
rect 9400 15200 13000 15300
rect 9500 15100 12900 15200
rect 9600 15000 12900 15100
rect 9700 14900 12800 15000
rect 9800 14800 12700 14900
rect 9900 14700 12600 14800
rect 10000 14600 12500 14700
rect 10200 14500 12300 14600
rect 10400 14400 12000 14500
rect 10600 14300 11700 14400
rect 5000 10500 6200 10600
rect 11200 10500 15800 10600
rect 18300 10500 22900 10600
rect 4900 10300 6300 10500
rect 10900 10400 16100 10500
rect 18000 10400 23200 10500
rect 10700 10300 16300 10400
rect 17800 10300 23400 10400
rect 4800 10200 6400 10300
rect 10600 10200 16400 10300
rect 17700 10200 23500 10300
rect 4700 10000 6500 10200
rect 10500 10100 16500 10200
rect 17600 10100 23600 10200
rect 4600 9800 6600 10000
rect 10400 9900 16600 10100
rect 17500 9900 23700 10100
rect 10300 9800 16700 9900
rect 4500 9700 6700 9800
rect 10300 9700 11700 9800
rect 15300 9700 16700 9800
rect 4400 9500 6800 9700
rect 10300 9600 11400 9700
rect 15600 9600 16700 9700
rect 17400 9800 23800 9900
rect 17400 9700 18800 9800
rect 22400 9700 23800 9800
rect 17400 9600 18500 9700
rect 22700 9600 23800 9700
rect 24400 9800 30500 10600
rect 4300 9400 5400 9500
rect 5800 9400 6900 9500
rect 4300 9300 5300 9400
rect 4200 9200 5300 9300
rect 5900 9300 6900 9400
rect 10200 9400 11200 9600
rect 15800 9400 16800 9600
rect 5900 9200 7000 9300
rect 4100 9000 5200 9200
rect 6000 9000 7100 9200
rect 10200 9100 11100 9400
rect 15900 9100 16800 9400
rect 4000 8900 5100 9000
rect 6100 8900 7200 9000
rect 4000 8800 5000 8900
rect 3900 8700 5000 8800
rect 6200 8800 7200 8900
rect 6200 8700 7300 8800
rect 3800 8500 4900 8700
rect 6300 8500 7400 8700
rect 3700 8400 4800 8500
rect 6400 8400 7500 8500
rect 3700 8300 4700 8400
rect 3600 8200 4700 8300
rect 6500 8300 7500 8400
rect 6500 8200 7600 8300
rect 3500 8000 4600 8200
rect 6600 8000 7700 8200
rect 3400 7900 4500 8000
rect 6700 7900 7800 8000
rect 3400 7800 4400 7900
rect 3300 7700 4400 7800
rect 6800 7800 7800 7900
rect 6800 7700 7900 7800
rect 3200 7500 4300 7700
rect 6900 7500 8000 7700
rect 3100 7400 4200 7500
rect 7000 7400 8100 7500
rect 3100 7300 4100 7400
rect 3000 7200 4100 7300
rect 7100 7300 8100 7400
rect 7100 7200 8200 7300
rect 2900 7000 4000 7200
rect 7200 7000 8300 7200
rect 2800 6900 3900 7000
rect 7300 6900 8400 7000
rect 2800 6800 3800 6900
rect 2700 6700 3800 6800
rect 7400 6800 8400 6900
rect 7400 6700 8500 6800
rect 2600 6500 3700 6700
rect 7500 6500 8600 6700
rect 2500 6300 3600 6500
rect 7600 6300 8700 6500
rect 2400 6200 8800 6300
rect 2300 6000 8900 6200
rect 10200 6000 11000 9100
rect 16000 8300 16800 9100
rect 17300 9400 18300 9600
rect 22900 9400 23900 9600
rect 17300 9100 18200 9400
rect 23000 9100 23900 9400
rect 17300 8300 18100 9100
rect 23100 8600 23900 9100
rect 23000 8400 23900 8600
rect 22900 8300 23800 8400
rect 22800 8200 23800 8300
rect 22600 8100 23800 8200
rect 22400 8000 23700 8100
rect 19600 7900 23700 8000
rect 24400 8000 25200 9800
rect 19600 7800 23600 7900
rect 19600 7700 23500 7800
rect 19600 7400 23300 7700
rect 19600 7300 23500 7400
rect 19600 7200 23600 7300
rect 24400 7200 30500 8000
rect 22600 7100 23700 7200
rect 22800 7000 23700 7100
rect 22900 6900 23800 7000
rect 16000 6000 16800 6800
rect 2200 5800 9000 6000
rect 2100 5700 9100 5800
rect 10200 5700 11100 6000
rect 15900 5700 16800 6000
rect 2000 5600 9200 5700
rect 2000 5500 3100 5600
rect 8000 5500 9200 5600
rect 10200 5500 11200 5700
rect 15800 5500 16800 5700
rect 17300 6000 18100 6800
rect 23000 6700 23800 6900
rect 23100 6000 23900 6700
rect 17300 5700 18200 6000
rect 23000 5700 23900 6000
rect 17300 5500 18300 5700
rect 22900 5500 23900 5700
rect 1900 5400 3000 5500
rect 8200 5400 9300 5500
rect 1900 5300 2900 5400
rect 1800 5200 2900 5300
rect 8300 5300 9300 5400
rect 10300 5400 11400 5500
rect 15600 5400 16700 5500
rect 10300 5300 11700 5400
rect 15300 5300 16700 5400
rect 8300 5200 9400 5300
rect 10300 5200 16700 5300
rect 17400 5400 18500 5500
rect 22700 5400 23800 5500
rect 17400 5300 18800 5400
rect 22400 5300 23800 5400
rect 17400 5200 23800 5300
rect 24400 5300 25200 7200
rect 1700 5000 2800 5200
rect 8400 5000 9500 5200
rect 10400 5000 16600 5200
rect 17500 5000 23700 5200
rect 1600 4900 2700 5000
rect 8500 4900 9600 5000
rect 10500 4900 16500 5000
rect 17600 4900 23600 5000
rect 1600 4800 2600 4900
rect 1500 4700 2600 4800
rect 8600 4800 9600 4900
rect 10600 4800 16400 4900
rect 17700 4800 23500 4900
rect 8600 4700 9700 4800
rect 10700 4700 16300 4800
rect 17800 4700 23400 4800
rect 1500 4500 2500 4700
rect 8700 4500 9700 4700
rect 10900 4600 16100 4700
rect 18000 4600 23200 4700
rect 11200 4500 15800 4600
rect 18300 4500 22900 4600
rect 24400 4500 30500 5300
<< comment >>
rect -100 32000 32100 32100
rect -100 0 0 32000
rect 32000 0 32100 32000
rect -100 -100 32100 0
<< end >>
