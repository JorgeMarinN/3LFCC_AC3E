magic
tech sky130A
magscale 1 2
timestamp 1667251862
<< metal1 >>
rect 2300 584600 16000 584800
rect 567796 584600 581496 584800
rect 2300 568890 2500 584600
rect 2300 568710 2310 568890
rect 2490 568710 2500 568890
rect 2300 568700 2500 568710
rect 4300 584300 16400 584500
rect 567396 584300 579496 584500
rect 4300 568890 4500 584300
rect 4300 568710 4310 568890
rect 4490 568710 4500 568890
rect 4300 568700 4500 568710
rect 6300 584000 16800 584200
rect 566996 584000 577496 584200
rect 6300 568890 6500 584000
rect 6300 568710 6310 568890
rect 6490 568710 6500 568890
rect 6300 568700 6500 568710
rect 8300 583700 17200 583900
rect 566596 583700 575496 583900
rect 8300 568890 8500 583700
rect 8300 568710 8310 568890
rect 8490 568710 8500 568890
rect 8300 568700 8500 568710
rect 575296 568890 575496 583700
rect 575296 568710 575306 568890
rect 575486 568710 575496 568890
rect 575296 568700 575496 568710
rect 577296 568890 577496 584000
rect 577296 568710 577306 568890
rect 577486 568710 577496 568890
rect 577296 568700 577496 568710
rect 579296 568890 579496 584300
rect 579296 568710 579306 568890
rect 579486 568710 579496 568890
rect 579296 568700 579496 568710
rect 581296 568890 581496 584600
rect 581296 568710 581306 568890
rect 581486 568710 581496 568890
rect 581296 568700 581496 568710
<< via1 >>
rect 2310 568710 2490 568890
rect 4310 568710 4490 568890
rect 6310 568710 6490 568890
rect 8310 568710 8490 568890
rect 575306 568710 575486 568890
rect 577306 568710 577486 568890
rect 579306 568710 579486 568890
rect 581306 568710 581486 568890
<< metal2 >>
rect 2300 568890 2500 568900
rect 2300 568710 2310 568890
rect 2490 568710 2500 568890
rect 2300 568700 2500 568710
rect 4300 568890 4500 568900
rect 4300 568710 4310 568890
rect 4490 568710 4500 568890
rect 4300 568700 4500 568710
rect 6300 568890 6500 568900
rect 6300 568710 6310 568890
rect 6490 568710 6500 568890
rect 6300 568700 6500 568710
rect 8300 568890 8500 568900
rect 8300 568710 8310 568890
rect 8490 568710 8500 568890
rect 8300 568700 8500 568710
rect 575296 568890 575496 568900
rect 575296 568710 575306 568890
rect 575486 568710 575496 568890
rect 575296 568700 575496 568710
rect 577296 568890 577496 568900
rect 577296 568710 577306 568890
rect 577486 568710 577496 568890
rect 577296 568700 577496 568710
rect 579296 568890 579496 568900
rect 579296 568710 579306 568890
rect 579486 568710 579496 568890
rect 579296 568700 579496 568710
rect 581296 568890 581496 568900
rect 581296 568710 581306 568890
rect 581486 568710 581496 568890
rect 581296 568700 581496 568710
<< via2 >>
rect 2310 568710 2490 568890
rect 4310 568710 4490 568890
rect 6310 568710 6490 568890
rect 8310 568710 8490 568890
rect 575306 568710 575486 568890
rect 577306 568710 577486 568890
rect 579306 568710 579486 568890
rect 581306 568710 581486 568890
<< metal3 >>
rect 2300 568890 2500 568900
rect 2300 568710 2310 568890
rect 2490 568710 2500 568890
rect 2300 379000 2500 568710
rect 4300 568890 4500 568900
rect 4300 568710 4310 568890
rect 4490 568710 4500 568890
rect 0 377800 4000 379000
rect 0 335300 4000 335758
rect 4300 335300 4500 568710
rect 0 335100 4500 335300
rect 6300 568890 6500 568900
rect 6300 568710 6310 568890
rect 6490 568710 6500 568890
rect 0 334558 4000 335100
rect 0 292100 4000 292536
rect 6300 292100 6500 568710
rect 0 291900 6500 292100
rect 8300 568890 8500 568900
rect 8300 568710 8310 568890
rect 8490 568710 8500 568890
rect 0 291336 4000 291900
rect 0 249000 4000 249514
rect 8300 249000 8500 568710
rect 9000 492000 11000 686000
rect 12000 582000 14000 702000
rect 68000 700000 125194 702300
rect 146000 702000 170600 702300
rect 175894 702000 181000 702300
rect 146000 700000 181000 702000
rect 217294 702000 222294 702300
rect 227594 702000 238000 702300
rect 217294 700000 238000 702000
rect 318994 702000 323994 702300
rect 329294 702000 362000 702300
rect 318994 700000 362000 702000
rect 413394 700000 472000 702300
rect 570000 582000 572000 702000
rect 12000 580000 16000 582000
rect 566000 580000 572000 582000
rect 573000 492000 575000 684000
rect 9000 490000 16000 492000
rect 566000 490000 575000 492000
rect 575296 568890 575496 568900
rect 575296 568710 575306 568890
rect 575486 568710 575496 568890
rect 575296 273000 575496 568710
rect 577296 568890 577496 568900
rect 577296 568710 577306 568890
rect 577486 568710 577496 568890
rect 577296 317400 577496 568710
rect 579296 568890 579496 568900
rect 579296 568710 579306 568890
rect 579486 568710 579496 568890
rect 579296 362600 579496 568710
rect 581296 568890 581496 568900
rect 581296 568710 581306 568890
rect 581486 568710 581496 568890
rect 581296 409524 581496 568710
rect 580000 408324 584000 409524
rect 580000 362600 584000 363101
rect 579296 362400 584000 362600
rect 580000 361901 584000 362400
rect 580000 317400 584000 317880
rect 577296 317200 584000 317400
rect 580000 316680 584000 317200
rect 580000 273000 584000 273458
rect 575296 272800 584000 273000
rect 580000 272258 584000 272800
rect 0 248800 8500 249000
rect 0 248314 4000 248800
<< metal4 >>
rect 68000 700000 125194 702300
rect 146000 702000 170600 702300
rect 175894 702000 181000 702300
rect 146000 700000 181000 702000
rect 217294 702000 222294 702300
rect 227594 702000 238000 702300
rect 217294 700000 238000 702000
rect 318994 702000 323994 702300
rect 329294 702000 362000 702300
rect 318994 700000 362000 702000
rect 413394 700000 472000 702300
<< metal5 >>
rect 68000 700000 125194 702300
rect 146000 702000 170600 702300
rect 175894 702000 181000 702300
rect 146000 700000 181000 702000
rect 217294 702000 222294 702300
rect 227594 702000 238000 702300
rect 217294 700000 238000 702000
rect 318994 702000 323994 702300
rect 329294 702000 362000 702300
rect 318994 700000 362000 702000
rect 413394 700000 472000 702300
<< comment >>
rect 28560 682200 88560 702200
rect 128560 682200 188560 702200
rect 228560 682200 288560 702200
rect 328560 682200 388560 702200
rect 428560 682200 488560 702200
rect 0 0 2000 2000
use interleaved  interleaved_0
timestamp 1667247273
transform 1 0 292560 0 1 251000
box -278240 0 277120 451200
<< end >>
