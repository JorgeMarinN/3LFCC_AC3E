magic
tech sky130A
magscale 1 2
timestamp 1665097055
<< nwell >>
rect -304 36844 3274 41092
<< mvpsubdiff >>
rect 3172 34952 3224 34976
rect -246 34904 -194 34928
rect 3172 33980 3224 34004
rect -246 33932 -194 33956
rect -166 32166 -142 32272
rect 3122 32166 3146 32272
<< mvnsubdiff >>
rect -44 40968 -14 41022
rect 2976 40968 3026 41022
rect 3152 39518 3206 39570
rect -238 39440 -184 39488
rect -186 38492 -184 39440
rect 3152 38570 3154 39518
rect 3152 38522 3206 38570
rect -238 38440 -184 38492
<< mvpsubdiffcont >>
rect -246 33956 -194 34904
rect 3172 34004 3224 34952
rect -142 32166 3122 32272
<< mvnsubdiffcont >>
rect -14 40968 2976 41022
rect -238 38492 -186 39440
rect 3154 38570 3206 39518
<< poly >>
rect -42 36358 18 36914
rect 116 36824 176 36916
rect 274 36824 334 36914
rect 116 36758 334 36824
rect 116 36358 176 36758
rect 274 36358 334 36758
rect 432 36824 492 36916
rect 590 36824 650 36914
rect 432 36758 650 36824
rect 432 36358 492 36758
rect 590 36358 650 36758
rect 748 36824 808 36916
rect 906 36824 966 36914
rect 748 36758 966 36824
rect 748 36358 808 36758
rect 906 36358 966 36758
rect 1064 36824 1124 36916
rect 1222 36824 1282 36914
rect 1064 36758 1282 36824
rect 1064 36358 1124 36758
rect 1222 36358 1282 36758
rect 1380 36824 1440 36916
rect 1538 36824 1598 36914
rect 1380 36758 1598 36824
rect 1380 36358 1440 36758
rect 1538 36358 1598 36758
rect 1696 36824 1756 36916
rect 1854 36824 1914 36914
rect 1696 36758 1914 36824
rect 1696 36358 1756 36758
rect 1854 36358 1914 36758
rect 2012 36824 2072 36916
rect 2170 36824 2230 36914
rect 2012 36758 2230 36824
rect 2012 36358 2072 36758
rect 2170 36358 2230 36758
rect 2328 36824 2388 36916
rect 2486 36824 2546 36914
rect 2328 36758 2546 36824
rect 2328 36358 2388 36758
rect 2486 36358 2546 36758
rect 2644 36824 2704 36916
rect 2802 36824 2862 36914
rect 2644 36758 2862 36824
rect 2644 36358 2704 36758
rect 2802 36358 2862 36758
rect 2960 36358 3020 36916
<< locali >>
rect -36 40968 -14 41022
rect 2976 40968 3018 41022
rect 3152 39518 3206 39562
rect -238 39440 -184 39480
rect -186 38492 -184 39440
rect 3152 38570 3154 39518
rect 3152 38530 3206 38570
rect -238 38448 -184 38492
rect 3172 34952 3224 34968
rect -246 34904 -194 34920
rect 3172 33988 3224 34004
rect -246 33940 -194 33956
rect -158 32166 -142 32272
rect 3122 32166 3138 32272
<< viali >>
rect -14 40968 2976 41022
rect -238 38492 -186 39440
rect 3154 38570 3206 39518
rect -142 32166 3122 32272
<< metal1 >>
rect -244 41022 3212 41032
rect -244 40968 -14 41022
rect 2976 40968 3212 41022
rect -244 40960 3212 40968
rect -244 39442 -180 40960
rect -110 40890 -76 40960
rect 206 40890 242 40960
rect 522 40890 558 40960
rect 838 40890 874 40960
rect 1154 40890 1190 40960
rect 1470 40890 1506 40960
rect 1786 40890 1822 40960
rect 2102 40890 2138 40960
rect 2418 40890 2454 40960
rect 2734 40890 2770 40960
rect 3050 40890 3086 40960
rect 3148 39518 3212 40960
rect -244 39440 -98 39442
rect -244 38492 -238 39440
rect -186 38492 -98 39440
rect 3082 38570 3154 39518
rect 3206 38570 3212 39518
rect 3082 38568 3212 38570
rect 3148 38558 3212 38568
rect -244 38480 -180 38492
rect -64 36758 -54 36824
rect 12 36758 22 36824
rect 50 36520 82 36914
rect 180 36758 190 36824
rect 256 36758 266 36824
rect 22 36454 32 36520
rect 98 36454 108 36520
rect 366 36518 398 36914
rect 496 36758 506 36824
rect 572 36758 582 36824
rect 682 36518 714 36914
rect 812 36758 822 36824
rect 888 36758 898 36824
rect 998 36518 1030 36914
rect 1128 36758 1138 36824
rect 1204 36758 1214 36824
rect 1314 36518 1346 36914
rect 1446 36758 1456 36824
rect 1522 36758 1532 36824
rect 1630 36518 1662 36914
rect 1762 36758 1772 36824
rect 1838 36758 1848 36824
rect 1946 36518 1978 36914
rect 2076 36758 2086 36824
rect 2152 36758 2162 36824
rect 2262 36518 2294 36914
rect 2392 36758 2402 36824
rect 2468 36758 2478 36824
rect 50 36358 82 36454
rect 340 36452 350 36518
rect 416 36452 426 36518
rect 656 36452 666 36518
rect 732 36452 742 36518
rect 974 36452 984 36518
rect 1050 36452 1060 36518
rect 1288 36452 1298 36518
rect 1364 36452 1374 36518
rect 1604 36452 1614 36518
rect 1680 36452 1690 36518
rect 1920 36452 1930 36518
rect 1996 36452 2006 36518
rect 2236 36452 2246 36518
rect 2312 36452 2322 36518
rect 2578 36516 2610 36914
rect 2710 36758 2720 36824
rect 2786 36758 2796 36824
rect 2894 36516 2926 36914
rect 2968 36758 2978 36824
rect 3044 36758 3054 36824
rect 366 36358 398 36452
rect 682 36358 714 36452
rect 998 36358 1030 36452
rect 1314 36358 1346 36452
rect 1630 36358 1662 36452
rect 1946 36358 1978 36452
rect 2262 36358 2294 36452
rect 2552 36450 2562 36516
rect 2628 36450 2638 36516
rect 2868 36450 2878 36516
rect 2944 36450 2954 36516
rect 2578 36358 2610 36450
rect 2894 36358 2926 36450
rect -246 33984 -90 34904
rect 3068 34024 3212 34954
rect 3068 34006 3224 34024
rect -248 33956 -90 33984
rect -248 32286 -194 33956
rect -108 32286 -74 32382
rect 206 32286 240 32384
rect 524 32286 558 32384
rect 838 32286 872 32384
rect 1156 32286 1190 32384
rect 1470 32286 1504 32384
rect 1788 32286 1822 32384
rect 2102 32286 2136 32384
rect 2420 32286 2454 32382
rect 2734 32286 2768 32382
rect 3052 32286 3086 32382
rect 3170 32286 3224 34006
rect -248 32272 3224 32286
rect -248 32166 -142 32272
rect 3122 32166 3224 32272
rect -248 32158 3224 32166
<< via1 >>
rect -54 36758 12 36824
rect 190 36758 256 36824
rect 32 36454 98 36520
rect 506 36758 572 36824
rect 822 36758 888 36824
rect 1138 36758 1204 36824
rect 1456 36758 1522 36824
rect 1772 36758 1838 36824
rect 2086 36758 2152 36824
rect 2402 36758 2468 36824
rect 350 36452 416 36518
rect 666 36452 732 36518
rect 984 36452 1050 36518
rect 1298 36452 1364 36518
rect 1614 36452 1680 36518
rect 1930 36452 1996 36518
rect 2246 36452 2312 36518
rect 2720 36758 2786 36824
rect 2978 36758 3044 36824
rect 2562 36450 2628 36516
rect 2878 36450 2944 36516
<< metal2 >>
rect -160 36824 3130 36840
rect -160 36758 -54 36824
rect 12 36758 190 36824
rect 256 36758 506 36824
rect 572 36758 822 36824
rect 888 36758 1138 36824
rect 1204 36758 1456 36824
rect 1522 36758 1772 36824
rect 1838 36758 2086 36824
rect 2152 36758 2402 36824
rect 2468 36758 2720 36824
rect 2786 36758 2978 36824
rect 3044 36758 3130 36824
rect -160 36740 3130 36758
rect -160 36520 3130 36536
rect -160 36454 32 36520
rect 98 36518 3130 36520
rect 98 36454 350 36518
rect -160 36452 350 36454
rect 416 36452 666 36518
rect 732 36452 984 36518
rect 1050 36452 1298 36518
rect 1364 36452 1614 36518
rect 1680 36452 1930 36518
rect 1996 36452 2246 36518
rect 2312 36516 3130 36518
rect 2312 36452 2562 36516
rect -160 36450 2562 36452
rect 2628 36450 2878 36516
rect 2944 36450 3130 36516
rect -160 36436 3130 36450
use cont_poly_min  cont_poly_min_0
timestamp 1663264347
transform 1 0 -21 0 1 36725
box -33 33 33 99
use cont_poly_min  cont_poly_min_2
timestamp 1663264347
transform 1 0 223 0 1 36725
box -33 33 33 99
use cont_poly_min  cont_poly_min_3
timestamp 1663264347
transform 1 0 539 0 1 36725
box -33 33 33 99
use cont_poly_min  cont_poly_min_4
timestamp 1663264347
transform 1 0 855 0 1 36725
box -33 33 33 99
use cont_poly_min  cont_poly_min_5
timestamp 1663264347
transform 1 0 1171 0 1 36725
box -33 33 33 99
use cont_poly_min  cont_poly_min_6
timestamp 1663264347
transform 1 0 1489 0 1 36725
box -33 33 33 99
use cont_poly_min  cont_poly_min_7
timestamp 1663264347
transform 1 0 1805 0 1 36725
box -33 33 33 99
use cont_poly_min  cont_poly_min_8
timestamp 1663264347
transform 1 0 2119 0 1 36725
box -33 33 33 99
use cont_poly_min  cont_poly_min_9
timestamp 1663264347
transform 1 0 2435 0 1 36725
box -33 33 33 99
use cont_poly_min  cont_poly_min_10
timestamp 1663264347
transform 1 0 2753 0 1 36725
box -33 33 33 99
use cont_poly_min  cont_poly_min_11
timestamp 1663264347
transform 1 0 3011 0 1 36725
box -33 33 33 99
use sky130_fd_pr__nfet_g5v0d10v5_PPR2BY  sky130_fd_pr__nfet_g5v0d10v5_PPR2BY_0
timestamp 1663359535
transform 1 0 1489 0 1 34364
box -1609 -2026 1609 2026
use sky130_fd_pr__pfet_g5v0d10v5_VJVCZ4  sky130_fd_pr__pfet_g5v0d10v5_VJVCZ4_0
timestamp 1663460437
transform 1 0 1489 0 1 38912
box -1675 -2066 1675 2066
<< labels >>
rlabel metal2 -160 36740 -54 36840 1 IN
rlabel metal2 2944 36436 3130 36536 1 OUT
<< end >>
