magic
tech sky130A
magscale 1 2
timestamp 1665425771
<< nwell >>
rect -200 8934 100 8936
rect -200 8930 3604 8934
rect -1924 6680 3604 8930
rect 26 4686 3604 6680
rect -1931 3092 -1321 3634
rect -910 2200 -272 2872
<< nmos >>
rect -1833 3785 -1803 3985
rect -1737 3785 -1707 3985
rect -1641 3785 -1611 3985
rect -1545 3785 -1515 3985
rect -1449 3785 -1419 3985
<< pmos >>
rect -1833 3334 -1803 3534
rect -1737 3334 -1707 3534
rect -1641 3334 -1611 3534
rect -1545 3334 -1515 3534
rect -1449 3334 -1419 3534
<< mvnmos >>
rect -1800 4320 -1700 6320
rect -1642 4320 -1542 6320
rect -1484 4320 -1384 6320
rect -1326 4320 -1226 6320
rect -1168 4320 -1068 6320
rect -1010 4320 -910 6320
rect -852 4320 -752 6320
rect -694 4320 -594 6320
rect -536 4320 -436 6320
rect -378 4320 -278 6320
rect -1098 3132 -998 3932
rect -940 3132 -840 3932
rect -782 3132 -682 3932
rect -484 3132 -384 3932
rect -326 3132 -226 3932
rect -168 3132 -68 3932
rect 268 206 368 4206
rect 426 206 526 4206
rect 584 206 684 4206
rect 742 206 842 4206
rect 900 206 1000 4206
rect 1058 206 1158 4206
rect 1216 206 1316 4206
rect 1374 206 1474 4206
rect 1532 206 1632 4206
rect 1690 206 1790 4206
rect 1848 206 1948 4206
rect 2006 206 2106 4206
rect 2164 206 2264 4206
rect 2322 206 2422 4206
rect 2480 206 2580 4206
rect 2638 206 2738 4206
rect 2796 206 2896 4206
rect 2954 206 3054 4206
rect 3112 206 3212 4206
rect 3270 206 3370 4206
<< mvpmos >>
rect -1800 6746 -1700 8746
rect -1642 6746 -1542 8746
rect -1484 6746 -1384 8746
rect -1326 6746 -1226 8746
rect -1168 6746 -1068 8746
rect -1010 6746 -910 8746
rect -852 6746 -752 8746
rect -694 6746 -594 8746
rect -536 6746 -436 8746
rect -378 6746 -278 8746
rect 268 4754 368 8754
rect 426 4754 526 8754
rect 584 4754 684 8754
rect 742 4754 842 8754
rect 900 4754 1000 8754
rect 1058 4754 1158 8754
rect 1216 4754 1316 8754
rect 1374 4754 1474 8754
rect 1532 4754 1632 8754
rect 1690 4754 1790 8754
rect 1848 4754 1948 8754
rect 2006 4754 2106 8754
rect 2164 4754 2264 8754
rect 2322 4754 2422 8754
rect 2480 4754 2580 8754
rect 2638 4754 2738 8754
rect 2796 4754 2896 8754
rect 2954 4754 3054 8754
rect 3112 4754 3212 8754
rect 3270 4754 3370 8754
rect -786 2372 -686 2772
rect -496 2372 -396 2772
<< ndiff >>
rect -1895 3973 -1833 3985
rect -1895 3797 -1883 3973
rect -1849 3797 -1833 3973
rect -1895 3785 -1833 3797
rect -1803 3973 -1737 3985
rect -1803 3797 -1787 3973
rect -1753 3797 -1737 3973
rect -1803 3785 -1737 3797
rect -1707 3973 -1641 3985
rect -1707 3797 -1691 3973
rect -1657 3797 -1641 3973
rect -1707 3785 -1641 3797
rect -1611 3973 -1545 3985
rect -1611 3797 -1595 3973
rect -1561 3797 -1545 3973
rect -1611 3785 -1545 3797
rect -1515 3973 -1449 3985
rect -1515 3797 -1499 3973
rect -1465 3797 -1449 3973
rect -1515 3785 -1449 3797
rect -1419 3973 -1357 3985
rect -1419 3797 -1403 3973
rect -1369 3797 -1357 3973
rect -1419 3785 -1357 3797
<< pdiff >>
rect -1895 3522 -1833 3534
rect -1895 3346 -1883 3522
rect -1849 3346 -1833 3522
rect -1895 3334 -1833 3346
rect -1803 3522 -1737 3534
rect -1803 3346 -1787 3522
rect -1753 3346 -1737 3522
rect -1803 3334 -1737 3346
rect -1707 3522 -1641 3534
rect -1707 3346 -1691 3522
rect -1657 3346 -1641 3522
rect -1707 3334 -1641 3346
rect -1611 3522 -1545 3534
rect -1611 3346 -1595 3522
rect -1561 3346 -1545 3522
rect -1611 3334 -1545 3346
rect -1515 3522 -1449 3534
rect -1515 3346 -1499 3522
rect -1465 3346 -1449 3522
rect -1515 3334 -1449 3346
rect -1419 3522 -1357 3534
rect -1419 3346 -1403 3522
rect -1369 3346 -1357 3522
rect -1419 3334 -1357 3346
<< mvndiff >>
rect -1858 6308 -1800 6320
rect -1858 4332 -1846 6308
rect -1812 4332 -1800 6308
rect -1858 4320 -1800 4332
rect -1700 6308 -1642 6320
rect -1700 4332 -1688 6308
rect -1654 4332 -1642 6308
rect -1700 4320 -1642 4332
rect -1542 6308 -1484 6320
rect -1542 4332 -1530 6308
rect -1496 4332 -1484 6308
rect -1542 4320 -1484 4332
rect -1384 6308 -1326 6320
rect -1384 4332 -1372 6308
rect -1338 4332 -1326 6308
rect -1384 4320 -1326 4332
rect -1226 6308 -1168 6320
rect -1226 4332 -1214 6308
rect -1180 4332 -1168 6308
rect -1226 4320 -1168 4332
rect -1068 6308 -1010 6320
rect -1068 4332 -1056 6308
rect -1022 4332 -1010 6308
rect -1068 4320 -1010 4332
rect -910 6308 -852 6320
rect -910 4332 -898 6308
rect -864 4332 -852 6308
rect -910 4320 -852 4332
rect -752 6308 -694 6320
rect -752 4332 -740 6308
rect -706 4332 -694 6308
rect -752 4320 -694 4332
rect -594 6308 -536 6320
rect -594 4332 -582 6308
rect -548 4332 -536 6308
rect -594 4320 -536 4332
rect -436 6308 -378 6320
rect -436 4332 -424 6308
rect -390 4332 -378 6308
rect -436 4320 -378 4332
rect -278 6308 -220 6320
rect -278 4332 -266 6308
rect -232 4332 -220 6308
rect -278 4320 -220 4332
rect 210 4194 268 4206
rect -1156 3920 -1098 3932
rect -1156 3144 -1144 3920
rect -1110 3144 -1098 3920
rect -1156 3132 -1098 3144
rect -998 3920 -940 3932
rect -998 3144 -986 3920
rect -952 3144 -940 3920
rect -998 3132 -940 3144
rect -840 3920 -782 3932
rect -840 3144 -828 3920
rect -794 3144 -782 3920
rect -840 3132 -782 3144
rect -682 3920 -624 3932
rect -682 3144 -670 3920
rect -636 3144 -624 3920
rect -682 3132 -624 3144
rect -542 3920 -484 3932
rect -542 3144 -530 3920
rect -496 3144 -484 3920
rect -542 3132 -484 3144
rect -384 3920 -326 3932
rect -384 3144 -372 3920
rect -338 3144 -326 3920
rect -384 3132 -326 3144
rect -226 3920 -168 3932
rect -226 3144 -214 3920
rect -180 3144 -168 3920
rect -226 3132 -168 3144
rect -68 3920 -10 3932
rect -68 3144 -56 3920
rect -22 3144 -10 3920
rect -68 3132 -10 3144
rect 210 218 222 4194
rect 256 218 268 4194
rect 210 206 268 218
rect 368 4194 426 4206
rect 368 218 380 4194
rect 414 218 426 4194
rect 368 206 426 218
rect 526 4194 584 4206
rect 526 218 538 4194
rect 572 218 584 4194
rect 526 206 584 218
rect 684 4194 742 4206
rect 684 218 696 4194
rect 730 218 742 4194
rect 684 206 742 218
rect 842 4194 900 4206
rect 842 218 854 4194
rect 888 218 900 4194
rect 842 206 900 218
rect 1000 4194 1058 4206
rect 1000 218 1012 4194
rect 1046 218 1058 4194
rect 1000 206 1058 218
rect 1158 4194 1216 4206
rect 1158 218 1170 4194
rect 1204 218 1216 4194
rect 1158 206 1216 218
rect 1316 4194 1374 4206
rect 1316 218 1328 4194
rect 1362 218 1374 4194
rect 1316 206 1374 218
rect 1474 4194 1532 4206
rect 1474 218 1486 4194
rect 1520 218 1532 4194
rect 1474 206 1532 218
rect 1632 4194 1690 4206
rect 1632 218 1644 4194
rect 1678 218 1690 4194
rect 1632 206 1690 218
rect 1790 4194 1848 4206
rect 1790 218 1802 4194
rect 1836 218 1848 4194
rect 1790 206 1848 218
rect 1948 4194 2006 4206
rect 1948 218 1960 4194
rect 1994 218 2006 4194
rect 1948 206 2006 218
rect 2106 4194 2164 4206
rect 2106 218 2118 4194
rect 2152 218 2164 4194
rect 2106 206 2164 218
rect 2264 4194 2322 4206
rect 2264 218 2276 4194
rect 2310 218 2322 4194
rect 2264 206 2322 218
rect 2422 4194 2480 4206
rect 2422 218 2434 4194
rect 2468 218 2480 4194
rect 2422 206 2480 218
rect 2580 4194 2638 4206
rect 2580 218 2592 4194
rect 2626 218 2638 4194
rect 2580 206 2638 218
rect 2738 4194 2796 4206
rect 2738 218 2750 4194
rect 2784 218 2796 4194
rect 2738 206 2796 218
rect 2896 4194 2954 4206
rect 2896 218 2908 4194
rect 2942 218 2954 4194
rect 2896 206 2954 218
rect 3054 4194 3112 4206
rect 3054 218 3066 4194
rect 3100 218 3112 4194
rect 3054 206 3112 218
rect 3212 4194 3270 4206
rect 3212 218 3224 4194
rect 3258 218 3270 4194
rect 3212 206 3270 218
rect 3370 4194 3428 4206
rect 3370 218 3382 4194
rect 3416 218 3428 4194
rect 3370 206 3428 218
<< mvpdiff >>
rect -1858 8734 -1800 8746
rect -1858 6758 -1846 8734
rect -1812 6758 -1800 8734
rect -1858 6746 -1800 6758
rect -1700 8734 -1642 8746
rect -1700 6758 -1688 8734
rect -1654 6758 -1642 8734
rect -1700 6746 -1642 6758
rect -1542 8734 -1484 8746
rect -1542 6758 -1530 8734
rect -1496 6758 -1484 8734
rect -1542 6746 -1484 6758
rect -1384 8734 -1326 8746
rect -1384 6758 -1372 8734
rect -1338 6758 -1326 8734
rect -1384 6746 -1326 6758
rect -1226 8734 -1168 8746
rect -1226 6758 -1214 8734
rect -1180 6758 -1168 8734
rect -1226 6746 -1168 6758
rect -1068 8734 -1010 8746
rect -1068 6758 -1056 8734
rect -1022 6758 -1010 8734
rect -1068 6746 -1010 6758
rect -910 8734 -852 8746
rect -910 6758 -898 8734
rect -864 6758 -852 8734
rect -910 6746 -852 6758
rect -752 8734 -694 8746
rect -752 6758 -740 8734
rect -706 6758 -694 8734
rect -752 6746 -694 6758
rect -594 8734 -536 8746
rect -594 6758 -582 8734
rect -548 6758 -536 8734
rect -594 6746 -536 6758
rect -436 8734 -378 8746
rect -436 6758 -424 8734
rect -390 6758 -378 8734
rect -436 6746 -378 6758
rect -278 8734 -220 8746
rect -278 6758 -266 8734
rect -232 6758 -220 8734
rect 210 8742 268 8754
rect -278 6746 -220 6758
rect 210 4766 222 8742
rect 256 4766 268 8742
rect 210 4754 268 4766
rect 368 8742 426 8754
rect 368 4766 380 8742
rect 414 4766 426 8742
rect 368 4754 426 4766
rect 526 8742 584 8754
rect 526 4766 538 8742
rect 572 4766 584 8742
rect 526 4754 584 4766
rect 684 8742 742 8754
rect 684 4766 696 8742
rect 730 4766 742 8742
rect 684 4754 742 4766
rect 842 8742 900 8754
rect 842 4766 854 8742
rect 888 4766 900 8742
rect 842 4754 900 4766
rect 1000 8742 1058 8754
rect 1000 4766 1012 8742
rect 1046 4766 1058 8742
rect 1000 4754 1058 4766
rect 1158 8742 1216 8754
rect 1158 4766 1170 8742
rect 1204 4766 1216 8742
rect 1158 4754 1216 4766
rect 1316 8742 1374 8754
rect 1316 4766 1328 8742
rect 1362 4766 1374 8742
rect 1316 4754 1374 4766
rect 1474 8742 1532 8754
rect 1474 4766 1486 8742
rect 1520 4766 1532 8742
rect 1474 4754 1532 4766
rect 1632 8742 1690 8754
rect 1632 4766 1644 8742
rect 1678 4766 1690 8742
rect 1632 4754 1690 4766
rect 1790 8742 1848 8754
rect 1790 4766 1802 8742
rect 1836 4766 1848 8742
rect 1790 4754 1848 4766
rect 1948 8742 2006 8754
rect 1948 4766 1960 8742
rect 1994 4766 2006 8742
rect 1948 4754 2006 4766
rect 2106 8742 2164 8754
rect 2106 4766 2118 8742
rect 2152 4766 2164 8742
rect 2106 4754 2164 4766
rect 2264 8742 2322 8754
rect 2264 4766 2276 8742
rect 2310 4766 2322 8742
rect 2264 4754 2322 4766
rect 2422 8742 2480 8754
rect 2422 4766 2434 8742
rect 2468 4766 2480 8742
rect 2422 4754 2480 4766
rect 2580 8742 2638 8754
rect 2580 4766 2592 8742
rect 2626 4766 2638 8742
rect 2580 4754 2638 4766
rect 2738 8742 2796 8754
rect 2738 4766 2750 8742
rect 2784 4766 2796 8742
rect 2738 4754 2796 4766
rect 2896 8742 2954 8754
rect 2896 4766 2908 8742
rect 2942 4766 2954 8742
rect 2896 4754 2954 4766
rect 3054 8742 3112 8754
rect 3054 4766 3066 8742
rect 3100 4766 3112 8742
rect 3054 4754 3112 4766
rect 3212 8742 3270 8754
rect 3212 4766 3224 8742
rect 3258 4766 3270 8742
rect 3212 4754 3270 4766
rect 3370 8742 3428 8754
rect 3370 4766 3382 8742
rect 3416 4766 3428 8742
rect 3370 4754 3428 4766
rect -844 2760 -786 2772
rect -844 2384 -832 2760
rect -798 2384 -786 2760
rect -844 2372 -786 2384
rect -686 2760 -628 2772
rect -686 2384 -674 2760
rect -640 2384 -628 2760
rect -686 2372 -628 2384
rect -554 2760 -496 2772
rect -554 2384 -542 2760
rect -508 2384 -496 2760
rect -554 2372 -496 2384
rect -396 2760 -338 2772
rect -396 2384 -384 2760
rect -350 2384 -338 2760
rect -396 2372 -338 2384
<< ndiffc >>
rect -1883 3797 -1849 3973
rect -1787 3797 -1753 3973
rect -1691 3797 -1657 3973
rect -1595 3797 -1561 3973
rect -1499 3797 -1465 3973
rect -1403 3797 -1369 3973
<< pdiffc >>
rect -1883 3346 -1849 3522
rect -1787 3346 -1753 3522
rect -1691 3346 -1657 3522
rect -1595 3346 -1561 3522
rect -1499 3346 -1465 3522
rect -1403 3346 -1369 3522
<< mvndiffc >>
rect -1846 4332 -1812 6308
rect -1688 4332 -1654 6308
rect -1530 4332 -1496 6308
rect -1372 4332 -1338 6308
rect -1214 4332 -1180 6308
rect -1056 4332 -1022 6308
rect -898 4332 -864 6308
rect -740 4332 -706 6308
rect -582 4332 -548 6308
rect -424 4332 -390 6308
rect -266 4332 -232 6308
rect -1144 3144 -1110 3920
rect -986 3144 -952 3920
rect -828 3144 -794 3920
rect -670 3144 -636 3920
rect -530 3144 -496 3920
rect -372 3144 -338 3920
rect -214 3144 -180 3920
rect -56 3144 -22 3920
rect 222 218 256 4194
rect 380 218 414 4194
rect 538 218 572 4194
rect 696 218 730 4194
rect 854 218 888 4194
rect 1012 218 1046 4194
rect 1170 218 1204 4194
rect 1328 218 1362 4194
rect 1486 218 1520 4194
rect 1644 218 1678 4194
rect 1802 218 1836 4194
rect 1960 218 1994 4194
rect 2118 218 2152 4194
rect 2276 218 2310 4194
rect 2434 218 2468 4194
rect 2592 218 2626 4194
rect 2750 218 2784 4194
rect 2908 218 2942 4194
rect 3066 218 3100 4194
rect 3224 218 3258 4194
rect 3382 218 3416 4194
<< mvpdiffc >>
rect -1846 6758 -1812 8734
rect -1688 6758 -1654 8734
rect -1530 6758 -1496 8734
rect -1372 6758 -1338 8734
rect -1214 6758 -1180 8734
rect -1056 6758 -1022 8734
rect -898 6758 -864 8734
rect -740 6758 -706 8734
rect -582 6758 -548 8734
rect -424 6758 -390 8734
rect -266 6758 -232 8734
rect 222 4766 256 8742
rect 380 4766 414 8742
rect 538 4766 572 8742
rect 696 4766 730 8742
rect 854 4766 888 8742
rect 1012 4766 1046 8742
rect 1170 4766 1204 8742
rect 1328 4766 1362 8742
rect 1486 4766 1520 8742
rect 1644 4766 1678 8742
rect 1802 4766 1836 8742
rect 1960 4766 1994 8742
rect 2118 4766 2152 8742
rect 2276 4766 2310 8742
rect 2434 4766 2468 8742
rect 2592 4766 2626 8742
rect 2750 4766 2784 8742
rect 2908 4766 2942 8742
rect 3066 4766 3100 8742
rect 3224 4766 3258 8742
rect 3382 4766 3416 8742
rect -832 2384 -798 2760
rect -674 2384 -640 2760
rect -542 2384 -508 2760
rect -384 2384 -350 2760
<< psubdiff >>
rect -1850 4043 -1826 4082
rect -1411 4043 -1387 4082
<< nsubdiff >>
rect -1888 3227 -1821 3261
rect -1432 3227 -1361 3261
<< mvpsubdiff >>
rect -1786 4160 -1762 4228
rect -324 4160 -220 4228
rect -1106 4016 -1082 4106
rect -82 4016 -58 4106
rect 84 2746 136 2770
rect 84 1774 136 1798
rect 3502 2794 3554 2818
rect 3502 1822 3554 1846
rect 164 8 188 114
rect 3452 8 3476 114
<< mvnsubdiff >>
rect -1780 8812 -1750 8864
rect -342 8812 -298 8864
rect 286 8810 316 8864
rect 3306 8810 3356 8864
rect 92 7282 146 7330
rect 144 6334 146 7282
rect 92 6282 146 6334
rect 3482 7360 3536 7412
rect 3482 6412 3484 7360
rect 3482 6364 3536 6412
rect -812 2266 -772 2308
rect -394 2266 -360 2308
<< psubdiffcont >>
rect -1826 4043 -1411 4082
<< nsubdiffcont >>
rect -1821 3227 -1432 3261
<< mvpsubdiffcont >>
rect -1762 4160 -324 4228
rect -1082 4016 -82 4106
rect 84 1798 136 2746
rect 3502 1846 3554 2794
rect 188 8 3452 114
<< mvnsubdiffcont >>
rect -1750 8812 -342 8864
rect 316 8810 3306 8864
rect 92 6334 144 7282
rect 3484 6412 3536 7360
rect -772 2266 -394 2308
<< poly >>
rect -1800 8746 -1700 8772
rect -1642 8746 -1542 8772
rect -1484 8746 -1384 8772
rect -1326 8746 -1226 8772
rect -1168 8746 -1068 8772
rect -1010 8746 -910 8772
rect -852 8746 -752 8772
rect -694 8746 -594 8772
rect -536 8746 -436 8772
rect -378 8746 -278 8772
rect 268 8754 368 8780
rect 426 8754 526 8780
rect 584 8754 684 8780
rect 742 8754 842 8780
rect 900 8754 1000 8780
rect 1058 8754 1158 8780
rect 1216 8754 1316 8780
rect 1374 8754 1474 8780
rect 1532 8754 1632 8780
rect 1690 8754 1790 8780
rect 1848 8754 1948 8780
rect 2006 8754 2106 8780
rect 2164 8754 2264 8780
rect 2322 8754 2422 8780
rect 2480 8754 2580 8780
rect 2638 8754 2738 8780
rect 2796 8754 2896 8780
rect 2954 8754 3054 8780
rect 3112 8754 3212 8780
rect 3270 8754 3370 8780
rect -1800 6720 -1700 6746
rect -1642 6720 -1542 6746
rect -1484 6720 -1384 6746
rect -1326 6720 -1226 6746
rect -1168 6720 -1068 6746
rect -1010 6720 -910 6746
rect -852 6720 -752 6746
rect -694 6720 -594 6746
rect -536 6720 -436 6746
rect -378 6720 -278 6746
rect -1780 6674 -1720 6720
rect -1622 6676 -1562 6720
rect -1464 6676 -1404 6720
rect -1784 6658 -1718 6674
rect -1784 6624 -1768 6658
rect -1734 6624 -1718 6658
rect -1784 6608 -1718 6624
rect -1622 6660 -1404 6676
rect -1622 6626 -1530 6660
rect -1496 6626 -1404 6660
rect -1622 6610 -1404 6626
rect -1622 6608 -1562 6610
rect -1464 6608 -1404 6610
rect -1306 6676 -1246 6720
rect -1148 6676 -1088 6720
rect -1306 6660 -1088 6676
rect -1306 6626 -1216 6660
rect -1182 6626 -1088 6660
rect -1306 6610 -1088 6626
rect -1306 6608 -1246 6610
rect -1148 6608 -1088 6610
rect -990 6674 -930 6720
rect -832 6674 -772 6720
rect -990 6658 -772 6674
rect -990 6624 -898 6658
rect -864 6624 -772 6658
rect -990 6608 -772 6624
rect -674 6674 -614 6720
rect -516 6674 -456 6720
rect -674 6658 -456 6674
rect -674 6624 -584 6658
rect -550 6624 -456 6658
rect -674 6608 -456 6624
rect -358 6674 -298 6720
rect -358 6658 -290 6674
rect -358 6624 -340 6658
rect -306 6624 -290 6658
rect -358 6608 -290 6624
rect -1780 6602 -1720 6608
rect -358 6602 -298 6608
rect -1780 6456 -1720 6462
rect -1784 6440 -1718 6456
rect -1784 6406 -1768 6440
rect -1734 6406 -1718 6440
rect -1784 6390 -1718 6406
rect -1622 6442 -1404 6458
rect -1622 6408 -1530 6442
rect -1496 6408 -1404 6442
rect -1622 6392 -1404 6408
rect -1780 6346 -1720 6390
rect -1622 6346 -1562 6392
rect -1464 6346 -1404 6392
rect -1306 6442 -1088 6458
rect -1306 6408 -1216 6442
rect -1182 6408 -1088 6442
rect -1306 6392 -1088 6408
rect -1306 6346 -1246 6392
rect -1148 6346 -1088 6392
rect -990 6456 -930 6458
rect -832 6456 -772 6458
rect -990 6440 -772 6456
rect -990 6406 -898 6440
rect -864 6406 -772 6440
rect -990 6390 -772 6406
rect -990 6346 -930 6390
rect -832 6346 -772 6390
rect -674 6456 -614 6458
rect -516 6456 -456 6458
rect -674 6440 -456 6456
rect -674 6406 -584 6440
rect -550 6406 -456 6440
rect -674 6390 -456 6406
rect -674 6346 -614 6390
rect -516 6346 -456 6390
rect -358 6456 -298 6462
rect -358 6440 -290 6456
rect -358 6406 -340 6440
rect -306 6406 -290 6440
rect -358 6390 -290 6406
rect -358 6346 -298 6390
rect -1800 6320 -1700 6346
rect -1642 6320 -1542 6346
rect -1484 6320 -1384 6346
rect -1326 6320 -1226 6346
rect -1168 6320 -1068 6346
rect -1010 6320 -910 6346
rect -852 6320 -752 6346
rect -694 6320 -594 6346
rect -536 6320 -436 6346
rect -378 6320 -278 6346
rect 268 4728 368 4754
rect 426 4728 526 4754
rect 584 4728 684 4754
rect 742 4728 842 4754
rect 900 4728 1000 4754
rect 1058 4728 1158 4754
rect 1216 4728 1316 4754
rect 1374 4728 1474 4754
rect 1532 4728 1632 4754
rect 1690 4728 1790 4754
rect 1848 4728 1948 4754
rect 2006 4728 2106 4754
rect 2164 4728 2264 4754
rect 2322 4728 2422 4754
rect 2480 4728 2580 4754
rect 2638 4728 2738 4754
rect 2796 4728 2896 4754
rect 2954 4728 3054 4754
rect 3112 4728 3212 4754
rect 3270 4728 3370 4754
rect 288 4666 348 4728
rect 276 4650 348 4666
rect 276 4616 292 4650
rect 326 4616 348 4650
rect 276 4600 348 4616
rect -1800 4294 -1700 4320
rect -1642 4294 -1542 4320
rect -1484 4294 -1384 4320
rect -1326 4294 -1226 4320
rect -1168 4294 -1068 4320
rect -1010 4294 -910 4320
rect -852 4294 -752 4320
rect -694 4294 -594 4320
rect -536 4294 -436 4320
rect -378 4294 -278 4320
rect 288 4232 348 4600
rect 446 4666 506 4728
rect 604 4666 664 4728
rect 446 4650 664 4666
rect 446 4616 536 4650
rect 570 4616 664 4650
rect 446 4600 664 4616
rect 446 4232 506 4600
rect 604 4232 664 4600
rect 762 4666 822 4728
rect 920 4666 980 4728
rect 762 4650 980 4666
rect 762 4616 852 4650
rect 886 4616 980 4650
rect 762 4600 980 4616
rect 762 4232 822 4600
rect 920 4232 980 4600
rect 1078 4666 1138 4728
rect 1236 4666 1296 4728
rect 1078 4650 1296 4666
rect 1078 4616 1168 4650
rect 1202 4616 1296 4650
rect 1078 4600 1296 4616
rect 1078 4232 1138 4600
rect 1236 4232 1296 4600
rect 1394 4666 1454 4728
rect 1552 4666 1612 4728
rect 1394 4650 1612 4666
rect 1394 4616 1484 4650
rect 1518 4616 1612 4650
rect 1394 4600 1612 4616
rect 1394 4232 1454 4600
rect 1552 4232 1612 4600
rect 1710 4666 1770 4728
rect 1868 4666 1928 4728
rect 1710 4650 1928 4666
rect 1710 4616 1802 4650
rect 1836 4616 1928 4650
rect 1710 4600 1928 4616
rect 1710 4232 1770 4600
rect 1868 4232 1928 4600
rect 2026 4666 2086 4728
rect 2184 4666 2244 4728
rect 2026 4650 2244 4666
rect 2026 4616 2118 4650
rect 2152 4616 2244 4650
rect 2026 4600 2244 4616
rect 2026 4232 2086 4600
rect 2184 4232 2244 4600
rect 2342 4666 2402 4728
rect 2500 4666 2560 4728
rect 2342 4650 2560 4666
rect 2342 4616 2432 4650
rect 2466 4616 2560 4650
rect 2342 4600 2560 4616
rect 2342 4232 2402 4600
rect 2500 4232 2560 4600
rect 2658 4666 2718 4728
rect 2816 4666 2876 4728
rect 2658 4650 2876 4666
rect 2658 4616 2748 4650
rect 2782 4616 2876 4650
rect 2658 4600 2876 4616
rect 2658 4232 2718 4600
rect 2816 4232 2876 4600
rect 2974 4666 3034 4728
rect 3132 4666 3192 4728
rect 2974 4650 3192 4666
rect 2974 4616 3066 4650
rect 3100 4616 3192 4650
rect 2974 4600 3192 4616
rect 2974 4232 3034 4600
rect 3132 4232 3192 4600
rect 3290 4666 3350 4728
rect 3290 4650 3374 4666
rect 3290 4616 3324 4650
rect 3358 4616 3374 4650
rect 3290 4600 3374 4616
rect 3290 4232 3350 4600
rect 268 4206 368 4232
rect 426 4206 526 4232
rect 584 4206 684 4232
rect 742 4206 842 4232
rect 900 4206 1000 4232
rect 1058 4206 1158 4232
rect 1216 4206 1316 4232
rect 1374 4206 1474 4232
rect 1532 4206 1632 4232
rect 1690 4206 1790 4232
rect 1848 4206 1948 4232
rect 2006 4206 2106 4232
rect 2164 4206 2264 4232
rect 2322 4206 2422 4232
rect 2480 4206 2580 4232
rect 2638 4206 2738 4232
rect 2796 4206 2896 4232
rect 2954 4206 3054 4232
rect 3112 4206 3212 4232
rect 3270 4206 3370 4232
rect -1833 3985 -1803 4011
rect -1737 3985 -1707 4011
rect -1641 3985 -1611 4011
rect -1545 3985 -1515 4011
rect -1449 3985 -1419 4011
rect -1098 3932 -998 3958
rect -940 3932 -840 3958
rect -782 3932 -682 3958
rect -484 3932 -384 3958
rect -326 3932 -226 3958
rect -168 3932 -68 3958
rect -1833 3634 -1803 3785
rect -1883 3618 -1803 3634
rect -1883 3584 -1867 3618
rect -1833 3584 -1803 3618
rect -1883 3568 -1803 3584
rect -1833 3534 -1803 3568
rect -1737 3634 -1707 3785
rect -1641 3634 -1611 3785
rect -1737 3618 -1611 3634
rect -1737 3584 -1691 3618
rect -1657 3584 -1611 3618
rect -1737 3568 -1611 3584
rect -1737 3534 -1707 3568
rect -1641 3534 -1611 3568
rect -1545 3631 -1515 3785
rect -1449 3631 -1419 3785
rect -1545 3615 -1419 3631
rect -1545 3581 -1499 3615
rect -1465 3581 -1419 3615
rect -1545 3565 -1419 3581
rect -1545 3534 -1515 3565
rect -1449 3534 -1419 3565
rect -1833 3308 -1803 3334
rect -1737 3303 -1707 3334
rect -1641 3308 -1611 3334
rect -1545 3303 -1515 3334
rect -1449 3308 -1419 3334
rect -1098 3106 -998 3132
rect -940 3106 -840 3132
rect -782 3106 -682 3132
rect -484 3106 -384 3132
rect -326 3106 -226 3132
rect -168 3106 -68 3132
rect -1080 3092 -1014 3106
rect -1080 3058 -1064 3092
rect -1030 3058 -1014 3092
rect -1080 3042 -1014 3058
rect -922 3094 -856 3106
rect -922 3060 -906 3094
rect -872 3060 -856 3094
rect -922 3044 -856 3060
rect -762 3094 -696 3106
rect -762 3060 -746 3094
rect -712 3060 -696 3094
rect -762 3044 -696 3060
rect -468 3094 -402 3106
rect -468 3060 -452 3094
rect -418 3060 -402 3094
rect -468 3044 -402 3060
rect -306 3094 -240 3106
rect -306 3060 -290 3094
rect -256 3060 -240 3094
rect -306 3044 -240 3060
rect -150 3094 -84 3106
rect -150 3060 -134 3094
rect -100 3060 -84 3094
rect -150 3044 -84 3060
rect -786 2853 -686 2869
rect -786 2819 -770 2853
rect -702 2819 -686 2853
rect -786 2772 -686 2819
rect -496 2853 -396 2869
rect -496 2819 -480 2853
rect -412 2819 -396 2853
rect -496 2772 -396 2819
rect -786 2346 -686 2372
rect -496 2346 -396 2372
rect 268 180 368 206
rect 426 180 526 206
rect 584 180 684 206
rect 742 180 842 206
rect 900 180 1000 206
rect 1058 180 1158 206
rect 1216 180 1316 206
rect 1374 180 1474 206
rect 1532 180 1632 206
rect 1690 180 1790 206
rect 1848 180 1948 206
rect 2006 180 2106 206
rect 2164 180 2264 206
rect 2322 180 2422 206
rect 2480 180 2580 206
rect 2638 180 2738 206
rect 2796 180 2896 206
rect 2954 180 3054 206
rect 3112 180 3212 206
rect 3270 180 3370 206
<< polycont >>
rect -1768 6624 -1734 6658
rect -1530 6626 -1496 6660
rect -1216 6626 -1182 6660
rect -898 6624 -864 6658
rect -584 6624 -550 6658
rect -340 6624 -306 6658
rect -1768 6406 -1734 6440
rect -1530 6408 -1496 6442
rect -1216 6408 -1182 6442
rect -898 6406 -864 6440
rect -584 6406 -550 6440
rect -340 6406 -306 6440
rect 292 4616 326 4650
rect 536 4616 570 4650
rect 852 4616 886 4650
rect 1168 4616 1202 4650
rect 1484 4616 1518 4650
rect 1802 4616 1836 4650
rect 2118 4616 2152 4650
rect 2432 4616 2466 4650
rect 2748 4616 2782 4650
rect 3066 4616 3100 4650
rect 3324 4616 3358 4650
rect -1867 3584 -1833 3618
rect -1691 3584 -1657 3618
rect -1499 3581 -1465 3615
rect -1064 3058 -1030 3092
rect -906 3060 -872 3094
rect -746 3060 -712 3094
rect -452 3060 -418 3094
rect -290 3060 -256 3094
rect -134 3060 -100 3094
rect -770 2819 -702 2853
rect -480 2819 -412 2853
<< locali >>
rect -1772 8812 -1750 8864
rect -342 8812 -306 8864
rect 294 8810 316 8864
rect 3306 8810 3348 8864
rect -1846 8734 -1812 8750
rect -1846 6742 -1812 6758
rect -1688 8734 -1654 8750
rect -1688 6742 -1654 6758
rect -1530 8734 -1496 8750
rect -1530 6742 -1496 6758
rect -1372 8734 -1338 8750
rect -1372 6742 -1338 6758
rect -1214 8734 -1180 8750
rect -1214 6742 -1180 6758
rect -1056 8734 -1022 8750
rect -1056 6742 -1022 6758
rect -898 8734 -864 8750
rect -898 6742 -864 6758
rect -740 8734 -706 8750
rect -740 6742 -706 6758
rect -582 8734 -548 8750
rect -582 6742 -548 6758
rect -424 8734 -390 8750
rect -424 6742 -390 6758
rect -266 8734 -232 8750
rect 222 8742 256 8758
rect -266 6742 -232 6758
rect 92 7282 146 7322
rect -1784 6624 -1768 6658
rect -1734 6624 -1718 6658
rect -1546 6626 -1530 6660
rect -1496 6626 -1480 6660
rect -1232 6626 -1216 6660
rect -1182 6626 -1166 6660
rect -914 6624 -898 6658
rect -864 6624 -848 6658
rect -600 6624 -584 6658
rect -550 6624 -534 6658
rect -356 6624 -340 6658
rect -306 6624 -290 6658
rect -1784 6406 -1768 6440
rect -1734 6406 -1718 6440
rect -1546 6408 -1530 6442
rect -1496 6408 -1480 6442
rect -1232 6408 -1216 6442
rect -1182 6408 -1166 6442
rect -914 6406 -898 6440
rect -864 6406 -848 6440
rect -600 6406 -584 6440
rect -550 6406 -534 6440
rect -356 6406 -340 6440
rect -306 6406 -290 6440
rect 144 6334 146 7282
rect -1846 6308 -1812 6324
rect -1846 4316 -1812 4332
rect -1688 6308 -1654 6324
rect -1688 4316 -1654 4332
rect -1530 6308 -1496 6324
rect -1530 4316 -1496 4332
rect -1372 6308 -1338 6324
rect -1372 4316 -1338 4332
rect -1214 6308 -1180 6324
rect -1214 4316 -1180 4332
rect -1056 6308 -1022 6324
rect -1056 4316 -1022 4332
rect -898 6308 -864 6324
rect -898 4316 -864 4332
rect -740 6308 -706 6324
rect -740 4316 -706 4332
rect -582 6308 -548 6324
rect -582 4316 -548 4332
rect -424 6308 -390 6324
rect -424 4316 -390 4332
rect -266 6308 -232 6324
rect 92 6290 146 6334
rect 222 4750 256 4766
rect 380 8742 414 8758
rect 380 4750 414 4766
rect 538 8742 572 8758
rect 538 4750 572 4766
rect 696 8742 730 8758
rect 696 4750 730 4766
rect 854 8742 888 8758
rect 854 4750 888 4766
rect 1012 8742 1046 8758
rect 1012 4750 1046 4766
rect 1170 8742 1204 8758
rect 1170 4750 1204 4766
rect 1328 8742 1362 8758
rect 1328 4750 1362 4766
rect 1486 8742 1520 8758
rect 1486 4750 1520 4766
rect 1644 8742 1678 8758
rect 1644 4750 1678 4766
rect 1802 8742 1836 8758
rect 1802 4750 1836 4766
rect 1960 8742 1994 8758
rect 1960 4750 1994 4766
rect 2118 8742 2152 8758
rect 2118 4750 2152 4766
rect 2276 8742 2310 8758
rect 2276 4750 2310 4766
rect 2434 8742 2468 8758
rect 2434 4750 2468 4766
rect 2592 8742 2626 8758
rect 2592 4750 2626 4766
rect 2750 8742 2784 8758
rect 2750 4750 2784 4766
rect 2908 8742 2942 8758
rect 2908 4750 2942 4766
rect 3066 8742 3100 8758
rect 3066 4750 3100 4766
rect 3224 8742 3258 8758
rect 3224 4750 3258 4766
rect 3382 8742 3416 8758
rect 3482 7360 3536 7404
rect 3482 6412 3484 7360
rect 3482 6372 3536 6412
rect 3382 4750 3416 4766
rect 276 4616 292 4650
rect 326 4616 342 4650
rect 520 4616 536 4650
rect 570 4616 586 4650
rect 836 4616 852 4650
rect 886 4616 902 4650
rect 1152 4616 1168 4650
rect 1202 4616 1218 4650
rect 1468 4616 1484 4650
rect 1518 4616 1534 4650
rect 1786 4616 1802 4650
rect 1836 4616 1852 4650
rect 2102 4616 2118 4650
rect 2152 4616 2168 4650
rect 2416 4616 2432 4650
rect 2466 4616 2482 4650
rect 2732 4616 2748 4650
rect 2782 4616 2798 4650
rect 3050 4616 3066 4650
rect 3100 4616 3116 4650
rect 3308 4616 3324 4650
rect 3358 4616 3374 4650
rect -266 4316 -232 4332
rect -1778 4160 -1762 4228
rect -324 4160 -308 4228
rect 222 4194 256 4210
rect -1098 4016 -1082 4106
rect -82 4016 -66 4106
rect -1883 3973 -1849 3989
rect -1883 3781 -1849 3797
rect -1787 3973 -1753 3989
rect -1787 3781 -1753 3797
rect -1691 3973 -1657 3989
rect -1691 3781 -1657 3797
rect -1595 3973 -1561 3989
rect -1595 3781 -1561 3797
rect -1499 3973 -1465 3989
rect -1499 3781 -1465 3797
rect -1403 3973 -1369 3989
rect -1403 3781 -1369 3797
rect -1144 3920 -1110 3936
rect -1883 3584 -1867 3618
rect -1833 3584 -1817 3618
rect -1707 3584 -1691 3618
rect -1657 3584 -1641 3618
rect -1515 3581 -1499 3615
rect -1465 3581 -1449 3615
rect -1883 3522 -1849 3538
rect -1883 3330 -1849 3346
rect -1787 3522 -1753 3538
rect -1787 3330 -1753 3346
rect -1691 3522 -1657 3538
rect -1691 3330 -1657 3346
rect -1595 3522 -1561 3538
rect -1595 3330 -1561 3346
rect -1499 3522 -1465 3538
rect -1499 3330 -1465 3346
rect -1403 3522 -1369 3538
rect -1403 3330 -1369 3346
rect -1144 3128 -1110 3144
rect -986 3920 -952 3936
rect -986 3128 -952 3144
rect -828 3920 -794 3936
rect -828 3128 -794 3144
rect -670 3920 -636 3936
rect -670 3128 -636 3144
rect -530 3920 -496 3936
rect -530 3128 -496 3144
rect -372 3920 -338 3936
rect -372 3128 -338 3144
rect -214 3920 -180 3936
rect -214 3128 -180 3144
rect -56 3920 -22 3936
rect -56 3128 -22 3144
rect -1080 3058 -1064 3092
rect -1030 3058 -1014 3092
rect -922 3060 -906 3094
rect -872 3060 -856 3094
rect -762 3060 -746 3094
rect -712 3060 -696 3094
rect -468 3060 -452 3094
rect -418 3060 -402 3094
rect -306 3060 -290 3094
rect -256 3060 -240 3094
rect -150 3060 -134 3094
rect -100 3060 -84 3094
rect -786 2819 -770 2853
rect -702 2819 -686 2853
rect -496 2819 -480 2853
rect -412 2819 -396 2853
rect -832 2760 -798 2776
rect -832 2368 -798 2384
rect -674 2760 -640 2776
rect -674 2368 -640 2384
rect -542 2760 -508 2776
rect -542 2368 -508 2384
rect -384 2760 -350 2776
rect -384 2368 -350 2384
rect 84 2746 136 2762
rect -804 2266 -772 2308
rect -394 2266 -368 2308
rect 84 1782 136 1798
rect 222 202 256 218
rect 380 4194 414 4210
rect 380 202 414 218
rect 538 4194 572 4210
rect 538 202 572 218
rect 696 4194 730 4210
rect 696 202 730 218
rect 854 4194 888 4210
rect 854 202 888 218
rect 1012 4194 1046 4210
rect 1012 202 1046 218
rect 1170 4194 1204 4210
rect 1170 202 1204 218
rect 1328 4194 1362 4210
rect 1328 202 1362 218
rect 1486 4194 1520 4210
rect 1486 202 1520 218
rect 1644 4194 1678 4210
rect 1644 202 1678 218
rect 1802 4194 1836 4210
rect 1802 202 1836 218
rect 1960 4194 1994 4210
rect 1960 202 1994 218
rect 2118 4194 2152 4210
rect 2118 202 2152 218
rect 2276 4194 2310 4210
rect 2276 202 2310 218
rect 2434 4194 2468 4210
rect 2434 202 2468 218
rect 2592 4194 2626 4210
rect 2592 202 2626 218
rect 2750 4194 2784 4210
rect 2750 202 2784 218
rect 2908 4194 2942 4210
rect 2908 202 2942 218
rect 3066 4194 3100 4210
rect 3066 202 3100 218
rect 3224 4194 3258 4210
rect 3224 202 3258 218
rect 3382 4194 3416 4210
rect 3502 2794 3554 2810
rect 3502 1830 3554 1846
rect 3382 202 3416 218
rect 172 8 188 114
rect 3452 8 3468 114
<< viali >>
rect -1750 8812 -342 8864
rect 316 8810 3306 8864
rect -1846 6758 -1812 8734
rect -1688 6758 -1654 8734
rect -1530 6758 -1496 8734
rect -1372 6758 -1338 8734
rect -1214 6758 -1180 8734
rect -1056 6758 -1022 8734
rect -898 6758 -864 8734
rect -740 6758 -706 8734
rect -582 6758 -548 8734
rect -424 6758 -390 8734
rect -266 6758 -232 8734
rect -1768 6624 -1734 6658
rect -1530 6626 -1496 6660
rect -1216 6626 -1182 6660
rect -898 6624 -864 6658
rect -584 6624 -550 6658
rect -340 6624 -306 6658
rect -1768 6406 -1734 6440
rect -1530 6408 -1496 6442
rect -1216 6408 -1182 6442
rect -898 6406 -864 6440
rect -584 6406 -550 6440
rect -340 6406 -306 6440
rect 92 6334 144 7282
rect -1846 4332 -1812 6308
rect -1688 4332 -1654 6308
rect -1530 4332 -1496 6308
rect -1372 4332 -1338 6308
rect -1214 4332 -1180 6308
rect -1056 4332 -1022 6308
rect -898 4332 -864 6308
rect -740 4332 -706 6308
rect -582 4332 -548 6308
rect -424 4332 -390 6308
rect -266 4332 -232 6308
rect 222 4766 256 8742
rect 380 4766 414 8742
rect 538 4766 572 8742
rect 696 4766 730 8742
rect 854 4766 888 8742
rect 1012 4766 1046 8742
rect 1170 4766 1204 8742
rect 1328 4766 1362 8742
rect 1486 4766 1520 8742
rect 1644 4766 1678 8742
rect 1802 4766 1836 8742
rect 1960 4766 1994 8742
rect 2118 4766 2152 8742
rect 2276 4766 2310 8742
rect 2434 4766 2468 8742
rect 2592 4766 2626 8742
rect 2750 4766 2784 8742
rect 2908 4766 2942 8742
rect 3066 4766 3100 8742
rect 3224 4766 3258 8742
rect 3382 4766 3416 8742
rect 3484 6412 3536 7360
rect 292 4616 326 4650
rect 536 4616 570 4650
rect 852 4616 886 4650
rect 1168 4616 1202 4650
rect 1484 4616 1518 4650
rect 1802 4616 1836 4650
rect 2118 4616 2152 4650
rect 2432 4616 2466 4650
rect 2748 4616 2782 4650
rect 3066 4616 3100 4650
rect 3324 4616 3358 4650
rect -1762 4162 -324 4228
rect -1891 4082 -1369 4086
rect -1891 4043 -1826 4082
rect -1826 4043 -1411 4082
rect -1411 4043 -1369 4082
rect -1891 4040 -1369 4043
rect -1082 4016 -82 4106
rect -1883 3797 -1849 3973
rect -1787 3797 -1753 3973
rect -1691 3797 -1657 3973
rect -1595 3797 -1561 3973
rect -1499 3797 -1465 3973
rect -1403 3797 -1369 3973
rect -1867 3584 -1833 3618
rect -1691 3584 -1657 3618
rect -1499 3581 -1465 3615
rect -1883 3346 -1849 3522
rect -1787 3346 -1753 3522
rect -1691 3346 -1657 3522
rect -1595 3346 -1561 3522
rect -1499 3346 -1465 3522
rect -1403 3346 -1369 3522
rect -1894 3261 -1359 3262
rect -1894 3227 -1821 3261
rect -1821 3227 -1432 3261
rect -1432 3227 -1359 3261
rect -1894 3226 -1359 3227
rect -1144 3144 -1110 3920
rect -986 3144 -952 3920
rect -828 3144 -794 3920
rect -670 3144 -636 3920
rect -530 3144 -496 3920
rect -372 3144 -338 3920
rect -214 3144 -180 3920
rect -56 3144 -22 3920
rect -1064 3058 -1030 3092
rect -906 3060 -872 3094
rect -746 3060 -712 3094
rect -452 3060 -418 3094
rect -290 3060 -256 3094
rect -134 3060 -100 3094
rect -770 2819 -702 2853
rect -480 2819 -412 2853
rect -832 2384 -798 2760
rect -674 2384 -640 2760
rect -542 2384 -508 2760
rect -384 2384 -350 2760
rect -772 2266 -394 2308
rect 222 218 256 4194
rect 380 218 414 4194
rect 538 218 572 4194
rect 696 218 730 4194
rect 854 218 888 4194
rect 1012 218 1046 4194
rect 1170 218 1204 4194
rect 1328 218 1362 4194
rect 1486 218 1520 4194
rect 1644 218 1678 4194
rect 1802 218 1836 4194
rect 1960 218 1994 4194
rect 2118 218 2152 4194
rect 2276 218 2310 4194
rect 2434 218 2468 4194
rect 2592 218 2626 4194
rect 2750 218 2784 4194
rect 2908 218 2942 4194
rect 3066 218 3100 4194
rect 3224 218 3258 4194
rect 3382 218 3416 4194
rect 188 8 3452 114
<< metal1 >>
rect -2436 8898 -2296 8900
rect -2436 8896 -1800 8898
rect -2436 8874 3274 8896
rect -2436 8864 3542 8874
rect -2436 8812 -1750 8864
rect -342 8812 316 8864
rect -2436 8810 316 8812
rect 3306 8810 3542 8864
rect -2436 8808 3542 8810
rect -2436 7738 -2296 8808
rect -1870 8806 3542 8808
rect -1846 8746 -1812 8806
rect -1530 8746 -1496 8806
rect -1214 8746 -1180 8806
rect -898 8746 -864 8806
rect -582 8746 -548 8806
rect -266 8746 -232 8806
rect 86 8802 3542 8806
rect -1852 8734 -1806 8746
rect -2436 7140 -2294 7738
rect -2434 2904 -2294 7140
rect -1852 6758 -1846 8734
rect -1812 6758 -1806 8734
rect -1852 6746 -1806 6758
rect -1694 8734 -1648 8746
rect -1694 6758 -1688 8734
rect -1654 6758 -1648 8734
rect -1694 6746 -1648 6758
rect -1536 8734 -1490 8746
rect -1536 6758 -1530 8734
rect -1496 6758 -1490 8734
rect -1536 6746 -1490 6758
rect -1378 8734 -1332 8746
rect -1378 6758 -1372 8734
rect -1338 6758 -1332 8734
rect -1378 6746 -1332 6758
rect -1220 8734 -1174 8746
rect -1220 6758 -1214 8734
rect -1180 6758 -1174 8734
rect -1220 6746 -1174 6758
rect -1062 8734 -1016 8746
rect -1062 6758 -1056 8734
rect -1022 6758 -1016 8734
rect -1062 6746 -1016 6758
rect -904 8734 -858 8746
rect -904 6758 -898 8734
rect -864 6758 -858 8734
rect -904 6746 -858 6758
rect -746 8734 -700 8746
rect -746 6758 -740 8734
rect -706 6758 -700 8734
rect -746 6746 -700 6758
rect -588 8734 -542 8746
rect -588 6758 -582 8734
rect -548 6758 -542 8734
rect -588 6746 -542 6758
rect -430 8734 -384 8746
rect -430 6758 -424 8734
rect -390 6758 -384 8734
rect -430 6746 -384 6758
rect -272 8734 -226 8746
rect -272 6758 -266 8734
rect -232 6758 -226 8734
rect -272 6746 -226 6758
rect 86 7284 150 8802
rect 220 8754 254 8802
rect 536 8754 572 8802
rect 852 8754 888 8802
rect 1168 8754 1204 8802
rect 1484 8754 1520 8802
rect 1800 8754 1836 8802
rect 2116 8754 2152 8802
rect 2432 8754 2468 8802
rect 2748 8754 2784 8802
rect 3064 8754 3100 8802
rect 3380 8754 3416 8802
rect 216 8742 262 8754
rect 216 7284 222 8742
rect 86 7282 222 7284
rect -2078 6694 -1938 6698
rect -2078 6594 -2058 6694
rect -1958 6594 -1938 6694
rect -1788 6616 -1778 6668
rect -1726 6616 -1716 6668
rect -2256 6472 -2116 6482
rect -2256 6372 -2238 6472
rect -2138 6372 -2116 6472
rect -2256 3652 -2116 6372
rect -2256 3552 -2238 3652
rect -2138 3552 -2116 3652
rect -2256 3538 -2116 3552
rect -2078 2998 -1938 6594
rect -1688 6558 -1654 6746
rect -1550 6616 -1540 6668
rect -1488 6616 -1478 6668
rect -1372 6558 -1338 6746
rect -1236 6616 -1226 6668
rect -1174 6616 -1164 6668
rect -1056 6558 -1022 6746
rect -918 6616 -908 6668
rect -856 6616 -846 6668
rect -740 6558 -706 6746
rect -604 6616 -594 6668
rect -542 6616 -532 6668
rect -424 6558 -390 6746
rect -360 6616 -350 6668
rect -298 6616 -288 6668
rect -116 6568 -106 6586
rect -1708 6506 -1698 6558
rect -1646 6506 -1636 6558
rect -1392 6506 -1382 6558
rect -1330 6506 -1320 6558
rect -1074 6506 -1064 6558
rect -1012 6506 -1002 6558
rect -758 6506 -748 6558
rect -696 6506 -686 6558
rect -442 6506 -432 6558
rect -380 6506 -370 6558
rect -1788 6398 -1778 6450
rect -1726 6398 -1716 6450
rect -1688 6320 -1654 6506
rect -1550 6398 -1540 6450
rect -1488 6398 -1478 6450
rect -1372 6320 -1338 6506
rect -1236 6398 -1226 6450
rect -1174 6398 -1164 6450
rect -1056 6320 -1022 6506
rect -918 6398 -908 6450
rect -856 6398 -846 6450
rect -740 6320 -706 6506
rect -604 6398 -594 6450
rect -542 6398 -532 6450
rect -424 6320 -390 6506
rect -122 6486 -106 6568
rect 0 6568 10 6586
rect 0 6486 18 6568
rect -360 6398 -350 6450
rect -298 6398 -288 6450
rect -1852 6308 -1806 6320
rect -1852 4332 -1846 6308
rect -1812 4332 -1806 6308
rect -1852 4320 -1806 4332
rect -1694 6308 -1648 6320
rect -1694 4332 -1688 6308
rect -1654 4332 -1648 6308
rect -1694 4320 -1648 4332
rect -1536 6308 -1490 6320
rect -1536 4332 -1530 6308
rect -1496 4332 -1490 6308
rect -1536 4320 -1490 4332
rect -1378 6308 -1332 6320
rect -1378 4332 -1372 6308
rect -1338 4332 -1332 6308
rect -1378 4320 -1332 4332
rect -1220 6308 -1174 6320
rect -1220 4332 -1214 6308
rect -1180 4332 -1174 6308
rect -1220 4320 -1174 4332
rect -1062 6308 -1016 6320
rect -1062 4332 -1056 6308
rect -1022 4332 -1016 6308
rect -1062 4320 -1016 4332
rect -904 6308 -858 6320
rect -904 4332 -898 6308
rect -864 4332 -858 6308
rect -904 4320 -858 4332
rect -746 6308 -700 6320
rect -746 4332 -740 6308
rect -706 4332 -700 6308
rect -746 4320 -700 4332
rect -588 6308 -542 6320
rect -588 4332 -582 6308
rect -548 4332 -542 6308
rect -588 4320 -542 4332
rect -430 6308 -384 6320
rect -430 4332 -424 6308
rect -390 4332 -384 6308
rect -430 4320 -384 4332
rect -272 6308 -226 6320
rect -272 4332 -266 6308
rect -232 4332 -226 6308
rect -122 4682 18 6486
rect 86 6334 92 7282
rect 144 6334 222 7282
rect 86 6322 150 6334
rect 216 4766 222 6334
rect 256 4766 262 8742
rect 216 4754 262 4766
rect 374 8742 420 8754
rect 374 4766 380 8742
rect 414 4766 420 8742
rect 374 4754 420 4766
rect 532 8742 578 8754
rect 532 4766 538 8742
rect 572 4766 578 8742
rect 532 4754 578 4766
rect 690 8742 736 8754
rect 690 4766 696 8742
rect 730 4766 736 8742
rect 690 4754 736 4766
rect 848 8742 894 8754
rect 848 4766 854 8742
rect 888 4766 894 8742
rect 848 4754 894 4766
rect 1006 8742 1052 8754
rect 1006 4766 1012 8742
rect 1046 4766 1052 8742
rect 1006 4754 1052 4766
rect 1164 8742 1210 8754
rect 1164 4766 1170 8742
rect 1204 4766 1210 8742
rect 1164 4754 1210 4766
rect 1322 8742 1368 8754
rect 1322 4766 1328 8742
rect 1362 4766 1368 8742
rect 1322 4754 1368 4766
rect 1480 8742 1526 8754
rect 1480 4766 1486 8742
rect 1520 4766 1526 8742
rect 1480 4754 1526 4766
rect 1638 8742 1684 8754
rect 1638 4766 1644 8742
rect 1678 4766 1684 8742
rect 1638 4754 1684 4766
rect 1796 8742 1842 8754
rect 1796 4766 1802 8742
rect 1836 4766 1842 8742
rect 1796 4754 1842 4766
rect 1954 8742 2000 8754
rect 1954 4766 1960 8742
rect 1994 4766 2000 8742
rect 1954 4754 2000 4766
rect 2112 8742 2158 8754
rect 2112 4766 2118 8742
rect 2152 4766 2158 8742
rect 2112 4754 2158 4766
rect 2270 8742 2316 8754
rect 2270 4766 2276 8742
rect 2310 4766 2316 8742
rect 2270 4754 2316 4766
rect 2428 8742 2474 8754
rect 2428 4766 2434 8742
rect 2468 4766 2474 8742
rect 2428 4754 2474 4766
rect 2586 8742 2632 8754
rect 2586 4766 2592 8742
rect 2626 4766 2632 8742
rect 2586 4754 2632 4766
rect 2744 8742 2790 8754
rect 2744 4766 2750 8742
rect 2784 4766 2790 8742
rect 2744 4754 2790 4766
rect 2902 8742 2948 8754
rect 2902 4766 2908 8742
rect 2942 4766 2948 8742
rect 2902 4754 2948 4766
rect 3060 8742 3106 8754
rect 3060 4766 3066 8742
rect 3100 4766 3106 8742
rect 3060 4754 3106 4766
rect 3218 8742 3264 8754
rect 3218 4766 3224 8742
rect 3258 4766 3264 8742
rect 3218 4754 3264 4766
rect 3376 8742 3422 8754
rect 3376 4766 3382 8742
rect 3416 7360 3422 8742
rect 3478 7360 3542 8802
rect 3416 6412 3484 7360
rect 3536 6412 3542 7360
rect 3416 6410 3542 6412
rect 3416 4766 3422 6410
rect 3478 6400 3542 6410
rect 3376 4754 3422 4766
rect -122 4582 -104 4682
rect 2 4582 18 4682
rect 266 4600 276 4666
rect 342 4600 352 4666
rect 380 4362 412 4754
rect 510 4600 520 4666
rect 586 4600 596 4666
rect -272 4320 -226 4332
rect -1846 4264 -1812 4320
rect -1530 4264 -1496 4320
rect -1214 4264 -1180 4320
rect -898 4264 -864 4320
rect -582 4264 -548 4320
rect -266 4264 -232 4320
rect 352 4296 362 4362
rect 428 4296 438 4362
rect 696 4360 728 4754
rect 826 4600 836 4666
rect 902 4600 912 4666
rect 1012 4360 1044 4754
rect 1142 4600 1152 4666
rect 1218 4600 1228 4666
rect 1328 4360 1360 4754
rect 1458 4600 1468 4666
rect 1534 4600 1544 4666
rect 1644 4360 1676 4754
rect 1776 4600 1786 4666
rect 1852 4600 1862 4666
rect 1960 4360 1992 4754
rect 2092 4600 2102 4666
rect 2168 4600 2178 4666
rect 2276 4360 2308 4754
rect 2406 4600 2416 4666
rect 2482 4600 2492 4666
rect 2592 4360 2624 4754
rect 2722 4600 2732 4666
rect 2798 4600 2808 4666
rect -1874 4228 160 4264
rect -1874 4162 -1762 4228
rect -324 4162 160 4228
rect 380 4206 412 4296
rect 670 4294 680 4360
rect 746 4294 756 4360
rect 986 4294 996 4360
rect 1062 4294 1072 4360
rect 1304 4294 1314 4360
rect 1380 4294 1390 4360
rect 1618 4294 1628 4360
rect 1694 4294 1704 4360
rect 1934 4294 1944 4360
rect 2010 4294 2020 4360
rect 2250 4294 2260 4360
rect 2326 4294 2336 4360
rect 2566 4294 2576 4360
rect 2642 4294 2652 4360
rect 2908 4358 2940 4754
rect 3040 4600 3050 4666
rect 3116 4600 3126 4666
rect 3224 4358 3256 4754
rect 3298 4600 3308 4666
rect 3374 4600 3384 4666
rect 696 4206 728 4294
rect 1012 4206 1044 4294
rect 1328 4206 1360 4294
rect 1644 4206 1676 4294
rect 1960 4206 1992 4294
rect 2276 4206 2308 4294
rect 2592 4206 2624 4294
rect 2882 4292 2892 4358
rect 2958 4292 2968 4358
rect 3198 4292 3208 4358
rect 3274 4292 3284 4358
rect 2908 4206 2940 4292
rect 3224 4206 3256 4292
rect -1874 4106 160 4162
rect -1874 4092 -1082 4106
rect -1903 4086 -1082 4092
rect -1903 4040 -1891 4086
rect -1369 4040 -1082 4086
rect -1903 4034 -1082 4040
rect -1883 3985 -1849 4034
rect -1691 3985 -1657 4034
rect -1499 3985 -1465 4034
rect -1150 4016 -1082 4034
rect -82 4016 160 4106
rect -1150 4010 160 4016
rect -1889 3973 -1843 3985
rect -1889 3797 -1883 3973
rect -1849 3797 -1843 3973
rect -1889 3785 -1843 3797
rect -1793 3973 -1747 3985
rect -1793 3797 -1787 3973
rect -1753 3797 -1747 3973
rect -1793 3785 -1747 3797
rect -1697 3973 -1651 3985
rect -1697 3797 -1691 3973
rect -1657 3797 -1651 3973
rect -1697 3785 -1651 3797
rect -1601 3973 -1555 3985
rect -1601 3797 -1595 3973
rect -1561 3797 -1555 3973
rect -1601 3785 -1555 3797
rect -1505 3973 -1459 3985
rect -1505 3797 -1499 3973
rect -1465 3797 -1459 3973
rect -1505 3785 -1459 3797
rect -1409 3973 -1363 3985
rect -1409 3797 -1403 3973
rect -1369 3797 -1363 3973
rect -1409 3785 -1363 3797
rect -1150 3920 -1104 4010
rect -1785 3757 -1755 3785
rect -1593 3757 -1563 3785
rect -1805 3705 -1795 3757
rect -1743 3705 -1733 3757
rect -1613 3705 -1603 3757
rect -1551 3705 -1541 3757
rect -1401 3756 -1371 3785
rect -1879 3618 -1821 3624
rect -1879 3617 -1867 3618
rect -1833 3617 -1821 3618
rect -1886 3565 -1876 3617
rect -1824 3565 -1814 3617
rect -1785 3534 -1755 3705
rect -1703 3618 -1645 3624
rect -1703 3616 -1691 3618
rect -1657 3616 -1645 3618
rect -1710 3564 -1700 3616
rect -1648 3564 -1638 3616
rect -1593 3534 -1563 3705
rect -1422 3704 -1412 3756
rect -1360 3704 -1350 3756
rect -1511 3615 -1453 3621
rect -1511 3614 -1499 3615
rect -1465 3614 -1453 3615
rect -1517 3562 -1507 3614
rect -1455 3562 -1445 3614
rect -1401 3534 -1371 3704
rect -1889 3522 -1843 3534
rect -1889 3346 -1883 3522
rect -1849 3346 -1843 3522
rect -1889 3334 -1843 3346
rect -1793 3522 -1747 3534
rect -1793 3346 -1787 3522
rect -1753 3346 -1747 3522
rect -1793 3334 -1747 3346
rect -1697 3522 -1651 3534
rect -1697 3346 -1691 3522
rect -1657 3346 -1651 3522
rect -1697 3334 -1651 3346
rect -1601 3522 -1555 3534
rect -1601 3346 -1595 3522
rect -1561 3346 -1555 3522
rect -1601 3334 -1555 3346
rect -1505 3522 -1459 3534
rect -1505 3346 -1499 3522
rect -1465 3346 -1459 3522
rect -1505 3334 -1459 3346
rect -1409 3522 -1363 3534
rect -1409 3346 -1403 3522
rect -1369 3346 -1363 3522
rect -1409 3334 -1363 3346
rect -1883 3270 -1849 3334
rect -1691 3270 -1657 3334
rect -1499 3270 -1465 3334
rect -1883 3268 -1318 3270
rect -1906 3262 -1318 3268
rect -1906 3226 -1894 3262
rect -1359 3226 -1318 3262
rect -1906 3220 -1318 3226
rect -1876 3184 -1318 3220
rect -1150 3144 -1144 3920
rect -1110 3144 -1104 3920
rect -1150 3132 -1104 3144
rect -992 3920 -946 3932
rect -992 3144 -986 3920
rect -952 3144 -946 3920
rect -992 3132 -946 3144
rect -834 3920 -788 4010
rect -654 3932 -622 3934
rect -834 3144 -828 3920
rect -794 3144 -788 3920
rect -834 3132 -788 3144
rect -676 3920 -622 3932
rect -676 3144 -670 3920
rect -636 3144 -622 3920
rect -676 3132 -622 3144
rect -536 3920 -490 4010
rect -536 3144 -530 3920
rect -496 3144 -490 3920
rect -536 3132 -490 3144
rect -378 3920 -332 3932
rect -378 3144 -372 3920
rect -338 3144 -332 3920
rect -378 3132 -332 3144
rect -220 3920 -174 4010
rect -220 3144 -214 3920
rect -180 3144 -174 3920
rect -220 3132 -174 3144
rect -62 3920 -16 3932
rect -62 3144 -56 3920
rect -22 3144 -16 3920
rect -62 3132 -16 3144
rect -1082 3058 -1072 3110
rect -1020 3058 -1010 3110
rect -1082 3056 -1010 3058
rect -1076 3052 -1018 3056
rect -982 2998 -952 3132
rect -924 3058 -914 3110
rect -862 3058 -852 3110
rect -766 3058 -756 3110
rect -704 3058 -694 3110
rect -918 3054 -860 3058
rect -758 3054 -700 3058
rect -654 2998 -622 3132
rect -472 3058 -462 3110
rect -410 3058 -400 3110
rect -464 3054 -406 3058
rect -2078 2944 -622 2998
rect -370 2956 -338 3132
rect -310 3058 -300 3110
rect -248 3058 -238 3110
rect -154 3058 -144 3110
rect -92 3058 -82 3110
rect -302 3054 -244 3058
rect -146 3054 -88 3058
rect -380 2946 -338 2956
rect -2446 2892 -2254 2904
rect -2446 2832 -2434 2892
rect -2374 2832 -2326 2892
rect -2266 2832 -2254 2892
rect -772 2864 -762 2916
rect -710 2864 -700 2916
rect -772 2859 -700 2864
rect -2446 2822 -2254 2832
rect -782 2853 -690 2859
rect -782 2819 -770 2853
rect -702 2819 -690 2853
rect -782 2813 -690 2819
rect -654 2854 -622 2944
rect -390 2894 -380 2946
rect -328 2936 -318 2946
rect -54 2936 -16 3132
rect -328 2902 -16 2936
rect -328 2894 -318 2902
rect -380 2882 -338 2894
rect -492 2854 -400 2859
rect -654 2853 -400 2854
rect -654 2819 -480 2853
rect -412 2819 -400 2853
rect -654 2818 -472 2819
rect -654 2772 -622 2818
rect -492 2813 -472 2818
rect -482 2792 -472 2813
rect -420 2813 -400 2819
rect -420 2792 -410 2813
rect -370 2772 -338 2882
rect -838 2760 -792 2772
rect -838 2384 -832 2760
rect -798 2384 -792 2760
rect -838 2372 -792 2384
rect -680 2760 -622 2772
rect -680 2384 -674 2760
rect -640 2384 -622 2760
rect -680 2372 -622 2384
rect -548 2760 -502 2772
rect -548 2384 -542 2760
rect -508 2384 -502 2760
rect -548 2372 -502 2384
rect -390 2760 -338 2772
rect -390 2384 -384 2760
rect -350 2384 -338 2760
rect -390 2372 -338 2384
rect 20 2746 160 4010
rect 216 4194 262 4206
rect 216 2746 222 4194
rect -832 2314 -798 2372
rect -542 2314 -508 2372
rect -832 2308 -766 2314
rect -706 2308 -620 2314
rect -560 2308 -466 2314
rect -406 2308 -352 2314
rect -832 2266 -772 2308
rect -394 2266 -352 2308
rect -832 2256 -766 2266
rect -776 2254 -766 2256
rect -706 2256 -620 2266
rect -706 2254 -696 2256
rect -630 2254 -620 2256
rect -560 2256 -466 2266
rect -560 2254 -550 2256
rect -476 2254 -466 2256
rect -406 2256 -352 2266
rect -406 2254 -396 2256
rect 20 1798 222 2746
rect 20 128 160 1798
rect 216 218 222 1798
rect 256 218 262 4194
rect 216 206 262 218
rect 374 4194 420 4206
rect 374 218 380 4194
rect 414 218 420 4194
rect 374 206 420 218
rect 532 4194 578 4206
rect 532 218 538 4194
rect 572 218 578 4194
rect 532 206 578 218
rect 690 4194 736 4206
rect 690 218 696 4194
rect 730 218 736 4194
rect 690 206 736 218
rect 848 4194 894 4206
rect 848 218 854 4194
rect 888 218 894 4194
rect 848 206 894 218
rect 1006 4194 1052 4206
rect 1006 218 1012 4194
rect 1046 218 1052 4194
rect 1006 206 1052 218
rect 1164 4194 1210 4206
rect 1164 218 1170 4194
rect 1204 218 1210 4194
rect 1164 206 1210 218
rect 1322 4194 1368 4206
rect 1322 218 1328 4194
rect 1362 218 1368 4194
rect 1322 206 1368 218
rect 1480 4194 1526 4206
rect 1480 218 1486 4194
rect 1520 218 1526 4194
rect 1480 206 1526 218
rect 1638 4194 1684 4206
rect 1638 218 1644 4194
rect 1678 218 1684 4194
rect 1638 206 1684 218
rect 1796 4194 1842 4206
rect 1796 218 1802 4194
rect 1836 218 1842 4194
rect 1796 206 1842 218
rect 1954 4194 2000 4206
rect 1954 218 1960 4194
rect 1994 218 2000 4194
rect 1954 206 2000 218
rect 2112 4194 2158 4206
rect 2112 218 2118 4194
rect 2152 218 2158 4194
rect 2112 206 2158 218
rect 2270 4194 2316 4206
rect 2270 218 2276 4194
rect 2310 218 2316 4194
rect 2270 206 2316 218
rect 2428 4194 2474 4206
rect 2428 218 2434 4194
rect 2468 218 2474 4194
rect 2428 206 2474 218
rect 2586 4194 2632 4206
rect 2586 218 2592 4194
rect 2626 218 2632 4194
rect 2586 206 2632 218
rect 2744 4194 2790 4206
rect 2744 218 2750 4194
rect 2784 218 2790 4194
rect 2744 206 2790 218
rect 2902 4194 2948 4206
rect 2902 218 2908 4194
rect 2942 218 2948 4194
rect 2902 206 2948 218
rect 3060 4194 3106 4206
rect 3060 218 3066 4194
rect 3100 218 3106 4194
rect 3060 206 3106 218
rect 3218 4194 3264 4206
rect 3218 218 3224 4194
rect 3258 218 3264 4194
rect 3218 206 3264 218
rect 3376 4194 3422 4206
rect 3376 218 3382 4194
rect 3416 2796 3422 4194
rect 3416 1866 3542 2796
rect 3416 1848 3554 1866
rect 3416 218 3422 1848
rect 3376 206 3422 218
rect 222 128 256 206
rect 536 128 570 206
rect 854 128 888 206
rect 1168 128 1202 206
rect 1486 128 1520 206
rect 1800 128 1834 206
rect 2118 128 2152 206
rect 2432 128 2466 206
rect 2750 128 2784 206
rect 3064 128 3098 206
rect 3382 128 3416 206
rect 3500 128 3554 1848
rect 20 114 3554 128
rect 20 8 188 114
rect 3452 8 3554 114
rect 20 0 3554 8
<< via1 >>
rect -2058 6594 -1958 6694
rect -1778 6658 -1726 6668
rect -1778 6624 -1768 6658
rect -1768 6624 -1734 6658
rect -1734 6624 -1726 6658
rect -1778 6616 -1726 6624
rect -2238 6372 -2138 6472
rect -2238 3552 -2138 3652
rect -1540 6660 -1488 6668
rect -1540 6626 -1530 6660
rect -1530 6626 -1496 6660
rect -1496 6626 -1488 6660
rect -1540 6616 -1488 6626
rect -1226 6660 -1174 6668
rect -1226 6626 -1216 6660
rect -1216 6626 -1182 6660
rect -1182 6626 -1174 6660
rect -1226 6616 -1174 6626
rect -908 6658 -856 6668
rect -908 6624 -898 6658
rect -898 6624 -864 6658
rect -864 6624 -856 6658
rect -908 6616 -856 6624
rect -594 6658 -542 6668
rect -594 6624 -584 6658
rect -584 6624 -550 6658
rect -550 6624 -542 6658
rect -594 6616 -542 6624
rect -350 6658 -298 6668
rect -350 6624 -340 6658
rect -340 6624 -306 6658
rect -306 6624 -298 6658
rect -350 6616 -298 6624
rect -1698 6506 -1646 6558
rect -1382 6506 -1330 6558
rect -1064 6506 -1012 6558
rect -748 6506 -696 6558
rect -432 6506 -380 6558
rect -1778 6440 -1726 6450
rect -1778 6406 -1768 6440
rect -1768 6406 -1734 6440
rect -1734 6406 -1726 6440
rect -1778 6398 -1726 6406
rect -1540 6442 -1488 6450
rect -1540 6408 -1530 6442
rect -1530 6408 -1496 6442
rect -1496 6408 -1488 6442
rect -1540 6398 -1488 6408
rect -1226 6442 -1174 6450
rect -1226 6408 -1216 6442
rect -1216 6408 -1182 6442
rect -1182 6408 -1174 6442
rect -1226 6398 -1174 6408
rect -908 6440 -856 6450
rect -908 6406 -898 6440
rect -898 6406 -864 6440
rect -864 6406 -856 6440
rect -908 6398 -856 6406
rect -594 6440 -542 6450
rect -594 6406 -584 6440
rect -584 6406 -550 6440
rect -550 6406 -542 6440
rect -594 6398 -542 6406
rect -106 6486 0 6586
rect -350 6440 -298 6450
rect -350 6406 -340 6440
rect -340 6406 -306 6440
rect -306 6406 -298 6440
rect -350 6398 -298 6406
rect -104 4582 2 4682
rect 276 4650 342 4666
rect 276 4616 292 4650
rect 292 4616 326 4650
rect 326 4616 342 4650
rect 276 4600 342 4616
rect 520 4650 586 4666
rect 520 4616 536 4650
rect 536 4616 570 4650
rect 570 4616 586 4650
rect 520 4600 586 4616
rect 362 4296 428 4362
rect 836 4650 902 4666
rect 836 4616 852 4650
rect 852 4616 886 4650
rect 886 4616 902 4650
rect 836 4600 902 4616
rect 1152 4650 1218 4666
rect 1152 4616 1168 4650
rect 1168 4616 1202 4650
rect 1202 4616 1218 4650
rect 1152 4600 1218 4616
rect 1468 4650 1534 4666
rect 1468 4616 1484 4650
rect 1484 4616 1518 4650
rect 1518 4616 1534 4650
rect 1468 4600 1534 4616
rect 1786 4650 1852 4666
rect 1786 4616 1802 4650
rect 1802 4616 1836 4650
rect 1836 4616 1852 4650
rect 1786 4600 1852 4616
rect 2102 4650 2168 4666
rect 2102 4616 2118 4650
rect 2118 4616 2152 4650
rect 2152 4616 2168 4650
rect 2102 4600 2168 4616
rect 2416 4650 2482 4666
rect 2416 4616 2432 4650
rect 2432 4616 2466 4650
rect 2466 4616 2482 4650
rect 2416 4600 2482 4616
rect 2732 4650 2798 4666
rect 2732 4616 2748 4650
rect 2748 4616 2782 4650
rect 2782 4616 2798 4650
rect 2732 4600 2798 4616
rect 680 4294 746 4360
rect 996 4294 1062 4360
rect 1314 4294 1380 4360
rect 1628 4294 1694 4360
rect 1944 4294 2010 4360
rect 2260 4294 2326 4360
rect 2576 4294 2642 4360
rect 3050 4650 3116 4666
rect 3050 4616 3066 4650
rect 3066 4616 3100 4650
rect 3100 4616 3116 4650
rect 3050 4600 3116 4616
rect 3308 4650 3374 4666
rect 3308 4616 3324 4650
rect 3324 4616 3358 4650
rect 3358 4616 3374 4650
rect 3308 4600 3374 4616
rect 2892 4292 2958 4358
rect 3208 4292 3274 4358
rect -1795 3705 -1743 3757
rect -1603 3705 -1551 3757
rect -1876 3584 -1867 3617
rect -1867 3584 -1833 3617
rect -1833 3584 -1824 3617
rect -1876 3565 -1824 3584
rect -1700 3584 -1691 3616
rect -1691 3584 -1657 3616
rect -1657 3584 -1648 3616
rect -1700 3564 -1648 3584
rect -1412 3704 -1360 3756
rect -1507 3581 -1499 3614
rect -1499 3581 -1465 3614
rect -1465 3581 -1455 3614
rect -1507 3562 -1455 3581
rect -1072 3092 -1020 3110
rect -1072 3058 -1064 3092
rect -1064 3058 -1030 3092
rect -1030 3058 -1020 3092
rect -914 3094 -862 3110
rect -914 3060 -906 3094
rect -906 3060 -872 3094
rect -872 3060 -862 3094
rect -914 3058 -862 3060
rect -756 3094 -704 3110
rect -756 3060 -746 3094
rect -746 3060 -712 3094
rect -712 3060 -704 3094
rect -756 3058 -704 3060
rect -462 3094 -410 3110
rect -462 3060 -452 3094
rect -452 3060 -418 3094
rect -418 3060 -410 3094
rect -462 3058 -410 3060
rect -300 3094 -248 3110
rect -300 3060 -290 3094
rect -290 3060 -256 3094
rect -256 3060 -248 3094
rect -300 3058 -248 3060
rect -144 3094 -92 3110
rect -144 3060 -134 3094
rect -134 3060 -100 3094
rect -100 3060 -92 3094
rect -144 3058 -92 3060
rect -2434 2832 -2374 2892
rect -2326 2832 -2266 2892
rect -762 2864 -710 2916
rect -380 2894 -328 2946
rect -472 2819 -420 2844
rect -472 2792 -420 2819
rect -766 2308 -706 2314
rect -620 2308 -560 2314
rect -466 2308 -406 2314
rect -766 2266 -706 2308
rect -620 2266 -560 2308
rect -466 2266 -406 2308
rect -766 2254 -706 2266
rect -620 2254 -560 2266
rect -466 2254 -406 2266
<< metal2 >>
rect -2058 6694 -1958 6704
rect -1958 6668 -156 6682
rect -1958 6616 -1778 6668
rect -1726 6616 -1540 6668
rect -1488 6616 -1226 6668
rect -1174 6616 -908 6668
rect -856 6616 -594 6668
rect -542 6616 -350 6668
rect -298 6616 -156 6668
rect -1958 6604 -156 6616
rect -1778 6602 -156 6604
rect -2058 6584 -1958 6594
rect -106 6586 0 6596
rect -1928 6558 -106 6572
rect -1928 6506 -1698 6558
rect -1646 6506 -1382 6558
rect -1330 6506 -1064 6558
rect -1012 6506 -748 6558
rect -696 6506 -432 6558
rect -380 6506 -106 6558
rect -1928 6492 -106 6506
rect -2238 6472 -2138 6482
rect -106 6476 0 6486
rect -2242 6384 -2238 6462
rect -2138 6450 -156 6462
rect -2138 6398 -1778 6450
rect -1726 6398 -1540 6450
rect -1488 6398 -1226 6450
rect -1174 6398 -908 6450
rect -856 6398 -594 6450
rect -542 6398 -350 6450
rect -298 6398 -156 6450
rect -2138 6384 -156 6398
rect -2238 6362 -2138 6372
rect -104 4682 2 4692
rect 2 4666 3460 4682
rect 2 4600 276 4666
rect 342 4600 520 4666
rect 586 4600 836 4666
rect 902 4600 1152 4666
rect 1218 4600 1468 4666
rect 1534 4600 1786 4666
rect 1852 4600 2102 4666
rect 2168 4600 2416 4666
rect 2482 4600 2732 4666
rect 2798 4600 3050 4666
rect 3116 4600 3308 4666
rect 3374 4600 3460 4666
rect 2 4582 3460 4600
rect -104 4572 2 4582
rect 170 4362 3460 4378
rect 170 4296 362 4362
rect 428 4360 3460 4362
rect 428 4296 680 4360
rect 170 4294 680 4296
rect 746 4294 996 4360
rect 1062 4294 1314 4360
rect 1380 4294 1628 4360
rect 1694 4294 1944 4360
rect 2010 4294 2260 4360
rect 2326 4294 2576 4360
rect 2642 4358 3460 4360
rect 2642 4294 2892 4358
rect 170 4292 2892 4294
rect 2958 4292 3208 4358
rect 3274 4292 3460 4358
rect 170 4278 3460 4292
rect -1795 3758 -1743 3767
rect -1603 3758 -1551 3767
rect -1412 3758 -1360 3766
rect -1897 3757 -1160 3758
rect -1897 3744 -1795 3757
rect -1932 3716 -1795 3744
rect -1897 3705 -1795 3716
rect -1743 3705 -1603 3757
rect -1551 3756 -1160 3757
rect -1551 3705 -1412 3756
rect -1795 3695 -1743 3705
rect -1603 3695 -1551 3705
rect -1360 3705 -1160 3756
rect -1412 3694 -1360 3704
rect -2238 3652 -2138 3658
rect -2138 3617 -1252 3628
rect -2138 3568 -1876 3617
rect -1824 3616 -1252 3617
rect -1824 3568 -1700 3616
rect -1876 3555 -1824 3565
rect -1648 3614 -1252 3616
rect -1648 3568 -1507 3614
rect -1700 3554 -1648 3564
rect -1455 3568 -1252 3614
rect -1507 3552 -1455 3562
rect -2238 3538 -2138 3552
rect -1312 3020 -1252 3568
rect -1220 3102 -1160 3705
rect -1072 3110 -1020 3120
rect -1220 3068 -1072 3102
rect -914 3110 -862 3120
rect -1020 3068 -914 3102
rect -1072 3048 -1020 3058
rect -756 3110 -704 3120
rect -862 3068 -756 3102
rect -914 3048 -862 3058
rect -462 3110 -410 3120
rect -704 3068 -694 3102
rect -756 3048 -704 3058
rect -462 3020 -410 3058
rect -300 3110 -248 3120
rect -300 3020 -248 3058
rect -144 3110 -92 3120
rect -144 3020 -92 3058
rect -1312 2986 -92 3020
rect -380 2946 -328 2956
rect -762 2916 -380 2936
rect -2446 2892 -2254 2904
rect -2446 2832 -2434 2892
rect -2374 2832 -2326 2892
rect -2266 2832 -906 2892
rect -710 2902 -380 2916
rect -380 2882 -328 2894
rect -762 2854 -710 2864
rect -2446 2822 -2254 2832
rect -948 2312 -906 2832
rect -496 2844 -272 2854
rect -496 2820 -472 2844
rect -420 2820 -272 2844
rect -472 2760 -420 2792
rect -766 2314 -706 2324
rect -948 2254 -766 2312
rect -620 2314 -560 2324
rect -706 2254 -620 2312
rect -466 2314 -406 2324
rect -560 2254 -466 2312
rect -406 2254 -322 2312
rect -928 2252 -322 2254
rect -766 2244 -706 2252
rect -620 2244 -560 2252
rect -466 2244 -406 2252
<< labels >>
rlabel metal1 -1876 3184 -1318 3270 1 VDD
rlabel metal1 -1870 8806 3274 8896 1 VH
rlabel metal1 -2256 3648 -2116 6372 1 IN
rlabel metal1 20 0 160 4264 1 GND
rlabel space 3274 4278 3460 4378 1 OUT
rlabel space 142 0 3496 8930 1 OUT
rlabel metal1 -1870 8864 -208 8870 1 stage_100_0/VH
rlabel metal2 -380 6492 -158 6572 1 stage_100_0/OUT
rlabel metal1 -1846 4154 -232 4160 1 stage_100_0/GND
rlabel space -1926 6602 -1778 6682 1 stage_100_0/A
rlabel metal2 -1926 6384 -1778 6462 1 stage_100_0/B
rlabel metal2 170 4582 276 4682 1 inv_400_0/IN
rlabel metal2 3274 4278 3460 4378 1 inv_400_0/OUT
rlabel metal1 -1903 4086 -1357 4092 5 inv_1_8_0/GND
rlabel metal2 -1360 3716 -1321 3744 5 inv_1_8_0/OUT
rlabel metal2 -1931 3576 -1876 3604 5 inv_1_8_0/IN
rlabel metal1 -1906 3220 -1347 3226 5 inv_1_8_0/VDD
rlabel metal2 -420 2820 -272 2854 5 cruzados_0/OUT
rlabel metal1 -832 2256 -352 2262 5 cruzados_0/VH
rlabel metal2 -1156 3068 -1072 3102 5 cruzados_0/IN1
rlabel metal2 -906 2986 -470 3020 5 cruzados_0/IN2
<< end >>
