magic
tech sky130A
timestamp 1668450285
<< metal5 >>
rect 3500 10000 6500 22500
rect 0 0 10000 10000
<< glass >>
rect 20 20 9980 9980
use stack30um_1_5  stack30um_1_5_0
timestamp 1668366526
transform 1 0 3500 0 1 19500
box 0 0 3000 3000
<< end >>
