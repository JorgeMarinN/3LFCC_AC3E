* NGSPICE file created from user_analog_project_wrapper.ext - technology: sky130A

.subckt unit_cap c2_30_30# c1_30_30# m3_0_0#
X0 c1_30_30# m3_0_0# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X1 c2_30_30# c1_30_30# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
.ends

.subckt stack_2um_1_5 m1_0_0#
R0 m1_0_0# m1_0_0# sky130_fd_pr__res_generic_m1 w=800000u l=0u
.ends

.subckt stack30um_1_5 m5_0_0#
Xstack_2um_1_5_40 m5_0_0# stack_2um_1_5
Xstack_2um_1_5_51 m5_0_0# stack_2um_1_5
Xstack_2um_1_5_50 m5_0_0# stack_2um_1_5
Xstack_2um_1_5_52 m5_0_0# stack_2um_1_5
Xstack_2um_1_5_41 m5_0_0# stack_2um_1_5
Xstack_2um_1_5_30 m5_0_0# stack_2um_1_5
Xstack_2um_1_5_20 m5_0_0# stack_2um_1_5
Xstack_2um_1_5_53 m5_0_0# stack_2um_1_5
Xstack_2um_1_5_42 m5_0_0# stack_2um_1_5
Xstack_2um_1_5_31 m5_0_0# stack_2um_1_5
Xstack_2um_1_5_10 m5_0_0# stack_2um_1_5
Xstack_2um_1_5_21 m5_0_0# stack_2um_1_5
Xstack_2um_1_5_54 m5_0_0# stack_2um_1_5
Xstack_2um_1_5_43 m5_0_0# stack_2um_1_5
Xstack_2um_1_5_32 m5_0_0# stack_2um_1_5
Xstack_2um_1_5_0 m5_0_0# stack_2um_1_5
Xstack_2um_1_5_55 m5_0_0# stack_2um_1_5
Xstack_2um_1_5_44 m5_0_0# stack_2um_1_5
Xstack_2um_1_5_33 m5_0_0# stack_2um_1_5
Xstack_2um_1_5_2 m5_0_0# stack_2um_1_5
Xstack_2um_1_5_1 m5_0_0# stack_2um_1_5
Xstack_2um_1_5_22 m5_0_0# stack_2um_1_5
Xstack_2um_1_5_11 m5_0_0# stack_2um_1_5
Xstack_2um_1_5_3 m5_0_0# stack_2um_1_5
Xstack_2um_1_5_23 m5_0_0# stack_2um_1_5
Xstack_2um_1_5_12 m5_0_0# stack_2um_1_5
Xstack_2um_1_5_34 m5_0_0# stack_2um_1_5
Xstack_2um_1_5_45 m5_0_0# stack_2um_1_5
Xstack_2um_1_5_24 m5_0_0# stack_2um_1_5
Xstack_2um_1_5_13 m5_0_0# stack_2um_1_5
Xstack_2um_1_5_35 m5_0_0# stack_2um_1_5
Xstack_2um_1_5_46 m5_0_0# stack_2um_1_5
Xstack_2um_1_5_4 m5_0_0# stack_2um_1_5
Xstack_2um_1_5_25 m5_0_0# stack_2um_1_5
Xstack_2um_1_5_14 m5_0_0# stack_2um_1_5
Xstack_2um_1_5_36 m5_0_0# stack_2um_1_5
Xstack_2um_1_5_47 m5_0_0# stack_2um_1_5
Xstack_2um_1_5_5 m5_0_0# stack_2um_1_5
Xstack_2um_1_5_48 m5_0_0# stack_2um_1_5
Xstack_2um_1_5_6 m5_0_0# stack_2um_1_5
Xstack_2um_1_5_38 m5_0_0# stack_2um_1_5
Xstack_2um_1_5_27 m5_0_0# stack_2um_1_5
Xstack_2um_1_5_49 m5_0_0# stack_2um_1_5
Xstack_2um_1_5_16 m5_0_0# stack_2um_1_5
Xstack_2um_1_5_37 m5_0_0# stack_2um_1_5
Xstack_2um_1_5_26 m5_0_0# stack_2um_1_5
Xstack_2um_1_5_15 m5_0_0# stack_2um_1_5
Xstack_2um_1_5_39 m5_0_0# stack_2um_1_5
Xstack_2um_1_5_28 m5_0_0# stack_2um_1_5
Xstack_2um_1_5_17 m5_0_0# stack_2um_1_5
Xstack_2um_1_5_7 m5_0_0# stack_2um_1_5
Xstack_2um_1_5_29 m5_0_0# stack_2um_1_5
Xstack_2um_1_5_18 m5_0_0# stack_2um_1_5
Xstack_2um_1_5_8 m5_0_0# stack_2um_1_5
Xstack_2um_1_5_9 m5_0_0# stack_2um_1_5
Xstack_2um_1_5_19 m5_0_0# stack_2um_1_5
.ends

.subckt power_pad_1_5 m5_0_0#
Xstack30um_1_5_29 m5_0_0# stack30um_1_5
Xstack30um_1_5_19 m5_0_0# stack30um_1_5
Xstack30um_1_5_18 m5_0_0# stack30um_1_5
Xstack30um_1_5_0 m5_0_0# stack30um_1_5
Xstack30um_1_5_1 m5_0_0# stack30um_1_5
Xstack30um_1_5_2 m5_0_0# stack30um_1_5
Xstack30um_1_5_3 m5_0_0# stack30um_1_5
Xstack30um_1_5_4 m5_0_0# stack30um_1_5
Xstack30um_1_5_5 m5_0_0# stack30um_1_5
Xstack30um_1_5_6 m5_0_0# stack30um_1_5
Xstack30um_1_5_8 m5_0_0# stack30um_1_5
Xstack30um_1_5_7 m5_0_0# stack30um_1_5
Xstack30um_1_5_9 m5_0_0# stack30um_1_5
Xstack30um_1_5_20 m5_0_0# stack30um_1_5
Xstack30um_1_5_21 m5_0_0# stack30um_1_5
Xstack30um_1_5_10 m5_0_0# stack30um_1_5
Xstack30um_1_5_11 m5_0_0# stack30um_1_5
Xstack30um_1_5_22 m5_0_0# stack30um_1_5
Xstack30um_1_5_23 m5_0_0# stack30um_1_5
Xstack30um_1_5_12 m5_0_0# stack30um_1_5
Xstack30um_1_5_24 m5_0_0# stack30um_1_5
Xstack30um_1_5_13 m5_0_0# stack30um_1_5
Xstack30um_1_5_14 m5_0_0# stack30um_1_5
Xstack30um_1_5_25 m5_0_0# stack30um_1_5
Xstack30um_1_5_26 m5_0_0# stack30um_1_5
Xstack30um_1_5_15 m5_0_0# stack30um_1_5
Xstack30um_1_5_27 m5_0_0# stack30um_1_5
Xstack30um_1_5_16 m5_0_0# stack30um_1_5
Xstack30um_1_5_17 m5_0_0# stack30um_1_5
Xstack30um_1_5_28 m5_0_0# stack30um_1_5
.ends

.subckt stack_2um_3_5 m3_0_0#
R0 m3_0_0# m3_0_0# sky130_fd_pr__res_generic_m3 w=800000u l=0u
.ends

.subckt stack30um_3_5 m5_0_0#
Xstack_2um_3_5_48 m5_0_0# stack_2um_3_5
Xstack_2um_3_5_6 m5_0_0# stack_2um_3_5
Xstack_2um_3_5_37 m5_0_0# stack_2um_3_5
Xstack_2um_3_5_26 m5_0_0# stack_2um_3_5
Xstack_2um_3_5_15 m5_0_0# stack_2um_3_5
Xstack_2um_3_5_38 m5_0_0# stack_2um_3_5
Xstack_2um_3_5_27 m5_0_0# stack_2um_3_5
Xstack_2um_3_5_49 m5_0_0# stack_2um_3_5
Xstack_2um_3_5_16 m5_0_0# stack_2um_3_5
Xstack_2um_3_5_7 m5_0_0# stack_2um_3_5
Xstack_2um_3_5_29 m5_0_0# stack_2um_3_5
Xstack_2um_3_5_18 m5_0_0# stack_2um_3_5
Xstack_2um_3_5_39 m5_0_0# stack_2um_3_5
Xstack_2um_3_5_28 m5_0_0# stack_2um_3_5
Xstack_2um_3_5_17 m5_0_0# stack_2um_3_5
Xstack_2um_3_5_8 m5_0_0# stack_2um_3_5
Xstack_2um_3_5_9 m5_0_0# stack_2um_3_5
Xstack_2um_3_5_19 m5_0_0# stack_2um_3_5
Xstack_2um_3_5_50 m5_0_0# stack_2um_3_5
Xstack_2um_3_5_40 m5_0_0# stack_2um_3_5
Xstack_2um_3_5_51 m5_0_0# stack_2um_3_5
Xstack_2um_3_5_20 m5_0_0# stack_2um_3_5
Xstack_2um_3_5_53 m5_0_0# stack_2um_3_5
Xstack_2um_3_5_42 m5_0_0# stack_2um_3_5
Xstack_2um_3_5_31 m5_0_0# stack_2um_3_5
Xstack_2um_3_5_52 m5_0_0# stack_2um_3_5
Xstack_2um_3_5_41 m5_0_0# stack_2um_3_5
Xstack_2um_3_5_30 m5_0_0# stack_2um_3_5
Xstack_2um_3_5_10 m5_0_0# stack_2um_3_5
Xstack_2um_3_5_21 m5_0_0# stack_2um_3_5
Xstack_2um_3_5_54 m5_0_0# stack_2um_3_5
Xstack_2um_3_5_43 m5_0_0# stack_2um_3_5
Xstack_2um_3_5_32 m5_0_0# stack_2um_3_5
Xstack_2um_3_5_0 m5_0_0# stack_2um_3_5
Xstack_2um_3_5_55 m5_0_0# stack_2um_3_5
Xstack_2um_3_5_44 m5_0_0# stack_2um_3_5
Xstack_2um_3_5_33 m5_0_0# stack_2um_3_5
Xstack_2um_3_5_1 m5_0_0# stack_2um_3_5
Xstack_2um_3_5_22 m5_0_0# stack_2um_3_5
Xstack_2um_3_5_11 m5_0_0# stack_2um_3_5
Xstack_2um_3_5_2 m5_0_0# stack_2um_3_5
Xstack_2um_3_5_23 m5_0_0# stack_2um_3_5
Xstack_2um_3_5_12 m5_0_0# stack_2um_3_5
Xstack_2um_3_5_34 m5_0_0# stack_2um_3_5
Xstack_2um_3_5_45 m5_0_0# stack_2um_3_5
Xstack_2um_3_5_3 m5_0_0# stack_2um_3_5
Xstack_2um_3_5_24 m5_0_0# stack_2um_3_5
Xstack_2um_3_5_13 m5_0_0# stack_2um_3_5
Xstack_2um_3_5_35 m5_0_0# stack_2um_3_5
Xstack_2um_3_5_46 m5_0_0# stack_2um_3_5
Xstack_2um_3_5_25 m5_0_0# stack_2um_3_5
Xstack_2um_3_5_14 m5_0_0# stack_2um_3_5
Xstack_2um_3_5_36 m5_0_0# stack_2um_3_5
Xstack_2um_3_5_47 m5_0_0# stack_2um_3_5
Xstack_2um_3_5_5 m5_0_0# stack_2um_3_5
Xstack_2um_3_5_4 m5_0_0# stack_2um_3_5
.ends

.subckt power_pad_3_5 m5_0_0#
Xstack30um_3_5_20 m5_0_0# stack30um_3_5
Xstack30um_3_5_21 m5_0_0# stack30um_3_5
Xstack30um_3_5_10 m5_0_0# stack30um_3_5
Xstack30um_3_5_23 m5_0_0# stack30um_3_5
Xstack30um_3_5_11 m5_0_0# stack30um_3_5
Xstack30um_3_5_22 m5_0_0# stack30um_3_5
Xstack30um_3_5_12 m5_0_0# stack30um_3_5
Xstack30um_3_5_24 m5_0_0# stack30um_3_5
Xstack30um_3_5_13 m5_0_0# stack30um_3_5
Xstack30um_3_5_14 m5_0_0# stack30um_3_5
Xstack30um_3_5_25 m5_0_0# stack30um_3_5
Xstack30um_3_5_26 m5_0_0# stack30um_3_5
Xstack30um_3_5_15 m5_0_0# stack30um_3_5
Xstack30um_3_5_27 m5_0_0# stack30um_3_5
Xstack30um_3_5_16 m5_0_0# stack30um_3_5
Xstack30um_3_5_17 m5_0_0# stack30um_3_5
Xstack30um_3_5_28 m5_0_0# stack30um_3_5
Xstack30um_3_5_29 m5_0_0# stack30um_3_5
Xstack30um_3_5_18 m5_0_0# stack30um_3_5
Xstack30um_3_5_19 m5_0_0# stack30um_3_5
Xstack30um_3_5_0 m5_0_0# stack30um_3_5
Xstack30um_3_5_2 m5_0_0# stack30um_3_5
Xstack30um_3_5_1 m5_0_0# stack30um_3_5
Xstack30um_3_5_3 m5_0_0# stack30um_3_5
Xstack30um_3_5_4 m5_0_0# stack30um_3_5
Xstack30um_3_5_5 m5_0_0# stack30um_3_5
Xstack30um_3_5_6 m5_0_0# stack30um_3_5
Xstack30um_3_5_7 m5_0_0# stack30um_3_5
Xstack30um_3_5_8 m5_0_0# stack30um_3_5
Xstack30um_3_5_9 m5_0_0# stack30um_3_5
.ends

.subckt nmos_drain a_0_212# dw_0_0# a_0_50# li_1022_1022# a_150_212# a_212_0# w_0_0#
X0 a_150_212# a_0_50# a_212_0# w_0_0# sky130_fd_pr__nfet_g5v0d10v5 ad=3.3792e+12p pd=3.668e+07u as=1.095e+12p ps=9.26e+06u w=4.38e+06u l=500000u
X1 a_150_212# a_0_50# a_0_212# w_0_0# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.095e+12p ps=9.26e+06u w=4.38e+06u l=500000u
.ends

.subckt nmos_source li_0_0# a_0_212# dw_0_0# a_0_50# a_212_0# w_0_0#
X0 w_0_0# a_0_50# a_212_0# w_0_0# sky130_fd_pr__nfet_g5v0d10v5 ad=1.15372e+13p pd=3.22e+07u as=1.095e+12p ps=9.26e+06u w=4.38e+06u l=500000u
X1 w_0_0# a_0_50# a_0_212# w_0_0# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.095e+12p ps=9.26e+06u w=4.38e+06u l=500000u
.ends

.subckt nmos_waffle_36x36 dw_n5900_n5900# a_8912_38400# a_n50_n50# a_112_3350# a_112_1150#
Xnmos_drain_7 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_543 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_458 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_576 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_403 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_521 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_436 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_554 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_469 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_414 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_510 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_425 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_565 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_447 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_532 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_9 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_drain_373 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_288 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_200 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_233 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_351 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_266 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_384 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_299 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_211 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_244 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_340 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_255 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_222 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_395 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_277 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_362 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_181 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_170 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_192 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_81 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_92 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_70 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_8 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_577 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_404 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_522 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_437 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_555 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_500 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_415 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_533 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_448 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_544 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_459 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_426 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_511 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_566 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_201 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_234 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_352 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_267 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_385 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_212 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_330 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_245 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_363 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_278 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_374 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_289 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_256 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_341 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_223 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_396 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_160 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_171 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_82 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_182 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_60 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_93 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_193 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_71 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_9 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_405 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_523 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_438 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_556 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_501 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_416 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_534 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_449 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_567 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_545 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_427 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_512 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_202 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_320 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_235 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_353 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_268 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_386 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_213 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_331 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_246 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_364 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_279 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_397 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_375 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_257 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_342 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_224 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_50 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_83 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_150 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_183 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_61 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_94 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_161 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_194 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_172 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_72 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_406 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_524 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_502 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_417 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_535 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_546 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_428 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_513 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_439 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_557 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_568 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_203 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_321 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_236 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_354 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_269 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_387 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_214 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_332 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_247 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_365 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_398 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_376 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_258 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_343 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_225 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_310 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_151 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_184 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_162 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_195 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_173 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_140 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_84 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_62 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_95 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_40 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_51 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_73 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_407 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_525 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_558 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_503 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_418 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_536 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_569 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_547 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_429 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_514 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_322 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_237 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_355 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_388 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_300 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_215 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_333 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_248 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_366 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_399 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_311 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_226 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_204 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_377 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_259 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_344 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_152 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_185 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_130 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_163 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_196 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_174 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_141 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_30 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_63 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_96 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_41 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_74 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_52 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_85 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_526 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_559 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_504 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_419 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_537 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_515 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_408 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_548 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_301 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_312 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_356 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_389 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_216 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_334 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_249 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_367 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_227 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_345 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_205 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_323 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_238 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_378 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_186 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_131 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_164 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_197 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_142 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_175 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_120 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_153 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_31 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_64 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_97 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_42 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_75 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_86 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_53 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_20 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_505 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_538 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_516 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_549 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_409 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_527 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_302 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_217 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_335 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_368 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_313 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_228 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_346 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_379 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_324 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_239 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_357 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_206 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_132 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_165 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_110 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_143 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_176 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_154 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_187 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_121 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_32 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_65 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_98 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_198 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_10 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_570 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_43 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_76 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_87 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_54 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_21 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_506 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_539 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_517 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_528 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_303 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_218 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_336 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_369 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_314 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_229 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_347 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_358 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_325 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_207 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_33 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_100 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_66 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_133 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_99 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_166 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_199 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_11 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_44 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_111 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_77 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_144 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_177 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_188 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_155 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_88 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_122 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_55 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_22 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_560 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_571 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_390 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_507 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_518 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_529 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_304 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_219 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_337 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_315 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_348 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_359 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_326 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_208 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_101 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_134 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_167 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_112 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_145 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_178 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_189 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_156 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_123 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_67 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_12 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_572 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_45 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_78 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_550 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_23 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_561 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_34 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_89 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_56 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_380 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_391 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_508 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_519 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_305 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_338 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_316 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_349 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_327 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_209 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_135 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_168 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_113 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_146 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_179 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_102 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_157 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_124 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_540 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_13 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_573 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_46 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_79 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_551 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_24 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_57 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_68 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_35 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_562 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_370 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_381 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_392 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_509 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_317 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_306 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_339 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_328 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_169 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_114 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_147 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_125 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_136 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_103 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_158 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_541 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_14 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_574 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_47 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_552 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_25 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_58 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_69 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_36 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_563 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_530 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_371 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_382 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_393 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_360 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_190 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_318 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_329 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_307 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_115 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_148 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_126 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_159 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_137 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_104 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_542 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_15 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_575 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_48 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_520 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_553 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_26 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_59 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_37 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_564 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_531 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_372 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_490 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_350 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_383 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_394 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_361 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_180 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_191 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_319 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_308 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_16 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_49 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_116 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_149 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_521 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_27 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_127 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_510 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_138 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_105 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_38 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_543 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_576 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_554 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_532 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_565 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_373 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_491 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_351 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_384 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_362 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_340 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_395 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_480 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_181 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_192 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_170 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_309 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_117 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_128 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_139 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_106 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_577 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_522 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_555 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_28 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_500 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_533 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_566 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_544 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_17 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_511 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_39 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_492 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_352 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_470 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_385 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_330 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_363 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_481 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_396 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_341 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_374 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_182 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_160 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_193 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_171 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_118 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_129 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_107 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_523 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_556 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_29 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_501 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_534 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_567 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_18 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_545 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_512 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_320 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_353 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_471 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_386 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_331 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_364 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_482 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_397 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_460 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_375 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_493 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_342 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_150 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_183 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_161 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_194 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_290 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_172 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_108 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_119 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_524 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_557 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_502 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_535 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_568 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_19 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_546 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_513 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_321 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_354 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_472 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_387 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_332 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_450 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_365 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_483 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_398 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_494 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_376 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_461 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_343 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_310 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_151 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_162 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_280 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_173 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_140 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_184 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_195 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_291 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_109 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_525 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_558 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_503 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_536 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_569 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_547 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_514 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_322 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_440 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_355 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_473 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_388 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_300 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_333 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_451 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_366 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_484 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_399 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_495 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_377 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_462 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_344 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_311 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_152 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_270 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_185 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_130 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_163 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_281 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_196 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_292 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_174 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_141 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_90 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_526 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_504 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_537 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_515 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_559 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_548 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_441 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_356 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_474 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_389 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_301 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_334 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_452 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_367 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_485 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_312 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_323 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_496 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_378 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_463 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_345 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_430 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_271 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_186 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_131 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_164 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_282 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_197 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_142 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_153 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_120 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_293 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_175 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_260 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_80 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_91 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_505 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_538 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_516 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_527 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_549 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_475 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_302 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_420 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_335 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_453 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_368 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_486 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_313 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_431 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_346 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_442 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_357 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_324 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_497 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_379 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_464 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_132 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_250 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_165 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_283 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_198 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_110 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_143 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_261 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_176 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_272 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_187 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_154 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_121 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_294 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_81 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_92 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_70 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_506 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_539 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_517 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_528 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_303 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_421 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_410 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_336 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_454 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_369 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_487 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_314 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_432 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_347 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_465 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_476 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_358 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_443 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_325 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_498 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_100 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_133 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_251 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_166 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_284 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_199 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_111 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_144 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_262 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_177 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_295 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_188 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_273 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_155 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_240 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_122 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_82 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_60 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_93 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_71 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_507 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_518 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_529 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_304 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_422 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_337 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_455 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_488 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_400 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_315 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_433 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_348 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_466 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_499 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_477 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_359 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_444 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_326 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_411 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_101 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_134 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_252 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_167 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_285 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_112 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_230 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_145 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_263 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_178 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_296 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_274 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_156 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_241 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_123 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_189 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_50 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_83 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_61 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_94 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_72 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_508 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_519 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_305 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_423 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_338 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_456 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_489 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_401 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_316 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_434 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_349 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_467 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_478 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_445 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_327 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_412 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_220 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_135 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_253 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_168 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_286 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_113 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_231 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_146 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_264 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_179 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_297 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_102 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_275 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_157 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_242 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_124 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_84 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_62 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_95 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_40 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_51 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_73 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_509 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_424 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_339 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_457 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_402 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_317 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_435 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_468 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_413 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_328 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_306 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_479 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_446 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_254 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_169 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_287 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_114 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_232 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_147 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_265 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_298 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_210 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_125 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_243 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_103 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_221 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_136 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_276 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_158 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_30 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_63 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_96 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_41 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_74 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_85 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_52 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_drain_458 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_403 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_318 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_436 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_469 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_414 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_329 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_447 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_307 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_425 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_288 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_200 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_115 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_233 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_148 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_266 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_299 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_211 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_126 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_244 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_159 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_277 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_222 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_137 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_255 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_104 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_31 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_64 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_97 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_42 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_75 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_86 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_53 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_20 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_490 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_404 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_319 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_415 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_426 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_308 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_437 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_448 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_459 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_201 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_116 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_234 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_149 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_267 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_212 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_127 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_245 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_278 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_256 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_289 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_138 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_223 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_105 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_32 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_10 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_21 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_491 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_65 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_98 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_43 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_76 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_87 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_54 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_480 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_405 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_438 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_416 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_449 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_427 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_309 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_202 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_117 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_235 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_268 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_213 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_128 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_246 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_279 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_257 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_139 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_224 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_106 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_33 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_492 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_66 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_99 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_470 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_11 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_44 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_77 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_88 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_55 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_481 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_22 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_drain_406 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_439 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_417 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_428 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_203 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_118 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_236 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_269 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_214 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_129 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_247 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_258 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_225 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_107 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_67 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_471 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_12 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_45 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_78 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_23 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_482 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_493 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_34 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_460 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_89 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_56 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_0 a_8912_38400# a_112_1150# dw_n5900_n5900# a_n50_n50# a_112_1150# a_8912_38400#
+ nmos_source
Xnmos_source_290 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_407 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_418 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_429 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_237 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_215 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_248 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_108 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_204 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_119 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_259 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_226 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_472 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_13 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_46 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_79 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_450 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_24 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_483 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_57 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_35 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_68 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_494 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_461 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_1 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_280 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_291 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_419 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_408 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_216 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_249 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_109 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_227 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_238 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_205 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_0 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_14 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_47 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_25 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_58 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_69 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_36 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_440 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_473 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_451 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_484 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_495 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_462 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_2 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_270 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_281 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_292 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_409 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_217 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_228 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_239 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_206 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_1 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_15 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_48 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_26 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_37 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_441 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_474 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_452 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_570 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_485 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_59 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_430 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_496 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_463 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_271 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_282 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_260 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_3 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_293 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_218 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_229 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_207 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_2 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_560 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_475 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_16 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_49 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_420 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_453 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_27 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_drain_571 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_486 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_431 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_464 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_442 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_38 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_497 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_4 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_drain_390 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_250 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_283 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_261 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_294 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_272 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_208 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_219 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_3 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_421 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_454 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_572 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_487 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_28 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_432 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_550 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_465 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_498 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_443 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_561 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_476 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_17 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_410 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_39 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_5 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_251 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_284 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_262 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_380 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_295 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_273 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_391 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_240 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_209 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_4 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_422 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_540 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_455 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_29 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_drain_573 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_488 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_400 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_433 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_551 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_466 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_499 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_477 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_562 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_18 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_444 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_411 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_6 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_252 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_370 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_285 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_230 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_263 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_381 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_296 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_392 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_274 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_241 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_5 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_401 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_19 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_drain_530 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_412 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_423 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_541 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_456 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_574 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_489 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_434 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_552 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_467 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_478 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_563 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_445 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_7 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_220 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_253 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_371 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_286 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_231 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_264 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_382 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_297 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_393 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_275 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_360 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_242 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_190 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_90 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_6 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_424 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_542 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_457 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_575 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_402 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_520 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_435 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_553 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_468 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_479 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_564 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_446 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_531 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_413 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_254 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_372 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_287 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_232 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_350 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_265 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_383 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_298 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_8 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350# a_8912_38400#
+ nmos_source
Xnmos_source_210 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_source_221 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_394 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_276 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_361 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_source_243 a_8912_38400# a_112_3350# dw_n5900_n5900# a_n50_n50# a_112_3350#
+ a_8912_38400# nmos_source
Xnmos_drain_180 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_191 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_80 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
Xnmos_drain_91 a_8912_38400# dw_n5900_n5900# a_n50_n50# a_112_3350# a_112_3350# a_8912_38400#
+ a_8912_38400# nmos_drain
X0 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=8.80377e+15p pd=2.05783e+10u as=3.48383e+15p ps=2.27266e+10u w=4.38e+06u l=500000u
X1 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X5 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X6 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X7 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X8 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X9 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X10 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X11 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X12 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X13 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X14 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X15 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X16 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X17 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X18 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X19 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X20 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X21 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X22 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X23 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X24 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X25 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X26 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X27 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X28 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X29 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X30 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X31 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X32 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X33 a_8912_38400# a_n50_n50# a_112_1150# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=8.1096e+12p ps=5.6365e+07u w=4.38e+06u l=500000u
X34 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X35 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X36 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X37 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X38 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X39 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X40 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X41 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X42 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X43 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X44 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X45 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X46 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X47 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X48 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X49 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X50 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X51 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X52 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X53 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X54 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X55 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X56 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X57 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X58 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X59 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X60 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X61 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X62 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X63 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X64 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X65 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X66 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X67 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X68 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X69 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X70 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X71 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X72 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X73 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X74 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X75 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X76 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X77 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X78 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X79 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X80 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X81 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X82 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X83 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X84 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X85 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X86 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X87 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X88 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X89 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X90 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X91 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X92 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X93 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X94 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X95 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X96 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X97 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X98 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X99 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X100 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X101 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X102 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X103 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X104 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X105 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X106 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X107 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X108 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X109 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X110 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X111 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X112 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X113 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X114 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X115 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X116 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X117 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X118 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X119 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X120 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X121 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X122 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X123 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X124 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X125 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X126 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X127 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X128 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X129 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X130 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X131 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X132 a_8912_38400# a_n50_n50# a_112_1150# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X133 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X134 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X135 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X136 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X137 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X138 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X139 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X140 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X141 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X142 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X143 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X144 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X145 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X146 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X147 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X148 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X149 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X150 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X151 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X152 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X153 a_112_1150# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X154 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X155 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X156 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X157 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X158 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X159 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X160 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X161 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X162 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X163 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X164 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X165 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X166 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X167 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X168 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X169 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X170 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X171 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X172 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X173 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X174 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X175 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X176 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X177 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X178 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X179 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X180 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X181 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X182 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X183 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X184 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X185 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X186 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X187 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X188 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X189 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X190 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X191 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X192 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X193 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X194 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X195 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X196 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X197 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X198 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X199 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X200 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X201 a_112_1150# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X202 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X203 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X204 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X205 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X206 a_112_3350# a_n50_n50# a_8912_38400# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X207 a_8912_38400# a_n50_n50# a_112_3350# a_8912_38400# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
.ends

.subckt pmos_source li_0_0# a_0_212# a_0_50# a_212_0# w_0_0#
X0 w_0_0# a_0_50# a_212_0# w_0_0# sky130_fd_pr__pfet_g5v0d10v5 ad=1.15372e+13p pd=3.22e+07u as=1.095e+12p ps=9.26e+06u w=4.38e+06u l=500000u
X1 w_0_0# a_0_50# a_0_212# w_0_0# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1.095e+12p ps=9.26e+06u w=4.38e+06u l=500000u
.ends

.subckt pmos_drain a_0_212# a_0_50# li_1022_1022# a_150_212# a_212_0# w_0_0#
X0 a_150_212# a_0_50# a_212_0# w_0_0# sky130_fd_pr__pfet_g5v0d10v5 ad=3.3792e+12p pd=3.668e+07u as=1.095e+12p ps=9.26e+06u w=4.38e+06u l=500000u
X1 a_150_212# a_0_50# a_0_212# w_0_0# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1.095e+12p ps=9.26e+06u w=4.38e+06u l=500000u
.ends

.subckt pmos_waffle_48x48 a_8912_51600# a_n50_n50# a_112_3350# a_112_1150#
Xpmos_source_50 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_72 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_94 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_83 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_61 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_71 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_93 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_82 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_60 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_807 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_829 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_818 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_800 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_822 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_833 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_855 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_811 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_866 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_844 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_615 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_877 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_899 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_626 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_648 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_604 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_888 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_659 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_637 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_118 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_129 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_107 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_641 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_685 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_663 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_696 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_674 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_652 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_630 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_401 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_412 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_434 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_478 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_456 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_489 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_467 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_445 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_423 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_990 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_482 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_231 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_253 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_460 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_493 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_471 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_242 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_220 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_275 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_297 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_286 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_264 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_290 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_40 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_95 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_51 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_73 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_84 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_62 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_72 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_50 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_61 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_94 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_83 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_808 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_819 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_823 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_801 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_845 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_867 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_878 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_856 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_834 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_812 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_889 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_616 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_638 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_649 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_627 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_605 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_119 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_108 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_620 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_413 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_642 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_435 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_664 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_686 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_697 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_675 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_653 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_424 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_631 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_402 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_457 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_479 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_468 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_446 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_991 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_980 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_450 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_210 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_232 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_461 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_254 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_276 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_483 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_494 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_265 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_472 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_221 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_243 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_298 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_287 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_280 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_291 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_41 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_30 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_63 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_96 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_74 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_52 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_85 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_40 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_73 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_95 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_51 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_84 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_62 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_809 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_802 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_824 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_617 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_846 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_868 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_879 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_857 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_835 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_606 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_813 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_639 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_628 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_109 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_621 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_632 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_610 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_643 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_436 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_665 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_458 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_687 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_414 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_698 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_469 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_676 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_447 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_654 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_425 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_403 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_992 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_970 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_981 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_440 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_462 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_484 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_473 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_451 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_211 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_233 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_255 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_277 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_299 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_288 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_495 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_266 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_244 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_222 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_200 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_270 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_281 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_292 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_20 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_42 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_64 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_53 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_31 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_86 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_97 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_75 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_41 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_63 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_74 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_96 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_52 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_30 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_85 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_803 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_825 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_814 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_618 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_869 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_847 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_858 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_629 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_836 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_607 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_666 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_600 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_622 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_644 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_655 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_633 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_611 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_459 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_688 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_415 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_437 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_699 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_677 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_448 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_426 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_404 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_960 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_982 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_993 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_971 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_201 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_463 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_485 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_441 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_474 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_496 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_452 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_430 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_256 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_278 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_212 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_234 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_267 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_289 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_245 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_223 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_790 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_271 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_293 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_282 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_260 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_21 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_43 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_87 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_65 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_98 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_76 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_54 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_32 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_10 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_20 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_64 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_42 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_86 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_97 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_75 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_53 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_31 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_804 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_826 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_848 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_837 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_815 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_619 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_859 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_608 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_689 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_601 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_623 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_645 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_667 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_678 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_656 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_612 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_634 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_416 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_438 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_449 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_405 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_427 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_961 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_983 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_994 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_972 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_950 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_202 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_431 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_224 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_453 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_486 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_464 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_442 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_213 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_420 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_497 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_475 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_257 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_279 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_235 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_268 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_246 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_780 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_791 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_250 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_272 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_294 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_283 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_261 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_22 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_44 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_66 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_88 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_99 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_77 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_55 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_33 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_11 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_21 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_43 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_54 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_32 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_10 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_65 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_87 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_98 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_76 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_827 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_849 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_805 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_838 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_816 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_609 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_1050 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_624 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_417 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_646 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_668 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_602 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_679 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_657 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_635 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_406 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_613 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_439 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_428 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_940 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_962 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_973 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_951 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_984 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_995 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_410 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_432 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_421 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_203 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_225 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_454 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_247 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_258 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_465 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_487 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_236 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_443 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_214 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_498 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_476 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_269 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_781 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_792 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_770 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_251 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_273 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_284 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_262 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_240 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_295 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_23 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_12 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_45 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_67 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_89 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_78 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_56 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_34 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_22 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_44 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_66 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_88 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_77 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_55 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_33 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_11 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_99 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_806 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_828 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_839 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_817 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_1051 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_1040 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_603 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_614 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_647 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_669 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_418 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_625 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_658 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_429 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_636 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_407 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_941 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_963 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_985 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_996 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_974 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_952 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_930 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_411 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_455 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_433 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_466 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_444 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_422 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_400 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_204 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_248 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_226 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_477 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_499 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_488 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_259 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_237 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_215 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_760 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_782 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_793 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_771 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_252 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_274 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_296 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_230 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_285 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_263 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_241 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_24 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_46 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_35 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_13 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_68 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_79 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_57 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_590 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_45 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_67 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_89 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_23 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_78 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_56 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_34 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_12 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_807 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_829 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_818 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_1030 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_1052 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_1041 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_615 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_637 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_648 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_626 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_604 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_408 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_419 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_659 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_942 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_964 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_986 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_920 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_997 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_975 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_953 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_931 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_412 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_434 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_456 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_478 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_489 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_467 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_445 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_423 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_401 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_205 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_227 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_249 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_238 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_216 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_990 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_761 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_783 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_794 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_772 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_750 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_275 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_297 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_231 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_253 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_286 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_264 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_242 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_220 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_25 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_69 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_47 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_58 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_14 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_36 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_580 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_591 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_68 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_46 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_24 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_79 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_57 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_35 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_13 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_808 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_819 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_1053 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_1031 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_1042 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_1020 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_616 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_638 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_649 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_627 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_605 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_409 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_921 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_910 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_965 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_987 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_943 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_998 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_976 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_954 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_932 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_413 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_206 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_435 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_457 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_479 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_468 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_446 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_424 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_402 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_228 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_239 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_217 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_762 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_991 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_740 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_980 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_751 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_784 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_773 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_795 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_210 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_232 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_221 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_298 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_254 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_276 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_287 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_265 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_243 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_26 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_48 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_59 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_37 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_15 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_570 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_592 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_581 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_25 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_36 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_14 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_47 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_69 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_58 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_809 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_1010 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_1032 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_1054 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_1043 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_1021 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_639 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_617 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_628 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_606 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_900 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_922 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_944 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_955 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_911 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_933 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_988 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_966 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_999 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_977 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_414 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_403 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_436 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_229 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_458 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_207 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_469 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_447 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_218 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_425 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_970 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_730 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_752 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_992 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_785 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_763 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_741 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_796 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_774 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_981 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_233 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_255 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_211 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_244 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_266 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_222 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_200 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_277 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_299 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_288 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_49 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_27 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_38 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_16 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_571 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_593 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_582 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_560 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_26 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_48 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_37 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_59 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_15 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_390 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_1011 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_1033 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_1022 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_1000 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_1055 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_1044 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_618 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_629 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_607 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_923 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_945 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_967 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_901 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_978 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_956 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_934 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_912 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_989 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_415 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_437 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_448 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_426 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_404 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_459 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_208 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_219 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_960 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_971 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_993 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_982 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_731 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_753 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_764 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_786 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_742 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_720 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_797 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_775 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_201 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_234 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_256 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_278 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_212 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_289 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_267 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_245 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_223 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_17 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_28 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_790 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_39 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_550 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_572 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_594 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_583 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_561 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_27 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_49 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_38 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_16 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_380 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_391 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_1034 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_1056 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_1012 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_1045 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_1023 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_1001 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_619 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_608 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_946 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_968 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_902 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_924 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_957 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_979 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_935 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_913 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_416 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_438 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_449 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_427 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_405 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_209 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_710 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_961 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_983 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_994 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_972 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_950 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_754 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_732 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_776 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_798 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_787 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_765 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_743 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_721 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_202 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_224 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_279 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_235 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_257 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_213 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_268 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_246 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_18 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_29 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_551 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_780 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_791 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_562 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_540 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_573 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_595 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_584 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_17 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_28 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_39 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_370 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_392 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_381 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_1057 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_1013 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_1035 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_1046 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_1024 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_1002 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_609 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_903 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_914 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_936 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_969 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_947 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_925 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_958 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_417 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_439 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_428 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_406 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_711 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_940 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_733 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_962 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_984 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_995 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_973 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_744 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_951 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_722 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_700 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_755 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_777 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_799 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_788 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_766 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_203 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_214 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_225 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_247 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_258 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_236 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_269 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_19 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_770 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_781 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_574 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_596 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_530 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_552 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_585 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_792 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_563 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_541 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_18 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_29 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_371 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_393 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_382 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_360 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_1014 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_1036 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_190 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_1047 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_1025 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_1003 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_915 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_937 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_926 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_904 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_948 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_959 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_418 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_429 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_407 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_941 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_952 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_930 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_712 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_734 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_963 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_756 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_985 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_778 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_996 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_767 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_974 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_745 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_723 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_701 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_789 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_204 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_226 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_248 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_237 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_215 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_259 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_760 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_782 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_793 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_771 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_597 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_531 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_553 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_575 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_586 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_564 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_542 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_520 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_19 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_590 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_394 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_350 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_372 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_383 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_361 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_1015 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_1004 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_180 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_1037 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_191 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_1026 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_1048 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_938 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_916 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_949 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_927 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_905 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_408 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_419 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_942 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_964 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_986 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_920 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_975 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_953 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_931 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_735 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_757 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_779 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_713 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_997 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_768 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_746 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_724 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_702 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_205 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_227 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_249 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_238 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_216 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_761 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_783 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_510 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_794 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_750 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_772 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_532 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_554 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_576 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_598 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_587 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_543 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_565 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_521 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_340 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_362 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_591 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_580 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_351 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_395 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_373 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_384 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_181 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_1005 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_1038 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_1016 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_192 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_170 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_1049 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_1027 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_917 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_939 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_928 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_906 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_409 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_965 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_987 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_921 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_943 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_998 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_976 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_954 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_932 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_910 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_758 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_714 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_736 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_769 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_747 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_725 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_703 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_206 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_228 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_239 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_217 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_500 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_522 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_762 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_784 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_533 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_740 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_511 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_795 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_773 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_544 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_751 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_555 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_577 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_599 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_588 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_566 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_341 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_570 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_363 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_592 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_385 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_374 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_581 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_352 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_330 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_396 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_160 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_182 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_1006 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_1017 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_1039 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_193 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_171 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_1028 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_918 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_929 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_907 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_900 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_988 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_922 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_715 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_944 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_966 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_999 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_977 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_955 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_726 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_933 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_704 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_911 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_737 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_759 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_748 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_229 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_207 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_218 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_730 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_741 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_752 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_501 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_523 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_785 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_578 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_534 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_556 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_763 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_512 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_796 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_567 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_774 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_545 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_589 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_593 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_571 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_582 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_560 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_320 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_342 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_386 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_364 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_397 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_375 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_353 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_331 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_390 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_183 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_1007 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_1029 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_161 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_1018 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_194 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_172 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_150 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_919 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_908 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_923 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_901 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_934 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_912 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_716 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_945 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_738 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_967 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_989 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_978 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_727 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_749 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_956 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_705 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_208 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_219 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_731 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_753 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_775 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_764 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_742 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_720 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_524 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_502 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_546 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_568 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_579 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_786 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_557 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_535 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_513 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_797 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_550 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_572 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_594 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_583 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_561 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_310 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_321 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_343 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_365 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_387 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_398 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_376 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_354 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_332 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_140 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_391 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_380 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_151 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_1008 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_162 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_184 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_1019 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_195 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_173 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_909 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_913 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_946 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_968 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_924 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_902 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_957 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_935 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_706 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_739 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_717 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_979 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_728 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_209 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_1050 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_710 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_732 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_754 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_776 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_787 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_765 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_743 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_721 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_798 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_503 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_525 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_547 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_569 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_558 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_536 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_514 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_551 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_344 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_573 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_595 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_300 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_322 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_584 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_562 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_333 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_540 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_311 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_366 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_388 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_399 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_377 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_355 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_1009 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_141 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_370 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_163 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_392 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_185 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_174 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_381 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_152 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_130 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_196 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_914 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_969 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_925 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_947 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_903 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_958 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_936 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_707 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_718 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_729 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_1040 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_1051 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_700 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_711 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_504 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_733 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_526 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_777 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_755 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_799 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_788 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_766 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_744 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_515 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_722 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_548 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_559 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_537 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_530 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_541 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_574 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_367 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_596 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_301 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_323 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_345 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_552 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_585 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_356 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_563 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_334 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_312 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_389 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_378 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_890 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_371 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_393 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_382 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_360 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_164 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_186 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_120 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_142 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_175 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_197 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_153 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_131 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_190 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_915 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_708 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_937 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_959 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_948 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_926 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_904 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_719 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_1030 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_1052 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_1041 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_712 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_723 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_701 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_505 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_734 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_527 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_756 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_549 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_778 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_789 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_767 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_538 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_745 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_516 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_531 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_553 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_575 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_564 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_520 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_542 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_597 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_302 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_324 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_346 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_368 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_379 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_586 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_357 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_313 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_335 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_891 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_880 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_110 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_394 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_372 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_350 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_383 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_361 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_132 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_165 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_187 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_143 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_121 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_198 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_176 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_154 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_180 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_191 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_916 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_905 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_709 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_938 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_949 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_927 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_1031 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_1053 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_1042 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_1020 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_735 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_757 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_713 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_746 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_724 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_702 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_528 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_779 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_506 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_768 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_539 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_517 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_532 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_554 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_576 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_598 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_510 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_587 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_565 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_543 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_521 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_303 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_325 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_347 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_369 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_358 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_336 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_314 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_892 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_870 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_881 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_111 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_340 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_133 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_362 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_373 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_395 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_351 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_122 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_100 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_384 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_155 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_166 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_188 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_144 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_199 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_177 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_181 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_192 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_170 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_0 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_917 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_939 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_928 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_906 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_1010 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_1032 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_1021 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_1054 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_1043 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_758 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_714 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_736 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_769 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_747 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_725 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_703 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_507 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_529 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_518 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_500 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_555 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_577 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_599 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_304 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_326 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_511 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_533 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_566 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_588 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_544 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_315 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_522 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_348 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_359 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_337 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_871 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_860 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_893 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_882 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_341 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_330 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_112 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_363 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_156 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_134 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_385 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_396 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_167 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_374 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_145 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_352 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_123 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_101 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_178 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_189 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_690 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_160 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_182 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_171 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_193 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_1 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_918 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_929 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_907 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_1011 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_1033 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_1055 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_1044 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_1022 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_1000 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_715 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_508 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_737 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_759 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_748 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_704 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_726 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_519 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_501 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_523 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_512 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_316 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_545 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_349 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_578 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_556 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_327 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_534 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_305 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_589 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_567 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_338 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_850 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_872 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_894 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_883 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_861 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_320 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_342 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_364 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_375 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_353 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_331 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_113 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_135 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_157 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_386 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_179 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_397 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_168 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_146 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_124 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_102 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_691 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_680 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_183 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_161 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_194 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_172 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_150 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_2 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_919 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_908 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_1034 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_1056 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_1012 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_1045 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_1023 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_1001 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_705 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_716 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_509 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_738 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_749 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_727 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_502 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_524 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_546 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_557 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_535 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_513 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_317 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_339 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_579 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_328 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_306 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_568 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_873 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_895 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_851 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_884 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_862 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_840 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_321 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_343 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_365 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_387 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_398 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_376 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_354 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_332 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_310 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_114 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_136 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_158 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_169 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_147 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_125 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_103 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_670 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_692 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_681 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_140 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_162 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_184 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_195 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_173 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_151 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_3 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_909 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_0 a_8912_51600# a_112_1150# a_n50_n50# a_112_1150# a_8912_51600# pmos_source
Xpmos_drain_1057 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_1013 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_1035 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_1046 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_1024 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_1002 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_739 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_717 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_728 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_706 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_503 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_547 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_525 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_569 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_558 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_536 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_514 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_318 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_329 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_307 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_830 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_896 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_852 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_874 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_885 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_863 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_841 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_344 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_366 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_388 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_300 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_115 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_322 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_399 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_377 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_355 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_333 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_104 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_311 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_137 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_159 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_148 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_126 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_660 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_671 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_693 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_682 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_141 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_130 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_163 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_185 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_196 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_152 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_174 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_4 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_490 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_1 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_1014 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_1003 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_1036 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_1047 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_1025 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_707 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_729 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_718 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_504 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_526 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_548 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_559 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_537 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_308 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_515 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_319 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_831 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_853 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_842 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_820 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_875 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_897 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_886 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_864 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_301 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_323 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_312 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_367 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_389 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_116 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_138 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_345 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_378 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_149 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_356 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_127 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_334 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_105 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_661 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_672 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_694 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_650 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_683 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_890 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_142 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_164 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_120 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_153 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_131 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_186 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_197 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_175 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_480 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_5 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_491 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_2 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_1015 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_1037 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_1048 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_1026 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_1004 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_708 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_719 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_505 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_527 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_549 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_538 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_309 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_516 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_854 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_876 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_810 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_832 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_865 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_887 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_843 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_821 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_898 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_302 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_324 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_346 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_357 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_335 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_313 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_117 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_139 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_368 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_379 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_128 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_106 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_891 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_880 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_662 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_640 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_684 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_695 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_673 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_651 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_110 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_132 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_187 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_143 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_165 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_121 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_198 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_176 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_154 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_481 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_6 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_492 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_470 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_3 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_1038 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_1016 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_1049 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_1027 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_1005 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_709 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_528 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_506 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_539 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_517 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_800 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_822 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_844 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_877 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_899 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_855 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_833 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_811 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_888 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_866 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_325 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_347 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_369 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_303 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_336 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_358 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_314 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_118 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_129 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_107 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_870 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_892 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_881 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_641 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_663 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_685 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_696 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_674 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_652 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_630 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_133 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_111 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_155 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_188 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_166 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_144 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_122 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_100 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_199 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_177 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_460 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_7 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_471 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_482 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_493 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_290 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_4 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_1006 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_1028 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_1039 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_1017 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_507 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_529 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_518 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_801 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_812 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_823 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_845 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_856 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_878 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_834 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_889 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_867 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_326 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_348 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_304 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_359 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_337 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_315 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_119 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_108 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_620 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_642 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_871 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_893 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_882 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_653 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_860 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_631 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_664 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_686 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_697 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_675 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_112 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_123 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_101 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_134 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_156 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_178 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_189 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_167 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_145 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_461 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_483 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_690 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_8 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_494 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_472 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_450 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_280 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_291 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_5 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_1007 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_1029 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_1018 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_508 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_519 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_802 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_824 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_835 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_813 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_846 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_868 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_879 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_857 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_305 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_316 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_109 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_327 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_349 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_338 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_850 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_861 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_643 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_872 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_665 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_894 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_687 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_621 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_676 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_883 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_654 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_632 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_610 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_698 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_113 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_135 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_146 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_124 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_102 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_179 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_157 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_168 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_691 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_680 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_440 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_462 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_484 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_9 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_495 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_451 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_473 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_270 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_281 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_292 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_6 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_1008 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_1019 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_90 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_509 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_803 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_825 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_847 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_869 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_858 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_836 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_814 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_317 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_339 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_328 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_306 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_873 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_851 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_884 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_862 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_840 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_666 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_895 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_688 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_600 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_622 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_644 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_699 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_677 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_655 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_633 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_611 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_114 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_136 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_158 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_169 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_147 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_125 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_103 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_670 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_692 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_681 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_430 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_463 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_485 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_441 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_496 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_474 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_452 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_271 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_260 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_293 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_282 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_7 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_1009 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_91 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_80 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_90 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_804 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_826 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_848 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_859 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_837 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_815 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_318 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_329 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_307 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_896 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_601 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_830 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_852 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_874 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_885 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_863 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_841 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_689 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_623 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_645 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_667 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_678 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_656 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_634 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_612 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_137 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_159 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_115 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_148 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_126 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_104 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_431 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_693 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_442 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_671 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_420 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_682 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_453 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_660 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_486 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_464 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_497 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_475 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_250 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_294 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_272 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_283 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_490 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_261 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_8 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_70 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_92 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_81 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_91 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_80 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_827 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_849 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_805 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_838 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_816 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_319 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_308 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_831 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_624 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_853 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_875 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_897 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_602 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_886 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_635 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_842 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_864 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_613 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_820 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_646 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_668 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_679 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_657 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_105 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_116 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_138 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_149 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_127 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_650 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_432 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_410 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_661 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_454 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_683 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_476 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_487 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_694 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_465 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_672 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_443 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_421 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_498 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_480 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_491 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_251 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_273 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_295 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_284 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_262 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_240 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_9 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_71 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_60 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_82 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_93 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_92 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_70 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_81 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_806 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_817 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_828 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_839 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_309 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_821 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_832 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_810 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_843 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_614 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_854 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_647 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_876 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_669 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_898 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_625 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_603 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_887 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_658 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_865 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_636 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_117 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_106 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_128 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_139 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_640 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_662 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_684 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_673 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_651 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_411 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_433 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_455 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_477 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_488 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_695 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_466 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_444 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_422 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_400 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_499 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_source_481 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_492 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_source_470 a_8912_51600# a_112_3350# a_n50_n50# a_112_3350# a_8912_51600# pmos_source
Xpmos_drain_252 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_274 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_296 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_230 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_285 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_263 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
Xpmos_drain_241 a_8912_51600# a_n50_n50# a_112_3350# a_112_3350# a_8912_51600# a_8912_51600#
+ pmos_drain
X0 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=6.25436e+15p pd=4.0771e+10u as=1.56894e+16p ps=3.65702e+10u w=4.38e+06u l=500000u
X1 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X5 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X6 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X7 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X8 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X9 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X10 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X11 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X12 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X13 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X14 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X15 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X16 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X17 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X18 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X19 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X20 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X21 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X22 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X23 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X24 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X25 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X26 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X27 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X28 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X29 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X30 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X31 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X32 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X33 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X34 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X35 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X36 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X37 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X38 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X39 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X40 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X41 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X42 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X43 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X44 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X45 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X46 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X47 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X48 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X49 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X50 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X51 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X52 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X53 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X54 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X55 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X56 a_8912_51600# a_n50_n50# a_112_1150# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.1096e+12p ps=5.6365e+07u w=4.38e+06u l=500000u
X57 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X58 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X59 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X60 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X61 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X62 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X63 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X64 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X65 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X66 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X67 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X68 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X69 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X70 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X71 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X72 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X73 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X74 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X75 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X76 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X77 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X78 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X79 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X80 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X81 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X82 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X83 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X84 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X85 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X86 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X87 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X88 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X89 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X90 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X91 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X92 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X93 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X94 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X95 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X96 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X97 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X98 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X99 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X100 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X101 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X102 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X103 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X104 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X105 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X106 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X107 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X108 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X109 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X110 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X111 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X112 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X113 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X114 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X115 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X116 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X117 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X118 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X119 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X120 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X121 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X122 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X123 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X124 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X125 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X126 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X127 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X128 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X129 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X130 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X131 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X132 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X133 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X134 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X135 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X136 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X137 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X138 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X139 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X140 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X141 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X142 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X143 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X144 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X145 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X146 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X147 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X148 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X149 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X150 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X151 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X152 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X153 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X154 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X155 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X156 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X157 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X158 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X159 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X160 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X161 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X162 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X163 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X164 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X165 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X166 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X167 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X168 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X169 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X170 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X171 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X172 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X173 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X174 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X175 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X176 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X177 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X178 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X179 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X180 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X181 a_8912_51600# a_n50_n50# a_112_1150# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X182 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X183 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X184 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X185 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X186 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X187 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X188 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X189 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X190 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X191 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X192 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X193 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X194 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X195 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X196 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X197 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X198 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X199 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X200 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X201 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X202 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X203 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X204 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X205 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X206 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X207 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X208 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X209 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X210 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X211 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X212 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X213 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X214 a_112_1150# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X215 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X216 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X217 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X218 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X219 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X220 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X221 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X222 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X223 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X224 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X225 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X226 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X227 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X228 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X229 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X230 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X231 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X232 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X233 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X234 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X235 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X236 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X237 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X238 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X239 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X240 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X241 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X242 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X243 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X244 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X245 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X246 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X247 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X248 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X249 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X250 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X251 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X252 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X253 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X254 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X255 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X256 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X257 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X258 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X259 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X260 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X261 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X262 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X263 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X264 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X265 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X266 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X267 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X268 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X269 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X270 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X271 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X272 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X273 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X274 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X275 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X276 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X277 a_112_3350# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X278 a_112_1150# a_n50_n50# a_8912_51600# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X279 a_8912_51600# a_n50_n50# a_112_3350# a_8912_51600# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
.ends

.subckt power_stage nmos_waffle_36x36_1/dw_n5900_n5900# VP nmos_waffle_36x36_0/dw_n5900_n5900#
+ s4 s3 s2 s1 fc2 VN out fc1 VSUBS
Xnmos_waffle_36x36_0 nmos_waffle_36x36_0/dw_n5900_n5900# VN s4 fc2 fc2 nmos_waffle_36x36
Xnmos_waffle_36x36_1 nmos_waffle_36x36_1/dw_n5900_n5900# fc2 s3 out out nmos_waffle_36x36
Xpmos_waffle_48x48_0 fc1 s2 out out pmos_waffle_48x48
Xpmos_waffle_48x48_1 VP s1 fc1 fc1 pmos_waffle_48x48
.ends

.subckt fc_pad m5_0_0#
Xstack30um_1_5_19 m5_0_0# stack30um_1_5
Xstack30um_1_5_18 m5_0_0# stack30um_1_5
Xstack30um_1_5_0 m5_0_0# stack30um_1_5
Xstack30um_1_5_1 m5_0_0# stack30um_1_5
Xstack30um_1_5_2 m5_0_0# stack30um_1_5
Xstack30um_1_5_3 m5_0_0# stack30um_1_5
Xstack30um_1_5_4 m5_0_0# stack30um_1_5
Xstack30um_1_5_5 m5_0_0# stack30um_1_5
Xstack30um_1_5_6 m5_0_0# stack30um_1_5
Xstack30um_1_5_8 m5_0_0# stack30um_1_5
Xstack30um_1_5_7 m5_0_0# stack30um_1_5
Xstack30um_1_5_9 m5_0_0# stack30um_1_5
Xstack30um_1_5_20 m5_0_0# stack30um_1_5
Xstack30um_1_5_10 m5_0_0# stack30um_1_5
Xstack30um_1_5_11 m5_0_0# stack30um_1_5
Xstack30um_1_5_12 m5_0_0# stack30um_1_5
Xstack30um_1_5_13 m5_0_0# stack30um_1_5
Xstack30um_1_5_14 m5_0_0# stack30um_1_5
Xstack30um_1_5_15 m5_0_0# stack30um_1_5
Xstack30um_1_5_16 m5_0_0# stack30um_1_5
Xstack30um_1_5_17 m5_0_0# stack30um_1_5
.ends

.subckt flying_cap m4_8380_242120# m5_8380_287100#
Xunit_cap_360 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_371 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_382 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_393 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1038 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1027 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1049 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1005 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1016 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1550 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1561 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1572 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1583 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1594 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_190 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2070 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2081 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2092 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1380 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1391 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_926 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_937 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_948 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_904 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_959 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_915 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_701 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_778 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_723 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_95 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_767 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_712 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_62 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_734 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_789 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_745 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_73 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_756 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_40 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1968 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1913 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1979 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1924 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1935 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1946 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1902 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1957 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_531 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_520 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_542 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_553 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_564 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_575 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_586 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_597 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1209 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1710 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1765 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1754 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1721 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1776 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1732 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1787 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1743 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1798 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_361 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_372 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_383 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_394 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_350 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1006 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1039 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1028 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1017 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2230 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1551 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1562 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1540 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1595 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1573 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1584 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_180 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_191 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2071 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1392 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2082 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2093 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1370 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1381 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2060 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_927 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_938 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_949 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_905 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_916 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_724 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_713 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_52 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_735 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_702 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_30 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_41 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_779 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_96 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_768 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_63 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_746 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_74 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_757 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1903 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1969 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1914 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1925 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1936 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1947 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1958 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_565 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_510 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_521 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_576 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_532 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_587 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_543 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_554 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_598 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1711 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1700 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1722 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1733 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1744 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1766 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1755 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1777 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1788 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1799 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_362 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_373 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_384 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_340 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_395 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_351 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1029 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1007 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1018 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2231 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1552 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2220 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1596 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1563 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1574 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1530 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1585 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1541 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_170 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_181 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_192 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2072 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1393 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2083 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1360 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1371 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2094 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2050 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1382 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2061 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_906 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_917 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_928 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_939 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1190 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_725 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_42 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_769 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_714 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_64 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_53 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_736 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_20 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_747 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_75 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_703 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_758 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1915 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1926 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1937 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1904 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1959 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1948 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_566 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_511 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_555 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_522 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_577 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_533 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_588 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_544 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_599 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_500 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1767 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1712 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1756 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1701 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1723 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1778 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1734 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1745 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1789 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_363 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_374 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_330 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_385 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_341 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_396 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_352 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1008 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1019 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2221 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2210 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2232 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1553 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1597 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1564 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1520 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1575 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1531 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1586 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1542 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_160 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_171 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_182 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_193 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2073 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2040 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2051 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2062 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1350 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1394 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2084 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1361 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1372 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2095 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1383 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_929 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_907 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_918 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1191 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1180 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_726 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_43 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_715 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_65 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_10 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_54 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_737 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_748 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_21 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_76 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_704 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_759 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1916 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1927 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1938 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1949 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1905 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_501 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_567 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_512 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_556 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_523 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_578 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_534 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_589 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_545 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1713 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1757 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1702 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1768 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1724 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1779 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1735 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1746 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_320 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_331 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_342 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_375 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_364 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_386 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_397 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_353 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1009 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2233 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2222 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1510 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2200 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2211 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1554 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1598 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1543 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1565 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1521 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1576 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1532 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1587 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_161 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_172 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_183 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_194 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1351 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2074 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2063 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1340 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2085 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2030 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1362 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2041 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2096 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2052 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1395 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1373 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1384 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_919 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_908 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1192 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1181 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1170 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_11 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_727 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_44 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_716 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_55 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_738 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_66 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_22 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_77 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_749 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_705 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1917 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1928 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1939 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1906 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_513 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_524 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_535 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_502 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_568 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_557 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_579 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_546 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1714 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1758 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1703 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1769 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1725 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1736 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1747 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_310 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_354 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_376 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_321 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_365 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_332 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_343 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_387 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_398 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2234 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1500 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2223 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1544 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1511 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1522 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2201 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1533 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2212 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1555 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1599 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1566 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1577 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1588 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_162 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_173 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_184 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_195 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2075 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2020 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2064 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1341 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2086 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2031 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1352 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1363 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2042 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2097 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1374 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2053 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1330 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1385 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1396 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_909 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1193 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1182 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1160 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1171 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_717 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_12 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_23 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_706 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_56 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_728 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_739 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_67 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_78 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1918 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1907 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1929 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_569 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_514 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_558 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_503 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_525 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_536 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_547 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1715 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1704 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1726 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1759 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1737 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1748 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_311 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_355 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_377 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_322 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_366 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_333 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_388 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_344 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_300 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_399 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2235 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1556 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1501 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2224 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1545 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1512 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1567 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1523 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1578 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2202 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1534 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2213 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1589 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_163 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_174 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_130 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_185 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_196 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2021 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2010 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2076 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1397 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1342 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2065 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2032 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1353 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1364 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2087 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1320 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2043 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2098 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1375 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2054 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1331 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1386 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1194 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1183 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1150 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1161 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1172 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_718 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_13 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_57 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_729 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_68 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_24 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_707 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_79 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1919 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1908 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_515 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_559 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_504 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_526 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_537 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_548 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1705 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1716 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1727 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1738 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1749 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_301 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_356 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_323 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_312 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_367 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_378 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_334 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_389 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_345 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_890 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2203 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1557 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1502 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2225 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1546 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1513 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1568 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1524 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1579 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1535 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2214 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_120 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_131 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_142 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_164 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_175 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_186 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_197 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2022 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2011 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2033 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1310 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2044 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2000 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2055 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2077 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1398 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1343 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2066 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1387 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1354 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1365 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2088 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2099 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1321 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1376 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1332 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1140 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1151 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1195 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1184 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1162 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1173 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xfc_pad_0 m5_8380_287100# fc_pad
Xunit_cap_719 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_58 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_14 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_69 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_25 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_708 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1909 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_516 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_505 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_527 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_538 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_549 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1706 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1717 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1728 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1739 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_302 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_324 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_313 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_357 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_368 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_379 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_335 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_346 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_880 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_891 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2226 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2204 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2215 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1558 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1503 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1547 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1514 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1569 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1525 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1536 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_165 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_110 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_121 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_176 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_132 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_143 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_198 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_187 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2078 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2023 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1344 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2067 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2012 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2034 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1300 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1311 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2089 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2045 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1322 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2001 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1333 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2056 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1399 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1388 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1355 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1366 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1377 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1141 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1185 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1130 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1152 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1163 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1174 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1196 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xfc_pad_1 m4_8380_242120# fc_pad
Xunit_cap_59 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_15 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_26 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_709 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_517 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_506 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_528 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_539 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1707 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1718 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1729 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_358 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_303 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_325 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_314 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_336 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_347 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_369 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_881 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_870 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_892 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2227 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1504 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1515 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1526 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2205 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2216 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1559 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1548 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1537 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_199 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_166 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_111 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_122 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_177 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_133 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_188 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_144 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2079 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2024 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1345 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2068 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2013 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1356 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1301 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1312 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2035 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1367 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2046 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1323 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2002 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1334 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2057 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1389 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1378 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1890 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1142 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1186 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1131 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1197 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1153 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1164 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1120 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1175 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_16 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_27 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_38 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_518 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_507 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_529 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1708 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1719 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_359 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_304 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_315 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_326 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_337 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_348 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_882 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_871 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_893 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_860 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1505 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2228 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1549 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1516 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1527 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2206 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1538 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2217 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_167 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_112 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_156 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_123 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_178 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_134 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_189 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_145 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_690 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2003 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2025 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1346 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2069 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2014 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1335 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1357 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1302 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1313 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2036 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1368 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2047 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1324 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1379 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2058 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1880 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1891 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1110 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1143 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1187 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1132 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1198 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1154 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1165 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1121 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1176 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_17 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_28 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_39 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_519 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_508 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1709 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_305 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_316 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_327 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_338 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_349 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_883 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_872 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_894 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_850 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_861 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1506 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2229 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1517 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1528 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2207 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1539 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2218 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_113 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_124 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_146 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_168 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_157 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_179 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_680 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_691 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2026 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2015 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2037 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2004 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1347 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1336 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1358 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1303 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1314 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1369 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2048 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1325 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2059 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1870 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1881 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1892 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1133 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1100 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1111 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1122 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1188 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1199 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1144 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1155 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1166 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1177 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_18 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_29 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_509 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_306 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_317 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_328 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_339 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_840 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_851 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_862 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_873 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_884 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_895 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2219 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2208 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1507 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1518 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1529 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_147 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_114 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_158 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_125 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_169 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_670 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_681 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_692 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2027 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2016 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1304 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2038 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1315 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1326 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2049 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2005 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1348 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1337 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1359 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1871 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1860 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1882 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1893 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1134 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1145 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1101 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1156 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1112 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1167 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1123 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1189 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1178 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1690 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_19 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_307 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_318 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_329 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_830 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_874 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_885 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_841 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_896 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_852 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_863 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1508 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2209 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1519 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_148 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_115 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_104 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_159 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_126 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_671 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_660 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_682 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_693 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1349 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2017 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1338 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2028 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1305 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2039 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1316 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1327 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2006 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1861 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1872 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1883 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1894 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1850 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_490 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1135 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1179 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1146 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1102 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1157 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1113 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1168 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1124 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1680 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1691 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_308 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_319 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_831 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_875 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_820 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_886 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_842 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_897 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_853 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_864 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1509 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_116 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_105 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_127 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_672 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_661 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_683 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_694 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_650 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2018 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1339 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2029 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1306 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1317 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1328 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2007 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1862 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1873 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1884 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1840 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1895 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1851 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_480 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_491 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1136 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1147 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1103 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1158 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1114 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1169 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1125 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1670 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1681 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1692 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2190 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_309 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_810 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_876 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_821 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_887 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_832 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_843 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_898 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_854 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_865 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_106 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_117 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_128 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_662 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_640 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_651 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_673 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_684 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_695 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2019 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2008 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1307 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1318 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1329 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1830 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1863 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1874 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1885 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1841 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1896 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1852 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_481 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_470 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_492 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1104 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1115 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1137 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1148 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1159 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1126 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1660 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1671 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1682 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1693 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2180 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2191 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1490 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_822 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_833 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_844 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_800 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_811 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_877 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_888 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_899 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_855 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_866 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_107 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_118 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_129 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_0 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_674 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_663 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_630 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_685 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_641 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_696 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_652 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1308 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2009 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1319 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1820 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1831 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1842 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1853 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1864 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1875 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1886 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1897 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_460 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_471 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_482 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_493 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1138 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1127 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1149 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1105 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1116 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1661 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1650 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1672 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1683 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1694 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_290 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2181 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2170 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1491 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2192 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1480 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_878 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_823 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_867 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_834 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_845 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_801 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_856 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_812 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_889 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_108 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_119 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_675 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_620 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_664 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_631 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_686 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_642 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_697 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_653 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1309 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1865 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1810 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1876 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1821 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1832 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1887 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1843 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1854 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1898 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_461 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_472 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_483 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_494 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_450 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1139 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1128 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1106 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1117 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1662 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1651 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1673 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1684 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1640 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1695 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_280 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_291 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2182 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2171 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2160 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1492 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2193 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1470 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1481 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_879 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_824 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_868 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_835 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_846 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_802 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_857 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_813 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_109 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_610 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_621 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_665 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_632 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_676 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_687 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_643 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_698 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_654 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1866 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1811 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1855 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1877 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1822 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1833 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1888 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1844 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1899 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1800 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_462 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_440 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_451 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_473 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_484 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_495 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1129 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1107 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1118 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1663 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1652 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1674 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1630 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1685 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1641 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1696 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_270 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_281 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_292 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2183 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2172 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1460 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2194 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1471 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2150 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2161 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1493 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1482 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1290 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_825 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_869 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_836 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_847 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_803 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_858 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_814 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_3 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_622 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_611 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_633 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_644 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_600 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_666 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_677 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_688 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_699 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_655 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1812 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1801 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1867 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1856 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1878 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1823 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1834 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1889 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1845 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_463 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_452 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_474 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_430 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_485 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_441 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_496 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1108 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1119 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1653 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1620 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1631 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1642 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1664 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1675 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1686 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1697 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_271 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_260 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_282 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_293 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1450 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2173 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1494 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2184 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1461 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2140 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2195 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1472 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2151 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1483 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2162 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1291 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1280 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_826 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_815 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_804 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_837 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_848 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_859 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_4 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_623 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_667 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_612 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_634 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_678 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_645 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_601 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_656 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_689 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1813 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1824 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1835 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1802 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1868 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1857 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1879 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1846 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_464 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_453 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_475 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_420 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_431 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_486 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_442 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_497 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1109 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1610 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1654 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1665 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1621 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1676 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1632 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1687 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1643 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1698 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_250 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_272 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_261 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_283 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_294 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2130 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2174 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1451 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1495 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1440 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2185 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1462 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2141 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2196 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1473 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2152 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1484 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2163 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1292 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1270 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1281 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_827 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_816 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_838 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_849 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_805 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_5 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_668 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_613 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_679 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_624 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_635 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_646 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_602 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_657 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1869 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1814 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1858 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1803 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1825 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1836 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1847 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_410 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_465 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_454 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_476 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_421 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_432 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_487 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_443 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_498 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1611 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1655 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1699 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1600 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1666 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1622 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1677 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1633 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1688 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1644 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_251 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_240 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_273 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_262 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_284 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_295 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2131 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2120 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2142 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2153 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2164 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2175 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1452 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1496 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1441 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2186 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1463 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2197 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1474 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1430 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1485 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1260 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1271 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1293 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1282 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_828 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_817 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_839 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_806 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1090 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_6 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_669 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_614 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_625 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_636 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_647 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_603 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_658 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1815 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1859 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1804 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1826 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1837 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1848 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_411 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_400 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_422 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_433 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_444 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_466 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_455 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_477 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_488 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_499 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1601 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1656 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1667 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1612 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1623 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1678 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1634 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1689 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1645 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_252 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_263 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_274 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_230 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_285 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_241 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_296 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1453 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2176 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2121 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1442 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2187 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2132 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2143 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1420 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2198 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1431 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2154 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2110 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2165 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1497 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1464 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1475 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1486 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1294 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1283 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1250 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1261 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1272 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_829 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_818 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_807 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1091 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1080 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_7 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_615 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_626 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_604 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_659 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_637 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_648 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1816 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1805 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1827 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1838 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1849 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_467 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_412 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_456 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_401 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_423 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_434 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_445 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_478 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_489 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_990 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1602 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1613 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1624 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1635 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1657 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1668 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1679 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1646 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_253 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_220 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_264 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_275 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_231 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_286 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_242 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_297 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1454 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2177 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2122 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1443 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2188 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2133 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1410 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1465 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2144 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1421 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1476 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2100 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2199 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2155 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1432 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1487 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2111 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2166 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1498 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1295 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1240 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1284 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1251 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1262 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1273 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_808 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_819 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1081 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1092 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1070 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_8 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_616 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_627 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_638 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_649 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_605 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1817 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1806 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1828 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1839 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_413 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_457 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_402 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_479 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_424 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_468 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_435 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_446 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_980 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_991 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1658 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1603 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1647 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1669 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1614 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1625 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1636 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_254 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_221 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_210 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_265 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_276 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_232 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_287 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_243 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_298 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2101 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2112 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1455 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2178 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2123 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1400 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1499 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2167 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1444 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2189 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2134 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1411 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1466 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2145 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1422 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1477 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2156 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1433 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1488 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1296 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1241 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1285 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1252 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1263 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1274 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1230 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_809 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1060 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1082 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1093 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1071 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_9 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_617 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_628 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_639 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_606 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1818 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1807 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1829 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_414 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_458 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_403 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_425 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_469 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_436 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_447 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_981 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_992 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_970 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1659 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1604 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1648 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1615 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1626 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1637 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_200 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_211 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_222 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_233 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_255 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_266 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_277 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_288 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_244 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_299 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1401 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2124 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2135 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2146 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2102 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2113 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2179 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2168 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1445 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1456 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1412 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1467 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1423 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1478 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2157 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1434 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1489 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1990 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1242 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1231 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1253 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1220 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1297 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1286 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1264 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1275 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1083 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1094 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1050 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1061 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1072 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_618 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_607 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_629 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1819 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1808 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_415 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_404 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_426 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_459 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_437 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_448 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_971 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_960 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_982 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_993 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1605 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1649 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1616 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1627 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1638 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_256 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_201 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_267 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_212 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_223 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_234 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_245 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_278 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_289 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_790 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1402 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2125 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2169 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2136 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1413 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1424 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2147 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2103 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2158 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1435 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2114 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1446 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1457 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1468 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1479 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1980 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1991 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1243 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1232 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1254 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1210 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1265 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1221 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1276 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1298 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1287 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1084 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1095 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1040 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1051 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1062 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1073 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_608 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_619 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1809 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_405 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_427 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_416 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_438 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_449 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_983 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_972 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_994 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_950 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_961 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1606 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1617 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1628 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1639 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_257 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_202 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_268 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_213 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_224 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_279 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_235 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_246 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_780 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_791 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1403 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2126 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1447 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2115 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2137 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1458 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1414 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1469 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2148 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1425 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2104 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2159 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1436 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1970 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1981 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1992 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1299 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1244 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1288 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1233 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1200 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1255 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1211 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1266 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1222 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1277 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1085 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1030 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1096 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1041 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1052 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1063 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1074 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_609 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_406 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_428 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_417 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_439 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_984 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_973 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_940 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_995 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_951 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_962 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1607 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1618 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1629 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_258 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_203 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_269 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_214 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_225 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_236 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_247 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_770 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_781 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_792 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2127 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1448 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2116 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2138 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1459 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1404 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1415 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2149 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1426 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2105 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1437 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1971 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1960 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1982 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1993 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1201 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1245 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1289 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1234 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1256 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1212 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1267 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1223 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1278 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1790 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1031 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1042 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1020 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1086 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1075 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1097 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1053 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1064 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_407 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_429 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_418 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_930 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_985 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_974 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_941 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_996 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_952 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_963 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1608 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1619 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_204 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_215 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_259 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_226 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_237 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_248 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_771 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_760 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_782 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_793 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2128 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2117 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2106 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1449 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1405 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1416 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2139 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1427 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1438 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1972 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1961 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1983 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1994 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1950 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_590 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1202 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1213 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1224 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1246 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1235 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1257 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1268 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1279 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1780 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1791 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1032 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1076 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1043 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1054 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1010 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1065 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1021 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1087 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1098 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_408 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_419 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_931 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_920 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_942 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_953 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_986 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_975 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_997 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_964 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1609 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_205 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_216 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_227 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_238 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_249 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_772 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_783 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_794 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_750 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_761 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2129 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2118 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1406 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1417 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2107 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1439 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1428 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1973 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1962 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1940 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1951 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1984 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1995 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_580 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_591 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1247 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1236 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1203 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1258 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1214 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1225 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1269 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1770 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1781 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1792 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1088 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1033 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1077 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1044 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1099 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1000 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1055 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1011 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1066 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1022 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_409 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_987 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_932 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_976 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_921 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_943 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_954 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_910 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_965 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_998 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_206 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_217 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_228 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_239 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_773 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_784 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_740 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_795 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_751 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_762 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_90 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2119 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1407 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1418 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1429 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2108 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1974 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1963 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1930 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1985 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1941 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1996 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1952 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_570 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_581 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_592 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1237 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1248 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1204 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1259 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1215 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1226 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1760 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1771 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1782 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1793 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1089 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1034 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1078 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1023 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1045 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1001 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1056 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1012 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1067 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1590 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_933 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_977 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_922 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_988 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_944 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_999 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_900 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_955 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_911 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_966 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_207 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_218 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_229 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_774 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_763 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_785 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_730 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_741 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_796 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_752 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_80 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_91 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1408 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1419 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2109 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1975 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1920 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1964 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1931 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1986 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1942 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1997 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1953 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_571 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_560 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_582 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_593 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1238 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1249 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1205 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1216 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1227 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1761 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1772 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1783 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1794 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1750 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_390 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1024 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1002 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1013 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1035 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1079 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1046 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1057 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1068 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1580 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1591 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_901 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_912 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_934 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_978 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_923 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_989 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_945 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_956 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_967 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_219 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_208 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_720 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_731 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_70 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_742 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_753 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_81 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_775 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_764 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_786 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_797 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_92 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1409 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1921 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1910 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1965 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1976 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1932 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1987 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1943 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1998 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1954 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_561 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_572 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_583 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_594 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_550 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1206 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1239 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1217 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1228 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1762 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1751 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1740 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1773 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1784 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1795 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_380 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_391 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1036 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1025 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1047 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1003 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1058 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1014 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1069 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1570 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1581 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1592 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2090 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_935 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_924 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_902 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_913 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_979 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_946 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_957 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_968 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_209 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_776 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_721 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_765 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_60 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_732 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_787 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_71 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_743 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_754 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_82 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_710 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_93 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_798 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1922 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1911 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1933 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1944 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1900 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1955 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1966 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1977 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1988 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1999 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_562 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_573 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_584 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_540 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_595 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_551 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1207 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1218 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1229 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1763 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1752 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1774 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1730 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1785 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1741 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1796 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_370 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_381 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_392 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1037 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1026 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1048 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1004 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1059 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1015 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1560 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1571 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1582 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1593 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2080 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_2091 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1390 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_925 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_936 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_947 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_903 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_958 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_914 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_969 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_777 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_722 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_94 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_766 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_711 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_61 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_733 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_788 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_72 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_744 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_799 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_700 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_755 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1923 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1967 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1912 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1978 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1934 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1945 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1901 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1956 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1989 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_563 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_530 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_574 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_585 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_541 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_596 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_552 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1208 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1219 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1764 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1753 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1720 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1775 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1731 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1786 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1742 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
Xunit_cap_1797 m5_8380_287100# m4_8380_242120# m5_8380_287100# unit_cap
.ends

.subckt converter power_stage_0/s4 power_stage_0/s3 power_stage_0/s2 power_stage_0/s1
+ power_stage_0/nmos_waffle_36x36_1/dw_n5900_n5900# power_stage_0/nmos_waffle_36x36_0/dw_n5900_n5900#
+ VSUBS power_stage_0/VN power_stage_0/fc1 power_stage_0/VP power_stage_0/out power_stage_0/fc2
Xpower_stage_0 power_stage_0/nmos_waffle_36x36_1/dw_n5900_n5900# power_stage_0/VP
+ power_stage_0/nmos_waffle_36x36_0/dw_n5900_n5900# power_stage_0/s4 power_stage_0/s3
+ power_stage_0/s2 power_stage_0/s1 power_stage_0/fc2 power_stage_0/VN power_stage_0/out
+ power_stage_0/fc1 VSUBS power_stage
Xflying_cap_0 power_stage_0/fc2 power_stage_0/fc1 flying_cap
.ends

.subckt level_shifter level_shifter_0/cruzados_0/VH level_shifter_0/inv_1_8_0/VDD
+ level_shifter_0/inv_400_0/OUT level_shifter_0/inv_1_8_0/GND level_shifter_0/cruzados_0/IN2
X0 a_1660_2346# level_shifter_0/cruzados_0/OUT level_shifter_0/cruzados_0/VH level_shifter_0/cruzados_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+11p pd=4.58e+06u as=8.236e+13p ps=5.7902e+08u w=2e+06u l=500000u
X1 level_shifter_0/inv_400_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/inv_1_8_0/GND level_shifter_0/inv_1_8_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=5.8e+13p pd=4.058e+08u as=8.584e+13p ps=6.0418e+08u w=2e+07u l=500000u
X2 level_shifter_0/inv_1_8_0/GND level_shifter_0/cruzados_0/IN2 level_shifter_0/inv_400_0/IN level_shifter_0/inv_1_8_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.45e+13p ps=1.029e+08u w=1e+07u l=500000u
X3 level_shifter_0/cruzados_0/VH level_shifter_0/inv_400_0/IN level_shifter_0/inv_400_0/OUT level_shifter_0/cruzados_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=5.8e+13p ps=4.058e+08u w=2e+07u l=500000u
X4 level_shifter_0/inv_400_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/cruzados_0/VH level_shifter_0/cruzados_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X5 level_shifter_0/inv_1_8_0/GND level_shifter_0/inv_400_0/IN level_shifter_0/inv_400_0/OUT level_shifter_0/inv_1_8_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X6 level_shifter_0/inv_400_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/inv_1_8_0/GND level_shifter_0/inv_1_8_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X7 level_shifter_0/cruzados_0/VH level_shifter_0/cruzados_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/cruzados_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1.45e+13p ps=1.029e+08u w=1e+07u l=500000u
X8 level_shifter_0/inv_400_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/cruzados_0/VH level_shifter_0/cruzados_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X9 level_shifter_0/inv_400_0/IN level_shifter_0/cruzados_0/OUT level_shifter_0/cruzados_0/VH level_shifter_0/cruzados_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+07u l=500000u
X10 level_shifter_0/cruzados_0/IN1 level_shifter_0/cruzados_0/IN2 level_shifter_0/inv_1_8_0/GND level_shifter_0/inv_1_8_0/GND sky130_fd_pr__nfet_01v8 ad=9.7e+11p pd=7.94e+06u as=9.7e+11p ps=7.94e+06u w=1e+06u l=150000u
X11 level_shifter_0/inv_400_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/inv_1_8_0/GND level_shifter_0/inv_1_8_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X12 level_shifter_0/inv_1_8_0/GND level_shifter_0/inv_400_0/IN level_shifter_0/inv_400_0/OUT level_shifter_0/inv_1_8_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X13 level_shifter_0/inv_1_8_0/GND level_shifter_0/inv_400_0/IN level_shifter_0/inv_400_0/OUT level_shifter_0/inv_1_8_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X14 level_shifter_0/inv_400_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/cruzados_0/VH level_shifter_0/cruzados_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X15 level_shifter_0/inv_400_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/inv_1_8_0/GND level_shifter_0/inv_1_8_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X16 level_shifter_0/inv_400_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/cruzados_0/VH level_shifter_0/cruzados_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X17 level_shifter_0/inv_1_8_0/GND level_shifter_0/cruzados_0/IN2 level_shifter_0/cruzados_0/IN1 level_shifter_0/inv_1_8_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 level_shifter_0/cruzados_0/VH level_shifter_0/cruzados_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/cruzados_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+07u l=500000u
X19 level_shifter_0/inv_400_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/cruzados_0/VH level_shifter_0/cruzados_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X20 level_shifter_0/cruzados_0/IN1 level_shifter_0/cruzados_0/IN2 level_shifter_0/inv_1_8_0/VDD level_shifter_0/inv_1_8_0/VDD sky130_fd_pr__pfet_01v8 ad=9.7e+11p pd=7.94e+06u as=9.7e+11p ps=7.94e+06u w=1e+06u l=150000u
X21 level_shifter_0/cruzados_0/OUT level_shifter_0/cruzados_0/IN1 level_shifter_0/inv_1_8_0/GND level_shifter_0/inv_1_8_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=2.32e+12p pd=1.716e+07u as=0p ps=0u w=4e+06u l=500000u
X22 level_shifter_0/inv_1_8_0/GND level_shifter_0/inv_400_0/IN level_shifter_0/inv_400_0/OUT level_shifter_0/inv_1_8_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X23 level_shifter_0/cruzados_0/VH level_shifter_0/inv_400_0/IN level_shifter_0/inv_400_0/OUT level_shifter_0/cruzados_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X24 level_shifter_0/inv_1_8_0/GND level_shifter_0/inv_400_0/IN level_shifter_0/inv_400_0/OUT level_shifter_0/inv_1_8_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X25 level_shifter_0/cruzados_0/IN1 level_shifter_0/cruzados_0/IN2 level_shifter_0/inv_1_8_0/VDD level_shifter_0/inv_1_8_0/VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 level_shifter_0/cruzados_0/VH level_shifter_0/inv_400_0/IN level_shifter_0/inv_400_0/OUT level_shifter_0/cruzados_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X27 level_shifter_0/cruzados_0/IN1 level_shifter_0/cruzados_0/IN2 level_shifter_0/inv_1_8_0/GND level_shifter_0/inv_1_8_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 level_shifter_0/inv_400_0/IN level_shifter_0/cruzados_0/IN2 level_shifter_0/inv_1_8_0/GND level_shifter_0/inv_1_8_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+07u l=500000u
X29 level_shifter_0/cruzados_0/VH level_shifter_0/inv_400_0/IN level_shifter_0/inv_400_0/OUT level_shifter_0/cruzados_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X30 level_shifter_0/inv_1_8_0/VDD level_shifter_0/cruzados_0/IN2 level_shifter_0/cruzados_0/IN1 level_shifter_0/inv_1_8_0/VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 level_shifter_0/inv_1_8_0/GND level_shifter_0/inv_400_0/IN level_shifter_0/inv_400_0/OUT level_shifter_0/inv_1_8_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X32 level_shifter_0/cruzados_0/OUT a_1660_2346# level_shifter_0/cruzados_0/VH level_shifter_0/cruzados_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X33 level_shifter_0/inv_400_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/inv_1_8_0/GND level_shifter_0/inv_1_8_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X34 level_shifter_0/inv_400_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/inv_1_8_0/GND level_shifter_0/inv_1_8_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X35 level_shifter_0/inv_400_0/IN level_shifter_0/cruzados_0/IN2 level_shifter_0/inv_1_8_0/GND level_shifter_0/inv_1_8_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+07u l=500000u
X36 level_shifter_0/inv_1_8_0/GND level_shifter_0/cruzados_0/IN2 level_shifter_0/inv_400_0/IN level_shifter_0/inv_1_8_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+07u l=500000u
X37 level_shifter_0/cruzados_0/OUT level_shifter_0/cruzados_0/IN1 level_shifter_0/inv_1_8_0/GND level_shifter_0/inv_1_8_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X38 level_shifter_0/inv_1_8_0/GND level_shifter_0/inv_400_0/IN level_shifter_0/inv_400_0/OUT level_shifter_0/inv_1_8_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X39 level_shifter_0/inv_400_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/inv_1_8_0/GND level_shifter_0/inv_1_8_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X40 level_shifter_0/inv_1_8_0/GND level_shifter_0/cruzados_0/IN2 a_1660_2346# level_shifter_0/inv_1_8_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=2.32e+12p ps=1.716e+07u w=4e+06u l=500000u
X41 level_shifter_0/inv_400_0/IN level_shifter_0/cruzados_0/OUT level_shifter_0/cruzados_0/VH level_shifter_0/cruzados_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+07u l=500000u
X42 level_shifter_0/inv_400_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/cruzados_0/VH level_shifter_0/cruzados_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X43 level_shifter_0/inv_400_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/cruzados_0/VH level_shifter_0/cruzados_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X44 level_shifter_0/inv_400_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/inv_1_8_0/GND level_shifter_0/inv_1_8_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X45 level_shifter_0/inv_1_8_0/GND level_shifter_0/cruzados_0/IN2 level_shifter_0/inv_400_0/IN level_shifter_0/inv_1_8_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+07u l=500000u
X46 level_shifter_0/inv_400_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/cruzados_0/VH level_shifter_0/cruzados_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X47 level_shifter_0/inv_1_8_0/GND level_shifter_0/cruzados_0/IN2 level_shifter_0/cruzados_0/IN1 level_shifter_0/inv_1_8_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X48 level_shifter_0/cruzados_0/IN1 level_shifter_0/cruzados_0/IN2 level_shifter_0/inv_1_8_0/VDD level_shifter_0/inv_1_8_0/VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X49 level_shifter_0/inv_1_8_0/GND level_shifter_0/inv_400_0/IN level_shifter_0/inv_400_0/OUT level_shifter_0/inv_1_8_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X50 level_shifter_0/inv_400_0/IN level_shifter_0/cruzados_0/OUT level_shifter_0/cruzados_0/VH level_shifter_0/cruzados_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+07u l=500000u
X51 level_shifter_0/cruzados_0/VH level_shifter_0/cruzados_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/cruzados_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+07u l=500000u
X52 level_shifter_0/inv_400_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/cruzados_0/VH level_shifter_0/cruzados_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X53 level_shifter_0/inv_400_0/IN level_shifter_0/cruzados_0/IN2 level_shifter_0/inv_1_8_0/GND level_shifter_0/inv_1_8_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+07u l=500000u
X54 level_shifter_0/inv_1_8_0/GND level_shifter_0/cruzados_0/IN2 level_shifter_0/inv_400_0/IN level_shifter_0/inv_1_8_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+07u l=500000u
X55 level_shifter_0/inv_400_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/cruzados_0/VH level_shifter_0/cruzados_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X56 level_shifter_0/cruzados_0/VH level_shifter_0/inv_400_0/IN level_shifter_0/inv_400_0/OUT level_shifter_0/cruzados_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X57 level_shifter_0/inv_1_8_0/GND level_shifter_0/cruzados_0/IN1 level_shifter_0/cruzados_0/OUT level_shifter_0/inv_1_8_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X58 level_shifter_0/cruzados_0/VH level_shifter_0/cruzados_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/cruzados_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+07u l=500000u
X59 a_1660_2346# level_shifter_0/cruzados_0/IN2 level_shifter_0/inv_1_8_0/GND level_shifter_0/inv_1_8_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X60 level_shifter_0/cruzados_0/VH level_shifter_0/inv_400_0/IN level_shifter_0/inv_400_0/OUT level_shifter_0/cruzados_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X61 level_shifter_0/inv_400_0/IN level_shifter_0/cruzados_0/IN2 level_shifter_0/inv_1_8_0/GND level_shifter_0/inv_1_8_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+07u l=500000u
X62 level_shifter_0/cruzados_0/VH level_shifter_0/inv_400_0/IN level_shifter_0/inv_400_0/OUT level_shifter_0/cruzados_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X63 level_shifter_0/inv_400_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/inv_1_8_0/GND level_shifter_0/inv_1_8_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X64 level_shifter_0/inv_400_0/IN level_shifter_0/cruzados_0/OUT level_shifter_0/cruzados_0/VH level_shifter_0/cruzados_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+07u l=500000u
X65 level_shifter_0/cruzados_0/VH level_shifter_0/inv_400_0/IN level_shifter_0/inv_400_0/OUT level_shifter_0/cruzados_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X66 level_shifter_0/inv_1_8_0/VDD level_shifter_0/cruzados_0/IN2 level_shifter_0/cruzados_0/IN1 level_shifter_0/inv_1_8_0/VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X67 level_shifter_0/cruzados_0/VH level_shifter_0/cruzados_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/cruzados_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+07u l=500000u
X68 level_shifter_0/cruzados_0/VH level_shifter_0/inv_400_0/IN level_shifter_0/inv_400_0/OUT level_shifter_0/cruzados_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X69 level_shifter_0/inv_400_0/OUT level_shifter_0/inv_400_0/IN level_shifter_0/inv_1_8_0/GND level_shifter_0/inv_1_8_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X70 level_shifter_0/inv_1_8_0/GND level_shifter_0/cruzados_0/IN2 level_shifter_0/inv_400_0/IN level_shifter_0/inv_1_8_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+07u l=500000u
X71 level_shifter_0/cruzados_0/VH level_shifter_0/inv_400_0/IN level_shifter_0/inv_400_0/OUT level_shifter_0/cruzados_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X72 level_shifter_0/cruzados_0/IN1 level_shifter_0/cruzados_0/IN2 level_shifter_0/inv_1_8_0/GND level_shifter_0/inv_1_8_0/GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X73 level_shifter_0/inv_1_8_0/GND level_shifter_0/inv_400_0/IN level_shifter_0/inv_400_0/OUT level_shifter_0/inv_1_8_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X74 level_shifter_0/inv_400_0/IN level_shifter_0/cruzados_0/OUT level_shifter_0/cruzados_0/VH level_shifter_0/cruzados_0/VH sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+07u l=500000u
X75 level_shifter_0/inv_400_0/IN level_shifter_0/cruzados_0/IN2 level_shifter_0/inv_1_8_0/GND level_shifter_0/inv_1_8_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+07u l=500000u
X76 a_1660_2346# level_shifter_0/cruzados_0/IN2 level_shifter_0/inv_1_8_0/GND level_shifter_0/inv_1_8_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X77 level_shifter_0/inv_1_8_0/GND level_shifter_0/inv_400_0/IN level_shifter_0/inv_400_0/OUT level_shifter_0/inv_1_8_0/GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
.ends

.subckt core D4 D2 D3 D1 converter_0/power_stage_0/nmos_waffle_36x36_1/dw_n5900_n5900#
+ converter_0/power_stage_0/VP VLS converter_0/power_stage_0/out converter_0/power_stage_0/nmos_waffle_36x36_0/dw_n5900_n5900#
+ converter_0/power_stage_0/fc1 VDD converter_0/power_stage_0/fc2 VSUBS
Xconverter_0 converter_0/power_stage_0/s4 converter_0/power_stage_0/s3 converter_0/power_stage_0/s2
+ converter_0/power_stage_0/s1 converter_0/power_stage_0/nmos_waffle_36x36_1/dw_n5900_n5900#
+ converter_0/power_stage_0/nmos_waffle_36x36_0/dw_n5900_n5900# VSUBS VSUBS converter_0/power_stage_0/fc1
+ converter_0/power_stage_0/VP converter_0/power_stage_0/out converter_0/power_stage_0/fc2
+ converter
Xlevel_shifter_0 VLS VDD converter_0/power_stage_0/s1 VSUBS D1 level_shifter
Xlevel_shifter_1 VLS VDD converter_0/power_stage_0/s2 VSUBS D2 level_shifter
Xlevel_shifter_2 VLS VDD converter_0/power_stage_0/s3 VSUBS D3 level_shifter
Xlevel_shifter_3 VLS VDD converter_0/power_stage_0/s4 VSUBS D4 level_shifter
.ends

.subckt interleaved core_1/VLS core_1/D4 core_1/D3 core_1/D2 core_1/D1 VH core_1/VDD
+ core_1/converter_0/power_stage_0/fc2 core_0/D4 core_0/D3 core_0/D2 core_0/D1 core_0/converter_0/power_stage_0/fc2
+ Vout2 Vout1 core_1/converter_0/power_stage_0/fc1 core_0/VLS core_0/converter_0/power_stage_0/fc1
+ GND
Xstack30um_1_5_29 Vout2 stack30um_1_5
Xstack30um_1_5_19 Vout1 stack30um_1_5
Xstack30um_1_5_18 Vout1 stack30um_1_5
Xpower_pad_1_5_0 GND power_pad_1_5
Xpower_pad_1_5_1 Vout1 power_pad_1_5
Xpower_pad_1_5_2 Vout2 power_pad_1_5
Xstack30um_1_5_0 GND stack30um_1_5
Xstack30um_1_5_1 GND stack30um_1_5
Xstack30um_1_5_2 GND stack30um_1_5
Xstack30um_1_5_3 GND stack30um_1_5
Xstack30um_1_5_4 GND stack30um_1_5
Xstack30um_1_5_5 GND stack30um_1_5
Xstack30um_1_5_6 GND stack30um_1_5
Xstack30um_1_5_8 GND stack30um_1_5
Xstack30um_1_5_7 GND stack30um_1_5
Xstack30um_1_5_9 GND stack30um_1_5
Xpower_pad_3_5_0 VH power_pad_3_5
Xpower_pad_3_5_1 VH power_pad_3_5
Xstack30um_1_5_40 Vout2 stack30um_1_5
Xstack30um_1_5_41 Vout2 stack30um_1_5
Xstack30um_1_5_30 Vout2 stack30um_1_5
Xstack30um_1_5_31 Vout2 stack30um_1_5
Xstack30um_1_5_32 Vout2 stack30um_1_5
Xstack30um_1_5_10 GND stack30um_1_5
Xstack30um_1_5_21 Vout1 stack30um_1_5
Xstack30um_1_5_20 Vout1 stack30um_1_5
Xstack30um_1_5_33 Vout2 stack30um_1_5
Xstack30um_1_5_11 GND stack30um_1_5
Xstack30um_1_5_22 Vout1 stack30um_1_5
Xstack30um_1_5_34 Vout2 stack30um_1_5
Xcore_0 core_0/D4 core_0/D2 core_0/D3 core_0/D1 VH VH core_0/VLS Vout1 VH core_0/converter_0/power_stage_0/fc1
+ core_1/VDD core_0/converter_0/power_stage_0/fc2 GND core
Xstack30um_1_5_12 GND stack30um_1_5
Xstack30um_1_5_23 Vout1 stack30um_1_5
Xcore_1 core_1/D4 core_1/D2 core_1/D3 core_1/D1 VH VH core_1/VLS Vout2 VH core_1/converter_0/power_stage_0/fc1
+ core_1/VDD core_1/converter_0/power_stage_0/fc2 GND core
Xstack30um_1_5_35 Vout2 stack30um_1_5
Xstack30um_1_5_13 GND stack30um_1_5
Xstack30um_1_5_24 Vout1 stack30um_1_5
Xstack30um_1_5_36 Vout2 stack30um_1_5
Xstack30um_1_5_14 GND stack30um_1_5
Xstack30um_1_5_25 Vout1 stack30um_1_5
Xstack30um_1_5_37 Vout2 stack30um_1_5
Xstack30um_1_5_26 Vout2 stack30um_1_5
Xstack30um_1_5_15 GND stack30um_1_5
Xstack30um_1_5_38 Vout2 stack30um_1_5
Xstack30um_1_5_27 Vout2 stack30um_1_5
Xstack30um_1_5_16 Vout1 stack30um_1_5
Xstack30um_1_5_39 Vout2 stack30um_1_5
Xstack30um_1_5_28 Vout2 stack30um_1_5
Xstack30um_1_5_17 Vout1 stack30um_1_5
.ends

.subckt calibration_pad m5_0_0#
Xstack30um_1_5_0 m5_0_0# stack30um_1_5
.ends

.subckt sky130_fd_pr__res_generic_po_KL3G6K a_n3000_n3540# a_n3000_3110#
R0 a_n3000_n3540# a_n3000_3110# sky130_fd_pr__res_generic_po w=3e+07u l=3.11e+07u
.ends

.subckt calibration
Xcalibration_pad_0 calibration_pad_0/m5_0_0# calibration_pad
Xsky130_fd_pr__res_generic_po_KL3G6K_0 calibration_pad_0/m5_0_0# calibration_pad_1/m5_0_0#
+ sky130_fd_pr__res_generic_po_KL3G6K
Xcalibration_pad_1 calibration_pad_1/m5_0_0# calibration_pad
.ends

.subckt inductors m3_0_80000# m3_0_123200# m3_0_36800# m3_0_15200# m3_1000_162000#
Xcalibration_pad_0 m1_407000_47000# calibration_pad
Xcalibration_pad_1 calibration_pad_1/m5_0_0# calibration_pad
Xcalibration_1 calibration
Xcalibration_0 calibration
R0 m3_0_123200# m3_0_80000# sky130_fd_pr__res_generic_m3 w=5e+06u l=1e+06u
R1 m3_0_36800# m3_0_15200# sky130_fd_pr__res_generic_m3 w=5e+06u l=1e+06u
.ends

.subckt topmodule inductors_0/m3_0_123200# VLS2 VLS1 VH_4 inductors_0/m3_1000_162000#
+ VH_3 FC2_1 VH_2 D8 D7 D6 D5 D4 D3 D2 inductors_0/m3_0_36800# FC2_1b D1 FC2_2b GND_2
+ interleaved_0/Vout1 inductors_0/m3_0_15200# FC1_1 interleaved_0/VH FC1_2 FC2_2 VDD
+ interleaved_0/Vout2 FC1_1b FC1_2b inductors_0/m3_0_80000# VSUBS
Xunit_cap_73 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_62 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_51 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_40 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_74 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_63 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_52 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_41 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_30 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_75 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_64 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_53 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_42 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_20 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_31 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_76 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_65 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_54 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_21 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_32 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_43 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_10 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_77 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_66 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_55 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_23 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_22 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_34 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_33 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_12 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_44 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_11 VSUBS interleaved_0/VH VSUBS unit_cap
Xinterleaved_0 VLS2 D8 D7 D6 D5 interleaved_0/VH VDD FC2_2 D4 D3 D2 D1 FC1_2 interleaved_0/Vout2
+ interleaved_0/Vout1 FC2_1 VLS1 FC1_1 VSUBS interleaved
Xunit_cap_78 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_68 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_67 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_57 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_56 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_79 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_35 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_24 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_13 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_45 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_46 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_69 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_58 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_36 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_25 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_14 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_47 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_59 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_37 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_26 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_15 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_48 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_38 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_27 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_16 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_49 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_39 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_28 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_17 VSUBS interleaved_0/VH VSUBS unit_cap
Xinductors_0 inductors_0/m3_0_80000# inductors_0/m3_0_123200# inductors_0/m3_0_36800#
+ inductors_0/m3_0_15200# inductors_0/m3_1000_162000# inductors
Xunit_cap_18 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_29 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_19 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_0 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_1 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_2 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_3 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_4 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_5 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_6 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_7 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_8 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_9 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_70 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_81 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_80 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_71 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_82 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_60 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_72 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_61 VSUBS interleaved_0/VH VSUBS unit_cap
Xunit_cap_50 VSUBS interleaved_0/VH VSUBS unit_cap
R0 interleaved_0/VH VH_2 sky130_fd_pr__res_generic_m3 w=2.6e+07u l=500000u
R1 VSUBS GND_2 sky130_fd_pr__res_generic_m3 w=8e+07u l=500000u
R2 FC1_2b FC1_2 sky130_fd_pr__res_generic_m3 w=5e+06u l=5e+06u
R3 interleaved_0/VH VH_3 sky130_fd_pr__res_generic_m3 w=2.6e+07u l=500000u
R4 FC2_1 FC2_1b sky130_fd_pr__res_generic_m3 w=5e+06u l=5e+06u
R5 interleaved_0/VH VH_4 sky130_fd_pr__res_generic_m3 w=2.6e+07u l=300000u
R6 FC1_1b FC1_1 sky130_fd_pr__res_generic_m3 w=5e+06u l=5e+06u
R7 FC2_2 FC2_2b sky130_fd_pr__res_generic_m3 w=5e+06u l=5e+06u
.ends

.subckt user_analog_project_wrapper gpio_analog[0] gpio_analog[10] gpio_analog[11]
+ gpio_analog[12] gpio_analog[13] gpio_analog[14] gpio_analog[15] gpio_analog[16]
+ gpio_analog[17] gpio_analog[1] gpio_analog[2] gpio_analog[3] gpio_analog[4] gpio_analog[5]
+ gpio_analog[6] gpio_analog[7] gpio_analog[8] gpio_analog[9] gpio_noesd[0] gpio_noesd[10]
+ gpio_noesd[11] gpio_noesd[12] gpio_noesd[13] gpio_noesd[14] gpio_noesd[15] gpio_noesd[16]
+ gpio_noesd[17] gpio_noesd[1] gpio_noesd[2] gpio_noesd[3] gpio_noesd[4] gpio_noesd[5]
+ gpio_noesd[6] gpio_noesd[7] gpio_noesd[8] gpio_noesd[9] io_analog[0] io_analog[10]
+ io_analog[1] io_analog[2] io_analog[3] io_analog[7] io_analog[8] io_analog[9] io_analog[4]
+ io_analog[5] io_analog[6] io_clamp_high[0] io_clamp_high[1] io_clamp_high[2] io_clamp_low[0]
+ io_clamp_low[1] io_clamp_low[2] io_in[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21]
+ io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_in[8] io_in[9] io_in_3v3[0] io_in_3v3[10] io_in_3v3[11] io_in_3v3[12]
+ io_in_3v3[13] io_in_3v3[14] io_in_3v3[15] io_in_3v3[16] io_in_3v3[17] io_in_3v3[18]
+ io_in_3v3[19] io_in_3v3[1] io_in_3v3[20] io_in_3v3[21] io_in_3v3[22] io_in_3v3[23]
+ io_in_3v3[24] io_in_3v3[25] io_in_3v3[26] io_in_3v3[2] io_in_3v3[3] io_in_3v3[4]
+ io_in_3v3[5] io_in_3v3[6] io_in_3v3[7] io_in_3v3[8] io_in_3v3[9] io_oeb[0] io_oeb[10]
+ io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18]
+ io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25]
+ io_oeb[26] io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8]
+ io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15]
+ io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22]
+ io_out[23] io_out[24] io_out[25] io_out[26] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100] la_data_in[101]
+ la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105] la_data_in[106]
+ la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110] la_data_in[111]
+ la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115] la_data_in[116]
+ la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120] la_data_in[121]
+ la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125] la_data_in[126]
+ la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15] la_data_in[16]
+ la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20] la_data_in[21]
+ la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26] la_data_in[27]
+ la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31] la_data_in[32]
+ la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37] la_data_in[38]
+ la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42] la_data_in[43]
+ la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48] la_data_in[49]
+ la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53] la_data_in[54]
+ la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59] la_data_in[5]
+ la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64] la_data_in[65]
+ la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6] la_data_in[70]
+ la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75] la_data_in[76]
+ la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80] la_data_in[81]
+ la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86] la_data_in[87]
+ la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91] la_data_in[92]
+ la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97] la_data_in[98]
+ la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101] la_data_out[102]
+ la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106] la_data_out[107]
+ la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110] la_data_out[111]
+ la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115] la_data_out[116]
+ la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11] la_data_out[120]
+ la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124] la_data_out[125]
+ la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24]
+ la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29]
+ la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34]
+ la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39]
+ la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44]
+ la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49]
+ la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54]
+ la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59]
+ la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[64]
+ la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68] la_data_out[69]
+ la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73] la_data_out[74]
+ la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78] la_data_out[79]
+ la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83] la_data_out[84]
+ la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88] la_data_out[89]
+ la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93] la_data_out[94]
+ la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98] la_data_out[99]
+ la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104]
+ la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109] la_oenb[10] la_oenb[110]
+ la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117]
+ la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121] la_oenb[122] la_oenb[123]
+ la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65]
+ la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6] la_oenb[70] la_oenb[71]
+ la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76] la_oenb[77] la_oenb[78]
+ la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84]
+ la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89] la_oenb[8] la_oenb[90]
+ la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97]
+ la_oenb[98] la_oenb[99] la_oenb[9] user_clock2 user_irq[0] user_irq[1] user_irq[2]
+ vccd1 vccd2 vdda1 vdda2 vssa1 vssa2 vssd1 vssd2 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0]
+ wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15]
+ wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20]
+ wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26]
+ wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31]
+ wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9]
+ wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13]
+ wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19]
+ wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24]
+ wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2]
+ wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6]
+ wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3]
+ wbs_stb_i wbs_we_i
Xtopmodule_0 gpio_noesd[14] vdda1 vdda2 io_analog[2] vssd2 io_analog[3] io_analog[1]
+ io_analog[7] io_in[10] io_in[9] io_in[8] io_in[7] io_in[17] io_in[18] io_in[19]
+ gpio_noesd[16] gpio_noesd[6] io_in[20] gpio_noesd[5] vssa1 io_analog[6] gpio_noesd[17]
+ io_analog[9] io_analog[8] io_analog[10] io_analog[0] vccd1 io_analog[4] gpio_noesd[7]
+ gpio_noesd[9] gpio_noesd[15] io_analog[5] topmodule
.ends

