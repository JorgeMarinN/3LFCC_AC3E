magic
tech sky130A
timestamp 1667913101
<< error_s >>
rect 25 1650 75 1657
rect 575 1650 625 1657
rect 660 1650 1090 1675
rect 1125 1650 1175 1657
rect 2 1212 4 1638
rect 265 1473 385 1485
rect 265 1377 277 1473
rect 373 1377 385 1473
rect 265 1365 385 1377
rect 815 1473 935 1485
rect 815 1377 827 1473
rect 923 1377 935 1473
rect 815 1365 935 1377
rect 1365 1473 1485 1485
rect 1365 1377 1377 1473
rect 1473 1377 1485 1473
rect 1365 1365 1485 1377
rect 1650 1125 1657 1175
rect 2 1096 17 1102
rect -15 654 0 671
rect 2 662 4 1088
rect 265 923 385 935
rect 265 827 277 923
rect 373 827 385 923
rect 265 815 385 827
rect 815 923 935 935
rect 815 827 827 923
rect 923 827 935 923
rect 815 815 935 827
rect 1365 923 1485 935
rect 1365 827 1377 923
rect 1473 827 1485 923
rect 1365 815 1485 827
rect 1650 689 1675 1090
rect 2 648 17 654
rect 1650 575 1657 625
rect 2 112 4 538
rect 265 373 385 385
rect 265 277 277 373
rect 373 277 385 373
rect 265 265 385 277
rect 815 373 935 385
rect 815 277 827 373
rect 923 277 935 373
rect 815 265 935 277
rect 1365 373 1485 385
rect 1365 277 1377 373
rect 1473 277 1485 373
rect 1365 265 1485 277
rect 1650 25 1657 75
rect 0 2 2 17
rect 112 2 538 4
rect 648 2 654 17
rect 662 2 1088 4
rect 1096 2 1102 17
rect 1212 2 1638 4
rect 0 0 17 2
use nmos_drain  nmos_drain_0
timestamp 1667912669
transform 1 0 550 0 1 0
box -15 0 575 575
use nmos_drain  nmos_drain_1
timestamp 1667912669
transform 1 0 0 0 1 550
box -15 0 575 575
use nmos_drain  nmos_drain_2
timestamp 1667912669
transform 1 0 1100 0 1 550
box -15 0 575 575
use nmos_drain  nmos_drain_3
timestamp 1667912669
transform 1 0 550 0 1 1100
box -15 0 575 575
use nmos_source  nmos_source_0
timestamp 1667912374
transform 1 0 0 0 1 0
box 0 0 557 557
use nmos_source  nmos_source_1
timestamp 1667912374
transform 1 0 550 0 1 550
box 0 0 557 557
use nmos_source  nmos_source_2
timestamp 1667912374
transform 1 0 0 0 1 1100
box 0 0 557 557
use nmos_source  nmos_source_3
timestamp 1667912374
transform 1 0 1100 0 1 0
box 0 0 557 557
use nmos_source  nmos_source_4
timestamp 1667912374
transform 1 0 1100 0 1 1100
box 0 0 557 557
<< end >>
