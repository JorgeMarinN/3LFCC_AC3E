magic
tech sky130A
timestamp 1667697191
<< metal4 >>
rect 0 30559 17840 30579
rect 0 27339 20 30559
rect 3240 30528 17840 30559
rect 3240 27370 14631 30528
rect 17789 27370 17840 30528
rect 3240 27339 17840 27370
rect 0 27319 17840 27339
<< via4 >>
rect 20 27339 3240 30559
rect 14631 27370 17789 30528
<< metal5 >>
rect 0 41900 50020 45160
rect 4860 37040 45160 40300
rect 0 30559 3260 30579
rect 0 27339 20 30559
rect 3240 27339 3260 30559
rect 0 27319 3260 27339
rect 4860 3260 8120 37040
rect 9720 32179 40300 35440
rect 9720 8120 12980 32179
rect 14580 30528 17840 30579
rect 14580 27370 14631 30528
rect 17789 27370 17840 30528
rect 14580 12980 17840 27370
rect 37039 12980 40300 32179
rect 14580 9720 40300 12980
rect 41900 8120 45160 37040
rect 9720 4860 45160 8120
rect 46760 3260 50020 41900
rect 4860 0 50020 3260
<< end >>
