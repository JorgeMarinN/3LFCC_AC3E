magic
tech sky130A
timestamp 1666566871
<< checkpaint >>
rect -1966 -1966 139166 209966
<< metal1 >>
rect 5050 41645 136600 41650
rect 5050 41555 5055 41645
rect 5145 41555 136600 41645
rect 5050 41550 136600 41555
rect 56750 41495 136800 41500
rect 56750 41405 56755 41495
rect 56845 41405 136800 41495
rect 56750 41400 136800 41405
rect 65750 41345 137000 41350
rect 65750 41255 65755 41345
rect 65845 41255 137000 41345
rect 65750 41250 137000 41255
rect 130950 41195 137200 41200
rect 130950 41105 130955 41195
rect 131045 41105 137200 41195
rect 130950 41100 137200 41105
rect 1000 41045 137200 41050
rect 1000 40855 4897 41045
rect 4930 40855 56597 41045
rect 56630 40855 65597 41045
rect 65630 40855 130797 41045
rect 130830 40855 137200 41045
rect 1000 40850 137200 40855
rect 1000 40795 137200 40800
rect 1000 40605 5335 40795
rect 5425 40605 57035 40795
rect 57125 40605 66035 40795
rect 66125 40605 131235 40795
rect 131325 40605 137200 40795
rect 1000 40600 137200 40605
rect 1000 37995 1500 40600
rect 2000 40350 137200 40550
rect 1000 37505 1005 37995
rect 1495 37505 1500 37995
rect 1000 37500 1500 37505
rect 135500 37995 136000 40350
rect 135500 37505 135505 37995
rect 135995 37505 136000 37995
rect 135500 37500 136000 37505
<< via1 >>
rect 5055 41555 5145 41645
rect 56755 41405 56845 41495
rect 65755 41255 65845 41345
rect 130955 41105 131045 41195
rect 4897 40855 4930 41045
rect 56597 40855 56630 41045
rect 65597 40855 65630 41045
rect 130797 40855 130830 41045
rect 5335 40605 5425 40795
rect 57035 40605 57125 40795
rect 66035 40605 66125 40795
rect 131235 40605 131325 40795
rect 4897 39906 4930 40136
rect 5335 39806 5425 40096
rect 56597 39906 56630 40136
rect 57035 39806 57125 40096
rect 65597 39906 65630 40136
rect 66035 39806 66125 40096
rect 130797 39906 130830 40136
rect 131235 39806 131325 40096
rect 1005 37505 1495 37995
rect 135505 37505 135995 37995
<< metal2 >>
rect 5050 41645 5150 41650
rect 5050 41555 5055 41645
rect 5145 41555 5150 41645
rect 4892 41045 4935 41050
rect 4892 40855 4897 41045
rect 4930 40855 4935 41045
rect 4892 40136 4935 40855
rect 5050 40266 5150 41555
rect 56750 41495 56850 41500
rect 56750 41405 56755 41495
rect 56845 41405 56850 41495
rect 56592 41045 56635 41050
rect 56592 40855 56597 41045
rect 56630 40855 56635 41045
rect 5330 40795 5430 40800
rect 5330 40605 5335 40795
rect 5425 40605 5430 40795
rect 4892 39906 4897 40136
rect 4930 39906 4935 40136
rect 4892 39901 4935 39906
rect 5330 40096 5430 40605
rect 5330 39806 5335 40096
rect 5425 39806 5430 40096
rect 56592 40136 56635 40855
rect 56750 40266 56850 41405
rect 65750 41345 65850 41350
rect 65750 41255 65755 41345
rect 65845 41255 65850 41345
rect 65592 41045 65635 41050
rect 65592 40855 65597 41045
rect 65630 40855 65635 41045
rect 57030 40795 57130 40800
rect 57030 40605 57035 40795
rect 57125 40605 57130 40795
rect 56592 39906 56597 40136
rect 56630 39906 56635 40136
rect 56592 39901 56635 39906
rect 57030 40096 57130 40605
rect 5330 39801 5430 39806
rect 57030 39806 57035 40096
rect 57125 39806 57130 40096
rect 65592 40136 65635 40855
rect 65750 40266 65850 41255
rect 130950 41195 131050 41200
rect 130950 41105 130955 41195
rect 131045 41105 131050 41195
rect 130792 41045 130835 41050
rect 130792 40855 130797 41045
rect 130830 40855 130835 41045
rect 66030 40795 66130 40800
rect 66030 40605 66035 40795
rect 66125 40605 66130 40795
rect 65592 39906 65597 40136
rect 65630 39906 65635 40136
rect 65592 39901 65635 39906
rect 66030 40096 66130 40605
rect 57030 39801 57130 39806
rect 66030 39806 66035 40096
rect 66125 39806 66130 40096
rect 130792 40136 130835 40855
rect 130950 40266 131050 41105
rect 131230 40795 131330 40800
rect 131230 40605 131235 40795
rect 131325 40605 131330 40795
rect 130792 39906 130797 40136
rect 130830 39906 130835 40136
rect 130792 39901 130835 39906
rect 131230 40096 131330 40605
rect 66030 39801 66130 39806
rect 131230 39806 131235 40096
rect 131325 39806 131330 40096
rect 131230 39801 131330 39806
rect 1000 37995 1500 38000
rect 1000 37505 1005 37995
rect 1495 37505 1500 37995
rect 1000 37500 1500 37505
rect 135500 37995 136000 38000
rect 135500 37505 135505 37995
rect 135995 37505 136000 37995
rect 135500 37500 136000 37505
rect 5347 34185 5647 37451
rect 5347 33515 5362 34185
rect 5632 33515 5647 34185
rect 5347 33500 5647 33515
rect 57047 34185 57347 37451
rect 57047 33515 57062 34185
rect 57332 33515 57347 34185
rect 57047 33500 57347 33515
rect 66047 34185 66347 37451
rect 66047 33515 66062 34185
rect 66332 33515 66347 34185
rect 66047 33500 66347 33515
rect 131247 34185 131547 37451
rect 131247 33515 131262 34185
rect 131532 33515 131547 34185
rect 131247 33500 131547 33515
<< via2 >>
rect 1005 37505 1495 37995
rect 135505 37505 135995 37995
rect 5362 33515 5632 34185
rect 57062 33515 57332 34185
rect 66062 33515 66332 34185
rect 131262 33515 131532 34185
<< metal3 >>
rect 1000 37995 1500 38000
rect 1000 37505 1005 37995
rect 1495 37505 1500 37995
rect 1000 31000 1500 37505
rect 135500 37995 136000 38000
rect 135500 37505 135505 37995
rect 135995 37505 136000 37995
rect 5347 34185 5647 37451
rect 5347 33515 5362 34185
rect 5632 33515 5647 34185
rect 5347 33500 5647 33515
rect 57047 34185 57347 37451
rect 57047 33515 57062 34185
rect 57332 33515 57347 34185
rect 57047 33500 57347 33515
rect 66047 34185 66347 37451
rect 66047 33515 66062 34185
rect 66332 33515 66347 34185
rect 66047 33500 66347 33515
rect 131247 34185 131547 37451
rect 131247 33515 131262 34185
rect 131532 33515 131547 34185
rect 131247 33500 131547 33515
rect 135500 31000 136000 37505
<< via3 >>
rect 5362 33515 5632 34185
rect 57062 33515 57332 34185
rect 66062 33515 66332 34185
rect 131262 33515 131532 34185
<< metal4 >>
rect 5347 34185 5647 37451
rect 5347 33515 5362 34185
rect 5632 33515 5647 34185
rect 5347 33500 5647 33515
rect 57047 34185 57347 37451
rect 57047 33515 57062 34185
rect 57332 33515 57347 34185
rect 57047 33500 57347 33515
rect 66047 34185 66347 37451
rect 66047 33515 66062 34185
rect 66332 33515 66347 34185
rect 66047 33500 66347 33515
rect 131247 34185 131547 37451
rect 131247 33515 131262 34185
rect 131532 33515 131547 34185
rect 131247 33500 131547 33515
<< via4 >>
rect 5362 33515 5632 34185
rect 57062 33515 57332 34185
rect 66062 33515 66332 34185
rect 131262 33515 131532 34185
<< metal5 >>
rect 5347 34185 5647 37451
rect 5347 33515 5362 34185
rect 5632 33515 5647 34185
rect 5347 33500 5647 33515
rect 57047 34185 57347 37451
rect 57047 33515 57062 34185
rect 57332 33515 57347 34185
rect 57047 33500 57347 33515
rect 66047 34185 66347 37451
rect 66047 33515 66062 34185
rect 66332 33515 66347 34185
rect 66047 33500 66347 33515
rect 131247 34185 131547 37451
rect 131247 33515 131262 34185
rect 131532 33515 131547 34185
rect 131247 33500 131547 33515
use converter  converter_0
timestamp 1666362992
transform 1 0 0 0 1 0
box 0 0 137200 208000
use level_shifter  level_shifter_0
timestamp 1666543010
transform 0 1 129200 -1 0 40426
box 0 0 3025 4468
use level_shifter  level_shifter_1
timestamp 1666543010
transform 0 1 64000 -1 0 40426
box 0 0 3025 4468
use level_shifter  level_shifter_2
timestamp 1666543010
transform 0 1 55000 -1 0 40426
box 0 0 3025 4468
use level_shifter  level_shifter_3
timestamp 1666543010
transform 0 1 3300 -1 0 40426
box 0 0 3025 4468
<< labels >>
rlabel metal1 137000 40850 137200 41050 7 VDD
rlabel metal1 137100 41100 137200 41200 7 D1
rlabel metal1 136900 41250 137000 41350 7 D2
rlabel metal1 136700 41400 136800 41500 7 D3
rlabel metal1 136500 41550 136600 41650 7 D1
<< end >>
