magic
tech sky130A
timestamp 1667571418
<< metal1 >>
rect 14280 351080 44280 351100
rect 14280 341120 14300 351080
rect 44260 341120 44280 351080
rect 14280 341100 44280 341120
rect 64280 351080 94280 351100
rect 64280 341120 64300 351080
rect 94260 341120 94280 351080
rect 64280 341100 94280 341120
rect 114280 351080 144280 351100
rect 114280 341120 114300 351080
rect 144260 341120 144280 351080
rect 114280 341100 144280 341120
rect 164280 351080 194280 351100
rect 164280 341120 164300 351080
rect 194260 341120 194280 351080
rect 164280 341100 194280 341120
rect 214280 351080 244280 351100
rect 214280 341120 214300 351080
rect 244260 341120 244280 351080
rect 214280 341100 244280 341120
rect 1500 293145 8000 293150
rect 1500 292855 1505 293145
rect 1795 292855 8000 293145
rect 1500 292850 8000 292855
rect 283000 293145 290500 293150
rect 283000 292855 290205 293145
rect 290495 292855 290500 293145
rect 283000 292850 290500 292855
rect 283000 292795 291100 292800
rect 283000 292555 290855 292795
rect 291095 292555 291100 292795
rect 283000 292550 291100 292555
rect 900 292495 8000 292500
rect 900 292405 905 292495
rect 995 292405 8000 292495
rect 900 292400 8000 292405
rect 283000 292495 291100 292500
rect 283000 292405 291005 292495
rect 291095 292405 291100 292495
rect 283000 292400 291100 292405
rect 1050 292345 8000 292350
rect 1050 292255 1055 292345
rect 1145 292255 8000 292345
rect 1050 292250 8000 292255
rect 283000 292345 290950 292350
rect 283000 292255 290855 292345
rect 290945 292255 290950 292345
rect 283000 292250 290950 292255
rect 1200 292195 8000 292200
rect 1200 292105 1205 292195
rect 1295 292105 8000 292195
rect 1200 292100 8000 292105
rect 283000 292195 290800 292200
rect 283000 292105 290705 292195
rect 290795 292105 290800 292195
rect 283000 292100 290800 292105
rect 1350 292045 8000 292050
rect 1350 291955 1355 292045
rect 1445 291955 8000 292045
rect 1350 291950 8000 291955
rect 283000 292045 290650 292050
rect 283000 291955 290555 292045
rect 290645 291955 290650 292045
rect 283000 291950 290650 291955
<< via1 >>
rect 14300 341120 44260 351080
rect 64300 341120 94260 351080
rect 114300 341120 144260 351080
rect 164300 341120 194260 351080
rect 214300 341120 244260 351080
rect 1505 292855 1795 293145
rect 290205 292855 290495 293145
rect 290855 292555 291095 292795
rect 905 292405 995 292495
rect 291005 292405 291095 292495
rect 1055 292255 1145 292345
rect 290855 292255 290945 292345
rect 1205 292105 1295 292195
rect 290705 292105 290795 292195
rect 1355 291955 1445 292045
rect 290555 291955 290645 292045
<< metal2 >>
rect 14280 351080 44280 351100
rect 14280 341120 14300 351080
rect 44260 341120 44280 351080
rect 14280 341100 44280 341120
rect 64280 351080 94280 351100
rect 64280 341120 64300 351080
rect 94260 341120 94280 351080
rect 64280 341100 94280 341120
rect 114280 351080 144280 351100
rect 114280 341120 114300 351080
rect 144260 341120 144280 351080
rect 114280 341100 144280 341120
rect 164280 351080 194280 351100
rect 164280 341120 164300 351080
rect 194260 341120 194280 351080
rect 164280 341100 194280 341120
rect 214280 351080 244280 351100
rect 214280 341120 214300 351080
rect 244260 341120 244280 351080
rect 214280 341100 244280 341120
rect 290850 322287 291100 322300
rect 290850 314897 290855 322287
rect 291095 314897 291100 322287
rect 1500 293145 1800 293150
rect 1500 292855 1505 293145
rect 1795 292855 1800 293145
rect 900 292495 1000 292500
rect 900 292405 905 292495
rect 995 292405 1000 292495
rect 900 124495 1000 292405
rect 1050 292345 1150 292350
rect 1050 292255 1055 292345
rect 1145 292255 1150 292345
rect 1050 146045 1150 292255
rect 1200 292195 1300 292200
rect 1200 292105 1205 292195
rect 1295 292105 1300 292195
rect 1200 167595 1300 292105
rect 1350 292045 1450 292050
rect 1350 291955 1355 292045
rect 1445 291955 1450 292045
rect 1350 189195 1450 291955
rect 1350 189105 1355 189195
rect 1445 189105 1450 189195
rect 1350 189100 1450 189105
rect 1200 167505 1205 167595
rect 1295 167505 1300 167595
rect 1200 167500 1300 167505
rect 1050 145955 1055 146045
rect 1145 145955 1150 146045
rect 1050 145950 1150 145955
rect 900 124405 905 124495
rect 995 124405 1000 124495
rect 900 124400 1000 124405
rect 1500 109839 1800 292855
rect 290200 293145 290500 293150
rect 290200 292855 290205 293145
rect 290495 292855 290500 293145
rect 290200 120010 290500 292855
rect 290850 292795 291100 314897
rect 290850 292555 290855 292795
rect 291095 292555 291100 292795
rect 290850 292550 291100 292555
rect 291000 292495 291100 292500
rect 291000 292405 291005 292495
rect 291095 292405 291100 292495
rect 290850 292345 290950 292350
rect 290850 292255 290855 292345
rect 290945 292255 290950 292345
rect 290700 292195 290800 292200
rect 290700 292105 290705 292195
rect 290795 292105 290800 292195
rect 290550 292045 290650 292050
rect 290550 291955 290555 292045
rect 290645 291955 290650 292045
rect 290550 204495 290650 291955
rect 290550 204405 290555 204495
rect 290645 204405 290650 204495
rect 290550 204400 290650 204405
rect 290700 181295 290800 292105
rect 290700 181205 290705 181295
rect 290795 181205 290800 181295
rect 290700 181200 290800 181205
rect 290850 158695 290950 292255
rect 290850 158605 290855 158695
rect 290945 158605 290950 158695
rect 290850 158600 290950 158605
rect 291000 136495 291100 292405
rect 291000 136405 291005 136495
rect 291095 136405 291100 136495
rect 291000 136400 291100 136405
rect 290200 112620 290205 120010
rect 290495 112620 290500 120010
rect 290200 112600 290500 112620
rect 1500 102449 1505 109839
rect 1795 102449 1800 109839
rect 1500 102400 1800 102449
<< via2 >>
rect 14300 341120 44260 351080
rect 64300 341120 94260 351080
rect 114300 341120 144260 351080
rect 164300 341120 194260 351080
rect 214300 341120 244260 351080
rect 290855 314897 291095 322287
rect 1355 189105 1445 189195
rect 1205 167505 1295 167595
rect 1055 145955 1145 146045
rect 905 124405 995 124495
rect 290555 204405 290645 204495
rect 290705 181205 290795 181295
rect 290855 158605 290945 158695
rect 291005 136405 291095 136495
rect 290205 112620 290495 120010
rect 1505 102449 1795 109839
<< metal3 >>
rect 8000 351000 11000 351200
rect 34000 351100 36600 351150
rect 73000 351100 85300 351150
rect 87947 351100 90500 351150
rect 7000 350000 11000 351000
rect 14280 351080 44280 351100
rect 800 340000 6500 342000
rect 5500 245000 6500 340000
rect 7000 289000 8000 350000
rect 14280 341120 14300 351080
rect 44260 341120 44280 351080
rect 14280 341100 44280 341120
rect 64280 351080 94280 351100
rect 64280 341120 64300 351080
rect 94260 341120 94280 351080
rect 108647 351000 111147 351150
rect 113797 351100 119000 351150
rect 113797 351080 144280 351100
rect 113797 351000 114300 351080
rect 108647 348000 114300 351000
rect 108647 347800 111600 348000
rect 114280 347800 114300 348000
rect 108647 344800 114300 347800
rect 64280 341100 94280 341120
rect 114280 341120 114300 344800
rect 144260 341120 144280 351080
rect 159497 351000 161997 351150
rect 164647 351100 181000 351150
rect 164280 351080 194280 351100
rect 164280 351000 164300 351080
rect 159497 348000 164300 351000
rect 159497 347800 162400 348000
rect 164280 347800 164300 348000
rect 159497 344800 164300 347800
rect 114280 341100 144280 341120
rect 164280 341120 164300 344800
rect 194260 341120 194280 351080
rect 164280 341100 194280 341120
rect 214280 351080 244280 351100
rect 214280 341120 214300 351080
rect 244260 341120 244280 351080
rect 214280 341100 244280 341120
rect 284000 289000 285000 351200
rect 285500 339000 291200 341000
rect 285500 245000 286500 339000
rect 290850 322287 291500 322292
rect 290850 314897 290855 322287
rect 291095 314897 291500 322287
rect 290850 314892 291500 314897
rect 5500 244000 8000 245000
rect 283000 244000 286500 245000
rect 290550 204495 292000 204700
rect 290550 204405 290555 204495
rect 290645 204405 292000 204495
rect 290550 204200 292000 204405
rect 0 189195 1450 189400
rect 0 189105 1355 189195
rect 1445 189105 1450 189195
rect 0 188900 1450 189105
rect 290700 181295 292000 181500
rect 290700 181205 290705 181295
rect 290795 181205 292000 181295
rect 290700 181000 292000 181205
rect 0 167595 1300 167800
rect 0 167505 1205 167595
rect 1295 167505 1300 167595
rect 0 167300 1300 167505
rect 290850 158695 292000 158900
rect 290850 158605 290855 158695
rect 290945 158605 292000 158695
rect 290850 158400 292000 158605
rect 0 146045 1150 146200
rect 0 145955 1055 146045
rect 1145 145955 1150 146045
rect 0 145700 1150 145955
rect 291000 136495 292000 136700
rect 291000 136405 291005 136495
rect 291095 136405 292000 136495
rect 291000 136200 292000 136405
rect 0 124495 1000 124700
rect 0 124405 905 124495
rect 995 124405 1000 124495
rect 0 124200 1000 124405
rect 290200 120010 291500 120015
rect 290200 112620 290205 120010
rect 290495 112620 291500 120010
rect 290200 112615 291500 112620
rect 500 109839 1800 109844
rect 500 102449 1505 109839
rect 1795 102449 1800 109839
rect 500 102444 1800 102449
<< rmetal3 >>
rect 60000 351100 62600 351150
rect 206600 351100 209200 351150
rect 232600 351100 235200 351150
<< via3 >>
rect 14300 341120 44260 351080
rect 64300 341120 94260 351080
rect 114300 341120 144260 351080
rect 164300 341120 194260 351080
rect 214300 341120 244260 351080
<< metal4 >>
rect 73000 351100 85300 351150
rect 87947 351100 90500 351150
rect 14280 351080 44280 351100
rect 14280 341120 14300 351080
rect 44260 341120 44280 351080
rect 14280 341100 44280 341120
rect 64280 351080 94280 351100
rect 64280 341120 64300 351080
rect 94260 341120 94280 351080
rect 108647 351000 111147 351150
rect 113797 351100 119000 351150
rect 113797 351080 144280 351100
rect 113797 351000 114300 351080
rect 108647 348000 114300 351000
rect 108647 347800 111600 348000
rect 114280 347800 114300 348000
rect 108647 344800 114300 347800
rect 64280 341100 94280 341120
rect 114280 341120 114300 344800
rect 144260 341120 144280 351080
rect 159497 351000 161997 351150
rect 164647 351100 181000 351150
rect 164280 351080 194280 351100
rect 164280 351000 164300 351080
rect 159497 348000 164300 351000
rect 159497 347800 162400 348000
rect 164280 347800 164300 348000
rect 159497 344800 164300 347800
rect 114280 341100 144280 341120
rect 164280 341120 164300 344800
rect 194260 341120 194280 351080
rect 164280 341100 194280 341120
rect 214280 351080 244280 351100
rect 214280 341120 214300 351080
rect 244260 341120 244280 351080
rect 214280 341100 244280 341120
<< via4 >>
rect 14300 341120 44260 351080
rect 64300 341120 94260 351080
rect 114300 341120 144260 351080
rect 164300 341120 194260 351080
rect 214300 341120 244260 351080
<< metal5 >>
rect 73000 351100 85300 351150
rect 87947 351100 90500 351150
rect 14280 351080 44280 351100
rect 14280 341120 14300 351080
rect 44260 341120 44280 351080
rect 14280 341100 44280 341120
rect 64280 351080 94280 351100
rect 64280 341120 64300 351080
rect 94260 341120 94280 351080
rect 108647 351000 111147 351150
rect 113797 351100 119000 351150
rect 113797 351080 144280 351100
rect 113797 351000 114300 351080
rect 108647 348000 114300 351000
rect 108647 347800 111600 348000
rect 114280 347800 114300 348000
rect 108647 344800 114300 347800
rect 64280 341100 94280 341120
rect 114280 341120 114300 344800
rect 144260 341120 144280 351080
rect 159497 351000 161997 351150
rect 164647 351100 181000 351150
rect 164280 351080 194280 351100
rect 164280 351000 164300 351080
rect 159497 348000 164300 351000
rect 159497 347800 162400 348000
rect 164280 347800 164300 348000
rect 159497 344800 164300 347800
rect 114280 341100 144280 341120
rect 164280 341120 164300 344800
rect 194260 341120 194280 351080
rect 164280 341100 194280 341120
rect 214280 351080 244280 351100
rect 214280 341120 214300 351080
rect 244260 341120 244280 351080
rect 214280 341100 244280 341120
<< glass >>
rect 14300 341120 44260 351080
rect 64300 341120 94260 351080
rect 114300 341120 144260 351080
rect 164300 341120 194260 351080
rect 214300 341120 244260 351080
rect 7460 268230 17420 290200
rect 274580 268230 284540 290200
rect 7460 223570 17420 245540
rect 274580 223570 284540 245540
<< comment >>
rect 0 0 1000 1000
use interleaved  interleaved_0
timestamp 1667562098
transform 1 0 146000 0 1 125500
box -138560 -1000 138560 225600
<< labels >>
rlabel metal3 0 124200 1000 124700 7 D1
rlabel metal3 0 145700 1150 146200 7 D2
rlabel metal3 0 167300 1300 167800 7 D3
rlabel metal3 0 188900 1450 189400 7 D4
rlabel metal3 291000 136200 292000 136700 3 D5
rlabel metal3 290850 158400 292000 158900 3 D6
rlabel metal3 290700 181000 292000 181500 3 D7
rlabel metal3 290550 204200 292000 204700 3 D8
rlabel metal3 500 102444 1800 109844 7 VLS1
rlabel metal3 290200 112615 291500 120015 3 VLS2
rlabel metal3 290850 314892 291500 322292 3 VDD
rlabel metal3 8000 350000 11000 351200 3 FC1_1
rlabel metal3 800 340000 6500 342000 1 FC1_2
rlabel metal3 284000 348000 285000 351000 3 FC2_1
rlabel metal3 285500 339000 291200 341000 1 FC2_2
<< end >>
