magic
tech sky130A
magscale 1 2
timestamp 1668450766
<< pwell >>
rect -3166 -3706 3166 3706
<< psubdiff >>
rect -3130 3636 -3034 3670
rect 3034 3636 3130 3670
rect -3130 3574 -3096 3636
rect 3096 3574 3130 3636
rect -3130 -3636 -3096 -3574
rect 3096 -3636 3130 -3574
rect -3130 -3670 -3034 -3636
rect 3034 -3670 3130 -3636
<< psubdiffcont >>
rect -3034 3636 3034 3670
rect -3130 -3574 -3096 3574
rect 3096 -3574 3130 3574
rect -3034 -3670 3034 -3636
<< poly >>
rect -3000 3524 3000 3540
rect -3000 3490 -2984 3524
rect 2984 3490 3000 3524
rect -3000 3110 3000 3490
rect -3000 -3490 3000 -3110
rect -3000 -3524 -2984 -3490
rect 2984 -3524 3000 -3490
rect -3000 -3540 3000 -3524
<< polycont >>
rect -2984 3490 2984 3524
rect -2984 -3524 2984 -3490
<< npolyres >>
rect -3000 -3110 3000 3110
<< locali >>
rect -3130 3636 -3034 3670
rect 3034 3636 3130 3670
rect -3130 3574 -3096 3636
rect 3096 3574 3130 3636
rect -3000 3490 -2984 3524
rect 2984 3490 3000 3524
rect -3000 -3524 -2984 -3490
rect 2984 -3524 3000 -3490
rect -3130 -3636 -3096 -3574
rect 3096 -3636 3130 -3574
rect -3130 -3670 -3034 -3636
rect 3034 -3670 3130 -3636
<< viali >>
rect -2984 3490 2984 3524
rect -2984 3127 2984 3490
rect -2984 -3490 2984 -3127
rect -2984 -3524 2984 -3490
<< metal1 >>
rect -2996 3524 2996 3530
rect -2996 3127 -2984 3524
rect 2984 3127 2996 3524
rect -2996 3121 2996 3127
rect -2996 -3127 2996 -3121
rect -2996 -3524 -2984 -3127
rect 2984 -3524 2996 -3127
rect -2996 -3530 2996 -3524
<< properties >>
string FIXED_BBOX -3113 -3653 3113 3653
string gencell sky130_fd_pr__res_generic_po
string library sky130
string parameters w 30 l 31.1 m 1 nx 1 wmin 0.330 lmin 1.650 rho 48.2 val 49.967 dummy 0 dw 0.0 term 0.0 sterm 0.0 caplen 0.4 snake 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 roverlap 0 endcov 100 full_metal 1 hv_guard 0 n_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
